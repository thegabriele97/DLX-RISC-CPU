
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ISSUE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ISSUE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA_IN : in 
         std_logic_vector (31 downto 0);  DRAM_DATA_OUT : out std_logic_vector 
         (31 downto 0);  DATA_SIZE : out std_logic_vector (1 downto 0);  
         DRAMRF_ADDRESS : out std_logic_vector (31 downto 0);  DRAMRF_ISSUE, 
         DRAMRF_READNOTWRITE : out std_logic;  DRAMRF_READY : in std_logic;  
         DRAMRF_DATA_IN : in std_logic_vector (31 downto 0);  DRAMRF_DATA_OUT :
         out std_logic_vector (31 downto 0);  DATA_SIZE_RF : out 
         std_logic_vector (1 downto 0);  OPCODE : out std_logic_vector (5 
         downto 0);  RS1, RS2, WS1 : out std_logic_vector (4 downto 0);  IRO, 
         PCO : out std_logic_vector (31 downto 0);  DIR_EN : out std_logic);

end DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port, 
      DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, 
      DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, 
      DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, 
      DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, 
      DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, 
      DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, 
      DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, 
      DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, 
      DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, 
      DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, 
      DRAM_ADDRESS_0_port, DRAM_ISSUE_port, DRAM_DATA_OUT_31_port, 
      DRAM_DATA_OUT_30_port, DRAM_DATA_OUT_29_port, DRAM_DATA_OUT_28_port, 
      DRAM_DATA_OUT_27_port, DRAM_DATA_OUT_26_port, DRAM_DATA_OUT_25_port, 
      DRAM_DATA_OUT_24_port, DRAM_DATA_OUT_23_port, DRAM_DATA_OUT_22_port, 
      DRAM_DATA_OUT_21_port, DRAM_DATA_OUT_20_port, DRAM_DATA_OUT_19_port, 
      DRAM_DATA_OUT_18_port, DRAM_DATA_OUT_17_port, DRAM_DATA_OUT_16_port, 
      DRAM_DATA_OUT_15_port, DRAM_DATA_OUT_14_port, DRAM_DATA_OUT_13_port, 
      DRAM_DATA_OUT_12_port, DRAM_DATA_OUT_11_port, DRAM_DATA_OUT_10_port, 
      DRAM_DATA_OUT_9_port, DRAM_DATA_OUT_8_port, DRAM_DATA_OUT_7_port, 
      DRAM_DATA_OUT_6_port, DRAM_DATA_OUT_5_port, DRAM_DATA_OUT_4_port, 
      DRAM_DATA_OUT_3_port, DRAM_DATA_OUT_2_port, DRAM_DATA_OUT_1_port, 
      DRAM_DATA_OUT_0_port, DATA_SIZE_1_port, DATA_SIZE_0_port, 
      DRAMRF_READNOTWRITE_port, OPCODE_5_port, OPCODE_4_port, OPCODE_3_port, 
      OPCODE_2_port, OPCODE_1_port, OPCODE_0_port, IRO_25_port, IRO_24_port, 
      IRO_23_port, IRO_22_port, IRO_21_port, IRO_20_port, IRO_19_port, 
      IRO_18_port, IRO_17_port, IRO_16_port, IRO_15_port, IRO_14_port, 
      IRO_13_port, IRO_12_port, IRO_11_port, IRO_10_port, IRO_9_port, 
      IRO_8_port, IRO_7_port, IRO_6_port, IRO_5_port, IRO_4_port, IRO_3_port, 
      IRO_2_port, IRO_1_port, IRO_0_port, i_RF_MEM_WM, i_EN2, i_S1, i_S2, 
      i_ALU_OP_4_port, i_ALU_OP_3_port, i_ALU_OP_1_port, i_ALU_OP_0_port, 
      i_SEL_ALU_SETCMP, i_SEL_LGET_1_port, i_SEL_LGET_0_port, i_DATAMEM_RM, 
      i_UNSIG_SIGN_N, i_EN3, i_ADD_WB_4_port, i_ADD_WB_3_port, i_ADD_WB_2_port,
      i_ADD_WB_1_port, i_ADD_WB_0_port, CU_I_n157, CU_I_n156, CU_I_n155, 
      CU_I_n154, CU_I_n153, CU_I_n152, CU_I_n151, CU_I_n148, CU_I_n147, 
      CU_I_n146, CU_I_n145, CU_I_n144, CU_I_n142, CU_I_n141, CU_I_n140, 
      CU_I_n139, CU_I_n138, CU_I_n137, CU_I_n136, CU_I_n135, CU_I_n134, 
      CU_I_n133, CU_I_n132, CU_I_n131, CU_I_n130, CU_I_n129, CU_I_n128, 
      CU_I_n127, CU_I_n126, CU_I_n118, CU_I_n114, CU_I_n113, CU_I_n112, 
      CU_I_n111, CU_I_n110, CU_I_n109, CU_I_n108, CU_I_n107, CU_I_n105, 
      CU_I_n104, CU_I_n103, CU_I_n102, CU_I_n101, CU_I_n99, CU_I_n98, CU_I_n71,
      CU_I_n58, CU_I_n22, CU_I_N50, CU_I_N49, DataPath_n3, DataPath_n2, 
      DataPath_i_PIPLIN_WRB2_0_port, DataPath_i_PIPLIN_WRB2_1_port, 
      DataPath_i_PIPLIN_WRB2_2_port, DataPath_i_PIPLIN_WRB2_3_port, 
      DataPath_i_PIPLIN_WRB2_4_port, DataPath_i_PIPLIN_WRB1_0_port, 
      DataPath_i_PIPLIN_WRB1_1_port, DataPath_i_PIPLIN_WRB1_2_port, 
      DataPath_i_PIPLIN_WRB1_3_port, DataPath_i_PIPLIN_WRB1_4_port, 
      DataPath_i_REG_MEM_ALUOUT_0_port, DataPath_i_REG_MEM_ALUOUT_1_port, 
      DataPath_i_REG_MEM_ALUOUT_2_port, DataPath_i_REG_MEM_ALUOUT_3_port, 
      DataPath_i_REG_MEM_ALUOUT_4_port, DataPath_i_REG_MEM_ALUOUT_5_port, 
      DataPath_i_REG_MEM_ALUOUT_6_port, DataPath_i_REG_MEM_ALUOUT_7_port, 
      DataPath_i_REG_MEM_ALUOUT_8_port, DataPath_i_REG_MEM_ALUOUT_9_port, 
      DataPath_i_REG_MEM_ALUOUT_10_port, DataPath_i_REG_MEM_ALUOUT_11_port, 
      DataPath_i_REG_MEM_ALUOUT_12_port, DataPath_i_REG_MEM_ALUOUT_13_port, 
      DataPath_i_REG_MEM_ALUOUT_14_port, DataPath_i_REG_MEM_ALUOUT_15_port, 
      DataPath_i_REG_MEM_ALUOUT_16_port, DataPath_i_REG_MEM_ALUOUT_17_port, 
      DataPath_i_REG_MEM_ALUOUT_18_port, DataPath_i_REG_MEM_ALUOUT_19_port, 
      DataPath_i_REG_MEM_ALUOUT_20_port, DataPath_i_REG_MEM_ALUOUT_21_port, 
      DataPath_i_REG_MEM_ALUOUT_22_port, DataPath_i_REG_MEM_ALUOUT_23_port, 
      DataPath_i_REG_MEM_ALUOUT_24_port, DataPath_i_REG_MEM_ALUOUT_25_port, 
      DataPath_i_REG_MEM_ALUOUT_26_port, DataPath_i_REG_MEM_ALUOUT_27_port, 
      DataPath_i_REG_MEM_ALUOUT_28_port, DataPath_i_REG_MEM_ALUOUT_29_port, 
      DataPath_i_REG_MEM_ALUOUT_30_port, DataPath_i_REG_MEM_ALUOUT_31_port, 
      DataPath_i_REG_LDSTR_OUT_0_port, DataPath_i_REG_LDSTR_OUT_1_port, 
      DataPath_i_REG_LDSTR_OUT_2_port, DataPath_i_REG_LDSTR_OUT_3_port, 
      DataPath_i_REG_LDSTR_OUT_4_port, DataPath_i_REG_LDSTR_OUT_5_port, 
      DataPath_i_REG_LDSTR_OUT_6_port, DataPath_i_REG_LDSTR_OUT_7_port, 
      DataPath_i_REG_LDSTR_OUT_8_port, DataPath_i_REG_LDSTR_OUT_9_port, 
      DataPath_i_REG_LDSTR_OUT_10_port, DataPath_i_REG_LDSTR_OUT_11_port, 
      DataPath_i_REG_LDSTR_OUT_12_port, DataPath_i_REG_LDSTR_OUT_13_port, 
      DataPath_i_REG_LDSTR_OUT_14_port, DataPath_i_REG_LDSTR_OUT_15_port, 
      DataPath_i_REG_LDSTR_OUT_16_port, DataPath_i_REG_LDSTR_OUT_17_port, 
      DataPath_i_REG_LDSTR_OUT_18_port, DataPath_i_REG_LDSTR_OUT_19_port, 
      DataPath_i_REG_LDSTR_OUT_20_port, DataPath_i_REG_LDSTR_OUT_21_port, 
      DataPath_i_REG_LDSTR_OUT_22_port, DataPath_i_REG_LDSTR_OUT_23_port, 
      DataPath_i_REG_LDSTR_OUT_24_port, DataPath_i_REG_LDSTR_OUT_25_port, 
      DataPath_i_REG_LDSTR_OUT_26_port, DataPath_i_REG_LDSTR_OUT_27_port, 
      DataPath_i_REG_LDSTR_OUT_28_port, DataPath_i_REG_LDSTR_OUT_29_port, 
      DataPath_i_REG_LDSTR_OUT_30_port, DataPath_i_REG_LDSTR_OUT_31_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_0_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_1_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_2_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_3_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_4_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_5_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_6_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_7_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_8_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_9_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_10_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_11_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_12_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_13_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_14_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_15_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_16_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_17_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_18_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_19_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_20_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_21_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_22_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_23_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_24_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_25_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_26_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_27_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_28_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_29_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_30_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_31_port, 
      DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_0_port, 
      DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_1_port, DataPath_i_ALU_OUT_0_port,
      DataPath_i_ALU_OUT_1_port, DataPath_i_ALU_OUT_2_port, 
      DataPath_i_ALU_OUT_3_port, DataPath_i_ALU_OUT_4_port, 
      DataPath_i_ALU_OUT_5_port, DataPath_i_ALU_OUT_6_port, 
      DataPath_i_ALU_OUT_7_port, DataPath_i_ALU_OUT_8_port, 
      DataPath_i_ALU_OUT_9_port, DataPath_i_ALU_OUT_10_port, 
      DataPath_i_ALU_OUT_11_port, DataPath_i_ALU_OUT_12_port, 
      DataPath_i_ALU_OUT_13_port, DataPath_i_ALU_OUT_14_port, 
      DataPath_i_ALU_OUT_15_port, DataPath_i_ALU_OUT_16_port, 
      DataPath_i_SETCMP_OUT_0_port, DataPath_i_LGET_0_port, 
      DataPath_i_LGET_1_port, DataPath_i_PIPLIN_IN2_0_port, 
      DataPath_i_PIPLIN_IN2_1_port, DataPath_i_PIPLIN_IN2_2_port, 
      DataPath_i_PIPLIN_IN2_3_port, DataPath_i_PIPLIN_IN2_4_port, 
      DataPath_i_PIPLIN_IN2_5_port, DataPath_i_PIPLIN_IN2_6_port, 
      DataPath_i_PIPLIN_IN2_7_port, DataPath_i_PIPLIN_IN2_8_port, 
      DataPath_i_PIPLIN_IN2_9_port, DataPath_i_PIPLIN_IN2_10_port, 
      DataPath_i_PIPLIN_IN2_11_port, DataPath_i_PIPLIN_IN2_12_port, 
      DataPath_i_PIPLIN_IN2_13_port, DataPath_i_PIPLIN_IN2_14_port, 
      DataPath_i_PIPLIN_IN2_15_port, DataPath_i_PIPLIN_IN2_16_port, 
      DataPath_i_PIPLIN_IN2_17_port, DataPath_i_PIPLIN_IN2_18_port, 
      DataPath_i_PIPLIN_IN2_19_port, DataPath_i_PIPLIN_IN2_20_port, 
      DataPath_i_PIPLIN_IN2_21_port, DataPath_i_PIPLIN_IN2_22_port, 
      DataPath_i_PIPLIN_IN2_23_port, DataPath_i_PIPLIN_IN2_24_port, 
      DataPath_i_PIPLIN_IN2_25_port, DataPath_i_PIPLIN_IN2_26_port, 
      DataPath_i_PIPLIN_IN2_27_port, DataPath_i_PIPLIN_IN2_28_port, 
      DataPath_i_PIPLIN_IN2_29_port, DataPath_i_PIPLIN_IN2_30_port, 
      DataPath_i_PIPLIN_IN2_31_port, DataPath_i_PIPLIN_IN1_0_port, 
      DataPath_i_PIPLIN_IN1_1_port, DataPath_i_PIPLIN_IN1_2_port, 
      DataPath_i_PIPLIN_IN1_3_port, DataPath_i_PIPLIN_IN1_4_port, 
      DataPath_i_PIPLIN_IN1_5_port, DataPath_i_PIPLIN_IN1_6_port, 
      DataPath_i_PIPLIN_IN1_7_port, DataPath_i_PIPLIN_IN1_8_port, 
      DataPath_i_PIPLIN_IN1_9_port, DataPath_i_PIPLIN_IN1_10_port, 
      DataPath_i_PIPLIN_IN1_11_port, DataPath_i_PIPLIN_IN1_12_port, 
      DataPath_i_PIPLIN_IN1_13_port, DataPath_i_PIPLIN_IN1_14_port, 
      DataPath_i_PIPLIN_IN1_15_port, DataPath_i_PIPLIN_IN1_16_port, 
      DataPath_i_PIPLIN_IN1_17_port, DataPath_i_PIPLIN_IN1_18_port, 
      DataPath_i_PIPLIN_IN1_19_port, DataPath_i_PIPLIN_IN1_20_port, 
      DataPath_i_PIPLIN_IN1_21_port, DataPath_i_PIPLIN_IN1_22_port, 
      DataPath_i_PIPLIN_IN1_23_port, DataPath_i_PIPLIN_IN1_24_port, 
      DataPath_i_PIPLIN_IN1_25_port, DataPath_i_PIPLIN_IN1_26_port, 
      DataPath_i_PIPLIN_IN1_27_port, DataPath_i_PIPLIN_IN1_28_port, 
      DataPath_i_PIPLIN_IN1_29_port, DataPath_i_PIPLIN_IN1_30_port, 
      DataPath_i_PIPLIN_IN1_31_port, DataPath_i_PIPLIN_B_0_port, 
      DataPath_i_PIPLIN_B_1_port, DataPath_i_PIPLIN_B_2_port, 
      DataPath_i_PIPLIN_B_3_port, DataPath_i_PIPLIN_B_4_port, 
      DataPath_i_PIPLIN_B_5_port, DataPath_i_PIPLIN_B_6_port, 
      DataPath_i_PIPLIN_B_7_port, DataPath_i_PIPLIN_B_8_port, 
      DataPath_i_PIPLIN_B_9_port, DataPath_i_PIPLIN_B_10_port, 
      DataPath_i_PIPLIN_B_11_port, DataPath_i_PIPLIN_B_12_port, 
      DataPath_i_PIPLIN_B_13_port, DataPath_i_PIPLIN_B_14_port, 
      DataPath_i_PIPLIN_B_15_port, DataPath_i_PIPLIN_B_16_port, 
      DataPath_i_PIPLIN_B_17_port, DataPath_i_PIPLIN_B_18_port, 
      DataPath_i_PIPLIN_B_19_port, DataPath_i_PIPLIN_B_20_port, 
      DataPath_i_PIPLIN_B_21_port, DataPath_i_PIPLIN_B_22_port, 
      DataPath_i_PIPLIN_B_23_port, DataPath_i_PIPLIN_B_24_port, 
      DataPath_i_PIPLIN_B_25_port, DataPath_i_PIPLIN_B_26_port, 
      DataPath_i_PIPLIN_B_27_port, DataPath_i_PIPLIN_B_28_port, 
      DataPath_i_PIPLIN_B_29_port, DataPath_i_PIPLIN_B_30_port, 
      DataPath_i_PIPLIN_B_31_port, DataPath_i_PIPLIN_A_0_port, 
      DataPath_i_PIPLIN_A_1_port, DataPath_i_PIPLIN_A_2_port, 
      DataPath_i_PIPLIN_A_3_port, DataPath_i_PIPLIN_A_4_port, 
      DataPath_i_PIPLIN_A_5_port, DataPath_i_PIPLIN_A_6_port, 
      DataPath_i_PIPLIN_A_7_port, DataPath_i_PIPLIN_A_8_port, 
      DataPath_i_PIPLIN_A_9_port, DataPath_i_PIPLIN_A_10_port, 
      DataPath_i_PIPLIN_A_11_port, DataPath_i_PIPLIN_A_12_port, 
      DataPath_i_PIPLIN_A_13_port, DataPath_i_PIPLIN_A_14_port, 
      DataPath_i_PIPLIN_A_15_port, DataPath_i_PIPLIN_A_16_port, 
      DataPath_i_PIPLIN_A_17_port, DataPath_i_PIPLIN_A_18_port, 
      DataPath_i_PIPLIN_A_19_port, DataPath_i_PIPLIN_A_20_port, 
      DataPath_i_PIPLIN_A_21_port, DataPath_i_PIPLIN_A_22_port, 
      DataPath_i_PIPLIN_A_23_port, DataPath_i_PIPLIN_A_24_port, 
      DataPath_i_PIPLIN_A_25_port, DataPath_i_PIPLIN_A_26_port, 
      DataPath_i_PIPLIN_A_27_port, DataPath_i_PIPLIN_A_28_port, 
      DataPath_i_PIPLIN_A_29_port, DataPath_i_PIPLIN_A_30_port, 
      DataPath_i_PIPLIN_A_31_port, DataPath_i_RF_BUS_FROM_RF_CU_0_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_1_port, DataPath_i_RF_BUS_FROM_RF_CU_2_port,
      DataPath_i_RF_BUS_FROM_RF_CU_3_port, DataPath_i_RF_BUS_FROM_RF_CU_4_port,
      DataPath_i_RF_BUS_FROM_RF_CU_5_port, DataPath_i_RF_BUS_FROM_RF_CU_6_port,
      DataPath_i_RF_BUS_FROM_RF_CU_7_port, DataPath_i_RF_BUS_FROM_RF_CU_8_port,
      DataPath_i_RF_BUS_FROM_RF_CU_9_port, DataPath_i_RF_BUS_FROM_RF_CU_10_port
      , DataPath_i_RF_BUS_FROM_RF_CU_11_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_12_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_13_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_14_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_15_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_16_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_17_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_18_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_19_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_20_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_21_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_22_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_23_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_24_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_25_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_26_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_27_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_28_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_29_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_30_port, 
      DataPath_i_RF_BUS_FROM_RF_CU_31_port, DataPath_i_DONE_FILL_EX, 
      DataPath_i_DONE_SPILL_EX, DataPath_i_WF, DataPath_RF_n10, DataPath_RF_n9,
      DataPath_RF_spill_address_0_port, DataPath_RF_spill_address_1_port, 
      DataPath_RF_spill_address_2_port, DataPath_RF_spill_address_3_port, 
      DataPath_RF_spill_address_ext_0_port, 
      DataPath_RF_spill_address_ext_1_port, 
      DataPath_RF_spill_address_ext_2_port, 
      DataPath_RF_spill_address_ext_3_port, 
      DataPath_RF_spill_address_ext_4_port, 
      DataPath_RF_spill_address_ext_5_port, 
      DataPath_RF_spill_address_ext_6_port, 
      DataPath_RF_spill_address_ext_7_port, 
      DataPath_RF_spill_address_ext_8_port, 
      DataPath_RF_spill_address_ext_9_port, 
      DataPath_RF_spill_address_ext_10_port, 
      DataPath_RF_spill_address_ext_11_port, 
      DataPath_RF_spill_address_ext_12_port, 
      DataPath_RF_spill_address_ext_13_port, 
      DataPath_RF_spill_address_ext_14_port, 
      DataPath_RF_spill_address_ext_15_port, 
      DataPath_RF_bus_sel_savedwin_data_0_port, 
      DataPath_RF_bus_sel_savedwin_data_1_port, 
      DataPath_RF_bus_sel_savedwin_data_2_port, 
      DataPath_RF_bus_sel_savedwin_data_3_port, 
      DataPath_RF_bus_sel_savedwin_data_4_port, 
      DataPath_RF_bus_sel_savedwin_data_5_port, 
      DataPath_RF_bus_sel_savedwin_data_6_port, 
      DataPath_RF_bus_sel_savedwin_data_7_port, 
      DataPath_RF_bus_sel_savedwin_data_8_port, 
      DataPath_RF_bus_sel_savedwin_data_9_port, 
      DataPath_RF_bus_sel_savedwin_data_10_port, 
      DataPath_RF_bus_sel_savedwin_data_11_port, 
      DataPath_RF_bus_sel_savedwin_data_12_port, 
      DataPath_RF_bus_sel_savedwin_data_13_port, 
      DataPath_RF_bus_sel_savedwin_data_14_port, 
      DataPath_RF_bus_sel_savedwin_data_15_port, 
      DataPath_RF_bus_sel_savedwin_data_16_port, 
      DataPath_RF_bus_sel_savedwin_data_17_port, 
      DataPath_RF_bus_sel_savedwin_data_18_port, 
      DataPath_RF_bus_sel_savedwin_data_19_port, 
      DataPath_RF_bus_sel_savedwin_data_20_port, 
      DataPath_RF_bus_sel_savedwin_data_21_port, 
      DataPath_RF_bus_sel_savedwin_data_22_port, 
      DataPath_RF_bus_sel_savedwin_data_23_port, 
      DataPath_RF_bus_sel_savedwin_data_24_port, 
      DataPath_RF_bus_sel_savedwin_data_25_port, 
      DataPath_RF_bus_sel_savedwin_data_26_port, 
      DataPath_RF_bus_sel_savedwin_data_27_port, 
      DataPath_RF_bus_sel_savedwin_data_28_port, 
      DataPath_RF_bus_sel_savedwin_data_29_port, 
      DataPath_RF_bus_sel_savedwin_data_30_port, 
      DataPath_RF_bus_sel_savedwin_data_31_port, 
      DataPath_RF_bus_sel_savedwin_data_32_port, 
      DataPath_RF_bus_sel_savedwin_data_33_port, 
      DataPath_RF_bus_sel_savedwin_data_34_port, 
      DataPath_RF_bus_sel_savedwin_data_35_port, 
      DataPath_RF_bus_sel_savedwin_data_36_port, 
      DataPath_RF_bus_sel_savedwin_data_37_port, 
      DataPath_RF_bus_sel_savedwin_data_38_port, 
      DataPath_RF_bus_sel_savedwin_data_39_port, 
      DataPath_RF_bus_sel_savedwin_data_40_port, 
      DataPath_RF_bus_sel_savedwin_data_41_port, 
      DataPath_RF_bus_sel_savedwin_data_42_port, 
      DataPath_RF_bus_sel_savedwin_data_43_port, 
      DataPath_RF_bus_sel_savedwin_data_44_port, 
      DataPath_RF_bus_sel_savedwin_data_45_port, 
      DataPath_RF_bus_sel_savedwin_data_46_port, 
      DataPath_RF_bus_sel_savedwin_data_47_port, 
      DataPath_RF_bus_sel_savedwin_data_48_port, 
      DataPath_RF_bus_sel_savedwin_data_49_port, 
      DataPath_RF_bus_sel_savedwin_data_50_port, 
      DataPath_RF_bus_sel_savedwin_data_51_port, 
      DataPath_RF_bus_sel_savedwin_data_52_port, 
      DataPath_RF_bus_sel_savedwin_data_53_port, 
      DataPath_RF_bus_sel_savedwin_data_54_port, 
      DataPath_RF_bus_sel_savedwin_data_55_port, 
      DataPath_RF_bus_sel_savedwin_data_56_port, 
      DataPath_RF_bus_sel_savedwin_data_57_port, 
      DataPath_RF_bus_sel_savedwin_data_58_port, 
      DataPath_RF_bus_sel_savedwin_data_59_port, 
      DataPath_RF_bus_sel_savedwin_data_60_port, 
      DataPath_RF_bus_sel_savedwin_data_61_port, 
      DataPath_RF_bus_sel_savedwin_data_62_port, 
      DataPath_RF_bus_sel_savedwin_data_63_port, 
      DataPath_RF_bus_sel_savedwin_data_64_port, 
      DataPath_RF_bus_sel_savedwin_data_65_port, 
      DataPath_RF_bus_sel_savedwin_data_66_port, 
      DataPath_RF_bus_sel_savedwin_data_67_port, 
      DataPath_RF_bus_sel_savedwin_data_68_port, 
      DataPath_RF_bus_sel_savedwin_data_69_port, 
      DataPath_RF_bus_sel_savedwin_data_70_port, 
      DataPath_RF_bus_sel_savedwin_data_71_port, 
      DataPath_RF_bus_sel_savedwin_data_72_port, 
      DataPath_RF_bus_sel_savedwin_data_73_port, 
      DataPath_RF_bus_sel_savedwin_data_74_port, 
      DataPath_RF_bus_sel_savedwin_data_75_port, 
      DataPath_RF_bus_sel_savedwin_data_76_port, 
      DataPath_RF_bus_sel_savedwin_data_77_port, 
      DataPath_RF_bus_sel_savedwin_data_78_port, 
      DataPath_RF_bus_sel_savedwin_data_79_port, 
      DataPath_RF_bus_sel_savedwin_data_80_port, 
      DataPath_RF_bus_sel_savedwin_data_81_port, 
      DataPath_RF_bus_sel_savedwin_data_82_port, 
      DataPath_RF_bus_sel_savedwin_data_83_port, 
      DataPath_RF_bus_sel_savedwin_data_84_port, 
      DataPath_RF_bus_sel_savedwin_data_85_port, 
      DataPath_RF_bus_sel_savedwin_data_86_port, 
      DataPath_RF_bus_sel_savedwin_data_87_port, 
      DataPath_RF_bus_sel_savedwin_data_88_port, 
      DataPath_RF_bus_sel_savedwin_data_89_port, 
      DataPath_RF_bus_sel_savedwin_data_90_port, 
      DataPath_RF_bus_sel_savedwin_data_91_port, 
      DataPath_RF_bus_sel_savedwin_data_92_port, 
      DataPath_RF_bus_sel_savedwin_data_93_port, 
      DataPath_RF_bus_sel_savedwin_data_94_port, 
      DataPath_RF_bus_sel_savedwin_data_95_port, 
      DataPath_RF_bus_sel_savedwin_data_96_port, 
      DataPath_RF_bus_sel_savedwin_data_97_port, 
      DataPath_RF_bus_sel_savedwin_data_98_port, 
      DataPath_RF_bus_sel_savedwin_data_99_port, 
      DataPath_RF_bus_sel_savedwin_data_100_port, 
      DataPath_RF_bus_sel_savedwin_data_101_port, 
      DataPath_RF_bus_sel_savedwin_data_102_port, 
      DataPath_RF_bus_sel_savedwin_data_103_port, 
      DataPath_RF_bus_sel_savedwin_data_104_port, 
      DataPath_RF_bus_sel_savedwin_data_105_port, 
      DataPath_RF_bus_sel_savedwin_data_106_port, 
      DataPath_RF_bus_sel_savedwin_data_107_port, 
      DataPath_RF_bus_sel_savedwin_data_108_port, 
      DataPath_RF_bus_sel_savedwin_data_109_port, 
      DataPath_RF_bus_sel_savedwin_data_110_port, 
      DataPath_RF_bus_sel_savedwin_data_111_port, 
      DataPath_RF_bus_sel_savedwin_data_112_port, 
      DataPath_RF_bus_sel_savedwin_data_113_port, 
      DataPath_RF_bus_sel_savedwin_data_114_port, 
      DataPath_RF_bus_sel_savedwin_data_115_port, 
      DataPath_RF_bus_sel_savedwin_data_116_port, 
      DataPath_RF_bus_sel_savedwin_data_117_port, 
      DataPath_RF_bus_sel_savedwin_data_118_port, 
      DataPath_RF_bus_sel_savedwin_data_119_port, 
      DataPath_RF_bus_sel_savedwin_data_120_port, 
      DataPath_RF_bus_sel_savedwin_data_121_port, 
      DataPath_RF_bus_sel_savedwin_data_122_port, 
      DataPath_RF_bus_sel_savedwin_data_123_port, 
      DataPath_RF_bus_sel_savedwin_data_124_port, 
      DataPath_RF_bus_sel_savedwin_data_125_port, 
      DataPath_RF_bus_sel_savedwin_data_126_port, 
      DataPath_RF_bus_sel_savedwin_data_127_port, 
      DataPath_RF_bus_sel_savedwin_data_128_port, 
      DataPath_RF_bus_sel_savedwin_data_129_port, 
      DataPath_RF_bus_sel_savedwin_data_130_port, 
      DataPath_RF_bus_sel_savedwin_data_131_port, 
      DataPath_RF_bus_sel_savedwin_data_132_port, 
      DataPath_RF_bus_sel_savedwin_data_133_port, 
      DataPath_RF_bus_sel_savedwin_data_134_port, 
      DataPath_RF_bus_sel_savedwin_data_135_port, 
      DataPath_RF_bus_sel_savedwin_data_136_port, 
      DataPath_RF_bus_sel_savedwin_data_137_port, 
      DataPath_RF_bus_sel_savedwin_data_138_port, 
      DataPath_RF_bus_sel_savedwin_data_139_port, 
      DataPath_RF_bus_sel_savedwin_data_140_port, 
      DataPath_RF_bus_sel_savedwin_data_141_port, 
      DataPath_RF_bus_sel_savedwin_data_142_port, 
      DataPath_RF_bus_sel_savedwin_data_143_port, 
      DataPath_RF_bus_sel_savedwin_data_144_port, 
      DataPath_RF_bus_sel_savedwin_data_145_port, 
      DataPath_RF_bus_sel_savedwin_data_146_port, 
      DataPath_RF_bus_sel_savedwin_data_147_port, 
      DataPath_RF_bus_sel_savedwin_data_148_port, 
      DataPath_RF_bus_sel_savedwin_data_149_port, 
      DataPath_RF_bus_sel_savedwin_data_150_port, 
      DataPath_RF_bus_sel_savedwin_data_151_port, 
      DataPath_RF_bus_sel_savedwin_data_152_port, 
      DataPath_RF_bus_sel_savedwin_data_153_port, 
      DataPath_RF_bus_sel_savedwin_data_154_port, 
      DataPath_RF_bus_sel_savedwin_data_155_port, 
      DataPath_RF_bus_sel_savedwin_data_156_port, 
      DataPath_RF_bus_sel_savedwin_data_157_port, 
      DataPath_RF_bus_sel_savedwin_data_158_port, 
      DataPath_RF_bus_sel_savedwin_data_159_port, 
      DataPath_RF_bus_sel_savedwin_data_160_port, 
      DataPath_RF_bus_sel_savedwin_data_161_port, 
      DataPath_RF_bus_sel_savedwin_data_162_port, 
      DataPath_RF_bus_sel_savedwin_data_163_port, 
      DataPath_RF_bus_sel_savedwin_data_164_port, 
      DataPath_RF_bus_sel_savedwin_data_165_port, 
      DataPath_RF_bus_sel_savedwin_data_166_port, 
      DataPath_RF_bus_sel_savedwin_data_167_port, 
      DataPath_RF_bus_sel_savedwin_data_168_port, 
      DataPath_RF_bus_sel_savedwin_data_169_port, 
      DataPath_RF_bus_sel_savedwin_data_170_port, 
      DataPath_RF_bus_sel_savedwin_data_171_port, 
      DataPath_RF_bus_sel_savedwin_data_172_port, 
      DataPath_RF_bus_sel_savedwin_data_173_port, 
      DataPath_RF_bus_sel_savedwin_data_174_port, 
      DataPath_RF_bus_sel_savedwin_data_175_port, 
      DataPath_RF_bus_sel_savedwin_data_176_port, 
      DataPath_RF_bus_sel_savedwin_data_177_port, 
      DataPath_RF_bus_sel_savedwin_data_178_port, 
      DataPath_RF_bus_sel_savedwin_data_179_port, 
      DataPath_RF_bus_sel_savedwin_data_180_port, 
      DataPath_RF_bus_sel_savedwin_data_181_port, 
      DataPath_RF_bus_sel_savedwin_data_182_port, 
      DataPath_RF_bus_sel_savedwin_data_183_port, 
      DataPath_RF_bus_sel_savedwin_data_184_port, 
      DataPath_RF_bus_sel_savedwin_data_185_port, 
      DataPath_RF_bus_sel_savedwin_data_186_port, 
      DataPath_RF_bus_sel_savedwin_data_187_port, 
      DataPath_RF_bus_sel_savedwin_data_188_port, 
      DataPath_RF_bus_sel_savedwin_data_189_port, 
      DataPath_RF_bus_sel_savedwin_data_190_port, 
      DataPath_RF_bus_sel_savedwin_data_191_port, 
      DataPath_RF_bus_sel_savedwin_data_192_port, 
      DataPath_RF_bus_sel_savedwin_data_193_port, 
      DataPath_RF_bus_sel_savedwin_data_194_port, 
      DataPath_RF_bus_sel_savedwin_data_195_port, 
      DataPath_RF_bus_sel_savedwin_data_196_port, 
      DataPath_RF_bus_sel_savedwin_data_197_port, 
      DataPath_RF_bus_sel_savedwin_data_198_port, 
      DataPath_RF_bus_sel_savedwin_data_199_port, 
      DataPath_RF_bus_sel_savedwin_data_200_port, 
      DataPath_RF_bus_sel_savedwin_data_201_port, 
      DataPath_RF_bus_sel_savedwin_data_202_port, 
      DataPath_RF_bus_sel_savedwin_data_203_port, 
      DataPath_RF_bus_sel_savedwin_data_204_port, 
      DataPath_RF_bus_sel_savedwin_data_205_port, 
      DataPath_RF_bus_sel_savedwin_data_206_port, 
      DataPath_RF_bus_sel_savedwin_data_207_port, 
      DataPath_RF_bus_sel_savedwin_data_208_port, 
      DataPath_RF_bus_sel_savedwin_data_209_port, 
      DataPath_RF_bus_sel_savedwin_data_210_port, 
      DataPath_RF_bus_sel_savedwin_data_211_port, 
      DataPath_RF_bus_sel_savedwin_data_212_port, 
      DataPath_RF_bus_sel_savedwin_data_213_port, 
      DataPath_RF_bus_sel_savedwin_data_214_port, 
      DataPath_RF_bus_sel_savedwin_data_215_port, 
      DataPath_RF_bus_sel_savedwin_data_216_port, 
      DataPath_RF_bus_sel_savedwin_data_217_port, 
      DataPath_RF_bus_sel_savedwin_data_218_port, 
      DataPath_RF_bus_sel_savedwin_data_219_port, 
      DataPath_RF_bus_sel_savedwin_data_220_port, 
      DataPath_RF_bus_sel_savedwin_data_221_port, 
      DataPath_RF_bus_sel_savedwin_data_222_port, 
      DataPath_RF_bus_sel_savedwin_data_223_port, 
      DataPath_RF_bus_sel_savedwin_data_224_port, 
      DataPath_RF_bus_sel_savedwin_data_225_port, 
      DataPath_RF_bus_sel_savedwin_data_226_port, 
      DataPath_RF_bus_sel_savedwin_data_227_port, 
      DataPath_RF_bus_sel_savedwin_data_228_port, 
      DataPath_RF_bus_sel_savedwin_data_229_port, 
      DataPath_RF_bus_sel_savedwin_data_230_port, 
      DataPath_RF_bus_sel_savedwin_data_231_port, 
      DataPath_RF_bus_sel_savedwin_data_232_port, 
      DataPath_RF_bus_sel_savedwin_data_233_port, 
      DataPath_RF_bus_sel_savedwin_data_234_port, 
      DataPath_RF_bus_sel_savedwin_data_235_port, 
      DataPath_RF_bus_sel_savedwin_data_236_port, 
      DataPath_RF_bus_sel_savedwin_data_237_port, 
      DataPath_RF_bus_sel_savedwin_data_238_port, 
      DataPath_RF_bus_sel_savedwin_data_239_port, 
      DataPath_RF_bus_sel_savedwin_data_240_port, 
      DataPath_RF_bus_sel_savedwin_data_241_port, 
      DataPath_RF_bus_sel_savedwin_data_242_port, 
      DataPath_RF_bus_sel_savedwin_data_243_port, 
      DataPath_RF_bus_sel_savedwin_data_244_port, 
      DataPath_RF_bus_sel_savedwin_data_245_port, 
      DataPath_RF_bus_sel_savedwin_data_246_port, 
      DataPath_RF_bus_sel_savedwin_data_247_port, 
      DataPath_RF_bus_sel_savedwin_data_248_port, 
      DataPath_RF_bus_sel_savedwin_data_249_port, 
      DataPath_RF_bus_sel_savedwin_data_250_port, 
      DataPath_RF_bus_sel_savedwin_data_251_port, 
      DataPath_RF_bus_sel_savedwin_data_252_port, 
      DataPath_RF_bus_sel_savedwin_data_253_port, 
      DataPath_RF_bus_sel_savedwin_data_254_port, 
      DataPath_RF_bus_sel_savedwin_data_255_port, 
      DataPath_RF_bus_sel_savedwin_data_256_port, 
      DataPath_RF_bus_sel_savedwin_data_257_port, 
      DataPath_RF_bus_sel_savedwin_data_258_port, 
      DataPath_RF_bus_sel_savedwin_data_259_port, 
      DataPath_RF_bus_sel_savedwin_data_260_port, 
      DataPath_RF_bus_sel_savedwin_data_261_port, 
      DataPath_RF_bus_sel_savedwin_data_262_port, 
      DataPath_RF_bus_sel_savedwin_data_263_port, 
      DataPath_RF_bus_sel_savedwin_data_264_port, 
      DataPath_RF_bus_sel_savedwin_data_265_port, 
      DataPath_RF_bus_sel_savedwin_data_266_port, 
      DataPath_RF_bus_sel_savedwin_data_267_port, 
      DataPath_RF_bus_sel_savedwin_data_268_port, 
      DataPath_RF_bus_sel_savedwin_data_269_port, 
      DataPath_RF_bus_sel_savedwin_data_270_port, 
      DataPath_RF_bus_sel_savedwin_data_271_port, 
      DataPath_RF_bus_sel_savedwin_data_272_port, 
      DataPath_RF_bus_sel_savedwin_data_273_port, 
      DataPath_RF_bus_sel_savedwin_data_274_port, 
      DataPath_RF_bus_sel_savedwin_data_275_port, 
      DataPath_RF_bus_sel_savedwin_data_276_port, 
      DataPath_RF_bus_sel_savedwin_data_277_port, 
      DataPath_RF_bus_sel_savedwin_data_278_port, 
      DataPath_RF_bus_sel_savedwin_data_279_port, 
      DataPath_RF_bus_sel_savedwin_data_280_port, 
      DataPath_RF_bus_sel_savedwin_data_281_port, 
      DataPath_RF_bus_sel_savedwin_data_282_port, 
      DataPath_RF_bus_sel_savedwin_data_283_port, 
      DataPath_RF_bus_sel_savedwin_data_284_port, 
      DataPath_RF_bus_sel_savedwin_data_285_port, 
      DataPath_RF_bus_sel_savedwin_data_286_port, 
      DataPath_RF_bus_sel_savedwin_data_287_port, 
      DataPath_RF_bus_sel_savedwin_data_288_port, 
      DataPath_RF_bus_sel_savedwin_data_289_port, 
      DataPath_RF_bus_sel_savedwin_data_290_port, 
      DataPath_RF_bus_sel_savedwin_data_291_port, 
      DataPath_RF_bus_sel_savedwin_data_292_port, 
      DataPath_RF_bus_sel_savedwin_data_293_port, 
      DataPath_RF_bus_sel_savedwin_data_294_port, 
      DataPath_RF_bus_sel_savedwin_data_295_port, 
      DataPath_RF_bus_sel_savedwin_data_296_port, 
      DataPath_RF_bus_sel_savedwin_data_297_port, 
      DataPath_RF_bus_sel_savedwin_data_298_port, 
      DataPath_RF_bus_sel_savedwin_data_299_port, 
      DataPath_RF_bus_sel_savedwin_data_300_port, 
      DataPath_RF_bus_sel_savedwin_data_301_port, 
      DataPath_RF_bus_sel_savedwin_data_302_port, 
      DataPath_RF_bus_sel_savedwin_data_303_port, 
      DataPath_RF_bus_sel_savedwin_data_304_port, 
      DataPath_RF_bus_sel_savedwin_data_305_port, 
      DataPath_RF_bus_sel_savedwin_data_306_port, 
      DataPath_RF_bus_sel_savedwin_data_307_port, 
      DataPath_RF_bus_sel_savedwin_data_308_port, 
      DataPath_RF_bus_sel_savedwin_data_309_port, 
      DataPath_RF_bus_sel_savedwin_data_310_port, 
      DataPath_RF_bus_sel_savedwin_data_311_port, 
      DataPath_RF_bus_sel_savedwin_data_312_port, 
      DataPath_RF_bus_sel_savedwin_data_313_port, 
      DataPath_RF_bus_sel_savedwin_data_314_port, 
      DataPath_RF_bus_sel_savedwin_data_315_port, 
      DataPath_RF_bus_sel_savedwin_data_316_port, 
      DataPath_RF_bus_sel_savedwin_data_317_port, 
      DataPath_RF_bus_sel_savedwin_data_318_port, 
      DataPath_RF_bus_sel_savedwin_data_319_port, 
      DataPath_RF_bus_sel_savedwin_data_320_port, 
      DataPath_RF_bus_sel_savedwin_data_321_port, 
      DataPath_RF_bus_sel_savedwin_data_322_port, 
      DataPath_RF_bus_sel_savedwin_data_323_port, 
      DataPath_RF_bus_sel_savedwin_data_324_port, 
      DataPath_RF_bus_sel_savedwin_data_325_port, 
      DataPath_RF_bus_sel_savedwin_data_326_port, 
      DataPath_RF_bus_sel_savedwin_data_327_port, 
      DataPath_RF_bus_sel_savedwin_data_328_port, 
      DataPath_RF_bus_sel_savedwin_data_329_port, 
      DataPath_RF_bus_sel_savedwin_data_330_port, 
      DataPath_RF_bus_sel_savedwin_data_331_port, 
      DataPath_RF_bus_sel_savedwin_data_332_port, 
      DataPath_RF_bus_sel_savedwin_data_333_port, 
      DataPath_RF_bus_sel_savedwin_data_334_port, 
      DataPath_RF_bus_sel_savedwin_data_335_port, 
      DataPath_RF_bus_sel_savedwin_data_336_port, 
      DataPath_RF_bus_sel_savedwin_data_337_port, 
      DataPath_RF_bus_sel_savedwin_data_338_port, 
      DataPath_RF_bus_sel_savedwin_data_339_port, 
      DataPath_RF_bus_sel_savedwin_data_340_port, 
      DataPath_RF_bus_sel_savedwin_data_341_port, 
      DataPath_RF_bus_sel_savedwin_data_342_port, 
      DataPath_RF_bus_sel_savedwin_data_343_port, 
      DataPath_RF_bus_sel_savedwin_data_344_port, 
      DataPath_RF_bus_sel_savedwin_data_345_port, 
      DataPath_RF_bus_sel_savedwin_data_346_port, 
      DataPath_RF_bus_sel_savedwin_data_347_port, 
      DataPath_RF_bus_sel_savedwin_data_348_port, 
      DataPath_RF_bus_sel_savedwin_data_349_port, 
      DataPath_RF_bus_sel_savedwin_data_350_port, 
      DataPath_RF_bus_sel_savedwin_data_351_port, 
      DataPath_RF_bus_sel_savedwin_data_352_port, 
      DataPath_RF_bus_sel_savedwin_data_353_port, 
      DataPath_RF_bus_sel_savedwin_data_354_port, 
      DataPath_RF_bus_sel_savedwin_data_355_port, 
      DataPath_RF_bus_sel_savedwin_data_356_port, 
      DataPath_RF_bus_sel_savedwin_data_357_port, 
      DataPath_RF_bus_sel_savedwin_data_358_port, 
      DataPath_RF_bus_sel_savedwin_data_359_port, 
      DataPath_RF_bus_sel_savedwin_data_360_port, 
      DataPath_RF_bus_sel_savedwin_data_361_port, 
      DataPath_RF_bus_sel_savedwin_data_362_port, 
      DataPath_RF_bus_sel_savedwin_data_363_port, 
      DataPath_RF_bus_sel_savedwin_data_364_port, 
      DataPath_RF_bus_sel_savedwin_data_365_port, 
      DataPath_RF_bus_sel_savedwin_data_366_port, 
      DataPath_RF_bus_sel_savedwin_data_367_port, 
      DataPath_RF_bus_sel_savedwin_data_368_port, 
      DataPath_RF_bus_sel_savedwin_data_369_port, 
      DataPath_RF_bus_sel_savedwin_data_370_port, 
      DataPath_RF_bus_sel_savedwin_data_371_port, 
      DataPath_RF_bus_sel_savedwin_data_372_port, 
      DataPath_RF_bus_sel_savedwin_data_373_port, 
      DataPath_RF_bus_sel_savedwin_data_374_port, 
      DataPath_RF_bus_sel_savedwin_data_375_port, 
      DataPath_RF_bus_sel_savedwin_data_376_port, 
      DataPath_RF_bus_sel_savedwin_data_377_port, 
      DataPath_RF_bus_sel_savedwin_data_378_port, 
      DataPath_RF_bus_sel_savedwin_data_379_port, 
      DataPath_RF_bus_sel_savedwin_data_380_port, 
      DataPath_RF_bus_sel_savedwin_data_381_port, 
      DataPath_RF_bus_sel_savedwin_data_382_port, 
      DataPath_RF_bus_sel_savedwin_data_383_port, 
      DataPath_RF_bus_sel_savedwin_data_384_port, 
      DataPath_RF_bus_sel_savedwin_data_385_port, 
      DataPath_RF_bus_sel_savedwin_data_386_port, 
      DataPath_RF_bus_sel_savedwin_data_387_port, 
      DataPath_RF_bus_sel_savedwin_data_388_port, 
      DataPath_RF_bus_sel_savedwin_data_389_port, 
      DataPath_RF_bus_sel_savedwin_data_390_port, 
      DataPath_RF_bus_sel_savedwin_data_391_port, 
      DataPath_RF_bus_sel_savedwin_data_392_port, 
      DataPath_RF_bus_sel_savedwin_data_393_port, 
      DataPath_RF_bus_sel_savedwin_data_394_port, 
      DataPath_RF_bus_sel_savedwin_data_395_port, 
      DataPath_RF_bus_sel_savedwin_data_396_port, 
      DataPath_RF_bus_sel_savedwin_data_397_port, 
      DataPath_RF_bus_sel_savedwin_data_398_port, 
      DataPath_RF_bus_sel_savedwin_data_399_port, 
      DataPath_RF_bus_sel_savedwin_data_400_port, 
      DataPath_RF_bus_sel_savedwin_data_401_port, 
      DataPath_RF_bus_sel_savedwin_data_402_port, 
      DataPath_RF_bus_sel_savedwin_data_403_port, 
      DataPath_RF_bus_sel_savedwin_data_404_port, 
      DataPath_RF_bus_sel_savedwin_data_405_port, 
      DataPath_RF_bus_sel_savedwin_data_406_port, 
      DataPath_RF_bus_sel_savedwin_data_407_port, 
      DataPath_RF_bus_sel_savedwin_data_408_port, 
      DataPath_RF_bus_sel_savedwin_data_409_port, 
      DataPath_RF_bus_sel_savedwin_data_410_port, 
      DataPath_RF_bus_sel_savedwin_data_411_port, 
      DataPath_RF_bus_sel_savedwin_data_412_port, 
      DataPath_RF_bus_sel_savedwin_data_413_port, 
      DataPath_RF_bus_sel_savedwin_data_414_port, 
      DataPath_RF_bus_sel_savedwin_data_415_port, 
      DataPath_RF_bus_sel_savedwin_data_416_port, 
      DataPath_RF_bus_sel_savedwin_data_417_port, 
      DataPath_RF_bus_sel_savedwin_data_418_port, 
      DataPath_RF_bus_sel_savedwin_data_419_port, 
      DataPath_RF_bus_sel_savedwin_data_420_port, 
      DataPath_RF_bus_sel_savedwin_data_421_port, 
      DataPath_RF_bus_sel_savedwin_data_422_port, 
      DataPath_RF_bus_sel_savedwin_data_423_port, 
      DataPath_RF_bus_sel_savedwin_data_424_port, 
      DataPath_RF_bus_sel_savedwin_data_425_port, 
      DataPath_RF_bus_sel_savedwin_data_426_port, 
      DataPath_RF_bus_sel_savedwin_data_427_port, 
      DataPath_RF_bus_sel_savedwin_data_428_port, 
      DataPath_RF_bus_sel_savedwin_data_429_port, 
      DataPath_RF_bus_sel_savedwin_data_430_port, 
      DataPath_RF_bus_sel_savedwin_data_431_port, 
      DataPath_RF_bus_sel_savedwin_data_432_port, 
      DataPath_RF_bus_sel_savedwin_data_433_port, 
      DataPath_RF_bus_sel_savedwin_data_434_port, 
      DataPath_RF_bus_sel_savedwin_data_435_port, 
      DataPath_RF_bus_sel_savedwin_data_436_port, 
      DataPath_RF_bus_sel_savedwin_data_437_port, 
      DataPath_RF_bus_sel_savedwin_data_438_port, 
      DataPath_RF_bus_sel_savedwin_data_439_port, 
      DataPath_RF_bus_sel_savedwin_data_440_port, 
      DataPath_RF_bus_sel_savedwin_data_441_port, 
      DataPath_RF_bus_sel_savedwin_data_442_port, 
      DataPath_RF_bus_sel_savedwin_data_443_port, 
      DataPath_RF_bus_sel_savedwin_data_444_port, 
      DataPath_RF_bus_sel_savedwin_data_445_port, 
      DataPath_RF_bus_sel_savedwin_data_446_port, 
      DataPath_RF_bus_sel_savedwin_data_447_port, 
      DataPath_RF_bus_sel_savedwin_data_448_port, 
      DataPath_RF_bus_sel_savedwin_data_449_port, 
      DataPath_RF_bus_sel_savedwin_data_450_port, 
      DataPath_RF_bus_sel_savedwin_data_451_port, 
      DataPath_RF_bus_sel_savedwin_data_452_port, 
      DataPath_RF_bus_sel_savedwin_data_453_port, 
      DataPath_RF_bus_sel_savedwin_data_454_port, 
      DataPath_RF_bus_sel_savedwin_data_455_port, 
      DataPath_RF_bus_sel_savedwin_data_456_port, 
      DataPath_RF_bus_sel_savedwin_data_457_port, 
      DataPath_RF_bus_sel_savedwin_data_458_port, 
      DataPath_RF_bus_sel_savedwin_data_459_port, 
      DataPath_RF_bus_sel_savedwin_data_460_port, 
      DataPath_RF_bus_sel_savedwin_data_461_port, 
      DataPath_RF_bus_sel_savedwin_data_462_port, 
      DataPath_RF_bus_sel_savedwin_data_463_port, 
      DataPath_RF_bus_sel_savedwin_data_464_port, 
      DataPath_RF_bus_sel_savedwin_data_465_port, 
      DataPath_RF_bus_sel_savedwin_data_466_port, 
      DataPath_RF_bus_sel_savedwin_data_467_port, 
      DataPath_RF_bus_sel_savedwin_data_468_port, 
      DataPath_RF_bus_sel_savedwin_data_469_port, 
      DataPath_RF_bus_sel_savedwin_data_470_port, 
      DataPath_RF_bus_sel_savedwin_data_471_port, 
      DataPath_RF_bus_sel_savedwin_data_472_port, 
      DataPath_RF_bus_sel_savedwin_data_473_port, 
      DataPath_RF_bus_sel_savedwin_data_474_port, 
      DataPath_RF_bus_sel_savedwin_data_475_port, 
      DataPath_RF_bus_sel_savedwin_data_476_port, 
      DataPath_RF_bus_sel_savedwin_data_477_port, 
      DataPath_RF_bus_sel_savedwin_data_478_port, 
      DataPath_RF_bus_sel_savedwin_data_479_port, 
      DataPath_RF_bus_sel_savedwin_data_480_port, 
      DataPath_RF_bus_sel_savedwin_data_481_port, 
      DataPath_RF_bus_sel_savedwin_data_482_port, 
      DataPath_RF_bus_sel_savedwin_data_483_port, 
      DataPath_RF_bus_sel_savedwin_data_484_port, 
      DataPath_RF_bus_sel_savedwin_data_485_port, 
      DataPath_RF_bus_sel_savedwin_data_486_port, 
      DataPath_RF_bus_sel_savedwin_data_487_port, 
      DataPath_RF_bus_sel_savedwin_data_488_port, 
      DataPath_RF_bus_sel_savedwin_data_489_port, 
      DataPath_RF_bus_sel_savedwin_data_490_port, 
      DataPath_RF_bus_sel_savedwin_data_491_port, 
      DataPath_RF_bus_sel_savedwin_data_492_port, 
      DataPath_RF_bus_sel_savedwin_data_493_port, 
      DataPath_RF_bus_sel_savedwin_data_494_port, 
      DataPath_RF_bus_sel_savedwin_data_495_port, 
      DataPath_RF_bus_sel_savedwin_data_496_port, 
      DataPath_RF_bus_sel_savedwin_data_497_port, 
      DataPath_RF_bus_sel_savedwin_data_498_port, 
      DataPath_RF_bus_sel_savedwin_data_499_port, 
      DataPath_RF_bus_sel_savedwin_data_500_port, 
      DataPath_RF_bus_sel_savedwin_data_501_port, 
      DataPath_RF_bus_sel_savedwin_data_502_port, 
      DataPath_RF_bus_sel_savedwin_data_503_port, 
      DataPath_RF_bus_sel_savedwin_data_504_port, 
      DataPath_RF_bus_sel_savedwin_data_505_port, 
      DataPath_RF_bus_sel_savedwin_data_506_port, 
      DataPath_RF_bus_sel_savedwin_data_507_port, 
      DataPath_RF_bus_sel_savedwin_data_508_port, 
      DataPath_RF_bus_sel_savedwin_data_509_port, 
      DataPath_RF_bus_sel_savedwin_data_510_port, 
      DataPath_RF_bus_sel_savedwin_data_511_port, DataPath_RF_next_swp_0_port, 
      DataPath_RF_next_swp_1_port, DataPath_RF_next_swp_2_port, 
      DataPath_RF_next_swp_3_port, DataPath_RF_next_swp_4_port, 
      DataPath_RF_c_swin_0_port, DataPath_RF_c_swin_1_port, 
      DataPath_RF_c_swin_2_port, DataPath_RF_c_swin_3_port, 
      DataPath_RF_c_swin_4_port, DataPath_RF_fill_address_ext_0_port, 
      DataPath_RF_fill_address_ext_1_port, DataPath_RF_fill_address_ext_2_port,
      DataPath_RF_fill_address_ext_3_port, DataPath_RF_fill_address_ext_4_port,
      DataPath_RF_fill_address_ext_5_port, DataPath_RF_fill_address_ext_6_port,
      DataPath_RF_fill_address_ext_7_port, DataPath_RF_fill_address_ext_8_port,
      DataPath_RF_fill_address_ext_9_port, DataPath_RF_fill_address_ext_10_port
      , DataPath_RF_fill_address_ext_11_port, 
      DataPath_RF_fill_address_ext_12_port, 
      DataPath_RF_fill_address_ext_13_port, 
      DataPath_RF_fill_address_ext_14_port, 
      DataPath_RF_fill_address_ext_15_port, DataPath_RF_dec_output_8_port, 
      DataPath_RF_dec_output_9_port, DataPath_RF_dec_output_10_port, 
      DataPath_RF_dec_output_11_port, DataPath_RF_dec_output_12_port, 
      DataPath_RF_dec_output_13_port, DataPath_RF_dec_output_14_port, 
      DataPath_RF_dec_output_15_port, DataPath_RF_dec_output_16_port, 
      DataPath_RF_dec_output_17_port, DataPath_RF_dec_output_18_port, 
      DataPath_RF_dec_output_19_port, DataPath_RF_dec_output_20_port, 
      DataPath_RF_dec_output_21_port, DataPath_RF_dec_output_22_port, 
      DataPath_RF_dec_output_23_port, DataPath_RF_dec_output_24_port, 
      DataPath_RF_dec_output_25_port, DataPath_RF_dec_output_26_port, 
      DataPath_RF_dec_output_27_port, DataPath_RF_dec_output_28_port, 
      DataPath_RF_dec_output_29_port, DataPath_RF_dec_output_30_port, 
      DataPath_RF_dec_output_31_port, DataPath_RF_internal_inloc_data_4_0_port,
      DataPath_RF_internal_inloc_data_4_1_port, 
      DataPath_RF_internal_inloc_data_4_2_port, 
      DataPath_RF_internal_inloc_data_4_3_port, 
      DataPath_RF_internal_inloc_data_4_4_port, 
      DataPath_RF_internal_inloc_data_4_5_port, 
      DataPath_RF_internal_inloc_data_4_6_port, 
      DataPath_RF_internal_inloc_data_4_7_port, 
      DataPath_RF_internal_inloc_data_4_8_port, 
      DataPath_RF_internal_inloc_data_4_9_port, 
      DataPath_RF_internal_inloc_data_4_10_port, 
      DataPath_RF_internal_inloc_data_4_11_port, 
      DataPath_RF_internal_inloc_data_4_12_port, 
      DataPath_RF_internal_inloc_data_4_13_port, 
      DataPath_RF_internal_inloc_data_4_14_port, 
      DataPath_RF_internal_inloc_data_4_15_port, 
      DataPath_RF_internal_inloc_data_4_16_port, 
      DataPath_RF_internal_inloc_data_4_17_port, 
      DataPath_RF_internal_inloc_data_4_18_port, 
      DataPath_RF_internal_inloc_data_4_19_port, 
      DataPath_RF_internal_inloc_data_4_20_port, 
      DataPath_RF_internal_inloc_data_4_21_port, 
      DataPath_RF_internal_inloc_data_4_22_port, 
      DataPath_RF_internal_inloc_data_4_23_port, 
      DataPath_RF_internal_inloc_data_4_24_port, 
      DataPath_RF_internal_inloc_data_4_25_port, 
      DataPath_RF_internal_inloc_data_4_26_port, 
      DataPath_RF_internal_inloc_data_4_27_port, 
      DataPath_RF_internal_inloc_data_4_28_port, 
      DataPath_RF_internal_inloc_data_4_29_port, 
      DataPath_RF_internal_inloc_data_4_30_port, 
      DataPath_RF_internal_inloc_data_4_31_port, 
      DataPath_RF_internal_inloc_data_3_0_port, 
      DataPath_RF_internal_inloc_data_3_1_port, 
      DataPath_RF_internal_inloc_data_3_2_port, 
      DataPath_RF_internal_inloc_data_3_3_port, 
      DataPath_RF_internal_inloc_data_3_4_port, 
      DataPath_RF_internal_inloc_data_3_5_port, 
      DataPath_RF_internal_inloc_data_3_6_port, 
      DataPath_RF_internal_inloc_data_3_7_port, 
      DataPath_RF_internal_inloc_data_3_8_port, 
      DataPath_RF_internal_inloc_data_3_9_port, 
      DataPath_RF_internal_inloc_data_3_10_port, 
      DataPath_RF_internal_inloc_data_3_11_port, 
      DataPath_RF_internal_inloc_data_3_12_port, 
      DataPath_RF_internal_inloc_data_3_13_port, 
      DataPath_RF_internal_inloc_data_3_14_port, 
      DataPath_RF_internal_inloc_data_3_15_port, 
      DataPath_RF_internal_inloc_data_3_16_port, 
      DataPath_RF_internal_inloc_data_3_17_port, 
      DataPath_RF_internal_inloc_data_3_18_port, 
      DataPath_RF_internal_inloc_data_3_19_port, 
      DataPath_RF_internal_inloc_data_3_20_port, 
      DataPath_RF_internal_inloc_data_3_21_port, 
      DataPath_RF_internal_inloc_data_3_22_port, 
      DataPath_RF_internal_inloc_data_3_23_port, 
      DataPath_RF_internal_inloc_data_3_24_port, 
      DataPath_RF_internal_inloc_data_3_25_port, 
      DataPath_RF_internal_inloc_data_3_26_port, 
      DataPath_RF_internal_inloc_data_3_27_port, 
      DataPath_RF_internal_inloc_data_3_28_port, 
      DataPath_RF_internal_inloc_data_3_29_port, 
      DataPath_RF_internal_inloc_data_3_30_port, 
      DataPath_RF_internal_inloc_data_3_31_port, 
      DataPath_RF_internal_inloc_data_2_0_port, 
      DataPath_RF_internal_inloc_data_2_1_port, 
      DataPath_RF_internal_inloc_data_2_2_port, 
      DataPath_RF_internal_inloc_data_2_3_port, 
      DataPath_RF_internal_inloc_data_2_4_port, 
      DataPath_RF_internal_inloc_data_2_5_port, 
      DataPath_RF_internal_inloc_data_2_6_port, 
      DataPath_RF_internal_inloc_data_2_7_port, 
      DataPath_RF_internal_inloc_data_2_8_port, 
      DataPath_RF_internal_inloc_data_2_9_port, 
      DataPath_RF_internal_inloc_data_2_10_port, 
      DataPath_RF_internal_inloc_data_2_11_port, 
      DataPath_RF_internal_inloc_data_2_12_port, 
      DataPath_RF_internal_inloc_data_2_13_port, 
      DataPath_RF_internal_inloc_data_2_14_port, 
      DataPath_RF_internal_inloc_data_2_15_port, 
      DataPath_RF_internal_inloc_data_2_16_port, 
      DataPath_RF_internal_inloc_data_2_17_port, 
      DataPath_RF_internal_inloc_data_2_18_port, 
      DataPath_RF_internal_inloc_data_2_19_port, 
      DataPath_RF_internal_inloc_data_2_20_port, 
      DataPath_RF_internal_inloc_data_2_21_port, 
      DataPath_RF_internal_inloc_data_2_22_port, 
      DataPath_RF_internal_inloc_data_2_23_port, 
      DataPath_RF_internal_inloc_data_2_24_port, 
      DataPath_RF_internal_inloc_data_2_25_port, 
      DataPath_RF_internal_inloc_data_2_26_port, 
      DataPath_RF_internal_inloc_data_2_27_port, 
      DataPath_RF_internal_inloc_data_2_28_port, 
      DataPath_RF_internal_inloc_data_2_29_port, 
      DataPath_RF_internal_inloc_data_2_30_port, 
      DataPath_RF_internal_inloc_data_2_31_port, 
      DataPath_RF_internal_inloc_data_1_0_port, 
      DataPath_RF_internal_inloc_data_1_1_port, 
      DataPath_RF_internal_inloc_data_1_2_port, 
      DataPath_RF_internal_inloc_data_1_3_port, 
      DataPath_RF_internal_inloc_data_1_4_port, 
      DataPath_RF_internal_inloc_data_1_5_port, 
      DataPath_RF_internal_inloc_data_1_6_port, 
      DataPath_RF_internal_inloc_data_1_7_port, 
      DataPath_RF_internal_inloc_data_1_8_port, 
      DataPath_RF_internal_inloc_data_1_9_port, 
      DataPath_RF_internal_inloc_data_1_10_port, 
      DataPath_RF_internal_inloc_data_1_11_port, 
      DataPath_RF_internal_inloc_data_1_12_port, 
      DataPath_RF_internal_inloc_data_1_13_port, 
      DataPath_RF_internal_inloc_data_1_14_port, 
      DataPath_RF_internal_inloc_data_1_15_port, 
      DataPath_RF_internal_inloc_data_1_16_port, 
      DataPath_RF_internal_inloc_data_1_17_port, 
      DataPath_RF_internal_inloc_data_1_18_port, 
      DataPath_RF_internal_inloc_data_1_19_port, 
      DataPath_RF_internal_inloc_data_1_20_port, 
      DataPath_RF_internal_inloc_data_1_21_port, 
      DataPath_RF_internal_inloc_data_1_22_port, 
      DataPath_RF_internal_inloc_data_1_23_port, 
      DataPath_RF_internal_inloc_data_1_24_port, 
      DataPath_RF_internal_inloc_data_1_25_port, 
      DataPath_RF_internal_inloc_data_1_26_port, 
      DataPath_RF_internal_inloc_data_1_27_port, 
      DataPath_RF_internal_inloc_data_1_28_port, 
      DataPath_RF_internal_inloc_data_1_29_port, 
      DataPath_RF_internal_inloc_data_1_30_port, 
      DataPath_RF_internal_inloc_data_1_31_port, 
      DataPath_RF_internal_inloc_data_0_0_port, 
      DataPath_RF_internal_inloc_data_0_1_port, 
      DataPath_RF_internal_inloc_data_0_2_port, 
      DataPath_RF_internal_inloc_data_0_3_port, 
      DataPath_RF_internal_inloc_data_0_4_port, 
      DataPath_RF_internal_inloc_data_0_5_port, 
      DataPath_RF_internal_inloc_data_0_6_port, 
      DataPath_RF_internal_inloc_data_0_7_port, 
      DataPath_RF_internal_inloc_data_0_8_port, 
      DataPath_RF_internal_inloc_data_0_9_port, 
      DataPath_RF_internal_inloc_data_0_10_port, 
      DataPath_RF_internal_inloc_data_0_11_port, 
      DataPath_RF_internal_inloc_data_0_12_port, 
      DataPath_RF_internal_inloc_data_0_13_port, 
      DataPath_RF_internal_inloc_data_0_14_port, 
      DataPath_RF_internal_inloc_data_0_15_port, 
      DataPath_RF_internal_inloc_data_0_16_port, 
      DataPath_RF_internal_inloc_data_0_17_port, 
      DataPath_RF_internal_inloc_data_0_18_port, 
      DataPath_RF_internal_inloc_data_0_19_port, 
      DataPath_RF_internal_inloc_data_0_20_port, 
      DataPath_RF_internal_inloc_data_0_21_port, 
      DataPath_RF_internal_inloc_data_0_22_port, 
      DataPath_RF_internal_inloc_data_0_23_port, 
      DataPath_RF_internal_inloc_data_0_24_port, 
      DataPath_RF_internal_inloc_data_0_25_port, 
      DataPath_RF_internal_inloc_data_0_26_port, 
      DataPath_RF_internal_inloc_data_0_27_port, 
      DataPath_RF_internal_inloc_data_0_28_port, 
      DataPath_RF_internal_inloc_data_0_29_port, 
      DataPath_RF_internal_inloc_data_0_30_port, 
      DataPath_RF_internal_inloc_data_0_31_port, 
      DataPath_RF_c_swin_masked_1bit_4_0_port, 
      DataPath_RF_c_swin_masked_1bit_3_0_port, 
      DataPath_RF_c_swin_masked_1bit_2_0_port, 
      DataPath_RF_c_swin_masked_1bit_1_0_port, 
      DataPath_RF_c_swin_masked_1bit_0_0_port, DataPath_RF_en_regi_8_port, 
      DataPath_RF_en_regi_9_port, DataPath_RF_en_regi_10_port, 
      DataPath_RF_en_regi_11_port, DataPath_RF_en_regi_12_port, 
      DataPath_RF_en_regi_13_port, DataPath_RF_en_regi_14_port, 
      DataPath_RF_en_regi_15_port, DataPath_RF_en_regi_16_port, 
      DataPath_RF_en_regi_17_port, DataPath_RF_en_regi_18_port, 
      DataPath_RF_en_regi_19_port, DataPath_RF_en_regi_20_port, 
      DataPath_RF_en_regi_21_port, DataPath_RF_en_regi_22_port, 
      DataPath_RF_en_regi_23_port, DataPath_RF_en_regi_24_port, 
      DataPath_RF_en_regi_25_port, DataPath_RF_en_regi_26_port, 
      DataPath_RF_en_regi_27_port, DataPath_RF_en_regi_28_port, 
      DataPath_RF_en_regi_29_port, DataPath_RF_en_regi_30_port, 
      DataPath_RF_en_regi_31_port, DataPath_RF_en_regi_32_port, 
      DataPath_RF_en_regi_33_port, DataPath_RF_en_regi_34_port, 
      DataPath_RF_en_regi_35_port, DataPath_RF_en_regi_36_port, 
      DataPath_RF_en_regi_37_port, DataPath_RF_en_regi_38_port, 
      DataPath_RF_en_regi_39_port, DataPath_RF_en_regi_40_port, 
      DataPath_RF_en_regi_41_port, DataPath_RF_en_regi_42_port, 
      DataPath_RF_en_regi_43_port, DataPath_RF_en_regi_44_port, 
      DataPath_RF_en_regi_45_port, DataPath_RF_en_regi_46_port, 
      DataPath_RF_en_regi_47_port, DataPath_RF_en_regi_48_port, 
      DataPath_RF_en_regi_49_port, DataPath_RF_en_regi_50_port, 
      DataPath_RF_en_regi_51_port, DataPath_RF_en_regi_52_port, 
      DataPath_RF_en_regi_53_port, DataPath_RF_en_regi_54_port, 
      DataPath_RF_en_regi_55_port, DataPath_RF_en_regi_56_port, 
      DataPath_RF_en_regi_57_port, DataPath_RF_en_regi_58_port, 
      DataPath_RF_en_regi_59_port, DataPath_RF_en_regi_60_port, 
      DataPath_RF_en_regi_61_port, DataPath_RF_en_regi_62_port, 
      DataPath_RF_en_regi_63_port, DataPath_RF_en_regi_64_port, 
      DataPath_RF_en_regi_65_port, DataPath_RF_en_regi_66_port, 
      DataPath_RF_en_regi_67_port, DataPath_RF_en_regi_68_port, 
      DataPath_RF_en_regi_69_port, DataPath_RF_en_regi_70_port, 
      DataPath_RF_en_regi_71_port, DataPath_RF_en_regi_72_port, 
      DataPath_RF_en_regi_73_port, DataPath_RF_en_regi_74_port, 
      DataPath_RF_en_regi_75_port, DataPath_RF_en_regi_76_port, 
      DataPath_RF_en_regi_77_port, DataPath_RF_en_regi_78_port, 
      DataPath_RF_en_regi_79_port, DataPath_RF_en_regi_80_port, 
      DataPath_RF_en_regi_81_port, DataPath_RF_en_regi_82_port, 
      DataPath_RF_en_regi_83_port, DataPath_RF_en_regi_84_port, 
      DataPath_RF_en_regi_85_port, DataPath_RF_en_regi_86_port, 
      DataPath_RF_en_regi_87_port, DataPath_RF_bus_reg_dataout_0_port, 
      DataPath_RF_bus_reg_dataout_1_port, DataPath_RF_bus_reg_dataout_2_port, 
      DataPath_RF_bus_reg_dataout_3_port, DataPath_RF_bus_reg_dataout_4_port, 
      DataPath_RF_bus_reg_dataout_5_port, DataPath_RF_bus_reg_dataout_6_port, 
      DataPath_RF_bus_reg_dataout_7_port, DataPath_RF_bus_reg_dataout_8_port, 
      DataPath_RF_bus_reg_dataout_9_port, DataPath_RF_bus_reg_dataout_10_port, 
      DataPath_RF_bus_reg_dataout_11_port, DataPath_RF_bus_reg_dataout_12_port,
      DataPath_RF_bus_reg_dataout_13_port, DataPath_RF_bus_reg_dataout_14_port,
      DataPath_RF_bus_reg_dataout_15_port, DataPath_RF_bus_reg_dataout_16_port,
      DataPath_RF_bus_reg_dataout_17_port, DataPath_RF_bus_reg_dataout_18_port,
      DataPath_RF_bus_reg_dataout_19_port, DataPath_RF_bus_reg_dataout_20_port,
      DataPath_RF_bus_reg_dataout_21_port, DataPath_RF_bus_reg_dataout_22_port,
      DataPath_RF_bus_reg_dataout_23_port, DataPath_RF_bus_reg_dataout_24_port,
      DataPath_RF_bus_reg_dataout_25_port, DataPath_RF_bus_reg_dataout_26_port,
      DataPath_RF_bus_reg_dataout_27_port, DataPath_RF_bus_reg_dataout_28_port,
      DataPath_RF_bus_reg_dataout_29_port, DataPath_RF_bus_reg_dataout_30_port,
      DataPath_RF_bus_reg_dataout_31_port, DataPath_RF_bus_reg_dataout_32_port,
      DataPath_RF_bus_reg_dataout_33_port, DataPath_RF_bus_reg_dataout_34_port,
      DataPath_RF_bus_reg_dataout_35_port, DataPath_RF_bus_reg_dataout_36_port,
      DataPath_RF_bus_reg_dataout_37_port, DataPath_RF_bus_reg_dataout_38_port,
      DataPath_RF_bus_reg_dataout_39_port, DataPath_RF_bus_reg_dataout_40_port,
      DataPath_RF_bus_reg_dataout_41_port, DataPath_RF_bus_reg_dataout_42_port,
      DataPath_RF_bus_reg_dataout_43_port, DataPath_RF_bus_reg_dataout_44_port,
      DataPath_RF_bus_reg_dataout_45_port, DataPath_RF_bus_reg_dataout_46_port,
      DataPath_RF_bus_reg_dataout_47_port, DataPath_RF_bus_reg_dataout_48_port,
      DataPath_RF_bus_reg_dataout_49_port, DataPath_RF_bus_reg_dataout_50_port,
      DataPath_RF_bus_reg_dataout_51_port, DataPath_RF_bus_reg_dataout_52_port,
      DataPath_RF_bus_reg_dataout_53_port, DataPath_RF_bus_reg_dataout_54_port,
      DataPath_RF_bus_reg_dataout_55_port, DataPath_RF_bus_reg_dataout_56_port,
      DataPath_RF_bus_reg_dataout_57_port, DataPath_RF_bus_reg_dataout_58_port,
      DataPath_RF_bus_reg_dataout_59_port, DataPath_RF_bus_reg_dataout_60_port,
      DataPath_RF_bus_reg_dataout_61_port, DataPath_RF_bus_reg_dataout_62_port,
      DataPath_RF_bus_reg_dataout_63_port, DataPath_RF_bus_reg_dataout_64_port,
      DataPath_RF_bus_reg_dataout_65_port, DataPath_RF_bus_reg_dataout_66_port,
      DataPath_RF_bus_reg_dataout_67_port, DataPath_RF_bus_reg_dataout_68_port,
      DataPath_RF_bus_reg_dataout_69_port, DataPath_RF_bus_reg_dataout_70_port,
      DataPath_RF_bus_reg_dataout_71_port, DataPath_RF_bus_reg_dataout_72_port,
      DataPath_RF_bus_reg_dataout_73_port, DataPath_RF_bus_reg_dataout_74_port,
      DataPath_RF_bus_reg_dataout_75_port, DataPath_RF_bus_reg_dataout_76_port,
      DataPath_RF_bus_reg_dataout_77_port, DataPath_RF_bus_reg_dataout_78_port,
      DataPath_RF_bus_reg_dataout_79_port, DataPath_RF_bus_reg_dataout_80_port,
      DataPath_RF_bus_reg_dataout_81_port, DataPath_RF_bus_reg_dataout_82_port,
      DataPath_RF_bus_reg_dataout_83_port, DataPath_RF_bus_reg_dataout_84_port,
      DataPath_RF_bus_reg_dataout_85_port, DataPath_RF_bus_reg_dataout_86_port,
      DataPath_RF_bus_reg_dataout_87_port, DataPath_RF_bus_reg_dataout_88_port,
      DataPath_RF_bus_reg_dataout_89_port, DataPath_RF_bus_reg_dataout_90_port,
      DataPath_RF_bus_reg_dataout_91_port, DataPath_RF_bus_reg_dataout_92_port,
      DataPath_RF_bus_reg_dataout_93_port, DataPath_RF_bus_reg_dataout_94_port,
      DataPath_RF_bus_reg_dataout_95_port, DataPath_RF_bus_reg_dataout_96_port,
      DataPath_RF_bus_reg_dataout_97_port, DataPath_RF_bus_reg_dataout_98_port,
      DataPath_RF_bus_reg_dataout_99_port, DataPath_RF_bus_reg_dataout_100_port
      , DataPath_RF_bus_reg_dataout_101_port, 
      DataPath_RF_bus_reg_dataout_102_port, 
      DataPath_RF_bus_reg_dataout_103_port, 
      DataPath_RF_bus_reg_dataout_104_port, 
      DataPath_RF_bus_reg_dataout_105_port, 
      DataPath_RF_bus_reg_dataout_106_port, 
      DataPath_RF_bus_reg_dataout_107_port, 
      DataPath_RF_bus_reg_dataout_108_port, 
      DataPath_RF_bus_reg_dataout_109_port, 
      DataPath_RF_bus_reg_dataout_110_port, 
      DataPath_RF_bus_reg_dataout_111_port, 
      DataPath_RF_bus_reg_dataout_112_port, 
      DataPath_RF_bus_reg_dataout_113_port, 
      DataPath_RF_bus_reg_dataout_114_port, 
      DataPath_RF_bus_reg_dataout_115_port, 
      DataPath_RF_bus_reg_dataout_116_port, 
      DataPath_RF_bus_reg_dataout_117_port, 
      DataPath_RF_bus_reg_dataout_118_port, 
      DataPath_RF_bus_reg_dataout_119_port, 
      DataPath_RF_bus_reg_dataout_120_port, 
      DataPath_RF_bus_reg_dataout_121_port, 
      DataPath_RF_bus_reg_dataout_122_port, 
      DataPath_RF_bus_reg_dataout_123_port, 
      DataPath_RF_bus_reg_dataout_124_port, 
      DataPath_RF_bus_reg_dataout_125_port, 
      DataPath_RF_bus_reg_dataout_126_port, 
      DataPath_RF_bus_reg_dataout_127_port, 
      DataPath_RF_bus_reg_dataout_128_port, 
      DataPath_RF_bus_reg_dataout_129_port, 
      DataPath_RF_bus_reg_dataout_130_port, 
      DataPath_RF_bus_reg_dataout_131_port, 
      DataPath_RF_bus_reg_dataout_132_port, 
      DataPath_RF_bus_reg_dataout_133_port, 
      DataPath_RF_bus_reg_dataout_134_port, 
      DataPath_RF_bus_reg_dataout_135_port, 
      DataPath_RF_bus_reg_dataout_136_port, 
      DataPath_RF_bus_reg_dataout_137_port, 
      DataPath_RF_bus_reg_dataout_138_port, 
      DataPath_RF_bus_reg_dataout_139_port, 
      DataPath_RF_bus_reg_dataout_140_port, 
      DataPath_RF_bus_reg_dataout_141_port, 
      DataPath_RF_bus_reg_dataout_142_port, 
      DataPath_RF_bus_reg_dataout_143_port, 
      DataPath_RF_bus_reg_dataout_144_port, 
      DataPath_RF_bus_reg_dataout_145_port, 
      DataPath_RF_bus_reg_dataout_146_port, 
      DataPath_RF_bus_reg_dataout_147_port, 
      DataPath_RF_bus_reg_dataout_148_port, 
      DataPath_RF_bus_reg_dataout_149_port, 
      DataPath_RF_bus_reg_dataout_150_port, 
      DataPath_RF_bus_reg_dataout_151_port, 
      DataPath_RF_bus_reg_dataout_152_port, 
      DataPath_RF_bus_reg_dataout_153_port, 
      DataPath_RF_bus_reg_dataout_154_port, 
      DataPath_RF_bus_reg_dataout_155_port, 
      DataPath_RF_bus_reg_dataout_156_port, 
      DataPath_RF_bus_reg_dataout_157_port, 
      DataPath_RF_bus_reg_dataout_158_port, 
      DataPath_RF_bus_reg_dataout_159_port, 
      DataPath_RF_bus_reg_dataout_160_port, 
      DataPath_RF_bus_reg_dataout_161_port, 
      DataPath_RF_bus_reg_dataout_162_port, 
      DataPath_RF_bus_reg_dataout_163_port, 
      DataPath_RF_bus_reg_dataout_164_port, 
      DataPath_RF_bus_reg_dataout_165_port, 
      DataPath_RF_bus_reg_dataout_166_port, 
      DataPath_RF_bus_reg_dataout_167_port, 
      DataPath_RF_bus_reg_dataout_168_port, 
      DataPath_RF_bus_reg_dataout_169_port, 
      DataPath_RF_bus_reg_dataout_170_port, 
      DataPath_RF_bus_reg_dataout_171_port, 
      DataPath_RF_bus_reg_dataout_172_port, 
      DataPath_RF_bus_reg_dataout_173_port, 
      DataPath_RF_bus_reg_dataout_174_port, 
      DataPath_RF_bus_reg_dataout_175_port, 
      DataPath_RF_bus_reg_dataout_176_port, 
      DataPath_RF_bus_reg_dataout_177_port, 
      DataPath_RF_bus_reg_dataout_178_port, 
      DataPath_RF_bus_reg_dataout_179_port, 
      DataPath_RF_bus_reg_dataout_180_port, 
      DataPath_RF_bus_reg_dataout_181_port, 
      DataPath_RF_bus_reg_dataout_182_port, 
      DataPath_RF_bus_reg_dataout_183_port, 
      DataPath_RF_bus_reg_dataout_184_port, 
      DataPath_RF_bus_reg_dataout_185_port, 
      DataPath_RF_bus_reg_dataout_186_port, 
      DataPath_RF_bus_reg_dataout_187_port, 
      DataPath_RF_bus_reg_dataout_188_port, 
      DataPath_RF_bus_reg_dataout_189_port, 
      DataPath_RF_bus_reg_dataout_190_port, 
      DataPath_RF_bus_reg_dataout_191_port, 
      DataPath_RF_bus_reg_dataout_192_port, 
      DataPath_RF_bus_reg_dataout_193_port, 
      DataPath_RF_bus_reg_dataout_194_port, 
      DataPath_RF_bus_reg_dataout_195_port, 
      DataPath_RF_bus_reg_dataout_196_port, 
      DataPath_RF_bus_reg_dataout_197_port, 
      DataPath_RF_bus_reg_dataout_198_port, 
      DataPath_RF_bus_reg_dataout_199_port, 
      DataPath_RF_bus_reg_dataout_200_port, 
      DataPath_RF_bus_reg_dataout_201_port, 
      DataPath_RF_bus_reg_dataout_202_port, 
      DataPath_RF_bus_reg_dataout_203_port, 
      DataPath_RF_bus_reg_dataout_204_port, 
      DataPath_RF_bus_reg_dataout_205_port, 
      DataPath_RF_bus_reg_dataout_206_port, 
      DataPath_RF_bus_reg_dataout_207_port, 
      DataPath_RF_bus_reg_dataout_208_port, 
      DataPath_RF_bus_reg_dataout_209_port, 
      DataPath_RF_bus_reg_dataout_210_port, 
      DataPath_RF_bus_reg_dataout_211_port, 
      DataPath_RF_bus_reg_dataout_212_port, 
      DataPath_RF_bus_reg_dataout_213_port, 
      DataPath_RF_bus_reg_dataout_214_port, 
      DataPath_RF_bus_reg_dataout_215_port, 
      DataPath_RF_bus_reg_dataout_216_port, 
      DataPath_RF_bus_reg_dataout_217_port, 
      DataPath_RF_bus_reg_dataout_218_port, 
      DataPath_RF_bus_reg_dataout_219_port, 
      DataPath_RF_bus_reg_dataout_220_port, 
      DataPath_RF_bus_reg_dataout_221_port, 
      DataPath_RF_bus_reg_dataout_222_port, 
      DataPath_RF_bus_reg_dataout_223_port, 
      DataPath_RF_bus_reg_dataout_224_port, 
      DataPath_RF_bus_reg_dataout_225_port, 
      DataPath_RF_bus_reg_dataout_226_port, 
      DataPath_RF_bus_reg_dataout_227_port, 
      DataPath_RF_bus_reg_dataout_228_port, 
      DataPath_RF_bus_reg_dataout_229_port, 
      DataPath_RF_bus_reg_dataout_230_port, 
      DataPath_RF_bus_reg_dataout_231_port, 
      DataPath_RF_bus_reg_dataout_232_port, 
      DataPath_RF_bus_reg_dataout_233_port, 
      DataPath_RF_bus_reg_dataout_234_port, 
      DataPath_RF_bus_reg_dataout_235_port, 
      DataPath_RF_bus_reg_dataout_236_port, 
      DataPath_RF_bus_reg_dataout_237_port, 
      DataPath_RF_bus_reg_dataout_238_port, 
      DataPath_RF_bus_reg_dataout_239_port, 
      DataPath_RF_bus_reg_dataout_240_port, 
      DataPath_RF_bus_reg_dataout_241_port, 
      DataPath_RF_bus_reg_dataout_242_port, 
      DataPath_RF_bus_reg_dataout_243_port, 
      DataPath_RF_bus_reg_dataout_244_port, 
      DataPath_RF_bus_reg_dataout_245_port, 
      DataPath_RF_bus_reg_dataout_246_port, 
      DataPath_RF_bus_reg_dataout_247_port, 
      DataPath_RF_bus_reg_dataout_248_port, 
      DataPath_RF_bus_reg_dataout_249_port, 
      DataPath_RF_bus_reg_dataout_250_port, 
      DataPath_RF_bus_reg_dataout_251_port, 
      DataPath_RF_bus_reg_dataout_252_port, 
      DataPath_RF_bus_reg_dataout_253_port, 
      DataPath_RF_bus_reg_dataout_254_port, 
      DataPath_RF_bus_reg_dataout_255_port, 
      DataPath_RF_bus_reg_dataout_256_port, 
      DataPath_RF_bus_reg_dataout_257_port, 
      DataPath_RF_bus_reg_dataout_258_port, 
      DataPath_RF_bus_reg_dataout_259_port, 
      DataPath_RF_bus_reg_dataout_260_port, 
      DataPath_RF_bus_reg_dataout_261_port, 
      DataPath_RF_bus_reg_dataout_262_port, 
      DataPath_RF_bus_reg_dataout_263_port, 
      DataPath_RF_bus_reg_dataout_264_port, 
      DataPath_RF_bus_reg_dataout_265_port, 
      DataPath_RF_bus_reg_dataout_266_port, 
      DataPath_RF_bus_reg_dataout_267_port, 
      DataPath_RF_bus_reg_dataout_268_port, 
      DataPath_RF_bus_reg_dataout_269_port, 
      DataPath_RF_bus_reg_dataout_270_port, 
      DataPath_RF_bus_reg_dataout_271_port, 
      DataPath_RF_bus_reg_dataout_272_port, 
      DataPath_RF_bus_reg_dataout_273_port, 
      DataPath_RF_bus_reg_dataout_274_port, 
      DataPath_RF_bus_reg_dataout_275_port, 
      DataPath_RF_bus_reg_dataout_276_port, 
      DataPath_RF_bus_reg_dataout_277_port, 
      DataPath_RF_bus_reg_dataout_278_port, 
      DataPath_RF_bus_reg_dataout_279_port, 
      DataPath_RF_bus_reg_dataout_280_port, 
      DataPath_RF_bus_reg_dataout_281_port, 
      DataPath_RF_bus_reg_dataout_282_port, 
      DataPath_RF_bus_reg_dataout_283_port, 
      DataPath_RF_bus_reg_dataout_284_port, 
      DataPath_RF_bus_reg_dataout_285_port, 
      DataPath_RF_bus_reg_dataout_286_port, 
      DataPath_RF_bus_reg_dataout_287_port, 
      DataPath_RF_bus_reg_dataout_288_port, 
      DataPath_RF_bus_reg_dataout_289_port, 
      DataPath_RF_bus_reg_dataout_290_port, 
      DataPath_RF_bus_reg_dataout_291_port, 
      DataPath_RF_bus_reg_dataout_292_port, 
      DataPath_RF_bus_reg_dataout_293_port, 
      DataPath_RF_bus_reg_dataout_294_port, 
      DataPath_RF_bus_reg_dataout_295_port, 
      DataPath_RF_bus_reg_dataout_296_port, 
      DataPath_RF_bus_reg_dataout_297_port, 
      DataPath_RF_bus_reg_dataout_298_port, 
      DataPath_RF_bus_reg_dataout_299_port, 
      DataPath_RF_bus_reg_dataout_300_port, 
      DataPath_RF_bus_reg_dataout_301_port, 
      DataPath_RF_bus_reg_dataout_302_port, 
      DataPath_RF_bus_reg_dataout_303_port, 
      DataPath_RF_bus_reg_dataout_304_port, 
      DataPath_RF_bus_reg_dataout_305_port, 
      DataPath_RF_bus_reg_dataout_306_port, 
      DataPath_RF_bus_reg_dataout_307_port, 
      DataPath_RF_bus_reg_dataout_308_port, 
      DataPath_RF_bus_reg_dataout_309_port, 
      DataPath_RF_bus_reg_dataout_310_port, 
      DataPath_RF_bus_reg_dataout_311_port, 
      DataPath_RF_bus_reg_dataout_312_port, 
      DataPath_RF_bus_reg_dataout_313_port, 
      DataPath_RF_bus_reg_dataout_314_port, 
      DataPath_RF_bus_reg_dataout_315_port, 
      DataPath_RF_bus_reg_dataout_316_port, 
      DataPath_RF_bus_reg_dataout_317_port, 
      DataPath_RF_bus_reg_dataout_318_port, 
      DataPath_RF_bus_reg_dataout_319_port, 
      DataPath_RF_bus_reg_dataout_320_port, 
      DataPath_RF_bus_reg_dataout_321_port, 
      DataPath_RF_bus_reg_dataout_322_port, 
      DataPath_RF_bus_reg_dataout_323_port, 
      DataPath_RF_bus_reg_dataout_324_port, 
      DataPath_RF_bus_reg_dataout_325_port, 
      DataPath_RF_bus_reg_dataout_326_port, 
      DataPath_RF_bus_reg_dataout_327_port, 
      DataPath_RF_bus_reg_dataout_328_port, 
      DataPath_RF_bus_reg_dataout_329_port, 
      DataPath_RF_bus_reg_dataout_330_port, 
      DataPath_RF_bus_reg_dataout_331_port, 
      DataPath_RF_bus_reg_dataout_332_port, 
      DataPath_RF_bus_reg_dataout_333_port, 
      DataPath_RF_bus_reg_dataout_334_port, 
      DataPath_RF_bus_reg_dataout_335_port, 
      DataPath_RF_bus_reg_dataout_336_port, 
      DataPath_RF_bus_reg_dataout_337_port, 
      DataPath_RF_bus_reg_dataout_338_port, 
      DataPath_RF_bus_reg_dataout_339_port, 
      DataPath_RF_bus_reg_dataout_340_port, 
      DataPath_RF_bus_reg_dataout_341_port, 
      DataPath_RF_bus_reg_dataout_342_port, 
      DataPath_RF_bus_reg_dataout_343_port, 
      DataPath_RF_bus_reg_dataout_344_port, 
      DataPath_RF_bus_reg_dataout_345_port, 
      DataPath_RF_bus_reg_dataout_346_port, 
      DataPath_RF_bus_reg_dataout_347_port, 
      DataPath_RF_bus_reg_dataout_348_port, 
      DataPath_RF_bus_reg_dataout_349_port, 
      DataPath_RF_bus_reg_dataout_350_port, 
      DataPath_RF_bus_reg_dataout_351_port, 
      DataPath_RF_bus_reg_dataout_352_port, 
      DataPath_RF_bus_reg_dataout_353_port, 
      DataPath_RF_bus_reg_dataout_354_port, 
      DataPath_RF_bus_reg_dataout_355_port, 
      DataPath_RF_bus_reg_dataout_356_port, 
      DataPath_RF_bus_reg_dataout_357_port, 
      DataPath_RF_bus_reg_dataout_358_port, 
      DataPath_RF_bus_reg_dataout_359_port, 
      DataPath_RF_bus_reg_dataout_360_port, 
      DataPath_RF_bus_reg_dataout_361_port, 
      DataPath_RF_bus_reg_dataout_362_port, 
      DataPath_RF_bus_reg_dataout_363_port, 
      DataPath_RF_bus_reg_dataout_364_port, 
      DataPath_RF_bus_reg_dataout_365_port, 
      DataPath_RF_bus_reg_dataout_366_port, 
      DataPath_RF_bus_reg_dataout_367_port, 
      DataPath_RF_bus_reg_dataout_368_port, 
      DataPath_RF_bus_reg_dataout_369_port, 
      DataPath_RF_bus_reg_dataout_370_port, 
      DataPath_RF_bus_reg_dataout_371_port, 
      DataPath_RF_bus_reg_dataout_372_port, 
      DataPath_RF_bus_reg_dataout_373_port, 
      DataPath_RF_bus_reg_dataout_374_port, 
      DataPath_RF_bus_reg_dataout_375_port, 
      DataPath_RF_bus_reg_dataout_376_port, 
      DataPath_RF_bus_reg_dataout_377_port, 
      DataPath_RF_bus_reg_dataout_378_port, 
      DataPath_RF_bus_reg_dataout_379_port, 
      DataPath_RF_bus_reg_dataout_380_port, 
      DataPath_RF_bus_reg_dataout_381_port, 
      DataPath_RF_bus_reg_dataout_382_port, 
      DataPath_RF_bus_reg_dataout_383_port, 
      DataPath_RF_bus_reg_dataout_384_port, 
      DataPath_RF_bus_reg_dataout_385_port, 
      DataPath_RF_bus_reg_dataout_386_port, 
      DataPath_RF_bus_reg_dataout_387_port, 
      DataPath_RF_bus_reg_dataout_388_port, 
      DataPath_RF_bus_reg_dataout_389_port, 
      DataPath_RF_bus_reg_dataout_390_port, 
      DataPath_RF_bus_reg_dataout_391_port, 
      DataPath_RF_bus_reg_dataout_392_port, 
      DataPath_RF_bus_reg_dataout_393_port, 
      DataPath_RF_bus_reg_dataout_394_port, 
      DataPath_RF_bus_reg_dataout_395_port, 
      DataPath_RF_bus_reg_dataout_396_port, 
      DataPath_RF_bus_reg_dataout_397_port, 
      DataPath_RF_bus_reg_dataout_398_port, 
      DataPath_RF_bus_reg_dataout_399_port, 
      DataPath_RF_bus_reg_dataout_400_port, 
      DataPath_RF_bus_reg_dataout_401_port, 
      DataPath_RF_bus_reg_dataout_402_port, 
      DataPath_RF_bus_reg_dataout_403_port, 
      DataPath_RF_bus_reg_dataout_404_port, 
      DataPath_RF_bus_reg_dataout_405_port, 
      DataPath_RF_bus_reg_dataout_406_port, 
      DataPath_RF_bus_reg_dataout_407_port, 
      DataPath_RF_bus_reg_dataout_408_port, 
      DataPath_RF_bus_reg_dataout_409_port, 
      DataPath_RF_bus_reg_dataout_410_port, 
      DataPath_RF_bus_reg_dataout_411_port, 
      DataPath_RF_bus_reg_dataout_412_port, 
      DataPath_RF_bus_reg_dataout_413_port, 
      DataPath_RF_bus_reg_dataout_414_port, 
      DataPath_RF_bus_reg_dataout_415_port, 
      DataPath_RF_bus_reg_dataout_416_port, 
      DataPath_RF_bus_reg_dataout_417_port, 
      DataPath_RF_bus_reg_dataout_418_port, 
      DataPath_RF_bus_reg_dataout_419_port, 
      DataPath_RF_bus_reg_dataout_420_port, 
      DataPath_RF_bus_reg_dataout_421_port, 
      DataPath_RF_bus_reg_dataout_422_port, 
      DataPath_RF_bus_reg_dataout_423_port, 
      DataPath_RF_bus_reg_dataout_424_port, 
      DataPath_RF_bus_reg_dataout_425_port, 
      DataPath_RF_bus_reg_dataout_426_port, 
      DataPath_RF_bus_reg_dataout_427_port, 
      DataPath_RF_bus_reg_dataout_428_port, 
      DataPath_RF_bus_reg_dataout_429_port, 
      DataPath_RF_bus_reg_dataout_430_port, 
      DataPath_RF_bus_reg_dataout_431_port, 
      DataPath_RF_bus_reg_dataout_432_port, 
      DataPath_RF_bus_reg_dataout_433_port, 
      DataPath_RF_bus_reg_dataout_434_port, 
      DataPath_RF_bus_reg_dataout_435_port, 
      DataPath_RF_bus_reg_dataout_436_port, 
      DataPath_RF_bus_reg_dataout_437_port, 
      DataPath_RF_bus_reg_dataout_438_port, 
      DataPath_RF_bus_reg_dataout_439_port, 
      DataPath_RF_bus_reg_dataout_440_port, 
      DataPath_RF_bus_reg_dataout_441_port, 
      DataPath_RF_bus_reg_dataout_442_port, 
      DataPath_RF_bus_reg_dataout_443_port, 
      DataPath_RF_bus_reg_dataout_444_port, 
      DataPath_RF_bus_reg_dataout_445_port, 
      DataPath_RF_bus_reg_dataout_446_port, 
      DataPath_RF_bus_reg_dataout_447_port, 
      DataPath_RF_bus_reg_dataout_448_port, 
      DataPath_RF_bus_reg_dataout_449_port, 
      DataPath_RF_bus_reg_dataout_450_port, 
      DataPath_RF_bus_reg_dataout_451_port, 
      DataPath_RF_bus_reg_dataout_452_port, 
      DataPath_RF_bus_reg_dataout_453_port, 
      DataPath_RF_bus_reg_dataout_454_port, 
      DataPath_RF_bus_reg_dataout_455_port, 
      DataPath_RF_bus_reg_dataout_456_port, 
      DataPath_RF_bus_reg_dataout_457_port, 
      DataPath_RF_bus_reg_dataout_458_port, 
      DataPath_RF_bus_reg_dataout_459_port, 
      DataPath_RF_bus_reg_dataout_460_port, 
      DataPath_RF_bus_reg_dataout_461_port, 
      DataPath_RF_bus_reg_dataout_462_port, 
      DataPath_RF_bus_reg_dataout_463_port, 
      DataPath_RF_bus_reg_dataout_464_port, 
      DataPath_RF_bus_reg_dataout_465_port, 
      DataPath_RF_bus_reg_dataout_466_port, 
      DataPath_RF_bus_reg_dataout_467_port, 
      DataPath_RF_bus_reg_dataout_468_port, 
      DataPath_RF_bus_reg_dataout_469_port, 
      DataPath_RF_bus_reg_dataout_470_port, 
      DataPath_RF_bus_reg_dataout_471_port, 
      DataPath_RF_bus_reg_dataout_472_port, 
      DataPath_RF_bus_reg_dataout_473_port, 
      DataPath_RF_bus_reg_dataout_474_port, 
      DataPath_RF_bus_reg_dataout_475_port, 
      DataPath_RF_bus_reg_dataout_476_port, 
      DataPath_RF_bus_reg_dataout_477_port, 
      DataPath_RF_bus_reg_dataout_478_port, 
      DataPath_RF_bus_reg_dataout_479_port, 
      DataPath_RF_bus_reg_dataout_480_port, 
      DataPath_RF_bus_reg_dataout_481_port, 
      DataPath_RF_bus_reg_dataout_482_port, 
      DataPath_RF_bus_reg_dataout_483_port, 
      DataPath_RF_bus_reg_dataout_484_port, 
      DataPath_RF_bus_reg_dataout_485_port, 
      DataPath_RF_bus_reg_dataout_486_port, 
      DataPath_RF_bus_reg_dataout_487_port, 
      DataPath_RF_bus_reg_dataout_488_port, 
      DataPath_RF_bus_reg_dataout_489_port, 
      DataPath_RF_bus_reg_dataout_490_port, 
      DataPath_RF_bus_reg_dataout_491_port, 
      DataPath_RF_bus_reg_dataout_492_port, 
      DataPath_RF_bus_reg_dataout_493_port, 
      DataPath_RF_bus_reg_dataout_494_port, 
      DataPath_RF_bus_reg_dataout_495_port, 
      DataPath_RF_bus_reg_dataout_496_port, 
      DataPath_RF_bus_reg_dataout_497_port, 
      DataPath_RF_bus_reg_dataout_498_port, 
      DataPath_RF_bus_reg_dataout_499_port, 
      DataPath_RF_bus_reg_dataout_500_port, 
      DataPath_RF_bus_reg_dataout_501_port, 
      DataPath_RF_bus_reg_dataout_502_port, 
      DataPath_RF_bus_reg_dataout_503_port, 
      DataPath_RF_bus_reg_dataout_504_port, 
      DataPath_RF_bus_reg_dataout_505_port, 
      DataPath_RF_bus_reg_dataout_506_port, 
      DataPath_RF_bus_reg_dataout_507_port, 
      DataPath_RF_bus_reg_dataout_508_port, 
      DataPath_RF_bus_reg_dataout_509_port, 
      DataPath_RF_bus_reg_dataout_510_port, 
      DataPath_RF_bus_reg_dataout_511_port, 
      DataPath_RF_bus_reg_dataout_512_port, 
      DataPath_RF_bus_reg_dataout_513_port, 
      DataPath_RF_bus_reg_dataout_514_port, 
      DataPath_RF_bus_reg_dataout_515_port, 
      DataPath_RF_bus_reg_dataout_516_port, 
      DataPath_RF_bus_reg_dataout_517_port, 
      DataPath_RF_bus_reg_dataout_518_port, 
      DataPath_RF_bus_reg_dataout_519_port, 
      DataPath_RF_bus_reg_dataout_520_port, 
      DataPath_RF_bus_reg_dataout_521_port, 
      DataPath_RF_bus_reg_dataout_522_port, 
      DataPath_RF_bus_reg_dataout_523_port, 
      DataPath_RF_bus_reg_dataout_524_port, 
      DataPath_RF_bus_reg_dataout_525_port, 
      DataPath_RF_bus_reg_dataout_526_port, 
      DataPath_RF_bus_reg_dataout_527_port, 
      DataPath_RF_bus_reg_dataout_528_port, 
      DataPath_RF_bus_reg_dataout_529_port, 
      DataPath_RF_bus_reg_dataout_530_port, 
      DataPath_RF_bus_reg_dataout_531_port, 
      DataPath_RF_bus_reg_dataout_532_port, 
      DataPath_RF_bus_reg_dataout_533_port, 
      DataPath_RF_bus_reg_dataout_534_port, 
      DataPath_RF_bus_reg_dataout_535_port, 
      DataPath_RF_bus_reg_dataout_536_port, 
      DataPath_RF_bus_reg_dataout_537_port, 
      DataPath_RF_bus_reg_dataout_538_port, 
      DataPath_RF_bus_reg_dataout_539_port, 
      DataPath_RF_bus_reg_dataout_540_port, 
      DataPath_RF_bus_reg_dataout_541_port, 
      DataPath_RF_bus_reg_dataout_542_port, 
      DataPath_RF_bus_reg_dataout_543_port, 
      DataPath_RF_bus_reg_dataout_544_port, 
      DataPath_RF_bus_reg_dataout_545_port, 
      DataPath_RF_bus_reg_dataout_546_port, 
      DataPath_RF_bus_reg_dataout_547_port, 
      DataPath_RF_bus_reg_dataout_548_port, 
      DataPath_RF_bus_reg_dataout_549_port, 
      DataPath_RF_bus_reg_dataout_550_port, 
      DataPath_RF_bus_reg_dataout_551_port, 
      DataPath_RF_bus_reg_dataout_552_port, 
      DataPath_RF_bus_reg_dataout_553_port, 
      DataPath_RF_bus_reg_dataout_554_port, 
      DataPath_RF_bus_reg_dataout_555_port, 
      DataPath_RF_bus_reg_dataout_556_port, 
      DataPath_RF_bus_reg_dataout_557_port, 
      DataPath_RF_bus_reg_dataout_558_port, 
      DataPath_RF_bus_reg_dataout_559_port, 
      DataPath_RF_bus_reg_dataout_560_port, 
      DataPath_RF_bus_reg_dataout_561_port, 
      DataPath_RF_bus_reg_dataout_562_port, 
      DataPath_RF_bus_reg_dataout_563_port, 
      DataPath_RF_bus_reg_dataout_564_port, 
      DataPath_RF_bus_reg_dataout_565_port, 
      DataPath_RF_bus_reg_dataout_566_port, 
      DataPath_RF_bus_reg_dataout_567_port, 
      DataPath_RF_bus_reg_dataout_568_port, 
      DataPath_RF_bus_reg_dataout_569_port, 
      DataPath_RF_bus_reg_dataout_570_port, 
      DataPath_RF_bus_reg_dataout_571_port, 
      DataPath_RF_bus_reg_dataout_572_port, 
      DataPath_RF_bus_reg_dataout_573_port, 
      DataPath_RF_bus_reg_dataout_574_port, 
      DataPath_RF_bus_reg_dataout_575_port, 
      DataPath_RF_bus_reg_dataout_576_port, 
      DataPath_RF_bus_reg_dataout_577_port, 
      DataPath_RF_bus_reg_dataout_578_port, 
      DataPath_RF_bus_reg_dataout_579_port, 
      DataPath_RF_bus_reg_dataout_580_port, 
      DataPath_RF_bus_reg_dataout_581_port, 
      DataPath_RF_bus_reg_dataout_582_port, 
      DataPath_RF_bus_reg_dataout_583_port, 
      DataPath_RF_bus_reg_dataout_584_port, 
      DataPath_RF_bus_reg_dataout_585_port, 
      DataPath_RF_bus_reg_dataout_586_port, 
      DataPath_RF_bus_reg_dataout_587_port, 
      DataPath_RF_bus_reg_dataout_588_port, 
      DataPath_RF_bus_reg_dataout_589_port, 
      DataPath_RF_bus_reg_dataout_590_port, 
      DataPath_RF_bus_reg_dataout_591_port, 
      DataPath_RF_bus_reg_dataout_592_port, 
      DataPath_RF_bus_reg_dataout_593_port, 
      DataPath_RF_bus_reg_dataout_594_port, 
      DataPath_RF_bus_reg_dataout_595_port, 
      DataPath_RF_bus_reg_dataout_596_port, 
      DataPath_RF_bus_reg_dataout_597_port, 
      DataPath_RF_bus_reg_dataout_598_port, 
      DataPath_RF_bus_reg_dataout_599_port, 
      DataPath_RF_bus_reg_dataout_600_port, 
      DataPath_RF_bus_reg_dataout_601_port, 
      DataPath_RF_bus_reg_dataout_602_port, 
      DataPath_RF_bus_reg_dataout_603_port, 
      DataPath_RF_bus_reg_dataout_604_port, 
      DataPath_RF_bus_reg_dataout_605_port, 
      DataPath_RF_bus_reg_dataout_606_port, 
      DataPath_RF_bus_reg_dataout_607_port, 
      DataPath_RF_bus_reg_dataout_608_port, 
      DataPath_RF_bus_reg_dataout_609_port, 
      DataPath_RF_bus_reg_dataout_610_port, 
      DataPath_RF_bus_reg_dataout_611_port, 
      DataPath_RF_bus_reg_dataout_612_port, 
      DataPath_RF_bus_reg_dataout_613_port, 
      DataPath_RF_bus_reg_dataout_614_port, 
      DataPath_RF_bus_reg_dataout_615_port, 
      DataPath_RF_bus_reg_dataout_616_port, 
      DataPath_RF_bus_reg_dataout_617_port, 
      DataPath_RF_bus_reg_dataout_618_port, 
      DataPath_RF_bus_reg_dataout_619_port, 
      DataPath_RF_bus_reg_dataout_620_port, 
      DataPath_RF_bus_reg_dataout_621_port, 
      DataPath_RF_bus_reg_dataout_622_port, 
      DataPath_RF_bus_reg_dataout_623_port, 
      DataPath_RF_bus_reg_dataout_624_port, 
      DataPath_RF_bus_reg_dataout_625_port, 
      DataPath_RF_bus_reg_dataout_626_port, 
      DataPath_RF_bus_reg_dataout_627_port, 
      DataPath_RF_bus_reg_dataout_628_port, 
      DataPath_RF_bus_reg_dataout_629_port, 
      DataPath_RF_bus_reg_dataout_630_port, 
      DataPath_RF_bus_reg_dataout_631_port, 
      DataPath_RF_bus_reg_dataout_632_port, 
      DataPath_RF_bus_reg_dataout_633_port, 
      DataPath_RF_bus_reg_dataout_634_port, 
      DataPath_RF_bus_reg_dataout_635_port, 
      DataPath_RF_bus_reg_dataout_636_port, 
      DataPath_RF_bus_reg_dataout_637_port, 
      DataPath_RF_bus_reg_dataout_638_port, 
      DataPath_RF_bus_reg_dataout_639_port, 
      DataPath_RF_bus_reg_dataout_640_port, 
      DataPath_RF_bus_reg_dataout_641_port, 
      DataPath_RF_bus_reg_dataout_642_port, 
      DataPath_RF_bus_reg_dataout_643_port, 
      DataPath_RF_bus_reg_dataout_644_port, 
      DataPath_RF_bus_reg_dataout_645_port, 
      DataPath_RF_bus_reg_dataout_646_port, 
      DataPath_RF_bus_reg_dataout_647_port, 
      DataPath_RF_bus_reg_dataout_648_port, 
      DataPath_RF_bus_reg_dataout_649_port, 
      DataPath_RF_bus_reg_dataout_650_port, 
      DataPath_RF_bus_reg_dataout_651_port, 
      DataPath_RF_bus_reg_dataout_652_port, 
      DataPath_RF_bus_reg_dataout_653_port, 
      DataPath_RF_bus_reg_dataout_654_port, 
      DataPath_RF_bus_reg_dataout_655_port, 
      DataPath_RF_bus_reg_dataout_656_port, 
      DataPath_RF_bus_reg_dataout_657_port, 
      DataPath_RF_bus_reg_dataout_658_port, 
      DataPath_RF_bus_reg_dataout_659_port, 
      DataPath_RF_bus_reg_dataout_660_port, 
      DataPath_RF_bus_reg_dataout_661_port, 
      DataPath_RF_bus_reg_dataout_662_port, 
      DataPath_RF_bus_reg_dataout_663_port, 
      DataPath_RF_bus_reg_dataout_664_port, 
      DataPath_RF_bus_reg_dataout_665_port, 
      DataPath_RF_bus_reg_dataout_666_port, 
      DataPath_RF_bus_reg_dataout_667_port, 
      DataPath_RF_bus_reg_dataout_668_port, 
      DataPath_RF_bus_reg_dataout_669_port, 
      DataPath_RF_bus_reg_dataout_670_port, 
      DataPath_RF_bus_reg_dataout_671_port, 
      DataPath_RF_bus_reg_dataout_672_port, 
      DataPath_RF_bus_reg_dataout_673_port, 
      DataPath_RF_bus_reg_dataout_674_port, 
      DataPath_RF_bus_reg_dataout_675_port, 
      DataPath_RF_bus_reg_dataout_676_port, 
      DataPath_RF_bus_reg_dataout_677_port, 
      DataPath_RF_bus_reg_dataout_678_port, 
      DataPath_RF_bus_reg_dataout_679_port, 
      DataPath_RF_bus_reg_dataout_680_port, 
      DataPath_RF_bus_reg_dataout_681_port, 
      DataPath_RF_bus_reg_dataout_682_port, 
      DataPath_RF_bus_reg_dataout_683_port, 
      DataPath_RF_bus_reg_dataout_684_port, 
      DataPath_RF_bus_reg_dataout_685_port, 
      DataPath_RF_bus_reg_dataout_686_port, 
      DataPath_RF_bus_reg_dataout_687_port, 
      DataPath_RF_bus_reg_dataout_688_port, 
      DataPath_RF_bus_reg_dataout_689_port, 
      DataPath_RF_bus_reg_dataout_690_port, 
      DataPath_RF_bus_reg_dataout_691_port, 
      DataPath_RF_bus_reg_dataout_692_port, 
      DataPath_RF_bus_reg_dataout_693_port, 
      DataPath_RF_bus_reg_dataout_694_port, 
      DataPath_RF_bus_reg_dataout_695_port, 
      DataPath_RF_bus_reg_dataout_696_port, 
      DataPath_RF_bus_reg_dataout_697_port, 
      DataPath_RF_bus_reg_dataout_698_port, 
      DataPath_RF_bus_reg_dataout_699_port, 
      DataPath_RF_bus_reg_dataout_700_port, 
      DataPath_RF_bus_reg_dataout_701_port, 
      DataPath_RF_bus_reg_dataout_702_port, 
      DataPath_RF_bus_reg_dataout_703_port, 
      DataPath_RF_bus_reg_dataout_704_port, 
      DataPath_RF_bus_reg_dataout_705_port, 
      DataPath_RF_bus_reg_dataout_706_port, 
      DataPath_RF_bus_reg_dataout_707_port, 
      DataPath_RF_bus_reg_dataout_708_port, 
      DataPath_RF_bus_reg_dataout_709_port, 
      DataPath_RF_bus_reg_dataout_710_port, 
      DataPath_RF_bus_reg_dataout_711_port, 
      DataPath_RF_bus_reg_dataout_712_port, 
      DataPath_RF_bus_reg_dataout_713_port, 
      DataPath_RF_bus_reg_dataout_714_port, 
      DataPath_RF_bus_reg_dataout_715_port, 
      DataPath_RF_bus_reg_dataout_716_port, 
      DataPath_RF_bus_reg_dataout_717_port, 
      DataPath_RF_bus_reg_dataout_718_port, 
      DataPath_RF_bus_reg_dataout_719_port, 
      DataPath_RF_bus_reg_dataout_720_port, 
      DataPath_RF_bus_reg_dataout_721_port, 
      DataPath_RF_bus_reg_dataout_722_port, 
      DataPath_RF_bus_reg_dataout_723_port, 
      DataPath_RF_bus_reg_dataout_724_port, 
      DataPath_RF_bus_reg_dataout_725_port, 
      DataPath_RF_bus_reg_dataout_726_port, 
      DataPath_RF_bus_reg_dataout_727_port, 
      DataPath_RF_bus_reg_dataout_728_port, 
      DataPath_RF_bus_reg_dataout_729_port, 
      DataPath_RF_bus_reg_dataout_730_port, 
      DataPath_RF_bus_reg_dataout_731_port, 
      DataPath_RF_bus_reg_dataout_732_port, 
      DataPath_RF_bus_reg_dataout_733_port, 
      DataPath_RF_bus_reg_dataout_734_port, 
      DataPath_RF_bus_reg_dataout_735_port, 
      DataPath_RF_bus_reg_dataout_736_port, 
      DataPath_RF_bus_reg_dataout_737_port, 
      DataPath_RF_bus_reg_dataout_738_port, 
      DataPath_RF_bus_reg_dataout_739_port, 
      DataPath_RF_bus_reg_dataout_740_port, 
      DataPath_RF_bus_reg_dataout_741_port, 
      DataPath_RF_bus_reg_dataout_742_port, 
      DataPath_RF_bus_reg_dataout_743_port, 
      DataPath_RF_bus_reg_dataout_744_port, 
      DataPath_RF_bus_reg_dataout_745_port, 
      DataPath_RF_bus_reg_dataout_746_port, 
      DataPath_RF_bus_reg_dataout_747_port, 
      DataPath_RF_bus_reg_dataout_748_port, 
      DataPath_RF_bus_reg_dataout_749_port, 
      DataPath_RF_bus_reg_dataout_750_port, 
      DataPath_RF_bus_reg_dataout_751_port, 
      DataPath_RF_bus_reg_dataout_752_port, 
      DataPath_RF_bus_reg_dataout_753_port, 
      DataPath_RF_bus_reg_dataout_754_port, 
      DataPath_RF_bus_reg_dataout_755_port, 
      DataPath_RF_bus_reg_dataout_756_port, 
      DataPath_RF_bus_reg_dataout_757_port, 
      DataPath_RF_bus_reg_dataout_758_port, 
      DataPath_RF_bus_reg_dataout_759_port, 
      DataPath_RF_bus_reg_dataout_760_port, 
      DataPath_RF_bus_reg_dataout_761_port, 
      DataPath_RF_bus_reg_dataout_762_port, 
      DataPath_RF_bus_reg_dataout_763_port, 
      DataPath_RF_bus_reg_dataout_764_port, 
      DataPath_RF_bus_reg_dataout_765_port, 
      DataPath_RF_bus_reg_dataout_766_port, 
      DataPath_RF_bus_reg_dataout_767_port, 
      DataPath_RF_bus_reg_dataout_768_port, 
      DataPath_RF_bus_reg_dataout_769_port, 
      DataPath_RF_bus_reg_dataout_770_port, 
      DataPath_RF_bus_reg_dataout_771_port, 
      DataPath_RF_bus_reg_dataout_772_port, 
      DataPath_RF_bus_reg_dataout_773_port, 
      DataPath_RF_bus_reg_dataout_774_port, 
      DataPath_RF_bus_reg_dataout_775_port, 
      DataPath_RF_bus_reg_dataout_776_port, 
      DataPath_RF_bus_reg_dataout_777_port, 
      DataPath_RF_bus_reg_dataout_778_port, 
      DataPath_RF_bus_reg_dataout_779_port, 
      DataPath_RF_bus_reg_dataout_780_port, 
      DataPath_RF_bus_reg_dataout_781_port, 
      DataPath_RF_bus_reg_dataout_782_port, 
      DataPath_RF_bus_reg_dataout_783_port, 
      DataPath_RF_bus_reg_dataout_784_port, 
      DataPath_RF_bus_reg_dataout_785_port, 
      DataPath_RF_bus_reg_dataout_786_port, 
      DataPath_RF_bus_reg_dataout_787_port, 
      DataPath_RF_bus_reg_dataout_788_port, 
      DataPath_RF_bus_reg_dataout_789_port, 
      DataPath_RF_bus_reg_dataout_790_port, 
      DataPath_RF_bus_reg_dataout_791_port, 
      DataPath_RF_bus_reg_dataout_792_port, 
      DataPath_RF_bus_reg_dataout_793_port, 
      DataPath_RF_bus_reg_dataout_794_port, 
      DataPath_RF_bus_reg_dataout_795_port, 
      DataPath_RF_bus_reg_dataout_796_port, 
      DataPath_RF_bus_reg_dataout_797_port, 
      DataPath_RF_bus_reg_dataout_798_port, 
      DataPath_RF_bus_reg_dataout_799_port, 
      DataPath_RF_bus_reg_dataout_800_port, 
      DataPath_RF_bus_reg_dataout_801_port, 
      DataPath_RF_bus_reg_dataout_802_port, 
      DataPath_RF_bus_reg_dataout_803_port, 
      DataPath_RF_bus_reg_dataout_804_port, 
      DataPath_RF_bus_reg_dataout_805_port, 
      DataPath_RF_bus_reg_dataout_806_port, 
      DataPath_RF_bus_reg_dataout_807_port, 
      DataPath_RF_bus_reg_dataout_808_port, 
      DataPath_RF_bus_reg_dataout_809_port, 
      DataPath_RF_bus_reg_dataout_810_port, 
      DataPath_RF_bus_reg_dataout_811_port, 
      DataPath_RF_bus_reg_dataout_812_port, 
      DataPath_RF_bus_reg_dataout_813_port, 
      DataPath_RF_bus_reg_dataout_814_port, 
      DataPath_RF_bus_reg_dataout_815_port, 
      DataPath_RF_bus_reg_dataout_816_port, 
      DataPath_RF_bus_reg_dataout_817_port, 
      DataPath_RF_bus_reg_dataout_818_port, 
      DataPath_RF_bus_reg_dataout_819_port, 
      DataPath_RF_bus_reg_dataout_820_port, 
      DataPath_RF_bus_reg_dataout_821_port, 
      DataPath_RF_bus_reg_dataout_822_port, 
      DataPath_RF_bus_reg_dataout_823_port, 
      DataPath_RF_bus_reg_dataout_824_port, 
      DataPath_RF_bus_reg_dataout_825_port, 
      DataPath_RF_bus_reg_dataout_826_port, 
      DataPath_RF_bus_reg_dataout_827_port, 
      DataPath_RF_bus_reg_dataout_828_port, 
      DataPath_RF_bus_reg_dataout_829_port, 
      DataPath_RF_bus_reg_dataout_830_port, 
      DataPath_RF_bus_reg_dataout_831_port, 
      DataPath_RF_bus_reg_dataout_832_port, 
      DataPath_RF_bus_reg_dataout_833_port, 
      DataPath_RF_bus_reg_dataout_834_port, 
      DataPath_RF_bus_reg_dataout_835_port, 
      DataPath_RF_bus_reg_dataout_836_port, 
      DataPath_RF_bus_reg_dataout_837_port, 
      DataPath_RF_bus_reg_dataout_838_port, 
      DataPath_RF_bus_reg_dataout_839_port, 
      DataPath_RF_bus_reg_dataout_840_port, 
      DataPath_RF_bus_reg_dataout_841_port, 
      DataPath_RF_bus_reg_dataout_842_port, 
      DataPath_RF_bus_reg_dataout_843_port, 
      DataPath_RF_bus_reg_dataout_844_port, 
      DataPath_RF_bus_reg_dataout_845_port, 
      DataPath_RF_bus_reg_dataout_846_port, 
      DataPath_RF_bus_reg_dataout_847_port, 
      DataPath_RF_bus_reg_dataout_848_port, 
      DataPath_RF_bus_reg_dataout_849_port, 
      DataPath_RF_bus_reg_dataout_850_port, 
      DataPath_RF_bus_reg_dataout_851_port, 
      DataPath_RF_bus_reg_dataout_852_port, 
      DataPath_RF_bus_reg_dataout_853_port, 
      DataPath_RF_bus_reg_dataout_854_port, 
      DataPath_RF_bus_reg_dataout_855_port, 
      DataPath_RF_bus_reg_dataout_856_port, 
      DataPath_RF_bus_reg_dataout_857_port, 
      DataPath_RF_bus_reg_dataout_858_port, 
      DataPath_RF_bus_reg_dataout_859_port, 
      DataPath_RF_bus_reg_dataout_860_port, 
      DataPath_RF_bus_reg_dataout_861_port, 
      DataPath_RF_bus_reg_dataout_862_port, 
      DataPath_RF_bus_reg_dataout_863_port, 
      DataPath_RF_bus_reg_dataout_864_port, 
      DataPath_RF_bus_reg_dataout_865_port, 
      DataPath_RF_bus_reg_dataout_866_port, 
      DataPath_RF_bus_reg_dataout_867_port, 
      DataPath_RF_bus_reg_dataout_868_port, 
      DataPath_RF_bus_reg_dataout_869_port, 
      DataPath_RF_bus_reg_dataout_870_port, 
      DataPath_RF_bus_reg_dataout_871_port, 
      DataPath_RF_bus_reg_dataout_872_port, 
      DataPath_RF_bus_reg_dataout_873_port, 
      DataPath_RF_bus_reg_dataout_874_port, 
      DataPath_RF_bus_reg_dataout_875_port, 
      DataPath_RF_bus_reg_dataout_876_port, 
      DataPath_RF_bus_reg_dataout_877_port, 
      DataPath_RF_bus_reg_dataout_878_port, 
      DataPath_RF_bus_reg_dataout_879_port, 
      DataPath_RF_bus_reg_dataout_880_port, 
      DataPath_RF_bus_reg_dataout_881_port, 
      DataPath_RF_bus_reg_dataout_882_port, 
      DataPath_RF_bus_reg_dataout_883_port, 
      DataPath_RF_bus_reg_dataout_884_port, 
      DataPath_RF_bus_reg_dataout_885_port, 
      DataPath_RF_bus_reg_dataout_886_port, 
      DataPath_RF_bus_reg_dataout_887_port, 
      DataPath_RF_bus_reg_dataout_888_port, 
      DataPath_RF_bus_reg_dataout_889_port, 
      DataPath_RF_bus_reg_dataout_890_port, 
      DataPath_RF_bus_reg_dataout_891_port, 
      DataPath_RF_bus_reg_dataout_892_port, 
      DataPath_RF_bus_reg_dataout_893_port, 
      DataPath_RF_bus_reg_dataout_894_port, 
      DataPath_RF_bus_reg_dataout_895_port, 
      DataPath_RF_bus_reg_dataout_896_port, 
      DataPath_RF_bus_reg_dataout_897_port, 
      DataPath_RF_bus_reg_dataout_898_port, 
      DataPath_RF_bus_reg_dataout_899_port, 
      DataPath_RF_bus_reg_dataout_900_port, 
      DataPath_RF_bus_reg_dataout_901_port, 
      DataPath_RF_bus_reg_dataout_902_port, 
      DataPath_RF_bus_reg_dataout_903_port, 
      DataPath_RF_bus_reg_dataout_904_port, 
      DataPath_RF_bus_reg_dataout_905_port, 
      DataPath_RF_bus_reg_dataout_906_port, 
      DataPath_RF_bus_reg_dataout_907_port, 
      DataPath_RF_bus_reg_dataout_908_port, 
      DataPath_RF_bus_reg_dataout_909_port, 
      DataPath_RF_bus_reg_dataout_910_port, 
      DataPath_RF_bus_reg_dataout_911_port, 
      DataPath_RF_bus_reg_dataout_912_port, 
      DataPath_RF_bus_reg_dataout_913_port, 
      DataPath_RF_bus_reg_dataout_914_port, 
      DataPath_RF_bus_reg_dataout_915_port, 
      DataPath_RF_bus_reg_dataout_916_port, 
      DataPath_RF_bus_reg_dataout_917_port, 
      DataPath_RF_bus_reg_dataout_918_port, 
      DataPath_RF_bus_reg_dataout_919_port, 
      DataPath_RF_bus_reg_dataout_920_port, 
      DataPath_RF_bus_reg_dataout_921_port, 
      DataPath_RF_bus_reg_dataout_922_port, 
      DataPath_RF_bus_reg_dataout_923_port, 
      DataPath_RF_bus_reg_dataout_924_port, 
      DataPath_RF_bus_reg_dataout_925_port, 
      DataPath_RF_bus_reg_dataout_926_port, 
      DataPath_RF_bus_reg_dataout_927_port, 
      DataPath_RF_bus_reg_dataout_928_port, 
      DataPath_RF_bus_reg_dataout_929_port, 
      DataPath_RF_bus_reg_dataout_930_port, 
      DataPath_RF_bus_reg_dataout_931_port, 
      DataPath_RF_bus_reg_dataout_932_port, 
      DataPath_RF_bus_reg_dataout_933_port, 
      DataPath_RF_bus_reg_dataout_934_port, 
      DataPath_RF_bus_reg_dataout_935_port, 
      DataPath_RF_bus_reg_dataout_936_port, 
      DataPath_RF_bus_reg_dataout_937_port, 
      DataPath_RF_bus_reg_dataout_938_port, 
      DataPath_RF_bus_reg_dataout_939_port, 
      DataPath_RF_bus_reg_dataout_940_port, 
      DataPath_RF_bus_reg_dataout_941_port, 
      DataPath_RF_bus_reg_dataout_942_port, 
      DataPath_RF_bus_reg_dataout_943_port, 
      DataPath_RF_bus_reg_dataout_944_port, 
      DataPath_RF_bus_reg_dataout_945_port, 
      DataPath_RF_bus_reg_dataout_946_port, 
      DataPath_RF_bus_reg_dataout_947_port, 
      DataPath_RF_bus_reg_dataout_948_port, 
      DataPath_RF_bus_reg_dataout_949_port, 
      DataPath_RF_bus_reg_dataout_950_port, 
      DataPath_RF_bus_reg_dataout_951_port, 
      DataPath_RF_bus_reg_dataout_952_port, 
      DataPath_RF_bus_reg_dataout_953_port, 
      DataPath_RF_bus_reg_dataout_954_port, 
      DataPath_RF_bus_reg_dataout_955_port, 
      DataPath_RF_bus_reg_dataout_956_port, 
      DataPath_RF_bus_reg_dataout_957_port, 
      DataPath_RF_bus_reg_dataout_958_port, 
      DataPath_RF_bus_reg_dataout_959_port, 
      DataPath_RF_bus_reg_dataout_960_port, 
      DataPath_RF_bus_reg_dataout_961_port, 
      DataPath_RF_bus_reg_dataout_962_port, 
      DataPath_RF_bus_reg_dataout_963_port, 
      DataPath_RF_bus_reg_dataout_964_port, 
      DataPath_RF_bus_reg_dataout_965_port, 
      DataPath_RF_bus_reg_dataout_966_port, 
      DataPath_RF_bus_reg_dataout_967_port, 
      DataPath_RF_bus_reg_dataout_968_port, 
      DataPath_RF_bus_reg_dataout_969_port, 
      DataPath_RF_bus_reg_dataout_970_port, 
      DataPath_RF_bus_reg_dataout_971_port, 
      DataPath_RF_bus_reg_dataout_972_port, 
      DataPath_RF_bus_reg_dataout_973_port, 
      DataPath_RF_bus_reg_dataout_974_port, 
      DataPath_RF_bus_reg_dataout_975_port, 
      DataPath_RF_bus_reg_dataout_976_port, 
      DataPath_RF_bus_reg_dataout_977_port, 
      DataPath_RF_bus_reg_dataout_978_port, 
      DataPath_RF_bus_reg_dataout_979_port, 
      DataPath_RF_bus_reg_dataout_980_port, 
      DataPath_RF_bus_reg_dataout_981_port, 
      DataPath_RF_bus_reg_dataout_982_port, 
      DataPath_RF_bus_reg_dataout_983_port, 
      DataPath_RF_bus_reg_dataout_984_port, 
      DataPath_RF_bus_reg_dataout_985_port, 
      DataPath_RF_bus_reg_dataout_986_port, 
      DataPath_RF_bus_reg_dataout_987_port, 
      DataPath_RF_bus_reg_dataout_988_port, 
      DataPath_RF_bus_reg_dataout_989_port, 
      DataPath_RF_bus_reg_dataout_990_port, 
      DataPath_RF_bus_reg_dataout_991_port, 
      DataPath_RF_bus_reg_dataout_992_port, 
      DataPath_RF_bus_reg_dataout_993_port, 
      DataPath_RF_bus_reg_dataout_994_port, 
      DataPath_RF_bus_reg_dataout_995_port, 
      DataPath_RF_bus_reg_dataout_996_port, 
      DataPath_RF_bus_reg_dataout_997_port, 
      DataPath_RF_bus_reg_dataout_998_port, 
      DataPath_RF_bus_reg_dataout_999_port, 
      DataPath_RF_bus_reg_dataout_1000_port, 
      DataPath_RF_bus_reg_dataout_1001_port, 
      DataPath_RF_bus_reg_dataout_1002_port, 
      DataPath_RF_bus_reg_dataout_1003_port, 
      DataPath_RF_bus_reg_dataout_1004_port, 
      DataPath_RF_bus_reg_dataout_1005_port, 
      DataPath_RF_bus_reg_dataout_1006_port, 
      DataPath_RF_bus_reg_dataout_1007_port, 
      DataPath_RF_bus_reg_dataout_1008_port, 
      DataPath_RF_bus_reg_dataout_1009_port, 
      DataPath_RF_bus_reg_dataout_1010_port, 
      DataPath_RF_bus_reg_dataout_1011_port, 
      DataPath_RF_bus_reg_dataout_1012_port, 
      DataPath_RF_bus_reg_dataout_1013_port, 
      DataPath_RF_bus_reg_dataout_1014_port, 
      DataPath_RF_bus_reg_dataout_1015_port, 
      DataPath_RF_bus_reg_dataout_1016_port, 
      DataPath_RF_bus_reg_dataout_1017_port, 
      DataPath_RF_bus_reg_dataout_1018_port, 
      DataPath_RF_bus_reg_dataout_1019_port, 
      DataPath_RF_bus_reg_dataout_1020_port, 
      DataPath_RF_bus_reg_dataout_1021_port, 
      DataPath_RF_bus_reg_dataout_1022_port, 
      DataPath_RF_bus_reg_dataout_1023_port, 
      DataPath_RF_bus_reg_dataout_1024_port, 
      DataPath_RF_bus_reg_dataout_1025_port, 
      DataPath_RF_bus_reg_dataout_1026_port, 
      DataPath_RF_bus_reg_dataout_1027_port, 
      DataPath_RF_bus_reg_dataout_1028_port, 
      DataPath_RF_bus_reg_dataout_1029_port, 
      DataPath_RF_bus_reg_dataout_1030_port, 
      DataPath_RF_bus_reg_dataout_1031_port, 
      DataPath_RF_bus_reg_dataout_1032_port, 
      DataPath_RF_bus_reg_dataout_1033_port, 
      DataPath_RF_bus_reg_dataout_1034_port, 
      DataPath_RF_bus_reg_dataout_1035_port, 
      DataPath_RF_bus_reg_dataout_1036_port, 
      DataPath_RF_bus_reg_dataout_1037_port, 
      DataPath_RF_bus_reg_dataout_1038_port, 
      DataPath_RF_bus_reg_dataout_1039_port, 
      DataPath_RF_bus_reg_dataout_1040_port, 
      DataPath_RF_bus_reg_dataout_1041_port, 
      DataPath_RF_bus_reg_dataout_1042_port, 
      DataPath_RF_bus_reg_dataout_1043_port, 
      DataPath_RF_bus_reg_dataout_1044_port, 
      DataPath_RF_bus_reg_dataout_1045_port, 
      DataPath_RF_bus_reg_dataout_1046_port, 
      DataPath_RF_bus_reg_dataout_1047_port, 
      DataPath_RF_bus_reg_dataout_1048_port, 
      DataPath_RF_bus_reg_dataout_1049_port, 
      DataPath_RF_bus_reg_dataout_1050_port, 
      DataPath_RF_bus_reg_dataout_1051_port, 
      DataPath_RF_bus_reg_dataout_1052_port, 
      DataPath_RF_bus_reg_dataout_1053_port, 
      DataPath_RF_bus_reg_dataout_1054_port, 
      DataPath_RF_bus_reg_dataout_1055_port, 
      DataPath_RF_bus_reg_dataout_1056_port, 
      DataPath_RF_bus_reg_dataout_1057_port, 
      DataPath_RF_bus_reg_dataout_1058_port, 
      DataPath_RF_bus_reg_dataout_1059_port, 
      DataPath_RF_bus_reg_dataout_1060_port, 
      DataPath_RF_bus_reg_dataout_1061_port, 
      DataPath_RF_bus_reg_dataout_1062_port, 
      DataPath_RF_bus_reg_dataout_1063_port, 
      DataPath_RF_bus_reg_dataout_1064_port, 
      DataPath_RF_bus_reg_dataout_1065_port, 
      DataPath_RF_bus_reg_dataout_1066_port, 
      DataPath_RF_bus_reg_dataout_1067_port, 
      DataPath_RF_bus_reg_dataout_1068_port, 
      DataPath_RF_bus_reg_dataout_1069_port, 
      DataPath_RF_bus_reg_dataout_1070_port, 
      DataPath_RF_bus_reg_dataout_1071_port, 
      DataPath_RF_bus_reg_dataout_1072_port, 
      DataPath_RF_bus_reg_dataout_1073_port, 
      DataPath_RF_bus_reg_dataout_1074_port, 
      DataPath_RF_bus_reg_dataout_1075_port, 
      DataPath_RF_bus_reg_dataout_1076_port, 
      DataPath_RF_bus_reg_dataout_1077_port, 
      DataPath_RF_bus_reg_dataout_1078_port, 
      DataPath_RF_bus_reg_dataout_1079_port, 
      DataPath_RF_bus_reg_dataout_1080_port, 
      DataPath_RF_bus_reg_dataout_1081_port, 
      DataPath_RF_bus_reg_dataout_1082_port, 
      DataPath_RF_bus_reg_dataout_1083_port, 
      DataPath_RF_bus_reg_dataout_1084_port, 
      DataPath_RF_bus_reg_dataout_1085_port, 
      DataPath_RF_bus_reg_dataout_1086_port, 
      DataPath_RF_bus_reg_dataout_1087_port, 
      DataPath_RF_bus_reg_dataout_1088_port, 
      DataPath_RF_bus_reg_dataout_1089_port, 
      DataPath_RF_bus_reg_dataout_1090_port, 
      DataPath_RF_bus_reg_dataout_1091_port, 
      DataPath_RF_bus_reg_dataout_1092_port, 
      DataPath_RF_bus_reg_dataout_1093_port, 
      DataPath_RF_bus_reg_dataout_1094_port, 
      DataPath_RF_bus_reg_dataout_1095_port, 
      DataPath_RF_bus_reg_dataout_1096_port, 
      DataPath_RF_bus_reg_dataout_1097_port, 
      DataPath_RF_bus_reg_dataout_1098_port, 
      DataPath_RF_bus_reg_dataout_1099_port, 
      DataPath_RF_bus_reg_dataout_1100_port, 
      DataPath_RF_bus_reg_dataout_1101_port, 
      DataPath_RF_bus_reg_dataout_1102_port, 
      DataPath_RF_bus_reg_dataout_1103_port, 
      DataPath_RF_bus_reg_dataout_1104_port, 
      DataPath_RF_bus_reg_dataout_1105_port, 
      DataPath_RF_bus_reg_dataout_1106_port, 
      DataPath_RF_bus_reg_dataout_1107_port, 
      DataPath_RF_bus_reg_dataout_1108_port, 
      DataPath_RF_bus_reg_dataout_1109_port, 
      DataPath_RF_bus_reg_dataout_1110_port, 
      DataPath_RF_bus_reg_dataout_1111_port, 
      DataPath_RF_bus_reg_dataout_1112_port, 
      DataPath_RF_bus_reg_dataout_1113_port, 
      DataPath_RF_bus_reg_dataout_1114_port, 
      DataPath_RF_bus_reg_dataout_1115_port, 
      DataPath_RF_bus_reg_dataout_1116_port, 
      DataPath_RF_bus_reg_dataout_1117_port, 
      DataPath_RF_bus_reg_dataout_1118_port, 
      DataPath_RF_bus_reg_dataout_1119_port, 
      DataPath_RF_bus_reg_dataout_1120_port, 
      DataPath_RF_bus_reg_dataout_1121_port, 
      DataPath_RF_bus_reg_dataout_1122_port, 
      DataPath_RF_bus_reg_dataout_1123_port, 
      DataPath_RF_bus_reg_dataout_1124_port, 
      DataPath_RF_bus_reg_dataout_1125_port, 
      DataPath_RF_bus_reg_dataout_1126_port, 
      DataPath_RF_bus_reg_dataout_1127_port, 
      DataPath_RF_bus_reg_dataout_1128_port, 
      DataPath_RF_bus_reg_dataout_1129_port, 
      DataPath_RF_bus_reg_dataout_1130_port, 
      DataPath_RF_bus_reg_dataout_1131_port, 
      DataPath_RF_bus_reg_dataout_1132_port, 
      DataPath_RF_bus_reg_dataout_1133_port, 
      DataPath_RF_bus_reg_dataout_1134_port, 
      DataPath_RF_bus_reg_dataout_1135_port, 
      DataPath_RF_bus_reg_dataout_1136_port, 
      DataPath_RF_bus_reg_dataout_1137_port, 
      DataPath_RF_bus_reg_dataout_1138_port, 
      DataPath_RF_bus_reg_dataout_1139_port, 
      DataPath_RF_bus_reg_dataout_1140_port, 
      DataPath_RF_bus_reg_dataout_1141_port, 
      DataPath_RF_bus_reg_dataout_1142_port, 
      DataPath_RF_bus_reg_dataout_1143_port, 
      DataPath_RF_bus_reg_dataout_1144_port, 
      DataPath_RF_bus_reg_dataout_1145_port, 
      DataPath_RF_bus_reg_dataout_1146_port, 
      DataPath_RF_bus_reg_dataout_1147_port, 
      DataPath_RF_bus_reg_dataout_1148_port, 
      DataPath_RF_bus_reg_dataout_1149_port, 
      DataPath_RF_bus_reg_dataout_1150_port, 
      DataPath_RF_bus_reg_dataout_1151_port, 
      DataPath_RF_bus_reg_dataout_1152_port, 
      DataPath_RF_bus_reg_dataout_1153_port, 
      DataPath_RF_bus_reg_dataout_1154_port, 
      DataPath_RF_bus_reg_dataout_1155_port, 
      DataPath_RF_bus_reg_dataout_1156_port, 
      DataPath_RF_bus_reg_dataout_1157_port, 
      DataPath_RF_bus_reg_dataout_1158_port, 
      DataPath_RF_bus_reg_dataout_1159_port, 
      DataPath_RF_bus_reg_dataout_1160_port, 
      DataPath_RF_bus_reg_dataout_1161_port, 
      DataPath_RF_bus_reg_dataout_1162_port, 
      DataPath_RF_bus_reg_dataout_1163_port, 
      DataPath_RF_bus_reg_dataout_1164_port, 
      DataPath_RF_bus_reg_dataout_1165_port, 
      DataPath_RF_bus_reg_dataout_1166_port, 
      DataPath_RF_bus_reg_dataout_1167_port, 
      DataPath_RF_bus_reg_dataout_1168_port, 
      DataPath_RF_bus_reg_dataout_1169_port, 
      DataPath_RF_bus_reg_dataout_1170_port, 
      DataPath_RF_bus_reg_dataout_1171_port, 
      DataPath_RF_bus_reg_dataout_1172_port, 
      DataPath_RF_bus_reg_dataout_1173_port, 
      DataPath_RF_bus_reg_dataout_1174_port, 
      DataPath_RF_bus_reg_dataout_1175_port, 
      DataPath_RF_bus_reg_dataout_1176_port, 
      DataPath_RF_bus_reg_dataout_1177_port, 
      DataPath_RF_bus_reg_dataout_1178_port, 
      DataPath_RF_bus_reg_dataout_1179_port, 
      DataPath_RF_bus_reg_dataout_1180_port, 
      DataPath_RF_bus_reg_dataout_1181_port, 
      DataPath_RF_bus_reg_dataout_1182_port, 
      DataPath_RF_bus_reg_dataout_1183_port, 
      DataPath_RF_bus_reg_dataout_1184_port, 
      DataPath_RF_bus_reg_dataout_1185_port, 
      DataPath_RF_bus_reg_dataout_1186_port, 
      DataPath_RF_bus_reg_dataout_1187_port, 
      DataPath_RF_bus_reg_dataout_1188_port, 
      DataPath_RF_bus_reg_dataout_1189_port, 
      DataPath_RF_bus_reg_dataout_1190_port, 
      DataPath_RF_bus_reg_dataout_1191_port, 
      DataPath_RF_bus_reg_dataout_1192_port, 
      DataPath_RF_bus_reg_dataout_1193_port, 
      DataPath_RF_bus_reg_dataout_1194_port, 
      DataPath_RF_bus_reg_dataout_1195_port, 
      DataPath_RF_bus_reg_dataout_1196_port, 
      DataPath_RF_bus_reg_dataout_1197_port, 
      DataPath_RF_bus_reg_dataout_1198_port, 
      DataPath_RF_bus_reg_dataout_1199_port, 
      DataPath_RF_bus_reg_dataout_1200_port, 
      DataPath_RF_bus_reg_dataout_1201_port, 
      DataPath_RF_bus_reg_dataout_1202_port, 
      DataPath_RF_bus_reg_dataout_1203_port, 
      DataPath_RF_bus_reg_dataout_1204_port, 
      DataPath_RF_bus_reg_dataout_1205_port, 
      DataPath_RF_bus_reg_dataout_1206_port, 
      DataPath_RF_bus_reg_dataout_1207_port, 
      DataPath_RF_bus_reg_dataout_1208_port, 
      DataPath_RF_bus_reg_dataout_1209_port, 
      DataPath_RF_bus_reg_dataout_1210_port, 
      DataPath_RF_bus_reg_dataout_1211_port, 
      DataPath_RF_bus_reg_dataout_1212_port, 
      DataPath_RF_bus_reg_dataout_1213_port, 
      DataPath_RF_bus_reg_dataout_1214_port, 
      DataPath_RF_bus_reg_dataout_1215_port, 
      DataPath_RF_bus_reg_dataout_1216_port, 
      DataPath_RF_bus_reg_dataout_1217_port, 
      DataPath_RF_bus_reg_dataout_1218_port, 
      DataPath_RF_bus_reg_dataout_1219_port, 
      DataPath_RF_bus_reg_dataout_1220_port, 
      DataPath_RF_bus_reg_dataout_1221_port, 
      DataPath_RF_bus_reg_dataout_1222_port, 
      DataPath_RF_bus_reg_dataout_1223_port, 
      DataPath_RF_bus_reg_dataout_1224_port, 
      DataPath_RF_bus_reg_dataout_1225_port, 
      DataPath_RF_bus_reg_dataout_1226_port, 
      DataPath_RF_bus_reg_dataout_1227_port, 
      DataPath_RF_bus_reg_dataout_1228_port, 
      DataPath_RF_bus_reg_dataout_1229_port, 
      DataPath_RF_bus_reg_dataout_1230_port, 
      DataPath_RF_bus_reg_dataout_1231_port, 
      DataPath_RF_bus_reg_dataout_1232_port, 
      DataPath_RF_bus_reg_dataout_1233_port, 
      DataPath_RF_bus_reg_dataout_1234_port, 
      DataPath_RF_bus_reg_dataout_1235_port, 
      DataPath_RF_bus_reg_dataout_1236_port, 
      DataPath_RF_bus_reg_dataout_1237_port, 
      DataPath_RF_bus_reg_dataout_1238_port, 
      DataPath_RF_bus_reg_dataout_1239_port, 
      DataPath_RF_bus_reg_dataout_1240_port, 
      DataPath_RF_bus_reg_dataout_1241_port, 
      DataPath_RF_bus_reg_dataout_1242_port, 
      DataPath_RF_bus_reg_dataout_1243_port, 
      DataPath_RF_bus_reg_dataout_1244_port, 
      DataPath_RF_bus_reg_dataout_1245_port, 
      DataPath_RF_bus_reg_dataout_1246_port, 
      DataPath_RF_bus_reg_dataout_1247_port, 
      DataPath_RF_bus_reg_dataout_1248_port, 
      DataPath_RF_bus_reg_dataout_1249_port, 
      DataPath_RF_bus_reg_dataout_1250_port, 
      DataPath_RF_bus_reg_dataout_1251_port, 
      DataPath_RF_bus_reg_dataout_1252_port, 
      DataPath_RF_bus_reg_dataout_1253_port, 
      DataPath_RF_bus_reg_dataout_1254_port, 
      DataPath_RF_bus_reg_dataout_1255_port, 
      DataPath_RF_bus_reg_dataout_1256_port, 
      DataPath_RF_bus_reg_dataout_1257_port, 
      DataPath_RF_bus_reg_dataout_1258_port, 
      DataPath_RF_bus_reg_dataout_1259_port, 
      DataPath_RF_bus_reg_dataout_1260_port, 
      DataPath_RF_bus_reg_dataout_1261_port, 
      DataPath_RF_bus_reg_dataout_1262_port, 
      DataPath_RF_bus_reg_dataout_1263_port, 
      DataPath_RF_bus_reg_dataout_1264_port, 
      DataPath_RF_bus_reg_dataout_1265_port, 
      DataPath_RF_bus_reg_dataout_1266_port, 
      DataPath_RF_bus_reg_dataout_1267_port, 
      DataPath_RF_bus_reg_dataout_1268_port, 
      DataPath_RF_bus_reg_dataout_1269_port, 
      DataPath_RF_bus_reg_dataout_1270_port, 
      DataPath_RF_bus_reg_dataout_1271_port, 
      DataPath_RF_bus_reg_dataout_1272_port, 
      DataPath_RF_bus_reg_dataout_1273_port, 
      DataPath_RF_bus_reg_dataout_1274_port, 
      DataPath_RF_bus_reg_dataout_1275_port, 
      DataPath_RF_bus_reg_dataout_1276_port, 
      DataPath_RF_bus_reg_dataout_1277_port, 
      DataPath_RF_bus_reg_dataout_1278_port, 
      DataPath_RF_bus_reg_dataout_1279_port, 
      DataPath_RF_bus_reg_dataout_1280_port, 
      DataPath_RF_bus_reg_dataout_1281_port, 
      DataPath_RF_bus_reg_dataout_1282_port, 
      DataPath_RF_bus_reg_dataout_1283_port, 
      DataPath_RF_bus_reg_dataout_1284_port, 
      DataPath_RF_bus_reg_dataout_1285_port, 
      DataPath_RF_bus_reg_dataout_1286_port, 
      DataPath_RF_bus_reg_dataout_1287_port, 
      DataPath_RF_bus_reg_dataout_1288_port, 
      DataPath_RF_bus_reg_dataout_1289_port, 
      DataPath_RF_bus_reg_dataout_1290_port, 
      DataPath_RF_bus_reg_dataout_1291_port, 
      DataPath_RF_bus_reg_dataout_1292_port, 
      DataPath_RF_bus_reg_dataout_1293_port, 
      DataPath_RF_bus_reg_dataout_1294_port, 
      DataPath_RF_bus_reg_dataout_1295_port, 
      DataPath_RF_bus_reg_dataout_1296_port, 
      DataPath_RF_bus_reg_dataout_1297_port, 
      DataPath_RF_bus_reg_dataout_1298_port, 
      DataPath_RF_bus_reg_dataout_1299_port, 
      DataPath_RF_bus_reg_dataout_1300_port, 
      DataPath_RF_bus_reg_dataout_1301_port, 
      DataPath_RF_bus_reg_dataout_1302_port, 
      DataPath_RF_bus_reg_dataout_1303_port, 
      DataPath_RF_bus_reg_dataout_1304_port, 
      DataPath_RF_bus_reg_dataout_1305_port, 
      DataPath_RF_bus_reg_dataout_1306_port, 
      DataPath_RF_bus_reg_dataout_1307_port, 
      DataPath_RF_bus_reg_dataout_1308_port, 
      DataPath_RF_bus_reg_dataout_1309_port, 
      DataPath_RF_bus_reg_dataout_1310_port, 
      DataPath_RF_bus_reg_dataout_1311_port, 
      DataPath_RF_bus_reg_dataout_1312_port, 
      DataPath_RF_bus_reg_dataout_1313_port, 
      DataPath_RF_bus_reg_dataout_1314_port, 
      DataPath_RF_bus_reg_dataout_1315_port, 
      DataPath_RF_bus_reg_dataout_1316_port, 
      DataPath_RF_bus_reg_dataout_1317_port, 
      DataPath_RF_bus_reg_dataout_1318_port, 
      DataPath_RF_bus_reg_dataout_1319_port, 
      DataPath_RF_bus_reg_dataout_1320_port, 
      DataPath_RF_bus_reg_dataout_1321_port, 
      DataPath_RF_bus_reg_dataout_1322_port, 
      DataPath_RF_bus_reg_dataout_1323_port, 
      DataPath_RF_bus_reg_dataout_1324_port, 
      DataPath_RF_bus_reg_dataout_1325_port, 
      DataPath_RF_bus_reg_dataout_1326_port, 
      DataPath_RF_bus_reg_dataout_1327_port, 
      DataPath_RF_bus_reg_dataout_1328_port, 
      DataPath_RF_bus_reg_dataout_1329_port, 
      DataPath_RF_bus_reg_dataout_1330_port, 
      DataPath_RF_bus_reg_dataout_1331_port, 
      DataPath_RF_bus_reg_dataout_1332_port, 
      DataPath_RF_bus_reg_dataout_1333_port, 
      DataPath_RF_bus_reg_dataout_1334_port, 
      DataPath_RF_bus_reg_dataout_1335_port, 
      DataPath_RF_bus_reg_dataout_1336_port, 
      DataPath_RF_bus_reg_dataout_1337_port, 
      DataPath_RF_bus_reg_dataout_1338_port, 
      DataPath_RF_bus_reg_dataout_1339_port, 
      DataPath_RF_bus_reg_dataout_1340_port, 
      DataPath_RF_bus_reg_dataout_1341_port, 
      DataPath_RF_bus_reg_dataout_1342_port, 
      DataPath_RF_bus_reg_dataout_1343_port, 
      DataPath_RF_bus_reg_dataout_1344_port, 
      DataPath_RF_bus_reg_dataout_1345_port, 
      DataPath_RF_bus_reg_dataout_1346_port, 
      DataPath_RF_bus_reg_dataout_1347_port, 
      DataPath_RF_bus_reg_dataout_1348_port, 
      DataPath_RF_bus_reg_dataout_1349_port, 
      DataPath_RF_bus_reg_dataout_1350_port, 
      DataPath_RF_bus_reg_dataout_1351_port, 
      DataPath_RF_bus_reg_dataout_1352_port, 
      DataPath_RF_bus_reg_dataout_1353_port, 
      DataPath_RF_bus_reg_dataout_1354_port, 
      DataPath_RF_bus_reg_dataout_1355_port, 
      DataPath_RF_bus_reg_dataout_1356_port, 
      DataPath_RF_bus_reg_dataout_1357_port, 
      DataPath_RF_bus_reg_dataout_1358_port, 
      DataPath_RF_bus_reg_dataout_1359_port, 
      DataPath_RF_bus_reg_dataout_1360_port, 
      DataPath_RF_bus_reg_dataout_1361_port, 
      DataPath_RF_bus_reg_dataout_1362_port, 
      DataPath_RF_bus_reg_dataout_1363_port, 
      DataPath_RF_bus_reg_dataout_1364_port, 
      DataPath_RF_bus_reg_dataout_1365_port, 
      DataPath_RF_bus_reg_dataout_1366_port, 
      DataPath_RF_bus_reg_dataout_1367_port, 
      DataPath_RF_bus_reg_dataout_1368_port, 
      DataPath_RF_bus_reg_dataout_1369_port, 
      DataPath_RF_bus_reg_dataout_1370_port, 
      DataPath_RF_bus_reg_dataout_1371_port, 
      DataPath_RF_bus_reg_dataout_1372_port, 
      DataPath_RF_bus_reg_dataout_1373_port, 
      DataPath_RF_bus_reg_dataout_1374_port, 
      DataPath_RF_bus_reg_dataout_1375_port, 
      DataPath_RF_bus_reg_dataout_1376_port, 
      DataPath_RF_bus_reg_dataout_1377_port, 
      DataPath_RF_bus_reg_dataout_1378_port, 
      DataPath_RF_bus_reg_dataout_1379_port, 
      DataPath_RF_bus_reg_dataout_1380_port, 
      DataPath_RF_bus_reg_dataout_1381_port, 
      DataPath_RF_bus_reg_dataout_1382_port, 
      DataPath_RF_bus_reg_dataout_1383_port, 
      DataPath_RF_bus_reg_dataout_1384_port, 
      DataPath_RF_bus_reg_dataout_1385_port, 
      DataPath_RF_bus_reg_dataout_1386_port, 
      DataPath_RF_bus_reg_dataout_1387_port, 
      DataPath_RF_bus_reg_dataout_1388_port, 
      DataPath_RF_bus_reg_dataout_1389_port, 
      DataPath_RF_bus_reg_dataout_1390_port, 
      DataPath_RF_bus_reg_dataout_1391_port, 
      DataPath_RF_bus_reg_dataout_1392_port, 
      DataPath_RF_bus_reg_dataout_1393_port, 
      DataPath_RF_bus_reg_dataout_1394_port, 
      DataPath_RF_bus_reg_dataout_1395_port, 
      DataPath_RF_bus_reg_dataout_1396_port, 
      DataPath_RF_bus_reg_dataout_1397_port, 
      DataPath_RF_bus_reg_dataout_1398_port, 
      DataPath_RF_bus_reg_dataout_1399_port, 
      DataPath_RF_bus_reg_dataout_1400_port, 
      DataPath_RF_bus_reg_dataout_1401_port, 
      DataPath_RF_bus_reg_dataout_1402_port, 
      DataPath_RF_bus_reg_dataout_1403_port, 
      DataPath_RF_bus_reg_dataout_1404_port, 
      DataPath_RF_bus_reg_dataout_1405_port, 
      DataPath_RF_bus_reg_dataout_1406_port, 
      DataPath_RF_bus_reg_dataout_1407_port, 
      DataPath_RF_bus_reg_dataout_1408_port, 
      DataPath_RF_bus_reg_dataout_1409_port, 
      DataPath_RF_bus_reg_dataout_1410_port, 
      DataPath_RF_bus_reg_dataout_1411_port, 
      DataPath_RF_bus_reg_dataout_1412_port, 
      DataPath_RF_bus_reg_dataout_1413_port, 
      DataPath_RF_bus_reg_dataout_1414_port, 
      DataPath_RF_bus_reg_dataout_1415_port, 
      DataPath_RF_bus_reg_dataout_1416_port, 
      DataPath_RF_bus_reg_dataout_1417_port, 
      DataPath_RF_bus_reg_dataout_1418_port, 
      DataPath_RF_bus_reg_dataout_1419_port, 
      DataPath_RF_bus_reg_dataout_1420_port, 
      DataPath_RF_bus_reg_dataout_1421_port, 
      DataPath_RF_bus_reg_dataout_1422_port, 
      DataPath_RF_bus_reg_dataout_1423_port, 
      DataPath_RF_bus_reg_dataout_1424_port, 
      DataPath_RF_bus_reg_dataout_1425_port, 
      DataPath_RF_bus_reg_dataout_1426_port, 
      DataPath_RF_bus_reg_dataout_1427_port, 
      DataPath_RF_bus_reg_dataout_1428_port, 
      DataPath_RF_bus_reg_dataout_1429_port, 
      DataPath_RF_bus_reg_dataout_1430_port, 
      DataPath_RF_bus_reg_dataout_1431_port, 
      DataPath_RF_bus_reg_dataout_1432_port, 
      DataPath_RF_bus_reg_dataout_1433_port, 
      DataPath_RF_bus_reg_dataout_1434_port, 
      DataPath_RF_bus_reg_dataout_1435_port, 
      DataPath_RF_bus_reg_dataout_1436_port, 
      DataPath_RF_bus_reg_dataout_1437_port, 
      DataPath_RF_bus_reg_dataout_1438_port, 
      DataPath_RF_bus_reg_dataout_1439_port, 
      DataPath_RF_bus_reg_dataout_1440_port, 
      DataPath_RF_bus_reg_dataout_1441_port, 
      DataPath_RF_bus_reg_dataout_1442_port, 
      DataPath_RF_bus_reg_dataout_1443_port, 
      DataPath_RF_bus_reg_dataout_1444_port, 
      DataPath_RF_bus_reg_dataout_1445_port, 
      DataPath_RF_bus_reg_dataout_1446_port, 
      DataPath_RF_bus_reg_dataout_1447_port, 
      DataPath_RF_bus_reg_dataout_1448_port, 
      DataPath_RF_bus_reg_dataout_1449_port, 
      DataPath_RF_bus_reg_dataout_1450_port, 
      DataPath_RF_bus_reg_dataout_1451_port, 
      DataPath_RF_bus_reg_dataout_1452_port, 
      DataPath_RF_bus_reg_dataout_1453_port, 
      DataPath_RF_bus_reg_dataout_1454_port, 
      DataPath_RF_bus_reg_dataout_1455_port, 
      DataPath_RF_bus_reg_dataout_1456_port, 
      DataPath_RF_bus_reg_dataout_1457_port, 
      DataPath_RF_bus_reg_dataout_1458_port, 
      DataPath_RF_bus_reg_dataout_1459_port, 
      DataPath_RF_bus_reg_dataout_1460_port, 
      DataPath_RF_bus_reg_dataout_1461_port, 
      DataPath_RF_bus_reg_dataout_1462_port, 
      DataPath_RF_bus_reg_dataout_1463_port, 
      DataPath_RF_bus_reg_dataout_1464_port, 
      DataPath_RF_bus_reg_dataout_1465_port, 
      DataPath_RF_bus_reg_dataout_1466_port, 
      DataPath_RF_bus_reg_dataout_1467_port, 
      DataPath_RF_bus_reg_dataout_1468_port, 
      DataPath_RF_bus_reg_dataout_1469_port, 
      DataPath_RF_bus_reg_dataout_1470_port, 
      DataPath_RF_bus_reg_dataout_1471_port, 
      DataPath_RF_bus_reg_dataout_1472_port, 
      DataPath_RF_bus_reg_dataout_1473_port, 
      DataPath_RF_bus_reg_dataout_1474_port, 
      DataPath_RF_bus_reg_dataout_1475_port, 
      DataPath_RF_bus_reg_dataout_1476_port, 
      DataPath_RF_bus_reg_dataout_1477_port, 
      DataPath_RF_bus_reg_dataout_1478_port, 
      DataPath_RF_bus_reg_dataout_1479_port, 
      DataPath_RF_bus_reg_dataout_1480_port, 
      DataPath_RF_bus_reg_dataout_1481_port, 
      DataPath_RF_bus_reg_dataout_1482_port, 
      DataPath_RF_bus_reg_dataout_1483_port, 
      DataPath_RF_bus_reg_dataout_1484_port, 
      DataPath_RF_bus_reg_dataout_1485_port, 
      DataPath_RF_bus_reg_dataout_1486_port, 
      DataPath_RF_bus_reg_dataout_1487_port, 
      DataPath_RF_bus_reg_dataout_1488_port, 
      DataPath_RF_bus_reg_dataout_1489_port, 
      DataPath_RF_bus_reg_dataout_1490_port, 
      DataPath_RF_bus_reg_dataout_1491_port, 
      DataPath_RF_bus_reg_dataout_1492_port, 
      DataPath_RF_bus_reg_dataout_1493_port, 
      DataPath_RF_bus_reg_dataout_1494_port, 
      DataPath_RF_bus_reg_dataout_1495_port, 
      DataPath_RF_bus_reg_dataout_1496_port, 
      DataPath_RF_bus_reg_dataout_1497_port, 
      DataPath_RF_bus_reg_dataout_1498_port, 
      DataPath_RF_bus_reg_dataout_1499_port, 
      DataPath_RF_bus_reg_dataout_1500_port, 
      DataPath_RF_bus_reg_dataout_1501_port, 
      DataPath_RF_bus_reg_dataout_1502_port, 
      DataPath_RF_bus_reg_dataout_1503_port, 
      DataPath_RF_bus_reg_dataout_1504_port, 
      DataPath_RF_bus_reg_dataout_1505_port, 
      DataPath_RF_bus_reg_dataout_1506_port, 
      DataPath_RF_bus_reg_dataout_1507_port, 
      DataPath_RF_bus_reg_dataout_1508_port, 
      DataPath_RF_bus_reg_dataout_1509_port, 
      DataPath_RF_bus_reg_dataout_1510_port, 
      DataPath_RF_bus_reg_dataout_1511_port, 
      DataPath_RF_bus_reg_dataout_1512_port, 
      DataPath_RF_bus_reg_dataout_1513_port, 
      DataPath_RF_bus_reg_dataout_1514_port, 
      DataPath_RF_bus_reg_dataout_1515_port, 
      DataPath_RF_bus_reg_dataout_1516_port, 
      DataPath_RF_bus_reg_dataout_1517_port, 
      DataPath_RF_bus_reg_dataout_1518_port, 
      DataPath_RF_bus_reg_dataout_1519_port, 
      DataPath_RF_bus_reg_dataout_1520_port, 
      DataPath_RF_bus_reg_dataout_1521_port, 
      DataPath_RF_bus_reg_dataout_1522_port, 
      DataPath_RF_bus_reg_dataout_1523_port, 
      DataPath_RF_bus_reg_dataout_1524_port, 
      DataPath_RF_bus_reg_dataout_1525_port, 
      DataPath_RF_bus_reg_dataout_1526_port, 
      DataPath_RF_bus_reg_dataout_1527_port, 
      DataPath_RF_bus_reg_dataout_1528_port, 
      DataPath_RF_bus_reg_dataout_1529_port, 
      DataPath_RF_bus_reg_dataout_1530_port, 
      DataPath_RF_bus_reg_dataout_1531_port, 
      DataPath_RF_bus_reg_dataout_1532_port, 
      DataPath_RF_bus_reg_dataout_1533_port, 
      DataPath_RF_bus_reg_dataout_1534_port, 
      DataPath_RF_bus_reg_dataout_1535_port, 
      DataPath_RF_bus_reg_dataout_1536_port, 
      DataPath_RF_bus_reg_dataout_1537_port, 
      DataPath_RF_bus_reg_dataout_1538_port, 
      DataPath_RF_bus_reg_dataout_1539_port, 
      DataPath_RF_bus_reg_dataout_1540_port, 
      DataPath_RF_bus_reg_dataout_1541_port, 
      DataPath_RF_bus_reg_dataout_1542_port, 
      DataPath_RF_bus_reg_dataout_1543_port, 
      DataPath_RF_bus_reg_dataout_1544_port, 
      DataPath_RF_bus_reg_dataout_1545_port, 
      DataPath_RF_bus_reg_dataout_1546_port, 
      DataPath_RF_bus_reg_dataout_1547_port, 
      DataPath_RF_bus_reg_dataout_1548_port, 
      DataPath_RF_bus_reg_dataout_1549_port, 
      DataPath_RF_bus_reg_dataout_1550_port, 
      DataPath_RF_bus_reg_dataout_1551_port, 
      DataPath_RF_bus_reg_dataout_1552_port, 
      DataPath_RF_bus_reg_dataout_1553_port, 
      DataPath_RF_bus_reg_dataout_1554_port, 
      DataPath_RF_bus_reg_dataout_1555_port, 
      DataPath_RF_bus_reg_dataout_1556_port, 
      DataPath_RF_bus_reg_dataout_1557_port, 
      DataPath_RF_bus_reg_dataout_1558_port, 
      DataPath_RF_bus_reg_dataout_1559_port, 
      DataPath_RF_bus_reg_dataout_1560_port, 
      DataPath_RF_bus_reg_dataout_1561_port, 
      DataPath_RF_bus_reg_dataout_1562_port, 
      DataPath_RF_bus_reg_dataout_1563_port, 
      DataPath_RF_bus_reg_dataout_1564_port, 
      DataPath_RF_bus_reg_dataout_1565_port, 
      DataPath_RF_bus_reg_dataout_1566_port, 
      DataPath_RF_bus_reg_dataout_1567_port, 
      DataPath_RF_bus_reg_dataout_1568_port, 
      DataPath_RF_bus_reg_dataout_1569_port, 
      DataPath_RF_bus_reg_dataout_1570_port, 
      DataPath_RF_bus_reg_dataout_1571_port, 
      DataPath_RF_bus_reg_dataout_1572_port, 
      DataPath_RF_bus_reg_dataout_1573_port, 
      DataPath_RF_bus_reg_dataout_1574_port, 
      DataPath_RF_bus_reg_dataout_1575_port, 
      DataPath_RF_bus_reg_dataout_1576_port, 
      DataPath_RF_bus_reg_dataout_1577_port, 
      DataPath_RF_bus_reg_dataout_1578_port, 
      DataPath_RF_bus_reg_dataout_1579_port, 
      DataPath_RF_bus_reg_dataout_1580_port, 
      DataPath_RF_bus_reg_dataout_1581_port, 
      DataPath_RF_bus_reg_dataout_1582_port, 
      DataPath_RF_bus_reg_dataout_1583_port, 
      DataPath_RF_bus_reg_dataout_1584_port, 
      DataPath_RF_bus_reg_dataout_1585_port, 
      DataPath_RF_bus_reg_dataout_1586_port, 
      DataPath_RF_bus_reg_dataout_1587_port, 
      DataPath_RF_bus_reg_dataout_1588_port, 
      DataPath_RF_bus_reg_dataout_1589_port, 
      DataPath_RF_bus_reg_dataout_1590_port, 
      DataPath_RF_bus_reg_dataout_1591_port, 
      DataPath_RF_bus_reg_dataout_1592_port, 
      DataPath_RF_bus_reg_dataout_1593_port, 
      DataPath_RF_bus_reg_dataout_1594_port, 
      DataPath_RF_bus_reg_dataout_1595_port, 
      DataPath_RF_bus_reg_dataout_1596_port, 
      DataPath_RF_bus_reg_dataout_1597_port, 
      DataPath_RF_bus_reg_dataout_1598_port, 
      DataPath_RF_bus_reg_dataout_1599_port, 
      DataPath_RF_bus_reg_dataout_1600_port, 
      DataPath_RF_bus_reg_dataout_1601_port, 
      DataPath_RF_bus_reg_dataout_1602_port, 
      DataPath_RF_bus_reg_dataout_1603_port, 
      DataPath_RF_bus_reg_dataout_1604_port, 
      DataPath_RF_bus_reg_dataout_1605_port, 
      DataPath_RF_bus_reg_dataout_1606_port, 
      DataPath_RF_bus_reg_dataout_1607_port, 
      DataPath_RF_bus_reg_dataout_1608_port, 
      DataPath_RF_bus_reg_dataout_1609_port, 
      DataPath_RF_bus_reg_dataout_1610_port, 
      DataPath_RF_bus_reg_dataout_1611_port, 
      DataPath_RF_bus_reg_dataout_1612_port, 
      DataPath_RF_bus_reg_dataout_1613_port, 
      DataPath_RF_bus_reg_dataout_1614_port, 
      DataPath_RF_bus_reg_dataout_1615_port, 
      DataPath_RF_bus_reg_dataout_1616_port, 
      DataPath_RF_bus_reg_dataout_1617_port, 
      DataPath_RF_bus_reg_dataout_1618_port, 
      DataPath_RF_bus_reg_dataout_1619_port, 
      DataPath_RF_bus_reg_dataout_1620_port, 
      DataPath_RF_bus_reg_dataout_1621_port, 
      DataPath_RF_bus_reg_dataout_1622_port, 
      DataPath_RF_bus_reg_dataout_1623_port, 
      DataPath_RF_bus_reg_dataout_1624_port, 
      DataPath_RF_bus_reg_dataout_1625_port, 
      DataPath_RF_bus_reg_dataout_1626_port, 
      DataPath_RF_bus_reg_dataout_1627_port, 
      DataPath_RF_bus_reg_dataout_1628_port, 
      DataPath_RF_bus_reg_dataout_1629_port, 
      DataPath_RF_bus_reg_dataout_1630_port, 
      DataPath_RF_bus_reg_dataout_1631_port, 
      DataPath_RF_bus_reg_dataout_1632_port, 
      DataPath_RF_bus_reg_dataout_1633_port, 
      DataPath_RF_bus_reg_dataout_1634_port, 
      DataPath_RF_bus_reg_dataout_1635_port, 
      DataPath_RF_bus_reg_dataout_1636_port, 
      DataPath_RF_bus_reg_dataout_1637_port, 
      DataPath_RF_bus_reg_dataout_1638_port, 
      DataPath_RF_bus_reg_dataout_1639_port, 
      DataPath_RF_bus_reg_dataout_1640_port, 
      DataPath_RF_bus_reg_dataout_1641_port, 
      DataPath_RF_bus_reg_dataout_1642_port, 
      DataPath_RF_bus_reg_dataout_1643_port, 
      DataPath_RF_bus_reg_dataout_1644_port, 
      DataPath_RF_bus_reg_dataout_1645_port, 
      DataPath_RF_bus_reg_dataout_1646_port, 
      DataPath_RF_bus_reg_dataout_1647_port, 
      DataPath_RF_bus_reg_dataout_1648_port, 
      DataPath_RF_bus_reg_dataout_1649_port, 
      DataPath_RF_bus_reg_dataout_1650_port, 
      DataPath_RF_bus_reg_dataout_1651_port, 
      DataPath_RF_bus_reg_dataout_1652_port, 
      DataPath_RF_bus_reg_dataout_1653_port, 
      DataPath_RF_bus_reg_dataout_1654_port, 
      DataPath_RF_bus_reg_dataout_1655_port, 
      DataPath_RF_bus_reg_dataout_1656_port, 
      DataPath_RF_bus_reg_dataout_1657_port, 
      DataPath_RF_bus_reg_dataout_1658_port, 
      DataPath_RF_bus_reg_dataout_1659_port, 
      DataPath_RF_bus_reg_dataout_1660_port, 
      DataPath_RF_bus_reg_dataout_1661_port, 
      DataPath_RF_bus_reg_dataout_1662_port, 
      DataPath_RF_bus_reg_dataout_1663_port, 
      DataPath_RF_bus_reg_dataout_1664_port, 
      DataPath_RF_bus_reg_dataout_1665_port, 
      DataPath_RF_bus_reg_dataout_1666_port, 
      DataPath_RF_bus_reg_dataout_1667_port, 
      DataPath_RF_bus_reg_dataout_1668_port, 
      DataPath_RF_bus_reg_dataout_1669_port, 
      DataPath_RF_bus_reg_dataout_1670_port, 
      DataPath_RF_bus_reg_dataout_1671_port, 
      DataPath_RF_bus_reg_dataout_1672_port, 
      DataPath_RF_bus_reg_dataout_1673_port, 
      DataPath_RF_bus_reg_dataout_1674_port, 
      DataPath_RF_bus_reg_dataout_1675_port, 
      DataPath_RF_bus_reg_dataout_1676_port, 
      DataPath_RF_bus_reg_dataout_1677_port, 
      DataPath_RF_bus_reg_dataout_1678_port, 
      DataPath_RF_bus_reg_dataout_1679_port, 
      DataPath_RF_bus_reg_dataout_1680_port, 
      DataPath_RF_bus_reg_dataout_1681_port, 
      DataPath_RF_bus_reg_dataout_1682_port, 
      DataPath_RF_bus_reg_dataout_1683_port, 
      DataPath_RF_bus_reg_dataout_1684_port, 
      DataPath_RF_bus_reg_dataout_1685_port, 
      DataPath_RF_bus_reg_dataout_1686_port, 
      DataPath_RF_bus_reg_dataout_1687_port, 
      DataPath_RF_bus_reg_dataout_1688_port, 
      DataPath_RF_bus_reg_dataout_1689_port, 
      DataPath_RF_bus_reg_dataout_1690_port, 
      DataPath_RF_bus_reg_dataout_1691_port, 
      DataPath_RF_bus_reg_dataout_1692_port, 
      DataPath_RF_bus_reg_dataout_1693_port, 
      DataPath_RF_bus_reg_dataout_1694_port, 
      DataPath_RF_bus_reg_dataout_1695_port, 
      DataPath_RF_bus_reg_dataout_1696_port, 
      DataPath_RF_bus_reg_dataout_1697_port, 
      DataPath_RF_bus_reg_dataout_1698_port, 
      DataPath_RF_bus_reg_dataout_1699_port, 
      DataPath_RF_bus_reg_dataout_1700_port, 
      DataPath_RF_bus_reg_dataout_1701_port, 
      DataPath_RF_bus_reg_dataout_1702_port, 
      DataPath_RF_bus_reg_dataout_1703_port, 
      DataPath_RF_bus_reg_dataout_1704_port, 
      DataPath_RF_bus_reg_dataout_1705_port, 
      DataPath_RF_bus_reg_dataout_1706_port, 
      DataPath_RF_bus_reg_dataout_1707_port, 
      DataPath_RF_bus_reg_dataout_1708_port, 
      DataPath_RF_bus_reg_dataout_1709_port, 
      DataPath_RF_bus_reg_dataout_1710_port, 
      DataPath_RF_bus_reg_dataout_1711_port, 
      DataPath_RF_bus_reg_dataout_1712_port, 
      DataPath_RF_bus_reg_dataout_1713_port, 
      DataPath_RF_bus_reg_dataout_1714_port, 
      DataPath_RF_bus_reg_dataout_1715_port, 
      DataPath_RF_bus_reg_dataout_1716_port, 
      DataPath_RF_bus_reg_dataout_1717_port, 
      DataPath_RF_bus_reg_dataout_1718_port, 
      DataPath_RF_bus_reg_dataout_1719_port, 
      DataPath_RF_bus_reg_dataout_1720_port, 
      DataPath_RF_bus_reg_dataout_1721_port, 
      DataPath_RF_bus_reg_dataout_1722_port, 
      DataPath_RF_bus_reg_dataout_1723_port, 
      DataPath_RF_bus_reg_dataout_1724_port, 
      DataPath_RF_bus_reg_dataout_1725_port, 
      DataPath_RF_bus_reg_dataout_1726_port, 
      DataPath_RF_bus_reg_dataout_1727_port, 
      DataPath_RF_bus_reg_dataout_1728_port, 
      DataPath_RF_bus_reg_dataout_1729_port, 
      DataPath_RF_bus_reg_dataout_1730_port, 
      DataPath_RF_bus_reg_dataout_1731_port, 
      DataPath_RF_bus_reg_dataout_1732_port, 
      DataPath_RF_bus_reg_dataout_1733_port, 
      DataPath_RF_bus_reg_dataout_1734_port, 
      DataPath_RF_bus_reg_dataout_1735_port, 
      DataPath_RF_bus_reg_dataout_1736_port, 
      DataPath_RF_bus_reg_dataout_1737_port, 
      DataPath_RF_bus_reg_dataout_1738_port, 
      DataPath_RF_bus_reg_dataout_1739_port, 
      DataPath_RF_bus_reg_dataout_1740_port, 
      DataPath_RF_bus_reg_dataout_1741_port, 
      DataPath_RF_bus_reg_dataout_1742_port, 
      DataPath_RF_bus_reg_dataout_1743_port, 
      DataPath_RF_bus_reg_dataout_1744_port, 
      DataPath_RF_bus_reg_dataout_1745_port, 
      DataPath_RF_bus_reg_dataout_1746_port, 
      DataPath_RF_bus_reg_dataout_1747_port, 
      DataPath_RF_bus_reg_dataout_1748_port, 
      DataPath_RF_bus_reg_dataout_1749_port, 
      DataPath_RF_bus_reg_dataout_1750_port, 
      DataPath_RF_bus_reg_dataout_1751_port, 
      DataPath_RF_bus_reg_dataout_1752_port, 
      DataPath_RF_bus_reg_dataout_1753_port, 
      DataPath_RF_bus_reg_dataout_1754_port, 
      DataPath_RF_bus_reg_dataout_1755_port, 
      DataPath_RF_bus_reg_dataout_1756_port, 
      DataPath_RF_bus_reg_dataout_1757_port, 
      DataPath_RF_bus_reg_dataout_1758_port, 
      DataPath_RF_bus_reg_dataout_1759_port, 
      DataPath_RF_bus_reg_dataout_1760_port, 
      DataPath_RF_bus_reg_dataout_1761_port, 
      DataPath_RF_bus_reg_dataout_1762_port, 
      DataPath_RF_bus_reg_dataout_1763_port, 
      DataPath_RF_bus_reg_dataout_1764_port, 
      DataPath_RF_bus_reg_dataout_1765_port, 
      DataPath_RF_bus_reg_dataout_1766_port, 
      DataPath_RF_bus_reg_dataout_1767_port, 
      DataPath_RF_bus_reg_dataout_1768_port, 
      DataPath_RF_bus_reg_dataout_1769_port, 
      DataPath_RF_bus_reg_dataout_1770_port, 
      DataPath_RF_bus_reg_dataout_1771_port, 
      DataPath_RF_bus_reg_dataout_1772_port, 
      DataPath_RF_bus_reg_dataout_1773_port, 
      DataPath_RF_bus_reg_dataout_1774_port, 
      DataPath_RF_bus_reg_dataout_1775_port, 
      DataPath_RF_bus_reg_dataout_1776_port, 
      DataPath_RF_bus_reg_dataout_1777_port, 
      DataPath_RF_bus_reg_dataout_1778_port, 
      DataPath_RF_bus_reg_dataout_1779_port, 
      DataPath_RF_bus_reg_dataout_1780_port, 
      DataPath_RF_bus_reg_dataout_1781_port, 
      DataPath_RF_bus_reg_dataout_1782_port, 
      DataPath_RF_bus_reg_dataout_1783_port, 
      DataPath_RF_bus_reg_dataout_1784_port, 
      DataPath_RF_bus_reg_dataout_1785_port, 
      DataPath_RF_bus_reg_dataout_1786_port, 
      DataPath_RF_bus_reg_dataout_1787_port, 
      DataPath_RF_bus_reg_dataout_1788_port, 
      DataPath_RF_bus_reg_dataout_1789_port, 
      DataPath_RF_bus_reg_dataout_1790_port, 
      DataPath_RF_bus_reg_dataout_1791_port, 
      DataPath_RF_bus_reg_dataout_1792_port, 
      DataPath_RF_bus_reg_dataout_1793_port, 
      DataPath_RF_bus_reg_dataout_1794_port, 
      DataPath_RF_bus_reg_dataout_1795_port, 
      DataPath_RF_bus_reg_dataout_1796_port, 
      DataPath_RF_bus_reg_dataout_1797_port, 
      DataPath_RF_bus_reg_dataout_1798_port, 
      DataPath_RF_bus_reg_dataout_1799_port, 
      DataPath_RF_bus_reg_dataout_1800_port, 
      DataPath_RF_bus_reg_dataout_1801_port, 
      DataPath_RF_bus_reg_dataout_1802_port, 
      DataPath_RF_bus_reg_dataout_1803_port, 
      DataPath_RF_bus_reg_dataout_1804_port, 
      DataPath_RF_bus_reg_dataout_1805_port, 
      DataPath_RF_bus_reg_dataout_1806_port, 
      DataPath_RF_bus_reg_dataout_1807_port, 
      DataPath_RF_bus_reg_dataout_1808_port, 
      DataPath_RF_bus_reg_dataout_1809_port, 
      DataPath_RF_bus_reg_dataout_1810_port, 
      DataPath_RF_bus_reg_dataout_1811_port, 
      DataPath_RF_bus_reg_dataout_1812_port, 
      DataPath_RF_bus_reg_dataout_1813_port, 
      DataPath_RF_bus_reg_dataout_1814_port, 
      DataPath_RF_bus_reg_dataout_1815_port, 
      DataPath_RF_bus_reg_dataout_1816_port, 
      DataPath_RF_bus_reg_dataout_1817_port, 
      DataPath_RF_bus_reg_dataout_1818_port, 
      DataPath_RF_bus_reg_dataout_1819_port, 
      DataPath_RF_bus_reg_dataout_1820_port, 
      DataPath_RF_bus_reg_dataout_1821_port, 
      DataPath_RF_bus_reg_dataout_1822_port, 
      DataPath_RF_bus_reg_dataout_1823_port, 
      DataPath_RF_bus_reg_dataout_1824_port, 
      DataPath_RF_bus_reg_dataout_1825_port, 
      DataPath_RF_bus_reg_dataout_1826_port, 
      DataPath_RF_bus_reg_dataout_1827_port, 
      DataPath_RF_bus_reg_dataout_1828_port, 
      DataPath_RF_bus_reg_dataout_1829_port, 
      DataPath_RF_bus_reg_dataout_1830_port, 
      DataPath_RF_bus_reg_dataout_1831_port, 
      DataPath_RF_bus_reg_dataout_1832_port, 
      DataPath_RF_bus_reg_dataout_1833_port, 
      DataPath_RF_bus_reg_dataout_1834_port, 
      DataPath_RF_bus_reg_dataout_1835_port, 
      DataPath_RF_bus_reg_dataout_1836_port, 
      DataPath_RF_bus_reg_dataout_1837_port, 
      DataPath_RF_bus_reg_dataout_1838_port, 
      DataPath_RF_bus_reg_dataout_1839_port, 
      DataPath_RF_bus_reg_dataout_1840_port, 
      DataPath_RF_bus_reg_dataout_1841_port, 
      DataPath_RF_bus_reg_dataout_1842_port, 
      DataPath_RF_bus_reg_dataout_1843_port, 
      DataPath_RF_bus_reg_dataout_1844_port, 
      DataPath_RF_bus_reg_dataout_1845_port, 
      DataPath_RF_bus_reg_dataout_1846_port, 
      DataPath_RF_bus_reg_dataout_1847_port, 
      DataPath_RF_bus_reg_dataout_1848_port, 
      DataPath_RF_bus_reg_dataout_1849_port, 
      DataPath_RF_bus_reg_dataout_1850_port, 
      DataPath_RF_bus_reg_dataout_1851_port, 
      DataPath_RF_bus_reg_dataout_1852_port, 
      DataPath_RF_bus_reg_dataout_1853_port, 
      DataPath_RF_bus_reg_dataout_1854_port, 
      DataPath_RF_bus_reg_dataout_1855_port, 
      DataPath_RF_bus_reg_dataout_1856_port, 
      DataPath_RF_bus_reg_dataout_1857_port, 
      DataPath_RF_bus_reg_dataout_1858_port, 
      DataPath_RF_bus_reg_dataout_1859_port, 
      DataPath_RF_bus_reg_dataout_1860_port, 
      DataPath_RF_bus_reg_dataout_1861_port, 
      DataPath_RF_bus_reg_dataout_1862_port, 
      DataPath_RF_bus_reg_dataout_1863_port, 
      DataPath_RF_bus_reg_dataout_1864_port, 
      DataPath_RF_bus_reg_dataout_1865_port, 
      DataPath_RF_bus_reg_dataout_1866_port, 
      DataPath_RF_bus_reg_dataout_1867_port, 
      DataPath_RF_bus_reg_dataout_1868_port, 
      DataPath_RF_bus_reg_dataout_1869_port, 
      DataPath_RF_bus_reg_dataout_1870_port, 
      DataPath_RF_bus_reg_dataout_1871_port, 
      DataPath_RF_bus_reg_dataout_1872_port, 
      DataPath_RF_bus_reg_dataout_1873_port, 
      DataPath_RF_bus_reg_dataout_1874_port, 
      DataPath_RF_bus_reg_dataout_1875_port, 
      DataPath_RF_bus_reg_dataout_1876_port, 
      DataPath_RF_bus_reg_dataout_1877_port, 
      DataPath_RF_bus_reg_dataout_1878_port, 
      DataPath_RF_bus_reg_dataout_1879_port, 
      DataPath_RF_bus_reg_dataout_1880_port, 
      DataPath_RF_bus_reg_dataout_1881_port, 
      DataPath_RF_bus_reg_dataout_1882_port, 
      DataPath_RF_bus_reg_dataout_1883_port, 
      DataPath_RF_bus_reg_dataout_1884_port, 
      DataPath_RF_bus_reg_dataout_1885_port, 
      DataPath_RF_bus_reg_dataout_1886_port, 
      DataPath_RF_bus_reg_dataout_1887_port, 
      DataPath_RF_bus_reg_dataout_1888_port, 
      DataPath_RF_bus_reg_dataout_1889_port, 
      DataPath_RF_bus_reg_dataout_1890_port, 
      DataPath_RF_bus_reg_dataout_1891_port, 
      DataPath_RF_bus_reg_dataout_1892_port, 
      DataPath_RF_bus_reg_dataout_1893_port, 
      DataPath_RF_bus_reg_dataout_1894_port, 
      DataPath_RF_bus_reg_dataout_1895_port, 
      DataPath_RF_bus_reg_dataout_1896_port, 
      DataPath_RF_bus_reg_dataout_1897_port, 
      DataPath_RF_bus_reg_dataout_1898_port, 
      DataPath_RF_bus_reg_dataout_1899_port, 
      DataPath_RF_bus_reg_dataout_1900_port, 
      DataPath_RF_bus_reg_dataout_1901_port, 
      DataPath_RF_bus_reg_dataout_1902_port, 
      DataPath_RF_bus_reg_dataout_1903_port, 
      DataPath_RF_bus_reg_dataout_1904_port, 
      DataPath_RF_bus_reg_dataout_1905_port, 
      DataPath_RF_bus_reg_dataout_1906_port, 
      DataPath_RF_bus_reg_dataout_1907_port, 
      DataPath_RF_bus_reg_dataout_1908_port, 
      DataPath_RF_bus_reg_dataout_1909_port, 
      DataPath_RF_bus_reg_dataout_1910_port, 
      DataPath_RF_bus_reg_dataout_1911_port, 
      DataPath_RF_bus_reg_dataout_1912_port, 
      DataPath_RF_bus_reg_dataout_1913_port, 
      DataPath_RF_bus_reg_dataout_1914_port, 
      DataPath_RF_bus_reg_dataout_1915_port, 
      DataPath_RF_bus_reg_dataout_1916_port, 
      DataPath_RF_bus_reg_dataout_1917_port, 
      DataPath_RF_bus_reg_dataout_1918_port, 
      DataPath_RF_bus_reg_dataout_1919_port, 
      DataPath_RF_bus_reg_dataout_1920_port, 
      DataPath_RF_bus_reg_dataout_1921_port, 
      DataPath_RF_bus_reg_dataout_1922_port, 
      DataPath_RF_bus_reg_dataout_1923_port, 
      DataPath_RF_bus_reg_dataout_1924_port, 
      DataPath_RF_bus_reg_dataout_1925_port, 
      DataPath_RF_bus_reg_dataout_1926_port, 
      DataPath_RF_bus_reg_dataout_1927_port, 
      DataPath_RF_bus_reg_dataout_1928_port, 
      DataPath_RF_bus_reg_dataout_1929_port, 
      DataPath_RF_bus_reg_dataout_1930_port, 
      DataPath_RF_bus_reg_dataout_1931_port, 
      DataPath_RF_bus_reg_dataout_1932_port, 
      DataPath_RF_bus_reg_dataout_1933_port, 
      DataPath_RF_bus_reg_dataout_1934_port, 
      DataPath_RF_bus_reg_dataout_1935_port, 
      DataPath_RF_bus_reg_dataout_1936_port, 
      DataPath_RF_bus_reg_dataout_1937_port, 
      DataPath_RF_bus_reg_dataout_1938_port, 
      DataPath_RF_bus_reg_dataout_1939_port, 
      DataPath_RF_bus_reg_dataout_1940_port, 
      DataPath_RF_bus_reg_dataout_1941_port, 
      DataPath_RF_bus_reg_dataout_1942_port, 
      DataPath_RF_bus_reg_dataout_1943_port, 
      DataPath_RF_bus_reg_dataout_1944_port, 
      DataPath_RF_bus_reg_dataout_1945_port, 
      DataPath_RF_bus_reg_dataout_1946_port, 
      DataPath_RF_bus_reg_dataout_1947_port, 
      DataPath_RF_bus_reg_dataout_1948_port, 
      DataPath_RF_bus_reg_dataout_1949_port, 
      DataPath_RF_bus_reg_dataout_1950_port, 
      DataPath_RF_bus_reg_dataout_1951_port, 
      DataPath_RF_bus_reg_dataout_1952_port, 
      DataPath_RF_bus_reg_dataout_1953_port, 
      DataPath_RF_bus_reg_dataout_1954_port, 
      DataPath_RF_bus_reg_dataout_1955_port, 
      DataPath_RF_bus_reg_dataout_1956_port, 
      DataPath_RF_bus_reg_dataout_1957_port, 
      DataPath_RF_bus_reg_dataout_1958_port, 
      DataPath_RF_bus_reg_dataout_1959_port, 
      DataPath_RF_bus_reg_dataout_1960_port, 
      DataPath_RF_bus_reg_dataout_1961_port, 
      DataPath_RF_bus_reg_dataout_1962_port, 
      DataPath_RF_bus_reg_dataout_1963_port, 
      DataPath_RF_bus_reg_dataout_1964_port, 
      DataPath_RF_bus_reg_dataout_1965_port, 
      DataPath_RF_bus_reg_dataout_1966_port, 
      DataPath_RF_bus_reg_dataout_1967_port, 
      DataPath_RF_bus_reg_dataout_1968_port, 
      DataPath_RF_bus_reg_dataout_1969_port, 
      DataPath_RF_bus_reg_dataout_1970_port, 
      DataPath_RF_bus_reg_dataout_1971_port, 
      DataPath_RF_bus_reg_dataout_1972_port, 
      DataPath_RF_bus_reg_dataout_1973_port, 
      DataPath_RF_bus_reg_dataout_1974_port, 
      DataPath_RF_bus_reg_dataout_1975_port, 
      DataPath_RF_bus_reg_dataout_1976_port, 
      DataPath_RF_bus_reg_dataout_1977_port, 
      DataPath_RF_bus_reg_dataout_1978_port, 
      DataPath_RF_bus_reg_dataout_1979_port, 
      DataPath_RF_bus_reg_dataout_1980_port, 
      DataPath_RF_bus_reg_dataout_1981_port, 
      DataPath_RF_bus_reg_dataout_1982_port, 
      DataPath_RF_bus_reg_dataout_1983_port, 
      DataPath_RF_bus_reg_dataout_1984_port, 
      DataPath_RF_bus_reg_dataout_1985_port, 
      DataPath_RF_bus_reg_dataout_1986_port, 
      DataPath_RF_bus_reg_dataout_1987_port, 
      DataPath_RF_bus_reg_dataout_1988_port, 
      DataPath_RF_bus_reg_dataout_1989_port, 
      DataPath_RF_bus_reg_dataout_1990_port, 
      DataPath_RF_bus_reg_dataout_1991_port, 
      DataPath_RF_bus_reg_dataout_1992_port, 
      DataPath_RF_bus_reg_dataout_1993_port, 
      DataPath_RF_bus_reg_dataout_1994_port, 
      DataPath_RF_bus_reg_dataout_1995_port, 
      DataPath_RF_bus_reg_dataout_1996_port, 
      DataPath_RF_bus_reg_dataout_1997_port, 
      DataPath_RF_bus_reg_dataout_1998_port, 
      DataPath_RF_bus_reg_dataout_1999_port, 
      DataPath_RF_bus_reg_dataout_2000_port, 
      DataPath_RF_bus_reg_dataout_2001_port, 
      DataPath_RF_bus_reg_dataout_2002_port, 
      DataPath_RF_bus_reg_dataout_2003_port, 
      DataPath_RF_bus_reg_dataout_2004_port, 
      DataPath_RF_bus_reg_dataout_2005_port, 
      DataPath_RF_bus_reg_dataout_2006_port, 
      DataPath_RF_bus_reg_dataout_2007_port, 
      DataPath_RF_bus_reg_dataout_2008_port, 
      DataPath_RF_bus_reg_dataout_2009_port, 
      DataPath_RF_bus_reg_dataout_2010_port, 
      DataPath_RF_bus_reg_dataout_2011_port, 
      DataPath_RF_bus_reg_dataout_2012_port, 
      DataPath_RF_bus_reg_dataout_2013_port, 
      DataPath_RF_bus_reg_dataout_2014_port, 
      DataPath_RF_bus_reg_dataout_2015_port, 
      DataPath_RF_bus_reg_dataout_2016_port, 
      DataPath_RF_bus_reg_dataout_2017_port, 
      DataPath_RF_bus_reg_dataout_2018_port, 
      DataPath_RF_bus_reg_dataout_2019_port, 
      DataPath_RF_bus_reg_dataout_2020_port, 
      DataPath_RF_bus_reg_dataout_2021_port, 
      DataPath_RF_bus_reg_dataout_2022_port, 
      DataPath_RF_bus_reg_dataout_2023_port, 
      DataPath_RF_bus_reg_dataout_2024_port, 
      DataPath_RF_bus_reg_dataout_2025_port, 
      DataPath_RF_bus_reg_dataout_2026_port, 
      DataPath_RF_bus_reg_dataout_2027_port, 
      DataPath_RF_bus_reg_dataout_2028_port, 
      DataPath_RF_bus_reg_dataout_2029_port, 
      DataPath_RF_bus_reg_dataout_2030_port, 
      DataPath_RF_bus_reg_dataout_2031_port, 
      DataPath_RF_bus_reg_dataout_2032_port, 
      DataPath_RF_bus_reg_dataout_2033_port, 
      DataPath_RF_bus_reg_dataout_2034_port, 
      DataPath_RF_bus_reg_dataout_2035_port, 
      DataPath_RF_bus_reg_dataout_2036_port, 
      DataPath_RF_bus_reg_dataout_2037_port, 
      DataPath_RF_bus_reg_dataout_2038_port, 
      DataPath_RF_bus_reg_dataout_2039_port, 
      DataPath_RF_bus_reg_dataout_2040_port, 
      DataPath_RF_bus_reg_dataout_2041_port, 
      DataPath_RF_bus_reg_dataout_2042_port, 
      DataPath_RF_bus_reg_dataout_2043_port, 
      DataPath_RF_bus_reg_dataout_2044_port, 
      DataPath_RF_bus_reg_dataout_2045_port, 
      DataPath_RF_bus_reg_dataout_2046_port, 
      DataPath_RF_bus_reg_dataout_2047_port, 
      DataPath_RF_bus_reg_dataout_2048_port, 
      DataPath_RF_bus_reg_dataout_2049_port, 
      DataPath_RF_bus_reg_dataout_2050_port, 
      DataPath_RF_bus_reg_dataout_2051_port, 
      DataPath_RF_bus_reg_dataout_2052_port, 
      DataPath_RF_bus_reg_dataout_2053_port, 
      DataPath_RF_bus_reg_dataout_2054_port, 
      DataPath_RF_bus_reg_dataout_2055_port, 
      DataPath_RF_bus_reg_dataout_2056_port, 
      DataPath_RF_bus_reg_dataout_2057_port, 
      DataPath_RF_bus_reg_dataout_2058_port, 
      DataPath_RF_bus_reg_dataout_2059_port, 
      DataPath_RF_bus_reg_dataout_2060_port, 
      DataPath_RF_bus_reg_dataout_2061_port, 
      DataPath_RF_bus_reg_dataout_2062_port, 
      DataPath_RF_bus_reg_dataout_2063_port, 
      DataPath_RF_bus_reg_dataout_2064_port, 
      DataPath_RF_bus_reg_dataout_2065_port, 
      DataPath_RF_bus_reg_dataout_2066_port, 
      DataPath_RF_bus_reg_dataout_2067_port, 
      DataPath_RF_bus_reg_dataout_2068_port, 
      DataPath_RF_bus_reg_dataout_2069_port, 
      DataPath_RF_bus_reg_dataout_2070_port, 
      DataPath_RF_bus_reg_dataout_2071_port, 
      DataPath_RF_bus_reg_dataout_2072_port, 
      DataPath_RF_bus_reg_dataout_2073_port, 
      DataPath_RF_bus_reg_dataout_2074_port, 
      DataPath_RF_bus_reg_dataout_2075_port, 
      DataPath_RF_bus_reg_dataout_2076_port, 
      DataPath_RF_bus_reg_dataout_2077_port, 
      DataPath_RF_bus_reg_dataout_2078_port, 
      DataPath_RF_bus_reg_dataout_2079_port, 
      DataPath_RF_bus_reg_dataout_2080_port, 
      DataPath_RF_bus_reg_dataout_2081_port, 
      DataPath_RF_bus_reg_dataout_2082_port, 
      DataPath_RF_bus_reg_dataout_2083_port, 
      DataPath_RF_bus_reg_dataout_2084_port, 
      DataPath_RF_bus_reg_dataout_2085_port, 
      DataPath_RF_bus_reg_dataout_2086_port, 
      DataPath_RF_bus_reg_dataout_2087_port, 
      DataPath_RF_bus_reg_dataout_2088_port, 
      DataPath_RF_bus_reg_dataout_2089_port, 
      DataPath_RF_bus_reg_dataout_2090_port, 
      DataPath_RF_bus_reg_dataout_2091_port, 
      DataPath_RF_bus_reg_dataout_2092_port, 
      DataPath_RF_bus_reg_dataout_2093_port, 
      DataPath_RF_bus_reg_dataout_2094_port, 
      DataPath_RF_bus_reg_dataout_2095_port, 
      DataPath_RF_bus_reg_dataout_2096_port, 
      DataPath_RF_bus_reg_dataout_2097_port, 
      DataPath_RF_bus_reg_dataout_2098_port, 
      DataPath_RF_bus_reg_dataout_2099_port, 
      DataPath_RF_bus_reg_dataout_2100_port, 
      DataPath_RF_bus_reg_dataout_2101_port, 
      DataPath_RF_bus_reg_dataout_2102_port, 
      DataPath_RF_bus_reg_dataout_2103_port, 
      DataPath_RF_bus_reg_dataout_2104_port, 
      DataPath_RF_bus_reg_dataout_2105_port, 
      DataPath_RF_bus_reg_dataout_2106_port, 
      DataPath_RF_bus_reg_dataout_2107_port, 
      DataPath_RF_bus_reg_dataout_2108_port, 
      DataPath_RF_bus_reg_dataout_2109_port, 
      DataPath_RF_bus_reg_dataout_2110_port, 
      DataPath_RF_bus_reg_dataout_2111_port, 
      DataPath_RF_bus_reg_dataout_2112_port, 
      DataPath_RF_bus_reg_dataout_2113_port, 
      DataPath_RF_bus_reg_dataout_2114_port, 
      DataPath_RF_bus_reg_dataout_2115_port, 
      DataPath_RF_bus_reg_dataout_2116_port, 
      DataPath_RF_bus_reg_dataout_2117_port, 
      DataPath_RF_bus_reg_dataout_2118_port, 
      DataPath_RF_bus_reg_dataout_2119_port, 
      DataPath_RF_bus_reg_dataout_2120_port, 
      DataPath_RF_bus_reg_dataout_2121_port, 
      DataPath_RF_bus_reg_dataout_2122_port, 
      DataPath_RF_bus_reg_dataout_2123_port, 
      DataPath_RF_bus_reg_dataout_2124_port, 
      DataPath_RF_bus_reg_dataout_2125_port, 
      DataPath_RF_bus_reg_dataout_2126_port, 
      DataPath_RF_bus_reg_dataout_2127_port, 
      DataPath_RF_bus_reg_dataout_2128_port, 
      DataPath_RF_bus_reg_dataout_2129_port, 
      DataPath_RF_bus_reg_dataout_2130_port, 
      DataPath_RF_bus_reg_dataout_2131_port, 
      DataPath_RF_bus_reg_dataout_2132_port, 
      DataPath_RF_bus_reg_dataout_2133_port, 
      DataPath_RF_bus_reg_dataout_2134_port, 
      DataPath_RF_bus_reg_dataout_2135_port, 
      DataPath_RF_bus_reg_dataout_2136_port, 
      DataPath_RF_bus_reg_dataout_2137_port, 
      DataPath_RF_bus_reg_dataout_2138_port, 
      DataPath_RF_bus_reg_dataout_2139_port, 
      DataPath_RF_bus_reg_dataout_2140_port, 
      DataPath_RF_bus_reg_dataout_2141_port, 
      DataPath_RF_bus_reg_dataout_2142_port, 
      DataPath_RF_bus_reg_dataout_2143_port, 
      DataPath_RF_bus_reg_dataout_2144_port, 
      DataPath_RF_bus_reg_dataout_2145_port, 
      DataPath_RF_bus_reg_dataout_2146_port, 
      DataPath_RF_bus_reg_dataout_2147_port, 
      DataPath_RF_bus_reg_dataout_2148_port, 
      DataPath_RF_bus_reg_dataout_2149_port, 
      DataPath_RF_bus_reg_dataout_2150_port, 
      DataPath_RF_bus_reg_dataout_2151_port, 
      DataPath_RF_bus_reg_dataout_2152_port, 
      DataPath_RF_bus_reg_dataout_2153_port, 
      DataPath_RF_bus_reg_dataout_2154_port, 
      DataPath_RF_bus_reg_dataout_2155_port, 
      DataPath_RF_bus_reg_dataout_2156_port, 
      DataPath_RF_bus_reg_dataout_2157_port, 
      DataPath_RF_bus_reg_dataout_2158_port, 
      DataPath_RF_bus_reg_dataout_2159_port, 
      DataPath_RF_bus_reg_dataout_2160_port, 
      DataPath_RF_bus_reg_dataout_2161_port, 
      DataPath_RF_bus_reg_dataout_2162_port, 
      DataPath_RF_bus_reg_dataout_2163_port, 
      DataPath_RF_bus_reg_dataout_2164_port, 
      DataPath_RF_bus_reg_dataout_2165_port, 
      DataPath_RF_bus_reg_dataout_2166_port, 
      DataPath_RF_bus_reg_dataout_2167_port, 
      DataPath_RF_bus_reg_dataout_2168_port, 
      DataPath_RF_bus_reg_dataout_2169_port, 
      DataPath_RF_bus_reg_dataout_2170_port, 
      DataPath_RF_bus_reg_dataout_2171_port, 
      DataPath_RF_bus_reg_dataout_2172_port, 
      DataPath_RF_bus_reg_dataout_2173_port, 
      DataPath_RF_bus_reg_dataout_2174_port, 
      DataPath_RF_bus_reg_dataout_2175_port, 
      DataPath_RF_bus_reg_dataout_2176_port, 
      DataPath_RF_bus_reg_dataout_2177_port, 
      DataPath_RF_bus_reg_dataout_2178_port, 
      DataPath_RF_bus_reg_dataout_2179_port, 
      DataPath_RF_bus_reg_dataout_2180_port, 
      DataPath_RF_bus_reg_dataout_2181_port, 
      DataPath_RF_bus_reg_dataout_2182_port, 
      DataPath_RF_bus_reg_dataout_2183_port, 
      DataPath_RF_bus_reg_dataout_2184_port, 
      DataPath_RF_bus_reg_dataout_2185_port, 
      DataPath_RF_bus_reg_dataout_2186_port, 
      DataPath_RF_bus_reg_dataout_2187_port, 
      DataPath_RF_bus_reg_dataout_2188_port, 
      DataPath_RF_bus_reg_dataout_2189_port, 
      DataPath_RF_bus_reg_dataout_2190_port, 
      DataPath_RF_bus_reg_dataout_2191_port, 
      DataPath_RF_bus_reg_dataout_2192_port, 
      DataPath_RF_bus_reg_dataout_2193_port, 
      DataPath_RF_bus_reg_dataout_2194_port, 
      DataPath_RF_bus_reg_dataout_2195_port, 
      DataPath_RF_bus_reg_dataout_2196_port, 
      DataPath_RF_bus_reg_dataout_2197_port, 
      DataPath_RF_bus_reg_dataout_2198_port, 
      DataPath_RF_bus_reg_dataout_2199_port, 
      DataPath_RF_bus_reg_dataout_2200_port, 
      DataPath_RF_bus_reg_dataout_2201_port, 
      DataPath_RF_bus_reg_dataout_2202_port, 
      DataPath_RF_bus_reg_dataout_2203_port, 
      DataPath_RF_bus_reg_dataout_2204_port, 
      DataPath_RF_bus_reg_dataout_2205_port, 
      DataPath_RF_bus_reg_dataout_2206_port, 
      DataPath_RF_bus_reg_dataout_2207_port, 
      DataPath_RF_bus_reg_dataout_2208_port, 
      DataPath_RF_bus_reg_dataout_2209_port, 
      DataPath_RF_bus_reg_dataout_2210_port, 
      DataPath_RF_bus_reg_dataout_2211_port, 
      DataPath_RF_bus_reg_dataout_2212_port, 
      DataPath_RF_bus_reg_dataout_2213_port, 
      DataPath_RF_bus_reg_dataout_2214_port, 
      DataPath_RF_bus_reg_dataout_2215_port, 
      DataPath_RF_bus_reg_dataout_2216_port, 
      DataPath_RF_bus_reg_dataout_2217_port, 
      DataPath_RF_bus_reg_dataout_2218_port, 
      DataPath_RF_bus_reg_dataout_2219_port, 
      DataPath_RF_bus_reg_dataout_2220_port, 
      DataPath_RF_bus_reg_dataout_2221_port, 
      DataPath_RF_bus_reg_dataout_2222_port, 
      DataPath_RF_bus_reg_dataout_2223_port, 
      DataPath_RF_bus_reg_dataout_2224_port, 
      DataPath_RF_bus_reg_dataout_2225_port, 
      DataPath_RF_bus_reg_dataout_2226_port, 
      DataPath_RF_bus_reg_dataout_2227_port, 
      DataPath_RF_bus_reg_dataout_2228_port, 
      DataPath_RF_bus_reg_dataout_2229_port, 
      DataPath_RF_bus_reg_dataout_2230_port, 
      DataPath_RF_bus_reg_dataout_2231_port, 
      DataPath_RF_bus_reg_dataout_2232_port, 
      DataPath_RF_bus_reg_dataout_2233_port, 
      DataPath_RF_bus_reg_dataout_2234_port, 
      DataPath_RF_bus_reg_dataout_2235_port, 
      DataPath_RF_bus_reg_dataout_2236_port, 
      DataPath_RF_bus_reg_dataout_2237_port, 
      DataPath_RF_bus_reg_dataout_2238_port, 
      DataPath_RF_bus_reg_dataout_2239_port, 
      DataPath_RF_bus_reg_dataout_2240_port, 
      DataPath_RF_bus_reg_dataout_2241_port, 
      DataPath_RF_bus_reg_dataout_2242_port, 
      DataPath_RF_bus_reg_dataout_2243_port, 
      DataPath_RF_bus_reg_dataout_2244_port, 
      DataPath_RF_bus_reg_dataout_2245_port, 
      DataPath_RF_bus_reg_dataout_2246_port, 
      DataPath_RF_bus_reg_dataout_2247_port, 
      DataPath_RF_bus_reg_dataout_2248_port, 
      DataPath_RF_bus_reg_dataout_2249_port, 
      DataPath_RF_bus_reg_dataout_2250_port, 
      DataPath_RF_bus_reg_dataout_2251_port, 
      DataPath_RF_bus_reg_dataout_2252_port, 
      DataPath_RF_bus_reg_dataout_2253_port, 
      DataPath_RF_bus_reg_dataout_2254_port, 
      DataPath_RF_bus_reg_dataout_2255_port, 
      DataPath_RF_bus_reg_dataout_2256_port, 
      DataPath_RF_bus_reg_dataout_2257_port, 
      DataPath_RF_bus_reg_dataout_2258_port, 
      DataPath_RF_bus_reg_dataout_2259_port, 
      DataPath_RF_bus_reg_dataout_2260_port, 
      DataPath_RF_bus_reg_dataout_2261_port, 
      DataPath_RF_bus_reg_dataout_2262_port, 
      DataPath_RF_bus_reg_dataout_2263_port, 
      DataPath_RF_bus_reg_dataout_2264_port, 
      DataPath_RF_bus_reg_dataout_2265_port, 
      DataPath_RF_bus_reg_dataout_2266_port, 
      DataPath_RF_bus_reg_dataout_2267_port, 
      DataPath_RF_bus_reg_dataout_2268_port, 
      DataPath_RF_bus_reg_dataout_2269_port, 
      DataPath_RF_bus_reg_dataout_2270_port, 
      DataPath_RF_bus_reg_dataout_2271_port, 
      DataPath_RF_bus_reg_dataout_2272_port, 
      DataPath_RF_bus_reg_dataout_2273_port, 
      DataPath_RF_bus_reg_dataout_2274_port, 
      DataPath_RF_bus_reg_dataout_2275_port, 
      DataPath_RF_bus_reg_dataout_2276_port, 
      DataPath_RF_bus_reg_dataout_2277_port, 
      DataPath_RF_bus_reg_dataout_2278_port, 
      DataPath_RF_bus_reg_dataout_2279_port, 
      DataPath_RF_bus_reg_dataout_2280_port, 
      DataPath_RF_bus_reg_dataout_2281_port, 
      DataPath_RF_bus_reg_dataout_2282_port, 
      DataPath_RF_bus_reg_dataout_2283_port, 
      DataPath_RF_bus_reg_dataout_2284_port, 
      DataPath_RF_bus_reg_dataout_2285_port, 
      DataPath_RF_bus_reg_dataout_2286_port, 
      DataPath_RF_bus_reg_dataout_2287_port, 
      DataPath_RF_bus_reg_dataout_2288_port, 
      DataPath_RF_bus_reg_dataout_2289_port, 
      DataPath_RF_bus_reg_dataout_2290_port, 
      DataPath_RF_bus_reg_dataout_2291_port, 
      DataPath_RF_bus_reg_dataout_2292_port, 
      DataPath_RF_bus_reg_dataout_2293_port, 
      DataPath_RF_bus_reg_dataout_2294_port, 
      DataPath_RF_bus_reg_dataout_2295_port, 
      DataPath_RF_bus_reg_dataout_2296_port, 
      DataPath_RF_bus_reg_dataout_2297_port, 
      DataPath_RF_bus_reg_dataout_2298_port, 
      DataPath_RF_bus_reg_dataout_2299_port, 
      DataPath_RF_bus_reg_dataout_2300_port, 
      DataPath_RF_bus_reg_dataout_2301_port, 
      DataPath_RF_bus_reg_dataout_2302_port, 
      DataPath_RF_bus_reg_dataout_2303_port, 
      DataPath_RF_bus_reg_dataout_2304_port, 
      DataPath_RF_bus_reg_dataout_2305_port, 
      DataPath_RF_bus_reg_dataout_2306_port, 
      DataPath_RF_bus_reg_dataout_2307_port, 
      DataPath_RF_bus_reg_dataout_2308_port, 
      DataPath_RF_bus_reg_dataout_2309_port, 
      DataPath_RF_bus_reg_dataout_2310_port, 
      DataPath_RF_bus_reg_dataout_2311_port, 
      DataPath_RF_bus_reg_dataout_2312_port, 
      DataPath_RF_bus_reg_dataout_2313_port, 
      DataPath_RF_bus_reg_dataout_2314_port, 
      DataPath_RF_bus_reg_dataout_2315_port, 
      DataPath_RF_bus_reg_dataout_2316_port, 
      DataPath_RF_bus_reg_dataout_2317_port, 
      DataPath_RF_bus_reg_dataout_2318_port, 
      DataPath_RF_bus_reg_dataout_2319_port, 
      DataPath_RF_bus_reg_dataout_2320_port, 
      DataPath_RF_bus_reg_dataout_2321_port, 
      DataPath_RF_bus_reg_dataout_2322_port, 
      DataPath_RF_bus_reg_dataout_2323_port, 
      DataPath_RF_bus_reg_dataout_2324_port, 
      DataPath_RF_bus_reg_dataout_2325_port, 
      DataPath_RF_bus_reg_dataout_2326_port, 
      DataPath_RF_bus_reg_dataout_2327_port, 
      DataPath_RF_bus_reg_dataout_2328_port, 
      DataPath_RF_bus_reg_dataout_2329_port, 
      DataPath_RF_bus_reg_dataout_2330_port, 
      DataPath_RF_bus_reg_dataout_2331_port, 
      DataPath_RF_bus_reg_dataout_2332_port, 
      DataPath_RF_bus_reg_dataout_2333_port, 
      DataPath_RF_bus_reg_dataout_2334_port, 
      DataPath_RF_bus_reg_dataout_2335_port, 
      DataPath_RF_bus_reg_dataout_2336_port, 
      DataPath_RF_bus_reg_dataout_2337_port, 
      DataPath_RF_bus_reg_dataout_2338_port, 
      DataPath_RF_bus_reg_dataout_2339_port, 
      DataPath_RF_bus_reg_dataout_2340_port, 
      DataPath_RF_bus_reg_dataout_2341_port, 
      DataPath_RF_bus_reg_dataout_2342_port, 
      DataPath_RF_bus_reg_dataout_2343_port, 
      DataPath_RF_bus_reg_dataout_2344_port, 
      DataPath_RF_bus_reg_dataout_2345_port, 
      DataPath_RF_bus_reg_dataout_2346_port, 
      DataPath_RF_bus_reg_dataout_2347_port, 
      DataPath_RF_bus_reg_dataout_2348_port, 
      DataPath_RF_bus_reg_dataout_2349_port, 
      DataPath_RF_bus_reg_dataout_2350_port, 
      DataPath_RF_bus_reg_dataout_2351_port, 
      DataPath_RF_bus_reg_dataout_2352_port, 
      DataPath_RF_bus_reg_dataout_2353_port, 
      DataPath_RF_bus_reg_dataout_2354_port, 
      DataPath_RF_bus_reg_dataout_2355_port, 
      DataPath_RF_bus_reg_dataout_2356_port, 
      DataPath_RF_bus_reg_dataout_2357_port, 
      DataPath_RF_bus_reg_dataout_2358_port, 
      DataPath_RF_bus_reg_dataout_2359_port, 
      DataPath_RF_bus_reg_dataout_2360_port, 
      DataPath_RF_bus_reg_dataout_2361_port, 
      DataPath_RF_bus_reg_dataout_2362_port, 
      DataPath_RF_bus_reg_dataout_2363_port, 
      DataPath_RF_bus_reg_dataout_2364_port, 
      DataPath_RF_bus_reg_dataout_2365_port, 
      DataPath_RF_bus_reg_dataout_2366_port, 
      DataPath_RF_bus_reg_dataout_2367_port, 
      DataPath_RF_bus_reg_dataout_2368_port, 
      DataPath_RF_bus_reg_dataout_2369_port, 
      DataPath_RF_bus_reg_dataout_2370_port, 
      DataPath_RF_bus_reg_dataout_2371_port, 
      DataPath_RF_bus_reg_dataout_2372_port, 
      DataPath_RF_bus_reg_dataout_2373_port, 
      DataPath_RF_bus_reg_dataout_2374_port, 
      DataPath_RF_bus_reg_dataout_2375_port, 
      DataPath_RF_bus_reg_dataout_2376_port, 
      DataPath_RF_bus_reg_dataout_2377_port, 
      DataPath_RF_bus_reg_dataout_2378_port, 
      DataPath_RF_bus_reg_dataout_2379_port, 
      DataPath_RF_bus_reg_dataout_2380_port, 
      DataPath_RF_bus_reg_dataout_2381_port, 
      DataPath_RF_bus_reg_dataout_2382_port, 
      DataPath_RF_bus_reg_dataout_2383_port, 
      DataPath_RF_bus_reg_dataout_2384_port, 
      DataPath_RF_bus_reg_dataout_2385_port, 
      DataPath_RF_bus_reg_dataout_2386_port, 
      DataPath_RF_bus_reg_dataout_2387_port, 
      DataPath_RF_bus_reg_dataout_2388_port, 
      DataPath_RF_bus_reg_dataout_2389_port, 
      DataPath_RF_bus_reg_dataout_2390_port, 
      DataPath_RF_bus_reg_dataout_2391_port, 
      DataPath_RF_bus_reg_dataout_2392_port, 
      DataPath_RF_bus_reg_dataout_2393_port, 
      DataPath_RF_bus_reg_dataout_2394_port, 
      DataPath_RF_bus_reg_dataout_2395_port, 
      DataPath_RF_bus_reg_dataout_2396_port, 
      DataPath_RF_bus_reg_dataout_2397_port, 
      DataPath_RF_bus_reg_dataout_2398_port, 
      DataPath_RF_bus_reg_dataout_2399_port, 
      DataPath_RF_bus_reg_dataout_2400_port, 
      DataPath_RF_bus_reg_dataout_2401_port, 
      DataPath_RF_bus_reg_dataout_2402_port, 
      DataPath_RF_bus_reg_dataout_2403_port, 
      DataPath_RF_bus_reg_dataout_2404_port, 
      DataPath_RF_bus_reg_dataout_2405_port, 
      DataPath_RF_bus_reg_dataout_2406_port, 
      DataPath_RF_bus_reg_dataout_2407_port, 
      DataPath_RF_bus_reg_dataout_2408_port, 
      DataPath_RF_bus_reg_dataout_2409_port, 
      DataPath_RF_bus_reg_dataout_2410_port, 
      DataPath_RF_bus_reg_dataout_2411_port, 
      DataPath_RF_bus_reg_dataout_2412_port, 
      DataPath_RF_bus_reg_dataout_2413_port, 
      DataPath_RF_bus_reg_dataout_2414_port, 
      DataPath_RF_bus_reg_dataout_2415_port, 
      DataPath_RF_bus_reg_dataout_2416_port, 
      DataPath_RF_bus_reg_dataout_2417_port, 
      DataPath_RF_bus_reg_dataout_2418_port, 
      DataPath_RF_bus_reg_dataout_2419_port, 
      DataPath_RF_bus_reg_dataout_2420_port, 
      DataPath_RF_bus_reg_dataout_2421_port, 
      DataPath_RF_bus_reg_dataout_2422_port, 
      DataPath_RF_bus_reg_dataout_2423_port, 
      DataPath_RF_bus_reg_dataout_2424_port, 
      DataPath_RF_bus_reg_dataout_2425_port, 
      DataPath_RF_bus_reg_dataout_2426_port, 
      DataPath_RF_bus_reg_dataout_2427_port, 
      DataPath_RF_bus_reg_dataout_2428_port, 
      DataPath_RF_bus_reg_dataout_2429_port, 
      DataPath_RF_bus_reg_dataout_2430_port, 
      DataPath_RF_bus_reg_dataout_2431_port, 
      DataPath_RF_bus_reg_dataout_2432_port, 
      DataPath_RF_bus_reg_dataout_2433_port, 
      DataPath_RF_bus_reg_dataout_2434_port, 
      DataPath_RF_bus_reg_dataout_2435_port, 
      DataPath_RF_bus_reg_dataout_2436_port, 
      DataPath_RF_bus_reg_dataout_2437_port, 
      DataPath_RF_bus_reg_dataout_2438_port, 
      DataPath_RF_bus_reg_dataout_2439_port, 
      DataPath_RF_bus_reg_dataout_2440_port, 
      DataPath_RF_bus_reg_dataout_2441_port, 
      DataPath_RF_bus_reg_dataout_2442_port, 
      DataPath_RF_bus_reg_dataout_2443_port, 
      DataPath_RF_bus_reg_dataout_2444_port, 
      DataPath_RF_bus_reg_dataout_2445_port, 
      DataPath_RF_bus_reg_dataout_2446_port, 
      DataPath_RF_bus_reg_dataout_2447_port, 
      DataPath_RF_bus_reg_dataout_2448_port, 
      DataPath_RF_bus_reg_dataout_2449_port, 
      DataPath_RF_bus_reg_dataout_2450_port, 
      DataPath_RF_bus_reg_dataout_2451_port, 
      DataPath_RF_bus_reg_dataout_2452_port, 
      DataPath_RF_bus_reg_dataout_2453_port, 
      DataPath_RF_bus_reg_dataout_2454_port, 
      DataPath_RF_bus_reg_dataout_2455_port, 
      DataPath_RF_bus_reg_dataout_2456_port, 
      DataPath_RF_bus_reg_dataout_2457_port, 
      DataPath_RF_bus_reg_dataout_2458_port, 
      DataPath_RF_bus_reg_dataout_2459_port, 
      DataPath_RF_bus_reg_dataout_2460_port, 
      DataPath_RF_bus_reg_dataout_2461_port, 
      DataPath_RF_bus_reg_dataout_2462_port, 
      DataPath_RF_bus_reg_dataout_2463_port, 
      DataPath_RF_bus_reg_dataout_2464_port, 
      DataPath_RF_bus_reg_dataout_2465_port, 
      DataPath_RF_bus_reg_dataout_2466_port, 
      DataPath_RF_bus_reg_dataout_2467_port, 
      DataPath_RF_bus_reg_dataout_2468_port, 
      DataPath_RF_bus_reg_dataout_2469_port, 
      DataPath_RF_bus_reg_dataout_2470_port, 
      DataPath_RF_bus_reg_dataout_2471_port, 
      DataPath_RF_bus_reg_dataout_2472_port, 
      DataPath_RF_bus_reg_dataout_2473_port, 
      DataPath_RF_bus_reg_dataout_2474_port, 
      DataPath_RF_bus_reg_dataout_2475_port, 
      DataPath_RF_bus_reg_dataout_2476_port, 
      DataPath_RF_bus_reg_dataout_2477_port, 
      DataPath_RF_bus_reg_dataout_2478_port, 
      DataPath_RF_bus_reg_dataout_2479_port, 
      DataPath_RF_bus_reg_dataout_2480_port, 
      DataPath_RF_bus_reg_dataout_2481_port, 
      DataPath_RF_bus_reg_dataout_2482_port, 
      DataPath_RF_bus_reg_dataout_2483_port, 
      DataPath_RF_bus_reg_dataout_2484_port, 
      DataPath_RF_bus_reg_dataout_2485_port, 
      DataPath_RF_bus_reg_dataout_2486_port, 
      DataPath_RF_bus_reg_dataout_2487_port, 
      DataPath_RF_bus_reg_dataout_2488_port, 
      DataPath_RF_bus_reg_dataout_2489_port, 
      DataPath_RF_bus_reg_dataout_2490_port, 
      DataPath_RF_bus_reg_dataout_2491_port, 
      DataPath_RF_bus_reg_dataout_2492_port, 
      DataPath_RF_bus_reg_dataout_2493_port, 
      DataPath_RF_bus_reg_dataout_2494_port, 
      DataPath_RF_bus_reg_dataout_2495_port, 
      DataPath_RF_bus_reg_dataout_2496_port, 
      DataPath_RF_bus_reg_dataout_2497_port, 
      DataPath_RF_bus_reg_dataout_2498_port, 
      DataPath_RF_bus_reg_dataout_2499_port, 
      DataPath_RF_bus_reg_dataout_2500_port, 
      DataPath_RF_bus_reg_dataout_2501_port, 
      DataPath_RF_bus_reg_dataout_2502_port, 
      DataPath_RF_bus_reg_dataout_2503_port, 
      DataPath_RF_bus_reg_dataout_2504_port, 
      DataPath_RF_bus_reg_dataout_2505_port, 
      DataPath_RF_bus_reg_dataout_2506_port, 
      DataPath_RF_bus_reg_dataout_2507_port, 
      DataPath_RF_bus_reg_dataout_2508_port, 
      DataPath_RF_bus_reg_dataout_2509_port, 
      DataPath_RF_bus_reg_dataout_2510_port, 
      DataPath_RF_bus_reg_dataout_2511_port, 
      DataPath_RF_bus_reg_dataout_2512_port, 
      DataPath_RF_bus_reg_dataout_2513_port, 
      DataPath_RF_bus_reg_dataout_2514_port, 
      DataPath_RF_bus_reg_dataout_2515_port, 
      DataPath_RF_bus_reg_dataout_2516_port, 
      DataPath_RF_bus_reg_dataout_2517_port, 
      DataPath_RF_bus_reg_dataout_2518_port, 
      DataPath_RF_bus_reg_dataout_2519_port, 
      DataPath_RF_bus_reg_dataout_2520_port, 
      DataPath_RF_bus_reg_dataout_2521_port, 
      DataPath_RF_bus_reg_dataout_2522_port, 
      DataPath_RF_bus_reg_dataout_2523_port, 
      DataPath_RF_bus_reg_dataout_2524_port, 
      DataPath_RF_bus_reg_dataout_2525_port, 
      DataPath_RF_bus_reg_dataout_2526_port, 
      DataPath_RF_bus_reg_dataout_2527_port, 
      DataPath_RF_bus_reg_dataout_2528_port, 
      DataPath_RF_bus_reg_dataout_2529_port, 
      DataPath_RF_bus_reg_dataout_2530_port, 
      DataPath_RF_bus_reg_dataout_2531_port, 
      DataPath_RF_bus_reg_dataout_2532_port, 
      DataPath_RF_bus_reg_dataout_2533_port, 
      DataPath_RF_bus_reg_dataout_2534_port, 
      DataPath_RF_bus_reg_dataout_2535_port, 
      DataPath_RF_bus_reg_dataout_2536_port, 
      DataPath_RF_bus_reg_dataout_2537_port, 
      DataPath_RF_bus_reg_dataout_2538_port, 
      DataPath_RF_bus_reg_dataout_2539_port, 
      DataPath_RF_bus_reg_dataout_2540_port, 
      DataPath_RF_bus_reg_dataout_2541_port, 
      DataPath_RF_bus_reg_dataout_2542_port, 
      DataPath_RF_bus_reg_dataout_2543_port, 
      DataPath_RF_bus_reg_dataout_2544_port, 
      DataPath_RF_bus_reg_dataout_2545_port, 
      DataPath_RF_bus_reg_dataout_2546_port, 
      DataPath_RF_bus_reg_dataout_2547_port, 
      DataPath_RF_bus_reg_dataout_2548_port, 
      DataPath_RF_bus_reg_dataout_2549_port, 
      DataPath_RF_bus_reg_dataout_2550_port, 
      DataPath_RF_bus_reg_dataout_2551_port, 
      DataPath_RF_bus_reg_dataout_2552_port, 
      DataPath_RF_bus_reg_dataout_2553_port, 
      DataPath_RF_bus_reg_dataout_2554_port, 
      DataPath_RF_bus_reg_dataout_2555_port, 
      DataPath_RF_bus_reg_dataout_2556_port, 
      DataPath_RF_bus_reg_dataout_2557_port, 
      DataPath_RF_bus_reg_dataout_2558_port, 
      DataPath_RF_bus_reg_dataout_2559_port, DataPath_RF_next_cwp_0_port, 
      DataPath_RF_next_cwp_1_port, DataPath_RF_next_cwp_2_port, 
      DataPath_RF_next_cwp_3_port, DataPath_RF_next_cwp_4_port, 
      DataPath_RF_c_win_0_port, DataPath_RF_c_win_1_port, 
      DataPath_RF_c_win_2_port, DataPath_RF_c_win_3_port, 
      DataPath_RF_c_win_4_port, DataPath_WRF_CUhw_n187, DataPath_WRF_CUhw_n186,
      DataPath_WRF_CUhw_n185, DataPath_WRF_CUhw_n184, DataPath_WRF_CUhw_n183, 
      DataPath_WRF_CUhw_n182, DataPath_WRF_CUhw_n181, DataPath_WRF_CUhw_n180, 
      DataPath_WRF_CUhw_n179, DataPath_WRF_CUhw_n178, DataPath_WRF_CUhw_n177, 
      DataPath_WRF_CUhw_n176, DataPath_WRF_CUhw_n175, DataPath_WRF_CUhw_n174, 
      DataPath_WRF_CUhw_n173, DataPath_WRF_CUhw_n172, DataPath_WRF_CUhw_n171, 
      DataPath_WRF_CUhw_n170, DataPath_WRF_CUhw_n169, DataPath_WRF_CUhw_n168, 
      DataPath_WRF_CUhw_n167, DataPath_WRF_CUhw_n166, DataPath_WRF_CUhw_n165, 
      DataPath_WRF_CUhw_n164, DataPath_WRF_CUhw_n163, DataPath_WRF_CUhw_n162, 
      DataPath_WRF_CUhw_n161, DataPath_WRF_CUhw_n160, DataPath_WRF_CUhw_n159, 
      DataPath_WRF_CUhw_n158, DataPath_WRF_CUhw_n157, DataPath_WRF_CUhw_n156, 
      DataPath_WRF_CUhw_n155, DataPath_WRF_CUhw_n154, DataPath_WRF_CUhw_n153, 
      DataPath_WRF_CUhw_n152, DataPath_WRF_CUhw_n150, DataPath_WRF_CUhw_n149, 
      DataPath_WRF_CUhw_n148, DataPath_WRF_CUhw_n147, DataPath_WRF_CUhw_n146, 
      DataPath_WRF_CUhw_n145, DataPath_WRF_CUhw_n144, DataPath_WRF_CUhw_n143, 
      DataPath_WRF_CUhw_n142, DataPath_WRF_CUhw_n141, DataPath_WRF_CUhw_n140, 
      DataPath_WRF_CUhw_n139, DataPath_WRF_CUhw_n138, DataPath_WRF_CUhw_n137, 
      DataPath_WRF_CUhw_n136, DataPath_WRF_CUhw_n135, DataPath_WRF_CUhw_n134, 
      DataPath_WRF_CUhw_n133, DataPath_WRF_CUhw_n132, DataPath_WRF_CUhw_n131, 
      DataPath_WRF_CUhw_n130, DataPath_WRF_CUhw_n129, DataPath_WRF_CUhw_n128, 
      DataPath_WRF_CUhw_n127, DataPath_WRF_CUhw_n126, DataPath_WRF_CUhw_n125, 
      DataPath_WRF_CUhw_n124, DataPath_WRF_CUhw_n123, DataPath_WRF_CUhw_n122, 
      DataPath_WRF_CUhw_n121, DataPath_WRF_CUhw_n120, DataPath_WRF_CUhw_n119, 
      DataPath_WRF_CUhw_n118, DataPath_WRF_CUhw_n117, DataPath_WRF_CUhw_n116, 
      DataPath_WRF_CUhw_n115, DataPath_WRF_CUhw_n114, DataPath_WRF_CUhw_n113, 
      DataPath_WRF_CUhw_n112, DataPath_WRF_CUhw_n73, DataPath_WRF_CUhw_n38, 
      DataPath_WRF_CUhw_n37, DataPath_WRF_CUhw_n36, DataPath_WRF_CUhw_n35, 
      DataPath_WRF_CUhw_n34, DataPath_WRF_CUhw_n33, DataPath_WRF_CUhw_n32, 
      DataPath_WRF_CUhw_n31, DataPath_WRF_CUhw_n30, DataPath_WRF_CUhw_n29, 
      DataPath_WRF_CUhw_n28, DataPath_WRF_CUhw_n27, DataPath_WRF_CUhw_n26, 
      DataPath_WRF_CUhw_n25, DataPath_WRF_CUhw_n24, DataPath_WRF_CUhw_n23, 
      DataPath_WRF_CUhw_n22, DataPath_WRF_CUhw_n21, DataPath_WRF_CUhw_n20, 
      DataPath_WRF_CUhw_n19, DataPath_WRF_CUhw_n18, DataPath_WRF_CUhw_n17, 
      DataPath_WRF_CUhw_n16, DataPath_WRF_CUhw_n15, DataPath_WRF_CUhw_n14, 
      DataPath_WRF_CUhw_n13, DataPath_WRF_CUhw_n12, DataPath_WRF_CUhw_n11, 
      DataPath_WRF_CUhw_n10, DataPath_WRF_CUhw_n9, DataPath_WRF_CUhw_n8, 
      DataPath_WRF_CUhw_n7, DataPath_WRF_CUhw_N217, DataPath_WRF_CUhw_N177_port
      , DataPath_WRF_CUhw_N176_port, DataPath_WRF_CUhw_N175_port, 
      DataPath_WRF_CUhw_N174_port, DataPath_WRF_CUhw_N173_port, 
      DataPath_WRF_CUhw_N172_port, DataPath_WRF_CUhw_N171_port, 
      DataPath_WRF_CUhw_N170_port, DataPath_WRF_CUhw_N169_port, 
      DataPath_WRF_CUhw_N168_port, DataPath_WRF_CUhw_N167_port, 
      DataPath_WRF_CUhw_N166_port, DataPath_WRF_CUhw_N165_port, 
      DataPath_WRF_CUhw_N164_port, DataPath_WRF_CUhw_N163_port, 
      DataPath_WRF_CUhw_N162_port, DataPath_WRF_CUhw_N161_port, 
      DataPath_WRF_CUhw_N160_port, DataPath_WRF_CUhw_N159_port, 
      DataPath_WRF_CUhw_N158_port, DataPath_WRF_CUhw_N157_port, 
      DataPath_WRF_CUhw_N156_port, DataPath_WRF_CUhw_N155_port, 
      DataPath_WRF_CUhw_N154_port, DataPath_WRF_CUhw_N153_port, 
      DataPath_WRF_CUhw_N152_port, DataPath_WRF_CUhw_N151, 
      DataPath_WRF_CUhw_N150_port, DataPath_WRF_CUhw_N149_port, 
      DataPath_WRF_CUhw_N148_port, DataPath_WRF_CUhw_N147_port, 
      DataPath_WRF_CUhw_N146_port, DataPath_WRF_CUhw_N145_port, 
      DataPath_WRF_CUhw_N144_port, DataPath_WRF_CUhw_N140_port, 
      DataPath_WRF_CUhw_N139_port, DataPath_WRF_CUhw_N138_port, 
      DataPath_WRF_CUhw_N137_port, DataPath_WRF_CUhw_N136_port, 
      DataPath_WRF_CUhw_N135_port, DataPath_WRF_CUhw_N134_port, 
      DataPath_WRF_CUhw_N133_port, DataPath_WRF_CUhw_N132_port, 
      DataPath_WRF_CUhw_N131_port, DataPath_WRF_CUhw_N130_port, 
      DataPath_WRF_CUhw_N129_port, DataPath_WRF_CUhw_N128_port, 
      DataPath_WRF_CUhw_N127_port, DataPath_WRF_CUhw_N126_port, 
      DataPath_WRF_CUhw_N125_port, DataPath_WRF_CUhw_N124_port, 
      DataPath_WRF_CUhw_N123_port, DataPath_WRF_CUhw_N122_port, 
      DataPath_WRF_CUhw_N121_port, DataPath_WRF_CUhw_N120_port, 
      DataPath_WRF_CUhw_N119_port, DataPath_WRF_CUhw_N118_port, 
      DataPath_WRF_CUhw_N117_port, DataPath_WRF_CUhw_N116_port, 
      DataPath_WRF_CUhw_N115_port, DataPath_WRF_CUhw_N114_port, 
      DataPath_WRF_CUhw_N113_port, DataPath_WRF_CUhw_N112_port, 
      DataPath_WRF_CUhw_N111, DataPath_WRF_CUhw_N109, 
      DataPath_WRF_CUhw_N26_port, DataPath_WRF_CUhw_curr_addr_1_port, 
      DataPath_WRF_CUhw_curr_addr_2_port, DataPath_WRF_CUhw_curr_addr_3_port, 
      DataPath_WRF_CUhw_curr_addr_4_port, DataPath_WRF_CUhw_curr_addr_5_port, 
      DataPath_WRF_CUhw_curr_addr_6_port, DataPath_WRF_CUhw_curr_addr_7_port, 
      DataPath_WRF_CUhw_curr_addr_8_port, DataPath_WRF_CUhw_curr_addr_9_port, 
      DataPath_WRF_CUhw_curr_addr_10_port, DataPath_WRF_CUhw_curr_addr_11_port,
      DataPath_WRF_CUhw_curr_addr_12_port, DataPath_WRF_CUhw_curr_addr_13_port,
      DataPath_WRF_CUhw_curr_addr_14_port, DataPath_WRF_CUhw_curr_addr_15_port,
      DataPath_WRF_CUhw_curr_addr_16_port, DataPath_WRF_CUhw_curr_addr_17_port,
      DataPath_WRF_CUhw_curr_addr_18_port, DataPath_WRF_CUhw_curr_addr_19_port,
      DataPath_WRF_CUhw_curr_addr_20_port, DataPath_WRF_CUhw_curr_addr_21_port,
      DataPath_WRF_CUhw_curr_addr_22_port, DataPath_WRF_CUhw_curr_addr_23_port,
      DataPath_WRF_CUhw_curr_addr_24_port, DataPath_WRF_CUhw_curr_addr_25_port,
      DataPath_WRF_CUhw_curr_addr_26_port, DataPath_WRF_CUhw_curr_addr_27_port,
      DataPath_WRF_CUhw_curr_addr_28_port, DataPath_WRF_CUhw_curr_addr_29_port,
      DataPath_WRF_CUhw_curr_addr_30_port, DataPath_WRF_CUhw_curr_addr_31_port,
      DataPath_WRF_CUhw_curr_state_0_port, DataPath_WRF_CUhw_curr_state_1_port,
      DataPath_SETCMP_n9, DataPath_SETCMP_n8, DataPath_SETCMP_n7, 
      DataPath_SETCMP_n6, DataPath_SETCMP_n5, DataPath_SETCMP_n4, 
      DataPath_ALUhw_i_Q_EXTENDED_76_port, DataPath_ALUhw_i_Q_EXTENDED_78_port,
      DataPath_ALUhw_i_Q_EXTENDED_79_port, DataPath_ALUhw_i_Q_EXTENDED_80_port,
      DataPath_ALUhw_i_Q_EXTENDED_96_port, DataPath_ALUhw_i_Q_EXTENDED_97_port,
      DataPath_ALUhw_i_Q_EXTENDED_98_port, DataPath_ALUhw_i_Q_EXTENDED_99_port,
      DataPath_ALUhw_i_Q_EXTENDED_100_port, 
      DataPath_ALUhw_i_Q_EXTENDED_101_port, 
      DataPath_ALUhw_i_Q_EXTENDED_102_port, 
      DataPath_ALUhw_i_Q_EXTENDED_103_port, 
      DataPath_ALUhw_i_Q_EXTENDED_104_port, 
      DataPath_ALUhw_i_Q_EXTENDED_105_port, 
      DataPath_ALUhw_i_Q_EXTENDED_106_port, 
      DataPath_ALUhw_i_Q_EXTENDED_107_port, 
      DataPath_ALUhw_i_Q_EXTENDED_108_port, 
      DataPath_ALUhw_i_Q_EXTENDED_109_port, 
      DataPath_ALUhw_i_Q_EXTENDED_110_port, 
      DataPath_ALUhw_i_Q_EXTENDED_111_port, 
      DataPath_ALUhw_i_Q_EXTENDED_112_port, DataPath_MEM_ADDR_MASK_n2, 
      DataPath_LDSTR_n86, DataPath_LDSTR_n85, DataPath_LDSTR_n84, 
      DataPath_LDSTR_n83, DataPath_LDSTR_n82, DataPath_LDSTR_n81, 
      DataPath_LDSTR_n80, DataPath_LDSTR_n79, DataPath_LDSTR_n78, 
      DataPath_LDSTR_n77, DataPath_LDSTR_n76, DataPath_LDSTR_n75, 
      DataPath_LDSTR_n74, DataPath_LDSTR_n73, DataPath_LDSTR_n72, 
      DataPath_LDSTR_n71, DataPath_LDSTR_n70, DataPath_LDSTR_n69, 
      DataPath_LDSTR_n68, DataPath_LDSTR_n67, DataPath_LDSTR_n66, 
      DataPath_LDSTR_n65, DataPath_LDSTR_n64, DataPath_LDSTR_n63, 
      DataPath_LDSTR_n62, DataPath_LDSTR_n61, DataPath_LDSTR_n60, 
      DataPath_LDSTR_n59, DataPath_LDSTR_n58, DataPath_LDSTR_n57, 
      DataPath_LDSTR_n56, DataPath_LDSTR_n55, DataPath_LDSTR_n54, 
      DataPath_LDSTR_n53, DataPath_LDSTR_n52, DataPath_LDSTR_n51, 
      DataPath_LDSTR_n50, DataPath_LDSTR_n49, DataPath_LDSTR_n48, 
      DataPath_LDSTR_n47, DataPath_LDSTR_n46, DataPath_LDSTR_n45, 
      DataPath_LDSTR_n44, DataPath_LDSTR_n43, DataPath_LDSTR_n42, 
      DataPath_LDSTR_n41, DataPath_LDSTR_n40, DataPath_LDSTR_n39, 
      DataPath_LDSTR_n38, DataPath_LDSTR_n37, DataPath_RF_CWP_n13, 
      DataPath_RF_MUX_SELINPUT_8_n65, DataPath_RF_MUX_SELINPUT_8_n64, 
      DataPath_RF_MUX_SELINPUT_8_n63, DataPath_RF_MUX_SELINPUT_8_n62, 
      DataPath_RF_MUX_SELINPUT_8_n61, DataPath_RF_MUX_SELINPUT_8_n60, 
      DataPath_RF_MUX_SELINPUT_8_n59, DataPath_RF_MUX_SELINPUT_8_n58, 
      DataPath_RF_MUX_SELINPUT_8_n57, DataPath_RF_MUX_SELINPUT_8_n56, 
      DataPath_RF_MUX_SELINPUT_8_n55, DataPath_RF_MUX_SELINPUT_8_n54, 
      DataPath_RF_MUX_SELINPUT_8_n53, DataPath_RF_MUX_SELINPUT_8_n52, 
      DataPath_RF_MUX_SELINPUT_8_n51, DataPath_RF_MUX_SELINPUT_8_n50, 
      DataPath_RF_MUX_SELINPUT_8_n49, DataPath_RF_MUX_SELINPUT_8_n48, 
      DataPath_RF_MUX_SELINPUT_8_n47, DataPath_RF_MUX_SELINPUT_8_n46, 
      DataPath_RF_MUX_SELINPUT_8_n45, DataPath_RF_MUX_SELINPUT_8_n44, 
      DataPath_RF_MUX_SELINPUT_8_n43, DataPath_RF_MUX_SELINPUT_8_n42, 
      DataPath_RF_MUX_SELINPUT_8_n41, DataPath_RF_MUX_SELINPUT_8_n40, 
      DataPath_RF_MUX_SELINPUT_8_n39, DataPath_RF_MUX_SELINPUT_8_n38, 
      DataPath_RF_MUX_SELINPUT_8_n37, DataPath_RF_MUX_SELINPUT_8_n36, 
      DataPath_RF_MUX_SELINPUT_8_n35, DataPath_RF_MUX_SELINPUT_8_n34, 
      DataPath_RF_DEC_n17, DataPath_RF_DEC_n16, DataPath_RF_DEC_n15, 
      DataPath_RF_DEC_n14, DataPath_RF_DEC_n13, DataPath_RF_DEC_n12, 
      DataPath_RF_DEC_n11, DataPath_RF_DEC_n10, DataPath_RF_DEC_n9, 
      DataPath_RF_DEC_n8, DataPath_RF_DEC_n7, DataPath_RF_SELBLOCK_INLOC_n1032,
      DataPath_RF_SELBLOCK_INLOC_n1031, DataPath_RF_SELBLOCK_INLOC_n1030, 
      DataPath_RF_SELBLOCK_INLOC_n1029, DataPath_RF_SELBLOCK_INLOC_n1028, 
      DataPath_RF_SELBLOCK_INLOC_n1027, DataPath_RF_SELBLOCK_INLOC_n1026, 
      DataPath_RF_SELBLOCK_INLOC_n1025, DataPath_RF_SELBLOCK_INLOC_n1024, 
      DataPath_RF_SELBLOCK_INLOC_n1023, DataPath_RF_SELBLOCK_INLOC_n1022, 
      DataPath_RF_SELBLOCK_INLOC_n1021, DataPath_RF_SELBLOCK_INLOC_n1020, 
      DataPath_RF_SELBLOCK_INLOC_n1019, DataPath_RF_SELBLOCK_INLOC_n1018, 
      DataPath_RF_SELBLOCK_INLOC_n1017, DataPath_RF_SELBLOCK_INLOC_n1016, 
      DataPath_RF_SELBLOCK_INLOC_n1015, DataPath_RF_SELBLOCK_INLOC_n1014, 
      DataPath_RF_SELBLOCK_INLOC_n1013, DataPath_RF_SELBLOCK_INLOC_n1012, 
      DataPath_RF_SELBLOCK_INLOC_n1011, DataPath_RF_SELBLOCK_INLOC_n1010, 
      DataPath_RF_SELBLOCK_INLOC_n1009, DataPath_RF_SELBLOCK_INLOC_n1008, 
      DataPath_RF_SELBLOCK_INLOC_n1007, DataPath_RF_SELBLOCK_INLOC_n1006, 
      DataPath_RF_SELBLOCK_INLOC_n1005, DataPath_RF_SELBLOCK_INLOC_n1004, 
      DataPath_RF_SELBLOCK_INLOC_n1003, DataPath_RF_SELBLOCK_INLOC_n1002, 
      DataPath_RF_SELBLOCK_INLOC_n1001, DataPath_RF_SELBLOCK_INLOC_n1000, 
      DataPath_RF_SELBLOCK_INLOC_n999, DataPath_RF_SELBLOCK_INLOC_n998, 
      DataPath_RF_SELBLOCK_INLOC_n997, DataPath_RF_SELBLOCK_INLOC_n996, 
      DataPath_RF_SELBLOCK_INLOC_n995, DataPath_RF_SELBLOCK_INLOC_n994, 
      DataPath_RF_SELBLOCK_INLOC_n993, DataPath_RF_SELBLOCK_INLOC_n992, 
      DataPath_RF_SELBLOCK_INLOC_n991, DataPath_RF_SELBLOCK_INLOC_n990, 
      DataPath_RF_SELBLOCK_INLOC_n989, DataPath_RF_SELBLOCK_INLOC_n988, 
      DataPath_RF_SELBLOCK_INLOC_n987, DataPath_RF_SELBLOCK_INLOC_n986, 
      DataPath_RF_SELBLOCK_INLOC_n985, DataPath_RF_SELBLOCK_INLOC_n984, 
      DataPath_RF_SELBLOCK_INLOC_n983, DataPath_RF_SELBLOCK_INLOC_n982, 
      DataPath_RF_SELBLOCK_INLOC_n981, DataPath_RF_SELBLOCK_INLOC_n980, 
      DataPath_RF_SELBLOCK_INLOC_n979, DataPath_RF_SELBLOCK_INLOC_n978, 
      DataPath_RF_SELBLOCK_INLOC_n977, DataPath_RF_SELBLOCK_INLOC_n976, 
      DataPath_RF_SELBLOCK_INLOC_n975, DataPath_RF_SELBLOCK_INLOC_n974, 
      DataPath_RF_SELBLOCK_INLOC_n973, DataPath_RF_SELBLOCK_INLOC_n972, 
      DataPath_RF_SELBLOCK_INLOC_n971, DataPath_RF_SELBLOCK_INLOC_n970, 
      DataPath_RF_SELBLOCK_INLOC_n969, DataPath_RF_SELBLOCK_INLOC_n968, 
      DataPath_RF_SELBLOCK_INLOC_n967, DataPath_RF_SELBLOCK_INLOC_n966, 
      DataPath_RF_SELBLOCK_INLOC_n965, DataPath_RF_SELBLOCK_INLOC_n964, 
      DataPath_RF_SELBLOCK_INLOC_n963, DataPath_RF_SELBLOCK_INLOC_n962, 
      DataPath_RF_SELBLOCK_INLOC_n961, DataPath_RF_SELBLOCK_INLOC_n960, 
      DataPath_RF_SELBLOCK_INLOC_n959, DataPath_RF_SELBLOCK_INLOC_n958, 
      DataPath_RF_SELBLOCK_INLOC_n957, DataPath_RF_SELBLOCK_INLOC_n956, 
      DataPath_RF_SELBLOCK_INLOC_n955, DataPath_RF_SELBLOCK_INLOC_n954, 
      DataPath_RF_SELBLOCK_INLOC_n953, DataPath_RF_SELBLOCK_INLOC_n952, 
      DataPath_RF_SELBLOCK_INLOC_n951, DataPath_RF_SELBLOCK_INLOC_n950, 
      DataPath_RF_SELBLOCK_INLOC_n949, DataPath_RF_SELBLOCK_INLOC_n948, 
      DataPath_RF_SELBLOCK_INLOC_n947, DataPath_RF_SELBLOCK_INLOC_n946, 
      DataPath_RF_SELBLOCK_INLOC_n945, DataPath_RF_SELBLOCK_INLOC_n944, 
      DataPath_RF_SELBLOCK_INLOC_n943, DataPath_RF_SELBLOCK_INLOC_n942, 
      DataPath_RF_SELBLOCK_INLOC_n941, DataPath_RF_SELBLOCK_INLOC_n940, 
      DataPath_RF_SELBLOCK_INLOC_n939, DataPath_RF_SELBLOCK_INLOC_n938, 
      DataPath_RF_SELBLOCK_INLOC_n937, DataPath_RF_SELBLOCK_INLOC_n936, 
      DataPath_RF_SELBLOCK_INLOC_n935, DataPath_RF_SELBLOCK_INLOC_n934, 
      DataPath_RF_SELBLOCK_INLOC_n933, DataPath_RF_SELBLOCK_INLOC_n932, 
      DataPath_RF_SELBLOCK_INLOC_n931, DataPath_RF_SELBLOCK_INLOC_n930, 
      DataPath_RF_SELBLOCK_INLOC_n929, DataPath_RF_SELBLOCK_INLOC_n928, 
      DataPath_RF_SELBLOCK_INLOC_n927, DataPath_RF_SELBLOCK_INLOC_n926, 
      DataPath_RF_SELBLOCK_INLOC_n925, DataPath_RF_SELBLOCK_INLOC_n924, 
      DataPath_RF_SELBLOCK_INLOC_n923, DataPath_RF_SELBLOCK_INLOC_n922, 
      DataPath_RF_SELBLOCK_INLOC_n921, DataPath_RF_SELBLOCK_INLOC_n920, 
      DataPath_RF_SELBLOCK_INLOC_n919, DataPath_RF_SELBLOCK_INLOC_n918, 
      DataPath_RF_SELBLOCK_INLOC_n917, DataPath_RF_SELBLOCK_INLOC_n916, 
      DataPath_RF_SELBLOCK_INLOC_n915, DataPath_RF_SELBLOCK_INLOC_n914, 
      DataPath_RF_SELBLOCK_INLOC_n913, DataPath_RF_SELBLOCK_INLOC_n912, 
      DataPath_RF_SELBLOCK_INLOC_n911, DataPath_RF_SELBLOCK_INLOC_n910, 
      DataPath_RF_SELBLOCK_INLOC_n909, DataPath_RF_SELBLOCK_INLOC_n908, 
      DataPath_RF_SELBLOCK_INLOC_n907, DataPath_RF_SELBLOCK_INLOC_n906, 
      DataPath_RF_SELBLOCK_INLOC_n905, DataPath_RF_SELBLOCK_INLOC_n904, 
      DataPath_RF_SELBLOCK_INLOC_n903, DataPath_RF_SELBLOCK_INLOC_n902, 
      DataPath_RF_SELBLOCK_INLOC_n901, DataPath_RF_SELBLOCK_INLOC_n900, 
      DataPath_RF_SELBLOCK_INLOC_n899, DataPath_RF_SELBLOCK_INLOC_n898, 
      DataPath_RF_SELBLOCK_INLOC_n897, DataPath_RF_SELBLOCK_INLOC_n896, 
      DataPath_RF_SELBLOCK_INLOC_n895, DataPath_RF_SELBLOCK_INLOC_n894, 
      DataPath_RF_SELBLOCK_INLOC_n893, DataPath_RF_SELBLOCK_INLOC_n892, 
      DataPath_RF_SELBLOCK_INLOC_n891, DataPath_RF_SELBLOCK_INLOC_n890, 
      DataPath_RF_SELBLOCK_INLOC_n889, DataPath_RF_SELBLOCK_INLOC_n888, 
      DataPath_RF_SELBLOCK_INLOC_n887, DataPath_RF_SELBLOCK_INLOC_n886, 
      DataPath_RF_SELBLOCK_INLOC_n885, DataPath_RF_SELBLOCK_INLOC_n884, 
      DataPath_RF_SELBLOCK_INLOC_n883, DataPath_RF_SELBLOCK_INLOC_n882, 
      DataPath_RF_SELBLOCK_INLOC_n881, DataPath_RF_SELBLOCK_INLOC_n880, 
      DataPath_RF_SELBLOCK_INLOC_n879, DataPath_RF_SELBLOCK_INLOC_n878, 
      DataPath_RF_SELBLOCK_INLOC_n877, DataPath_RF_SELBLOCK_INLOC_n876, 
      DataPath_RF_SELBLOCK_INLOC_n875, DataPath_RF_SELBLOCK_INLOC_n874, 
      DataPath_RF_SELBLOCK_INLOC_n873, DataPath_RF_SELBLOCK_INLOC_n872, 
      DataPath_RF_SELBLOCK_INLOC_n871, DataPath_RF_SELBLOCK_INLOC_n870, 
      DataPath_RF_SELBLOCK_INLOC_n869, DataPath_RF_SELBLOCK_INLOC_n868, 
      DataPath_RF_SELBLOCK_INLOC_n867, DataPath_RF_SELBLOCK_INLOC_n866, 
      DataPath_RF_SELBLOCK_INLOC_n865, DataPath_RF_SELBLOCK_INLOC_n864, 
      DataPath_RF_SELBLOCK_INLOC_n863, DataPath_RF_SELBLOCK_INLOC_n862, 
      DataPath_RF_SELBLOCK_INLOC_n861, DataPath_RF_SELBLOCK_INLOC_n860, 
      DataPath_RF_SELBLOCK_INLOC_n859, DataPath_RF_SELBLOCK_INLOC_n858, 
      DataPath_RF_SELBLOCK_INLOC_n857, DataPath_RF_SELBLOCK_INLOC_n856, 
      DataPath_RF_SELBLOCK_INLOC_n855, DataPath_RF_SELBLOCK_INLOC_n854, 
      DataPath_RF_SELBLOCK_INLOC_n853, DataPath_RF_SELBLOCK_INLOC_n852, 
      DataPath_RF_SELBLOCK_INLOC_n851, DataPath_RF_SELBLOCK_INLOC_n850, 
      DataPath_RF_SELBLOCK_INLOC_n849, DataPath_RF_SELBLOCK_INLOC_n848, 
      DataPath_RF_SELBLOCK_INLOC_n847, DataPath_RF_SELBLOCK_INLOC_n846, 
      DataPath_RF_SELBLOCK_INLOC_n845, DataPath_RF_SELBLOCK_INLOC_n844, 
      DataPath_RF_SELBLOCK_INLOC_n843, DataPath_RF_SELBLOCK_INLOC_n842, 
      DataPath_RF_SELBLOCK_INLOC_n841, DataPath_RF_SELBLOCK_INLOC_n840, 
      DataPath_RF_SELBLOCK_INLOC_n839, DataPath_RF_SELBLOCK_INLOC_n838, 
      DataPath_RF_SELBLOCK_INLOC_n837, DataPath_RF_SELBLOCK_INLOC_n836, 
      DataPath_RF_SELBLOCK_INLOC_n835, DataPath_RF_SELBLOCK_INLOC_n834, 
      DataPath_RF_SELBLOCK_INLOC_n833, DataPath_RF_SELBLOCK_INLOC_n832, 
      DataPath_RF_SELBLOCK_INLOC_n831, DataPath_RF_SELBLOCK_INLOC_n830, 
      DataPath_RF_SELBLOCK_INLOC_n829, DataPath_RF_SELBLOCK_INLOC_n828, 
      DataPath_RF_SELBLOCK_INLOC_n827, DataPath_RF_SELBLOCK_INLOC_n826, 
      DataPath_RF_SELBLOCK_INLOC_n825, DataPath_RF_SELBLOCK_INLOC_n824, 
      DataPath_RF_SELBLOCK_INLOC_n823, DataPath_RF_SELBLOCK_INLOC_n822, 
      DataPath_RF_SELBLOCK_INLOC_n821, DataPath_RF_SELBLOCK_INLOC_n820, 
      DataPath_RF_SELBLOCK_INLOC_n819, DataPath_RF_SELBLOCK_INLOC_n818, 
      DataPath_RF_SELBLOCK_INLOC_n817, DataPath_RF_SELBLOCK_INLOC_n816, 
      DataPath_RF_SELBLOCK_INLOC_n815, DataPath_RF_SELBLOCK_INLOC_n814, 
      DataPath_RF_SELBLOCK_INLOC_n813, DataPath_RF_SELBLOCK_INLOC_n812, 
      DataPath_RF_SELBLOCK_INLOC_n811, DataPath_RF_SELBLOCK_INLOC_n810, 
      DataPath_RF_SELBLOCK_INLOC_n809, DataPath_RF_SELBLOCK_INLOC_n808, 
      DataPath_RF_SELBLOCK_INLOC_n807, DataPath_RF_SELBLOCK_INLOC_n806, 
      DataPath_RF_SELBLOCK_INLOC_n805, DataPath_RF_SELBLOCK_INLOC_n804, 
      DataPath_RF_SELBLOCK_INLOC_n803, DataPath_RF_SELBLOCK_INLOC_n802, 
      DataPath_RF_SELBLOCK_INLOC_n801, DataPath_RF_SELBLOCK_INLOC_n800, 
      DataPath_RF_SELBLOCK_INLOC_n799, DataPath_RF_SELBLOCK_INLOC_n798, 
      DataPath_RF_SELBLOCK_INLOC_n797, DataPath_RF_SELBLOCK_INLOC_n796, 
      DataPath_RF_SELBLOCK_INLOC_n795, DataPath_RF_SELBLOCK_INLOC_n794, 
      DataPath_RF_SELBLOCK_INLOC_n793, DataPath_RF_SELBLOCK_INLOC_n792, 
      DataPath_RF_SELBLOCK_INLOC_n791, DataPath_RF_SELBLOCK_INLOC_n790, 
      DataPath_RF_SELBLOCK_INLOC_n789, DataPath_RF_SELBLOCK_INLOC_n788, 
      DataPath_RF_SELBLOCK_INLOC_n787, DataPath_RF_SELBLOCK_INLOC_n786, 
      DataPath_RF_SELBLOCK_INLOC_n785, DataPath_RF_SELBLOCK_INLOC_n784, 
      DataPath_RF_SELBLOCK_INLOC_n783, DataPath_RF_SELBLOCK_INLOC_n782, 
      DataPath_RF_SELBLOCK_INLOC_n781, DataPath_RF_SELBLOCK_INLOC_n780, 
      DataPath_RF_SELBLOCK_INLOC_n779, DataPath_RF_SELBLOCK_INLOC_n778, 
      DataPath_RF_SELBLOCK_INLOC_n777, DataPath_RF_SELBLOCK_INLOC_n776, 
      DataPath_RF_SELBLOCK_INLOC_n775, DataPath_RF_SELBLOCK_INLOC_n774, 
      DataPath_RF_SELBLOCK_INLOC_n773, DataPath_RF_SELBLOCK_INLOC_n772, 
      DataPath_RF_SELBLOCK_INLOC_n771, DataPath_RF_SELBLOCK_INLOC_n770, 
      DataPath_RF_SELBLOCK_INLOC_n769, DataPath_RF_SELBLOCK_INLOC_n768, 
      DataPath_RF_SELBLOCK_INLOC_n767, DataPath_RF_SELBLOCK_INLOC_n766, 
      DataPath_RF_SELBLOCK_INLOC_n765, DataPath_RF_SELBLOCK_INLOC_n764, 
      DataPath_RF_SELBLOCK_INLOC_n763, DataPath_RF_SELBLOCK_INLOC_n762, 
      DataPath_RF_SELBLOCK_INLOC_n761, DataPath_RF_SELBLOCK_INLOC_n760, 
      DataPath_RF_SELBLOCK_INLOC_n759, DataPath_RF_SELBLOCK_INLOC_n758, 
      DataPath_RF_SELBLOCK_INLOC_n757, DataPath_RF_SELBLOCK_INLOC_n756, 
      DataPath_RF_SELBLOCK_INLOC_n755, DataPath_RF_SELBLOCK_INLOC_n754, 
      DataPath_RF_SELBLOCK_INLOC_n753, DataPath_RF_SELBLOCK_INLOC_n752, 
      DataPath_RF_SELBLOCK_INLOC_n751, DataPath_RF_SELBLOCK_INLOC_n750, 
      DataPath_RF_SELBLOCK_INLOC_n749, DataPath_RF_SELBLOCK_INLOC_n748, 
      DataPath_RF_SELBLOCK_INLOC_n747, DataPath_RF_SELBLOCK_INLOC_n746, 
      DataPath_RF_SELBLOCK_INLOC_n745, DataPath_RF_SELBLOCK_INLOC_n744, 
      DataPath_RF_SELBLOCK_INLOC_n743, DataPath_RF_SELBLOCK_INLOC_n742, 
      DataPath_RF_SELBLOCK_INLOC_n741, DataPath_RF_SELBLOCK_INLOC_n740, 
      DataPath_RF_SELBLOCK_INLOC_n739, DataPath_RF_SELBLOCK_INLOC_n738, 
      DataPath_RF_SELBLOCK_INLOC_n737, DataPath_RF_SELBLOCK_INLOC_n736, 
      DataPath_RF_SELBLOCK_INLOC_n735, DataPath_RF_SELBLOCK_INLOC_n734, 
      DataPath_RF_SELBLOCK_INLOC_n733, DataPath_RF_SELBLOCK_INLOC_n732, 
      DataPath_RF_SELBLOCK_INLOC_n731, DataPath_RF_SELBLOCK_INLOC_n730, 
      DataPath_RF_SELBLOCK_INLOC_n729, DataPath_RF_SELBLOCK_INLOC_n728, 
      DataPath_RF_SELBLOCK_INLOC_n727, DataPath_RF_SELBLOCK_INLOC_n726, 
      DataPath_RF_SELBLOCK_INLOC_n725, DataPath_RF_SELBLOCK_INLOC_n724, 
      DataPath_RF_SELBLOCK_INLOC_n723, DataPath_RF_SELBLOCK_INLOC_n722, 
      DataPath_RF_SELBLOCK_INLOC_n721, DataPath_RF_SELBLOCK_INLOC_n720, 
      DataPath_RF_SELBLOCK_INLOC_n719, DataPath_RF_SELBLOCK_INLOC_n718, 
      DataPath_RF_SELBLOCK_INLOC_n717, DataPath_RF_SELBLOCK_INLOC_n716, 
      DataPath_RF_SELBLOCK_INLOC_n715, DataPath_RF_SELBLOCK_INLOC_n714, 
      DataPath_RF_SELBLOCK_INLOC_n713, DataPath_RF_SELBLOCK_INLOC_n712, 
      DataPath_RF_SELBLOCK_INLOC_n711, DataPath_RF_SELBLOCK_INLOC_n710, 
      DataPath_RF_SELBLOCK_INLOC_n709, DataPath_RF_SELBLOCK_INLOC_n708, 
      DataPath_RF_SELBLOCK_INLOC_n707, DataPath_RF_SELBLOCK_INLOC_n706, 
      DataPath_RF_SELBLOCK_INLOC_n705, DataPath_RF_SELBLOCK_INLOC_n704, 
      DataPath_RF_SELBLOCK_INLOC_n703, DataPath_RF_SELBLOCK_INLOC_n702, 
      DataPath_RF_SELBLOCK_INLOC_n701, DataPath_RF_SELBLOCK_INLOC_n700, 
      DataPath_RF_SELBLOCK_INLOC_n699, DataPath_RF_SELBLOCK_INLOC_n698, 
      DataPath_RF_SELBLOCK_INLOC_n697, DataPath_RF_SELBLOCK_INLOC_n696, 
      DataPath_RF_SELBLOCK_INLOC_n695, DataPath_RF_SELBLOCK_INLOC_n694, 
      DataPath_RF_SELBLOCK_INLOC_n693, DataPath_RF_SELBLOCK_INLOC_n692, 
      DataPath_RF_SELBLOCK_INLOC_n691, DataPath_RF_SELBLOCK_INLOC_n690, 
      DataPath_RF_SELBLOCK_INLOC_n689, DataPath_RF_SELBLOCK_INLOC_n688, 
      DataPath_RF_SELBLOCK_INLOC_n687, DataPath_RF_SELBLOCK_INLOC_n686, 
      DataPath_RF_SELBLOCK_INLOC_n685, DataPath_RF_SELBLOCK_INLOC_n684, 
      DataPath_RF_SELBLOCK_INLOC_n683, DataPath_RF_SELBLOCK_INLOC_n682, 
      DataPath_RF_SELBLOCK_INLOC_n681, DataPath_RF_SELBLOCK_INLOC_n680, 
      DataPath_RF_SELBLOCK_INLOC_n679, DataPath_RF_SELBLOCK_INLOC_n678, 
      DataPath_RF_SELBLOCK_INLOC_n677, DataPath_RF_SELBLOCK_INLOC_n676, 
      DataPath_RF_SELBLOCK_INLOC_n675, DataPath_RF_SELBLOCK_INLOC_n674, 
      DataPath_RF_SELBLOCK_INLOC_n673, DataPath_RF_SELBLOCK_INLOC_n672, 
      DataPath_RF_SELBLOCK_INLOC_n671, DataPath_RF_SELBLOCK_INLOC_n670, 
      DataPath_RF_SELBLOCK_INLOC_n669, DataPath_RF_SELBLOCK_INLOC_n668, 
      DataPath_RF_SELBLOCK_INLOC_n667, DataPath_RF_SELBLOCK_INLOC_n666, 
      DataPath_RF_SELBLOCK_INLOC_n665, DataPath_RF_SELBLOCK_INLOC_n664, 
      DataPath_RF_SELBLOCK_INLOC_n663, DataPath_RF_SELBLOCK_INLOC_n662, 
      DataPath_RF_SELBLOCK_INLOC_n661, DataPath_RF_SELBLOCK_INLOC_n660, 
      DataPath_RF_SELBLOCK_INLOC_n659, DataPath_RF_SELBLOCK_INLOC_n658, 
      DataPath_RF_SELBLOCK_INLOC_n657, DataPath_RF_SELBLOCK_INLOC_n656, 
      DataPath_RF_SELBLOCK_INLOC_n655, DataPath_RF_SELBLOCK_INLOC_n654, 
      DataPath_RF_SELBLOCK_INLOC_n653, DataPath_RF_SELBLOCK_INLOC_n652, 
      DataPath_RF_SELBLOCK_INLOC_n651, DataPath_RF_SELBLOCK_INLOC_n650, 
      DataPath_RF_SELBLOCK_INLOC_n649, DataPath_RF_SELBLOCK_INLOC_n648, 
      DataPath_RF_SELBLOCK_INLOC_n647, DataPath_RF_SELBLOCK_INLOC_n646, 
      DataPath_RF_SELBLOCK_INLOC_n645, DataPath_RF_SELBLOCK_INLOC_n644, 
      DataPath_RF_SELBLOCK_INLOC_n643, DataPath_RF_SELBLOCK_INLOC_n642, 
      DataPath_RF_SELBLOCK_INLOC_n641, DataPath_RF_SELBLOCK_INLOC_n640, 
      DataPath_RF_SELBLOCK_INLOC_n639, DataPath_RF_SELBLOCK_INLOC_n638, 
      DataPath_RF_SELBLOCK_INLOC_n637, DataPath_RF_SELBLOCK_INLOC_n636, 
      DataPath_RF_SELBLOCK_INLOC_n635, DataPath_RF_SELBLOCK_INLOC_n634, 
      DataPath_RF_SELBLOCK_INLOC_n633, DataPath_RF_SELBLOCK_INLOC_n632, 
      DataPath_RF_SELBLOCK_INLOC_n631, DataPath_RF_SELBLOCK_INLOC_n630, 
      DataPath_RF_SELBLOCK_INLOC_n629, DataPath_RF_SELBLOCK_INLOC_n628, 
      DataPath_RF_SELBLOCK_INLOC_n627, DataPath_RF_SELBLOCK_INLOC_n626, 
      DataPath_RF_SELBLOCK_INLOC_n625, DataPath_RF_SELBLOCK_INLOC_n624, 
      DataPath_RF_SELBLOCK_INLOC_n623, DataPath_RF_SELBLOCK_INLOC_n622, 
      DataPath_RF_SELBLOCK_INLOC_n621, DataPath_RF_SELBLOCK_INLOC_n620, 
      DataPath_RF_SELBLOCK_INLOC_n619, DataPath_RF_SELBLOCK_INLOC_n618, 
      DataPath_RF_SELBLOCK_INLOC_n617, DataPath_RF_SELBLOCK_INLOC_n616, 
      DataPath_RF_SELBLOCK_INLOC_n615, DataPath_RF_SELBLOCK_INLOC_n614, 
      DataPath_RF_SELBLOCK_INLOC_n613, DataPath_RF_SELBLOCK_INLOC_n612, 
      DataPath_RF_SELBLOCK_INLOC_n611, DataPath_RF_SELBLOCK_INLOC_n610, 
      DataPath_RF_SELBLOCK_INLOC_n609, DataPath_RF_SELBLOCK_INLOC_n608, 
      DataPath_RF_SELBLOCK_INLOC_n607, DataPath_RF_SELBLOCK_INLOC_n606, 
      DataPath_RF_SELBLOCK_INLOC_n605, DataPath_RF_SELBLOCK_INLOC_n604, 
      DataPath_RF_SELBLOCK_INLOC_n603, DataPath_RF_SELBLOCK_INLOC_n602, 
      DataPath_RF_SELBLOCK_INLOC_n601, DataPath_RF_SELBLOCK_INLOC_n600, 
      DataPath_RF_SELBLOCK_INLOC_n599, DataPath_RF_SELBLOCK_INLOC_n598, 
      DataPath_RF_SELBLOCK_INLOC_n597, DataPath_RF_SELBLOCK_INLOC_n596, 
      DataPath_RF_SELBLOCK_INLOC_n595, DataPath_RF_SELBLOCK_INLOC_n594, 
      DataPath_RF_SELBLOCK_INLOC_n593, DataPath_RF_SELBLOCK_INLOC_n592, 
      DataPath_RF_SELBLOCK_INLOC_n591, DataPath_RF_SELBLOCK_INLOC_n590, 
      DataPath_RF_SELBLOCK_INLOC_n589, DataPath_RF_SELBLOCK_INLOC_n588, 
      DataPath_RF_SELBLOCK_INLOC_n587, DataPath_RF_SELBLOCK_INLOC_n586, 
      DataPath_RF_SELBLOCK_INLOC_n585, DataPath_RF_SELBLOCK_INLOC_n584, 
      DataPath_RF_SELBLOCK_INLOC_n583, DataPath_RF_SELBLOCK_INLOC_n582, 
      DataPath_RF_SELBLOCK_INLOC_n581, DataPath_RF_SELBLOCK_INLOC_n580, 
      DataPath_RF_SELBLOCK_INLOC_n579, DataPath_RF_SELBLOCK_INLOC_n578, 
      DataPath_RF_SELBLOCK_INLOC_n577, DataPath_RF_SELBLOCK_INLOC_n576, 
      DataPath_RF_SELBLOCK_INLOC_n575, DataPath_RF_SELBLOCK_INLOC_n574, 
      DataPath_RF_SELBLOCK_INLOC_n573, DataPath_RF_SELBLOCK_INLOC_n572, 
      DataPath_RF_SELBLOCK_INLOC_n571, DataPath_RF_SELBLOCK_INLOC_n570, 
      DataPath_RF_SELBLOCK_INLOC_n569, DataPath_RF_SELBLOCK_INLOC_n568, 
      DataPath_RF_SELBLOCK_INLOC_n567, DataPath_RF_SELBLOCK_INLOC_n566, 
      DataPath_RF_SELBLOCK_INLOC_n565, DataPath_RF_SELBLOCK_INLOC_n564, 
      DataPath_RF_SELBLOCK_INLOC_n563, DataPath_RF_SELBLOCK_INLOC_n562, 
      DataPath_RF_SELBLOCK_INLOC_n561, DataPath_RF_SELBLOCK_INLOC_n560, 
      DataPath_RF_SELBLOCK_INLOC_n559, DataPath_RF_SELBLOCK_INLOC_n558, 
      DataPath_RF_SELBLOCK_INLOC_n557, DataPath_RF_SELBLOCK_INLOC_n556, 
      DataPath_RF_SELBLOCK_INLOC_n555, DataPath_RF_SELBLOCK_INLOC_n554, 
      DataPath_RF_SELBLOCK_INLOC_n553, DataPath_RF_SELBLOCK_INLOC_n552, 
      DataPath_RF_SELBLOCK_INLOC_n551, DataPath_RF_SELBLOCK_INLOC_n550, 
      DataPath_RF_SELBLOCK_INLOC_n549, DataPath_RF_SELBLOCK_INLOC_n548, 
      DataPath_RF_SELBLOCK_INLOC_n547, DataPath_RF_SELBLOCK_INLOC_n546, 
      DataPath_RF_SELBLOCK_INLOC_n545, DataPath_RF_SELBLOCK_INLOC_n544, 
      DataPath_RF_SELBLOCK_INLOC_n543, DataPath_RF_SELBLOCK_INLOC_n542, 
      DataPath_RF_SELBLOCK_INLOC_n541, DataPath_RF_SELBLOCK_INLOC_n540, 
      DataPath_RF_SELBLOCK_INLOC_n539, DataPath_RF_SELBLOCK_INLOC_n538, 
      DataPath_RF_SELBLOCK_INLOC_n537, DataPath_RF_SELBLOCK_INLOC_n536, 
      DataPath_RF_SELBLOCK_INLOC_n535, DataPath_RF_SELBLOCK_INLOC_n534, 
      DataPath_RF_SELBLOCK_INLOC_n533, DataPath_RF_SELBLOCK_INLOC_n532, 
      DataPath_RF_SELBLOCK_INLOC_n531, DataPath_RF_SELBLOCK_INLOC_n530, 
      DataPath_RF_SELBLOCK_INLOC_n529, DataPath_RF_SELBLOCK_INLOC_n528, 
      DataPath_RF_SELBLOCK_INLOC_n527, DataPath_RF_SELBLOCK_INLOC_n526, 
      DataPath_RF_SELBLOCK_INLOC_n525, DataPath_RF_SELBLOCK_INLOC_n524, 
      DataPath_RF_SELBLOCK_INLOC_n523, DataPath_RF_SELBLOCK_INLOC_n522, 
      DataPath_RF_SELBLOCK_INLOC_n521, DataPath_RF_SELBLOCK_INLOC_n520, 
      DataPath_RF_SELBLOCK_INLOC_n519, DataPath_RF_SELBLOCK_INLOC_n518, 
      DataPath_RF_SELBLOCK_INLOC_n517, DataPath_RF_SELBLOCK_INLOC_n516, 
      DataPath_RF_SELBLOCK_INLOC_n515, DataPath_RF_SELBLOCK_INLOC_n514, 
      DataPath_RF_SELBLOCK_INLOC_n513, DataPath_RF_SELBLOCK_INLOC_n512, 
      DataPath_RF_SELBLOCK_INLOC_n511, DataPath_RF_SELBLOCK_INLOC_n510, 
      DataPath_RF_SELBLOCK_INLOC_n509, DataPath_RF_SELBLOCK_INLOC_n508, 
      DataPath_RF_SELBLOCK_INLOC_n507, DataPath_RF_SELBLOCK_INLOC_n506, 
      DataPath_RF_SELBLOCK_INLOC_n505, DataPath_RF_SELBLOCK_INLOC_n504, 
      DataPath_RF_SELBLOCK_INLOC_n503, DataPath_RF_SELBLOCK_INLOC_n502, 
      DataPath_RF_SELBLOCK_INLOC_n501, DataPath_RF_SELBLOCK_INLOC_n500, 
      DataPath_RF_SELBLOCK_INLOC_n499, DataPath_RF_SELBLOCK_INLOC_n498, 
      DataPath_RF_SELBLOCK_INLOC_n497, DataPath_RF_SELBLOCK_INLOC_n496, 
      DataPath_RF_SELBLOCK_INLOC_n495, DataPath_RF_SELBLOCK_INLOC_n494, 
      DataPath_RF_SELBLOCK_INLOC_n493, DataPath_RF_SELBLOCK_INLOC_n492, 
      DataPath_RF_SELBLOCK_INLOC_n491, DataPath_RF_SELBLOCK_INLOC_n490, 
      DataPath_RF_SELBLOCK_INLOC_n489, DataPath_RF_SELBLOCK_INLOC_n488, 
      DataPath_RF_SELBLOCK_INLOC_n487, DataPath_RF_SELBLOCK_INLOC_n486, 
      DataPath_RF_SELBLOCK_INLOC_n485, DataPath_RF_SELBLOCK_INLOC_n484, 
      DataPath_RF_SELBLOCK_INLOC_n483, DataPath_RF_SELBLOCK_INLOC_n482, 
      DataPath_RF_SELBLOCK_INLOC_n481, DataPath_RF_SELBLOCK_INLOC_n480, 
      DataPath_RF_SELBLOCK_INLOC_n479, DataPath_RF_SELBLOCK_INLOC_n478, 
      DataPath_RF_SELBLOCK_INLOC_n477, DataPath_RF_SELBLOCK_INLOC_n476, 
      DataPath_RF_SELBLOCK_INLOC_n475, DataPath_RF_SELBLOCK_INLOC_n474, 
      DataPath_RF_SELBLOCK_INLOC_n473, DataPath_RF_SELBLOCK_INLOC_n472, 
      DataPath_RF_SELBLOCK_INLOC_n471, DataPath_RF_SELBLOCK_INLOC_n470, 
      DataPath_RF_SELBLOCK_INLOC_n469, DataPath_RF_SELBLOCK_INLOC_n468, 
      DataPath_RF_SELBLOCK_INLOC_n467, DataPath_RF_SELBLOCK_INLOC_n466, 
      DataPath_RF_SELBLOCK_INLOC_n465, DataPath_RF_SELBLOCK_INLOC_n464, 
      DataPath_RF_SELBLOCK_INLOC_n463, DataPath_RF_SELBLOCK_INLOC_n462, 
      DataPath_RF_SELBLOCK_INLOC_n461, DataPath_RF_SELBLOCK_INLOC_n460, 
      DataPath_RF_SELBLOCK_INLOC_n459, DataPath_RF_SELBLOCK_INLOC_n458, 
      DataPath_RF_SELBLOCK_INLOC_n457, DataPath_RF_SELBLOCK_INLOC_n456, 
      DataPath_RF_SELBLOCK_INLOC_n455, DataPath_RF_SELBLOCK_INLOC_n454, 
      DataPath_RF_SELBLOCK_INLOC_n453, DataPath_RF_SELBLOCK_INLOC_n452, 
      DataPath_RF_SELBLOCK_INLOC_n451, DataPath_RF_SELBLOCK_INLOC_n450, 
      DataPath_RF_SELBLOCK_INLOC_n449, DataPath_RF_SELBLOCK_INLOC_n448, 
      DataPath_RF_SELBLOCK_INLOC_n447, DataPath_RF_SELBLOCK_INLOC_n446, 
      DataPath_RF_SELBLOCK_INLOC_n445, DataPath_RF_SELBLOCK_INLOC_n444, 
      DataPath_RF_SELBLOCK_INLOC_n443, DataPath_RF_SELBLOCK_INLOC_n442, 
      DataPath_RF_SELBLOCK_INLOC_n441, DataPath_RF_SELBLOCK_INLOC_n440, 
      DataPath_RF_SELBLOCK_INLOC_n439, DataPath_RF_SELBLOCK_INLOC_n438, 
      DataPath_RF_SELBLOCK_INLOC_n437, DataPath_RF_SELBLOCK_INLOC_n436, 
      DataPath_RF_SELBLOCK_INLOC_n435, DataPath_RF_SELBLOCK_INLOC_n434, 
      DataPath_RF_SELBLOCK_INLOC_n433, DataPath_RF_SELBLOCK_INLOC_n432, 
      DataPath_RF_SELBLOCK_INLOC_n431, DataPath_RF_SELBLOCK_INLOC_n430, 
      DataPath_RF_SELBLOCK_INLOC_n429, DataPath_RF_SELBLOCK_INLOC_n428, 
      DataPath_RF_SELBLOCK_INLOC_n427, DataPath_RF_SELBLOCK_INLOC_n426, 
      DataPath_RF_SELBLOCK_INLOC_n425, DataPath_RF_SELBLOCK_INLOC_n424, 
      DataPath_RF_SELBLOCK_INLOC_n423, DataPath_RF_SELBLOCK_INLOC_n422, 
      DataPath_RF_SELBLOCK_INLOC_n421, DataPath_RF_SELBLOCK_INLOC_n420, 
      DataPath_RF_SELBLOCK_INLOC_n419, DataPath_RF_SELBLOCK_INLOC_n418, 
      DataPath_RF_SELBLOCK_INLOC_n417, DataPath_RF_SELBLOCK_INLOC_n416, 
      DataPath_RF_SELBLOCK_INLOC_n415, DataPath_RF_SELBLOCK_INLOC_n414, 
      DataPath_RF_SELBLOCK_INLOC_n413, DataPath_RF_SELBLOCK_INLOC_n412, 
      DataPath_RF_SELBLOCK_INLOC_n411, DataPath_RF_SELBLOCK_INLOC_n410, 
      DataPath_RF_SELBLOCK_INLOC_n409, DataPath_RF_SELBLOCK_INLOC_n408, 
      DataPath_RF_SELBLOCK_INLOC_n407, DataPath_RF_SELBLOCK_INLOC_n406, 
      DataPath_RF_SELBLOCK_INLOC_n405, DataPath_RF_SELBLOCK_INLOC_n404, 
      DataPath_RF_SELBLOCK_INLOC_n403, DataPath_RF_SELBLOCK_INLOC_n402, 
      DataPath_RF_SELBLOCK_INLOC_n401, DataPath_RF_SELBLOCK_INLOC_n400, 
      DataPath_RF_SELBLOCK_INLOC_n399, DataPath_RF_SELBLOCK_INLOC_n398, 
      DataPath_RF_SELBLOCK_INLOC_n397, DataPath_RF_SELBLOCK_INLOC_n396, 
      DataPath_RF_SELBLOCK_INLOC_n395, DataPath_RF_SELBLOCK_INLOC_n394, 
      DataPath_RF_SELBLOCK_INLOC_n393, DataPath_RF_SELBLOCK_INLOC_n392, 
      DataPath_RF_SELBLOCK_INLOC_n391, DataPath_RF_SELBLOCK_INLOC_n390, 
      DataPath_RF_SELBLOCK_INLOC_n389, DataPath_RF_SELBLOCK_INLOC_n388, 
      DataPath_RF_SELBLOCK_INLOC_n387, DataPath_RF_SELBLOCK_INLOC_n386, 
      DataPath_RF_SELBLOCK_INLOC_n385, DataPath_RF_SELBLOCK_INLOC_n384, 
      DataPath_RF_SELBLOCK_INLOC_n383, DataPath_RF_SELBLOCK_INLOC_n382, 
      DataPath_RF_SELBLOCK_INLOC_n381, DataPath_RF_SELBLOCK_INLOC_n380, 
      DataPath_RF_SELBLOCK_INLOC_n379, DataPath_RF_SELBLOCK_INLOC_n378, 
      DataPath_RF_SELBLOCK_INLOC_n377, DataPath_RF_SELBLOCK_INLOC_n376, 
      DataPath_RF_SELBLOCK_INLOC_n375, DataPath_RF_SELBLOCK_INLOC_n374, 
      DataPath_RF_SELBLOCK_INLOC_n373, DataPath_RF_SELBLOCK_INLOC_n372, 
      DataPath_RF_SELBLOCK_INLOC_n371, DataPath_RF_SELBLOCK_INLOC_n370, 
      DataPath_RF_SELBLOCK_INLOC_n369, DataPath_RF_SELBLOCK_INLOC_n368, 
      DataPath_RF_SELBLOCK_INLOC_n367, DataPath_RF_SELBLOCK_INLOC_n366, 
      DataPath_RF_SELBLOCK_INLOC_n365, DataPath_RF_SELBLOCK_INLOC_n364, 
      DataPath_RF_SELBLOCK_INLOC_n363, DataPath_RF_SELBLOCK_INLOC_n362, 
      DataPath_RF_SELBLOCK_INLOC_n361, DataPath_RF_SELBLOCK_INLOC_n360, 
      DataPath_RF_SELBLOCK_INLOC_n359, DataPath_RF_SELBLOCK_INLOC_n358, 
      DataPath_RF_SELBLOCK_INLOC_n357, DataPath_RF_SELBLOCK_INLOC_n356, 
      DataPath_RF_SELBLOCK_INLOC_n355, DataPath_RF_SELBLOCK_INLOC_n354, 
      DataPath_RF_SELBLOCK_INLOC_n353, DataPath_RF_SELBLOCK_INLOC_n352, 
      DataPath_RF_SELBLOCK_INLOC_n351, DataPath_RF_SELBLOCK_INLOC_n350, 
      DataPath_RF_SELBLOCK_INLOC_n349, DataPath_RF_SELBLOCK_INLOC_n348, 
      DataPath_RF_SELBLOCK_INLOC_n347, DataPath_RF_SELBLOCK_INLOC_n346, 
      DataPath_RF_SELBLOCK_INLOC_n345, DataPath_RF_SELBLOCK_INLOC_n344, 
      DataPath_RF_SELBLOCK_INLOC_n343, DataPath_RF_SELBLOCK_INLOC_n342, 
      DataPath_RF_SELBLOCK_INLOC_n341, DataPath_RF_SELBLOCK_INLOC_n340, 
      DataPath_RF_SELBLOCK_INLOC_n339, DataPath_RF_SELBLOCK_INLOC_n338, 
      DataPath_RF_SELBLOCK_INLOC_n337, DataPath_RF_SELBLOCK_INLOC_n336, 
      DataPath_RF_SELBLOCK_INLOC_n335, DataPath_RF_SELBLOCK_INLOC_n334, 
      DataPath_RF_SELBLOCK_INLOC_n333, DataPath_RF_SELBLOCK_INLOC_n332, 
      DataPath_RF_SELBLOCK_INLOC_n331, DataPath_RF_SELBLOCK_INLOC_n330, 
      DataPath_RF_SELBLOCK_INLOC_n329, DataPath_RF_SELBLOCK_INLOC_n328, 
      DataPath_RF_SELBLOCK_INLOC_n327, DataPath_RF_SELBLOCK_INLOC_n326, 
      DataPath_RF_SELBLOCK_INLOC_n325, DataPath_RF_SELBLOCK_INLOC_n324, 
      DataPath_RF_SELBLOCK_INLOC_n323, DataPath_RF_SELBLOCK_INLOC_n322, 
      DataPath_RF_SELBLOCK_INLOC_n321, DataPath_RF_SELBLOCK_INLOC_n320, 
      DataPath_RF_SELBLOCK_INLOC_n319, DataPath_RF_SELBLOCK_INLOC_n318, 
      DataPath_RF_SELBLOCK_INLOC_n317, DataPath_RF_SELBLOCK_INLOC_n316, 
      DataPath_RF_SELBLOCK_INLOC_n315, DataPath_RF_SELBLOCK_INLOC_n314, 
      DataPath_RF_SELBLOCK_INLOC_n313, DataPath_RF_SELBLOCK_INLOC_n312, 
      DataPath_RF_SELBLOCK_INLOC_n311, DataPath_RF_SELBLOCK_INLOC_n310, 
      DataPath_RF_SELBLOCK_INLOC_n309, DataPath_RF_SELBLOCK_INLOC_n308, 
      DataPath_RF_SELBLOCK_INLOC_n307, DataPath_RF_SELBLOCK_INLOC_n306, 
      DataPath_RF_SELBLOCK_INLOC_n305, DataPath_RF_SELBLOCK_INLOC_n304, 
      DataPath_RF_SELBLOCK_INLOC_n303, DataPath_RF_SELBLOCK_INLOC_n302, 
      DataPath_RF_SELBLOCK_INLOC_n301, DataPath_RF_SELBLOCK_INLOC_n300, 
      DataPath_RF_SELBLOCK_INLOC_n299, DataPath_RF_SELBLOCK_INLOC_n298, 
      DataPath_RF_SELBLOCK_INLOC_n297, DataPath_RF_SELBLOCK_INLOC_n296, 
      DataPath_RF_SELBLOCK_INLOC_n295, DataPath_RF_SELBLOCK_INLOC_n294, 
      DataPath_RF_SELBLOCK_INLOC_n293, DataPath_RF_SELBLOCK_INLOC_n292, 
      DataPath_RF_SELBLOCK_INLOC_n291, DataPath_RF_SELBLOCK_INLOC_n290, 
      DataPath_RF_SELBLOCK_INLOC_n289, DataPath_RF_SELBLOCK_INLOC_n288, 
      DataPath_RF_SELBLOCK_INLOC_n287, DataPath_RF_SELBLOCK_INLOC_n286, 
      DataPath_RF_SELBLOCK_INLOC_n285, DataPath_RF_SELBLOCK_INLOC_n284, 
      DataPath_RF_SELBLOCK_INLOC_n283, DataPath_RF_SELBLOCK_INLOC_n282, 
      DataPath_RF_SELBLOCK_INLOC_n281, DataPath_RF_SELBLOCK_INLOC_n280, 
      DataPath_RF_SELBLOCK_INLOC_n279, DataPath_RF_SELBLOCK_INLOC_n278, 
      DataPath_RF_SELBLOCK_INLOC_n277, DataPath_RF_SELBLOCK_INLOC_n276, 
      DataPath_RF_SELBLOCK_INLOC_n275, DataPath_RF_SELBLOCK_INLOC_n274, 
      DataPath_RF_SELBLOCK_INLOC_n273, DataPath_RF_SELBLOCK_INLOC_n272, 
      DataPath_RF_SELBLOCK_INLOC_n271, DataPath_RF_SELBLOCK_INLOC_n270, 
      DataPath_RF_SELBLOCK_INLOC_n269, DataPath_RF_SELBLOCK_INLOC_n268, 
      DataPath_RF_SELBLOCK_INLOC_n267, DataPath_RF_SELBLOCK_INLOC_n266, 
      DataPath_RF_SELBLOCK_INLOC_n265, DataPath_RF_SELBLOCK_INLOC_n264, 
      DataPath_RF_SELBLOCK_INLOC_n263, DataPath_RF_SELBLOCK_INLOC_n262, 
      DataPath_RF_SELBLOCK_INLOC_n261, DataPath_RF_SELBLOCK_INLOC_n260, 
      DataPath_RF_SELBLOCK_INLOC_n259, DataPath_RF_SELBLOCK_INLOC_n258, 
      DataPath_RF_SELBLOCK_INLOC_n257, DataPath_RF_SELBLOCK_INLOC_n256, 
      DataPath_RF_SELBLOCK_INLOC_n255, DataPath_RF_SELBLOCK_INLOC_n254, 
      DataPath_RF_SELBLOCK_INLOC_n253, DataPath_RF_SELBLOCK_INLOC_n252, 
      DataPath_RF_SELBLOCK_INLOC_n251, DataPath_RF_SELBLOCK_INLOC_n250, 
      DataPath_RF_SELBLOCK_INLOC_n249, DataPath_RF_SELBLOCK_INLOC_n248, 
      DataPath_RF_SELBLOCK_INLOC_n247, DataPath_RF_SELBLOCK_INLOC_n246, 
      DataPath_RF_SELBLOCK_INLOC_n245, DataPath_RF_SELBLOCK_INLOC_n244, 
      DataPath_RF_SELBLOCK_INLOC_n243, DataPath_RF_SELBLOCK_INLOC_n242, 
      DataPath_RF_SELBLOCK_INLOC_n241, DataPath_RF_SELBLOCK_INLOC_n240, 
      DataPath_RF_SELBLOCK_INLOC_n239, DataPath_RF_SELBLOCK_INLOC_n238, 
      DataPath_RF_SELBLOCK_INLOC_n237, DataPath_RF_SELBLOCK_INLOC_n236, 
      DataPath_RF_SELBLOCK_INLOC_n235, DataPath_RF_SELBLOCK_INLOC_n234, 
      DataPath_RF_SELBLOCK_INLOC_n233, DataPath_RF_SELBLOCK_INLOC_n232, 
      DataPath_RF_SELBLOCK_INLOC_n231, DataPath_RF_SELBLOCK_INLOC_n230, 
      DataPath_RF_SELBLOCK_INLOC_n229, DataPath_RF_SELBLOCK_INLOC_n228, 
      DataPath_RF_SELBLOCK_INLOC_n227, DataPath_RF_SELBLOCK_INLOC_n226, 
      DataPath_RF_SELBLOCK_INLOC_n225, DataPath_RF_SELBLOCK_INLOC_n224, 
      DataPath_RF_SELBLOCK_INLOC_n223, DataPath_RF_SELBLOCK_INLOC_n222, 
      DataPath_RF_SELBLOCK_INLOC_n221, DataPath_RF_SELBLOCK_INLOC_n220, 
      DataPath_RF_SELBLOCK_INLOC_n219, DataPath_RF_SELBLOCK_INLOC_n218, 
      DataPath_RF_SELBLOCK_INLOC_n217, DataPath_RF_SELBLOCK_INLOC_n216, 
      DataPath_RF_SELBLOCK_INLOC_n215, DataPath_RF_SELBLOCK_INLOC_n214, 
      DataPath_RF_SELBLOCK_INLOC_n213, DataPath_RF_SELBLOCK_INLOC_n212, 
      DataPath_RF_SELBLOCK_INLOC_n211, DataPath_RF_SELBLOCK_INLOC_n210, 
      DataPath_RF_SELBLOCK_INLOC_n209, DataPath_RF_SELBLOCK_INLOC_n208, 
      DataPath_RF_SELBLOCK_INLOC_n207, DataPath_RF_SELBLOCK_INLOC_n206, 
      DataPath_RF_SELBLOCK_INLOC_n205, DataPath_RF_SELBLOCK_INLOC_n204, 
      DataPath_RF_SELBLOCK_INLOC_n203, DataPath_RF_SELBLOCK_INLOC_n202, 
      DataPath_RF_SELBLOCK_INLOC_n201, DataPath_RF_SELBLOCK_INLOC_n200, 
      DataPath_RF_SELBLOCK_INLOC_n199, DataPath_RF_SELBLOCK_INLOC_n198, 
      DataPath_RF_SELBLOCK_INLOC_n197, DataPath_RF_SELBLOCK_INLOC_n196, 
      DataPath_RF_SELBLOCK_INLOC_n195, DataPath_RF_SELBLOCK_INLOC_n194, 
      DataPath_RF_SELBLOCK_INLOC_n193, DataPath_RF_SELBLOCK_INLOC_n192, 
      DataPath_RF_SELBLOCK_INLOC_n191, DataPath_RF_SELBLOCK_INLOC_n190, 
      DataPath_RF_SELBLOCK_INLOC_n189, DataPath_RF_SELBLOCK_INLOC_n188, 
      DataPath_RF_SELBLOCK_INLOC_n187, DataPath_RF_SELBLOCK_INLOC_n186, 
      DataPath_RF_SELBLOCK_INLOC_n185, DataPath_RF_SELBLOCK_INLOC_n184, 
      DataPath_RF_SELBLOCK_INLOC_n183, DataPath_RF_SELBLOCK_INLOC_n182, 
      DataPath_RF_SELBLOCK_INLOC_n181, DataPath_RF_SELBLOCK_INLOC_n180, 
      DataPath_RF_SELBLOCK_INLOC_n179, DataPath_RF_SELBLOCK_INLOC_n178, 
      DataPath_RF_SELBLOCK_INLOC_n177, DataPath_RF_SELBLOCK_INLOC_n176, 
      DataPath_RF_SELBLOCK_INLOC_n175, DataPath_RF_SELBLOCK_INLOC_n174, 
      DataPath_RF_SELBLOCK_INLOC_n173, DataPath_RF_SELBLOCK_INLOC_n172, 
      DataPath_RF_SELBLOCK_INLOC_n171, DataPath_RF_SELBLOCK_INLOC_n170, 
      DataPath_RF_SELBLOCK_INLOC_n169, DataPath_RF_SELBLOCK_INLOC_n168, 
      DataPath_RF_SELBLOCK_INLOC_n167, DataPath_RF_SELBLOCK_INLOC_n166, 
      DataPath_RF_SELBLOCK_INLOC_n165, DataPath_RF_SELBLOCK_INLOC_n164, 
      DataPath_RF_SELBLOCK_INLOC_n163, DataPath_RF_SELBLOCK_INLOC_n162, 
      DataPath_RF_SELBLOCK_INLOC_n161, DataPath_RF_SELBLOCK_INLOC_n160, 
      DataPath_RF_SELBLOCK_INLOC_n159, DataPath_RF_SELBLOCK_INLOC_n158, 
      DataPath_RF_SELBLOCK_INLOC_n157, DataPath_RF_SELBLOCK_INLOC_n156, 
      DataPath_RF_SELBLOCK_INLOC_n155, DataPath_RF_SELBLOCK_INLOC_n154, 
      DataPath_RF_SELBLOCK_INLOC_n153, DataPath_RF_SELBLOCK_INLOC_n152, 
      DataPath_RF_SELBLOCK_INLOC_n151, DataPath_RF_SELBLOCK_INLOC_n150, 
      DataPath_RF_SELBLOCK_INLOC_n149, DataPath_RF_SELBLOCK_INLOC_n148, 
      DataPath_RF_SELBLOCK_INLOC_n147, DataPath_RF_SELBLOCK_INLOC_n146, 
      DataPath_RF_SELBLOCK_INLOC_n145, DataPath_RF_SELBLOCK_INLOC_n144, 
      DataPath_RF_SELBLOCK_INLOC_n143, DataPath_RF_SELBLOCK_INLOC_n142, 
      DataPath_RF_SELBLOCK_INLOC_n141, DataPath_RF_SELBLOCK_INLOC_n140, 
      DataPath_RF_SELBLOCK_INLOC_n139, DataPath_RF_SELBLOCK_INLOC_n138, 
      DataPath_RF_SELBLOCK_INLOC_n137, DataPath_RF_SELBLOCK_INLOC_n136, 
      DataPath_RF_SELBLOCK_INLOC_n135, DataPath_RF_SELBLOCK_INLOC_n134, 
      DataPath_RF_SELBLOCK_INLOC_n133, DataPath_RF_SELBLOCK_INLOC_n132, 
      DataPath_RF_SELBLOCK_INLOC_n131, DataPath_RF_SELBLOCK_INLOC_n130, 
      DataPath_RF_SELBLOCK_INLOC_n129, DataPath_RF_SELBLOCK_INLOC_n128, 
      DataPath_RF_SELBLOCK_INLOC_n127, DataPath_RF_SELBLOCK_INLOC_n126, 
      DataPath_RF_SELBLOCK_INLOC_n125, DataPath_RF_SELBLOCK_INLOC_n124, 
      DataPath_RF_SELBLOCK_INLOC_n123, DataPath_RF_SELBLOCK_INLOC_n122, 
      DataPath_RF_SELBLOCK_INLOC_n121, DataPath_RF_SELBLOCK_INLOC_n120, 
      DataPath_RF_SELBLOCK_INLOC_n119, DataPath_RF_SELBLOCK_INLOC_n118, 
      DataPath_RF_SELBLOCK_INLOC_n117, DataPath_RF_SELBLOCK_INLOC_n116, 
      DataPath_RF_SELBLOCK_INLOC_n115, DataPath_RF_SELBLOCK_INLOC_n114, 
      DataPath_RF_SELBLOCK_INLOC_n113, DataPath_RF_SELBLOCK_INLOC_n112, 
      DataPath_RF_SELBLOCK_INLOC_n111, DataPath_RF_SELBLOCK_INLOC_n110, 
      DataPath_RF_SELBLOCK_INLOC_n109, DataPath_RF_SELBLOCK_INLOC_n108, 
      DataPath_RF_SELBLOCK_INLOC_n107, DataPath_RF_SELBLOCK_INLOC_n106, 
      DataPath_RF_SELBLOCK_INLOC_n105, DataPath_RF_SELBLOCK_INLOC_n104, 
      DataPath_RF_SELBLOCK_INLOC_n103, DataPath_RF_SELBLOCK_INLOC_n102, 
      DataPath_RF_SELBLOCK_INLOC_n101, DataPath_RF_SELBLOCK_INLOC_n100, 
      DataPath_RF_SELBLOCK_INLOC_n99, DataPath_RF_SELBLOCK_INLOC_n98, 
      DataPath_RF_SELBLOCK_INLOC_n97, DataPath_RF_SELBLOCK_INLOC_n96, 
      DataPath_RF_SELBLOCK_INLOC_n95, DataPath_RF_SELBLOCK_INLOC_n94, 
      DataPath_RF_SELBLOCK_INLOC_n93, DataPath_RF_SELBLOCK_INLOC_n92, 
      DataPath_RF_SELBLOCK_INLOC_n91, DataPath_RF_SELBLOCK_INLOC_n90, 
      DataPath_RF_SELBLOCK_INLOC_n89, DataPath_RF_SELBLOCK_INLOC_n88, 
      DataPath_RF_SELBLOCK_INLOC_n87, DataPath_RF_SELBLOCK_INLOC_n86, 
      DataPath_RF_SELBLOCK_INLOC_n85, DataPath_RF_SELBLOCK_INLOC_n84, 
      DataPath_RF_SELBLOCK_INLOC_n83, DataPath_RF_SELBLOCK_INLOC_n82, 
      DataPath_RF_SELBLOCK_INLOC_n81, DataPath_RF_SELBLOCK_INLOC_n80, 
      DataPath_RF_SELBLOCK_INLOC_n79, DataPath_RF_SELBLOCK_INLOC_n78, 
      DataPath_RF_SELBLOCK_INLOC_n77, DataPath_RF_SELBLOCK_INLOC_n76, 
      DataPath_RF_SELBLOCK_INLOC_n75, DataPath_RF_SELBLOCK_INLOC_n74, 
      DataPath_RF_SELBLOCK_INLOC_n73, DataPath_RF_SELBLOCK_INLOC_n72, 
      DataPath_RF_SELBLOCK_INLOC_n71, DataPath_RF_SELBLOCK_INLOC_n70, 
      DataPath_RF_SELBLOCK_INLOC_n69, DataPath_RF_SELBLOCK_INLOC_n68, 
      DataPath_RF_SELBLOCK_INLOC_n67, DataPath_RF_SELBLOCK_INLOC_n66, 
      DataPath_RF_SELBLOCK_INLOC_n65, DataPath_RF_SELBLOCK_INLOC_n64, 
      DataPath_RF_SELBLOCK_INLOC_n63, DataPath_RF_SELBLOCK_INLOC_n62, 
      DataPath_RF_SELBLOCK_INLOC_n61, DataPath_RF_SELBLOCK_INLOC_n60, 
      DataPath_RF_SELBLOCK_INLOC_n59, DataPath_RF_SELBLOCK_INLOC_n58, 
      DataPath_RF_SELBLOCK_INLOC_n57, DataPath_RF_SELBLOCK_INLOC_n56, 
      DataPath_RF_SELBLOCK_INLOC_n55, DataPath_RF_SELBLOCK_INLOC_n54, 
      DataPath_RF_SELBLOCK_INLOC_n53, DataPath_RF_SELBLOCK_INLOC_n52, 
      DataPath_RF_SELBLOCK_INLOC_n51, DataPath_RF_SELBLOCK_INLOC_n50, 
      DataPath_RF_SELBLOCK_INLOC_n49, DataPath_RF_SELBLOCK_INLOC_n48, 
      DataPath_RF_SELBLOCK_INLOC_n47, DataPath_RF_SELBLOCK_INLOC_n46, 
      DataPath_RF_SELBLOCK_INLOC_n45, DataPath_RF_SELBLOCK_INLOC_n44, 
      DataPath_RF_SELBLOCK_INLOC_n43, DataPath_RF_SELBLOCK_INLOC_n42, 
      DataPath_RF_SELBLOCK_INLOC_n41, DataPath_RF_SELBLOCK_INLOC_n40, 
      DataPath_RF_SELBLOCK_INLOC_n39, DataPath_RF_SELBLOCK_INLOC_n38, 
      DataPath_RF_SELBLOCK_INLOC_n37, DataPath_RF_SELBLOCK_INLOC_n36, 
      DataPath_RF_SELBLOCK_INLOC_n35, DataPath_RF_SELBLOCK_INLOC_n34, 
      DataPath_RF_SELBLOCK_INLOC_n33, DataPath_RF_SELBLOCK_INLOC_n32, 
      DataPath_RF_SELBLOCK_INLOC_n31, DataPath_RF_SELBLOCK_INLOC_n30, 
      DataPath_RF_SELBLOCK_INLOC_n29, DataPath_RF_SELBLOCK_INLOC_n28, 
      DataPath_RF_SELBLOCK_INLOC_n27, DataPath_RF_SELBLOCK_INLOC_n26, 
      DataPath_RF_SELBLOCK_INLOC_n25, DataPath_RF_SELBLOCK_INLOC_n24, 
      DataPath_RF_SELBLOCK_INLOC_n23, DataPath_RF_SELBLOCK_INLOC_n22, 
      DataPath_RF_SELBLOCK_INLOC_n21, DataPath_RF_SELBLOCK_INLOC_n20, 
      DataPath_RF_SELBLOCK_INLOC_n19, DataPath_RF_SELBLOCK_INLOC_n18, 
      DataPath_RF_SELBLOCK_INLOC_n17, DataPath_RF_SELBLOCK_INLOC_n16, 
      DataPath_RF_SELBLOCK_INLOC_n15, DataPath_RF_SELBLOCK_INLOC_n14, 
      DataPath_RF_SELBLOCK_INLOC_n13, DataPath_RF_SELBLOCK_INLOC_n12, 
      DataPath_RF_SELBLOCK_INLOC_n11, DataPath_RF_SELBLOCK_INLOC_n10, 
      DataPath_RF_SELBLOCK_INLOC_n9, DataPath_RF_SELBLOCK_INLOC_n8, 
      DataPath_RF_SELBLOCK_INLOC_n7, DataPath_RF_SELBLOCK_INLOC_n6, 
      DataPath_RF_SELBLOCK_INLOC_n5, DataPath_RF_SELBLOCK_INLOC_n4, 
      DataPath_RF_PUSH_ADDRGEN_n54, DataPath_RF_PUSH_ADDRGEN_n53, 
      DataPath_RF_PUSH_ADDRGEN_n52, DataPath_RF_PUSH_ADDRGEN_n51, 
      DataPath_RF_PUSH_ADDRGEN_n50, DataPath_RF_PUSH_ADDRGEN_n49, 
      DataPath_RF_PUSH_ADDRGEN_n48, DataPath_RF_PUSH_ADDRGEN_n47, 
      DataPath_RF_PUSH_ADDRGEN_n46, DataPath_RF_PUSH_ADDRGEN_n45, 
      DataPath_RF_PUSH_ADDRGEN_n44, DataPath_RF_PUSH_ADDRGEN_n43, 
      DataPath_RF_PUSH_ADDRGEN_n42, DataPath_RF_PUSH_ADDRGEN_n41, 
      DataPath_RF_PUSH_ADDRGEN_n40, DataPath_RF_PUSH_ADDRGEN_n39, 
      DataPath_RF_PUSH_ADDRGEN_n38, DataPath_RF_PUSH_ADDRGEN_n37, 
      DataPath_RF_PUSH_ADDRGEN_n36, DataPath_RF_PUSH_ADDRGEN_n35, 
      DataPath_RF_PUSH_ADDRGEN_n34, DataPath_RF_PUSH_ADDRGEN_n33, 
      DataPath_RF_PUSH_ADDRGEN_n32, DataPath_RF_PUSH_ADDRGEN_n31, 
      DataPath_RF_PUSH_ADDRGEN_n30, DataPath_RF_PUSH_ADDRGEN_n29, 
      DataPath_RF_PUSH_ADDRGEN_n28, DataPath_RF_PUSH_ADDRGEN_n27, 
      DataPath_RF_PUSH_ADDRGEN_n26, DataPath_RF_PUSH_ADDRGEN_n22, 
      DataPath_RF_PUSH_ADDRGEN_n20, DataPath_RF_PUSH_ADDRGEN_n18, 
      DataPath_RF_PUSH_ADDRGEN_n17, DataPath_RF_PUSH_ADDRGEN_n16, 
      DataPath_RF_PUSH_ADDRGEN_n15, DataPath_RF_PUSH_ADDRGEN_n14, 
      DataPath_RF_PUSH_ADDRGEN_n13, DataPath_RF_PUSH_ADDRGEN_n12, 
      DataPath_RF_PUSH_ADDRGEN_n11, DataPath_RF_PUSH_ADDRGEN_n10, 
      DataPath_RF_PUSH_ADDRGEN_n9, DataPath_RF_PUSH_ADDRGEN_n8, 
      DataPath_RF_PUSH_ADDRGEN_n7, DataPath_RF_PUSH_ADDRGEN_n6, 
      DataPath_RF_PUSH_ADDRGEN_n5, DataPath_RF_PUSH_ADDRGEN_n4, 
      DataPath_RF_PUSH_ADDRGEN_n1, DataPath_RF_PUSH_ADDRGEN_N61, 
      DataPath_RF_PUSH_ADDRGEN_N60, DataPath_RF_PUSH_ADDRGEN_N59, 
      DataPath_RF_PUSH_ADDRGEN_N58, DataPath_RF_PUSH_ADDRGEN_N57, 
      DataPath_RF_PUSH_ADDRGEN_N56, DataPath_RF_PUSH_ADDRGEN_N55, 
      DataPath_RF_PUSH_ADDRGEN_N54_port, DataPath_RF_PUSH_ADDRGEN_N53_port, 
      DataPath_RF_PUSH_ADDRGEN_N52_port, DataPath_RF_PUSH_ADDRGEN_N51_port, 
      DataPath_RF_PUSH_ADDRGEN_N50_port, DataPath_RF_PUSH_ADDRGEN_N49_port, 
      DataPath_RF_PUSH_ADDRGEN_N48_port, DataPath_RF_PUSH_ADDRGEN_N47_port, 
      DataPath_RF_PUSH_ADDRGEN_N46_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_state_1_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, DataPath_RF_SPILLADDR_ENC_n34
      , DataPath_RF_SPILLADDR_ENC_n33, DataPath_RF_SPILLADDR_ENC_n32, 
      DataPath_RF_SPILLADDR_ENC_n31, DataPath_RF_SPILLADDR_ENC_n30, 
      DataPath_RF_SPILLADDR_ENC_n29, DataPath_RF_SPILLADDR_ENC_n28, 
      DataPath_RF_SPILLADDR_ENC_n27, DataPath_RF_SPILLADDR_ENC_n26, 
      DataPath_RF_SPILLADDR_ENC_n25, DataPath_RF_SPILLADDR_ENC_n24, 
      DataPath_RF_SPILLADDR_ENC_n23, DataPath_RF_SPILLADDR_ENC_n22, 
      DataPath_RF_SPILLADDR_ENC_n21, DataPath_RF_SPILLADDR_ENC_n20, 
      DataPath_RF_SPILLADDR_ENC_n19, DataPath_RF_SPILLADDR_ENC_n18, 
      DataPath_RF_SPILLADDR_ENC_n17, DataPath_RF_SPILLADDR_ENC_n16, 
      DataPath_RF_SPILLADDR_ENC_n15, DataPath_RF_SPILLADDR_ENC_n14, 
      DataPath_RF_SPILLADDR_ENC_n13, DataPath_RF_SPILLADDR_ENC_n12, 
      DataPath_RF_RDPORT_SPILL_n347, DataPath_RF_RDPORT_SPILL_n346, 
      DataPath_RF_RDPORT_SPILL_n345, DataPath_RF_RDPORT_SPILL_n344, 
      DataPath_RF_RDPORT_SPILL_n343, DataPath_RF_RDPORT_SPILL_n342, 
      DataPath_RF_RDPORT_SPILL_n341, DataPath_RF_RDPORT_SPILL_n340, 
      DataPath_RF_RDPORT_SPILL_n339, DataPath_RF_RDPORT_SPILL_n338, 
      DataPath_RF_RDPORT_SPILL_n337, DataPath_RF_RDPORT_SPILL_n336, 
      DataPath_RF_RDPORT_SPILL_n335, DataPath_RF_RDPORT_SPILL_n334, 
      DataPath_RF_RDPORT_SPILL_n333, DataPath_RF_RDPORT_SPILL_n332, 
      DataPath_RF_RDPORT_SPILL_n331, DataPath_RF_RDPORT_SPILL_n330, 
      DataPath_RF_RDPORT_SPILL_n329, DataPath_RF_RDPORT_SPILL_n328, 
      DataPath_RF_RDPORT_SPILL_n327, DataPath_RF_RDPORT_SPILL_n326, 
      DataPath_RF_RDPORT_SPILL_n325, DataPath_RF_RDPORT_SPILL_n324, 
      DataPath_RF_RDPORT_SPILL_n323, DataPath_RF_RDPORT_SPILL_n322, 
      DataPath_RF_RDPORT_SPILL_n321, DataPath_RF_RDPORT_SPILL_n320, 
      DataPath_RF_RDPORT_SPILL_n319, DataPath_RF_RDPORT_SPILL_n318, 
      DataPath_RF_RDPORT_SPILL_n317, DataPath_RF_RDPORT_SPILL_n316, 
      DataPath_RF_RDPORT_SPILL_n315, DataPath_RF_RDPORT_SPILL_n314, 
      DataPath_RF_RDPORT_SPILL_n313, DataPath_RF_RDPORT_SPILL_n312, 
      DataPath_RF_RDPORT_SPILL_n311, DataPath_RF_RDPORT_SPILL_n310, 
      DataPath_RF_RDPORT_SPILL_n309, DataPath_RF_RDPORT_SPILL_n308, 
      DataPath_RF_RDPORT_SPILL_n307, DataPath_RF_RDPORT_SPILL_n306, 
      DataPath_RF_RDPORT_SPILL_n305, DataPath_RF_RDPORT_SPILL_n304, 
      DataPath_RF_RDPORT_SPILL_n303, DataPath_RF_RDPORT_SPILL_n302, 
      DataPath_RF_RDPORT_SPILL_n301, DataPath_RF_RDPORT_SPILL_n300, 
      DataPath_RF_RDPORT_SPILL_n299, DataPath_RF_RDPORT_SPILL_n298, 
      DataPath_RF_RDPORT_SPILL_n297, DataPath_RF_RDPORT_SPILL_n296, 
      DataPath_RF_RDPORT_SPILL_n295, DataPath_RF_RDPORT_SPILL_n294, 
      DataPath_RF_RDPORT_SPILL_n293, DataPath_RF_RDPORT_SPILL_n292, 
      DataPath_RF_RDPORT_SPILL_n291, DataPath_RF_RDPORT_SPILL_n290, 
      DataPath_RF_RDPORT_SPILL_n289, DataPath_RF_RDPORT_SPILL_n288, 
      DataPath_RF_RDPORT_SPILL_n287, DataPath_RF_RDPORT_SPILL_n286, 
      DataPath_RF_RDPORT_SPILL_n285, DataPath_RF_RDPORT_SPILL_n284, 
      DataPath_RF_RDPORT_SPILL_n283, DataPath_RF_RDPORT_SPILL_n282, 
      DataPath_RF_RDPORT_SPILL_n281, DataPath_RF_RDPORT_SPILL_n280, 
      DataPath_RF_RDPORT_SPILL_n279, DataPath_RF_RDPORT_SPILL_n278, 
      DataPath_RF_RDPORT_SPILL_n277, DataPath_RF_RDPORT_SPILL_n276, 
      DataPath_RF_RDPORT_SPILL_n275, DataPath_RF_RDPORT_SPILL_n274, 
      DataPath_RF_RDPORT_SPILL_n273, DataPath_RF_RDPORT_SPILL_n272, 
      DataPath_RF_RDPORT_SPILL_n271, DataPath_RF_RDPORT_SPILL_n270, 
      DataPath_RF_RDPORT_SPILL_n269, DataPath_RF_RDPORT_SPILL_n268, 
      DataPath_RF_RDPORT_SPILL_n267, DataPath_RF_RDPORT_SPILL_n266, 
      DataPath_RF_RDPORT_SPILL_n265, DataPath_RF_RDPORT_SPILL_n264, 
      DataPath_RF_RDPORT_SPILL_n263, DataPath_RF_RDPORT_SPILL_n262, 
      DataPath_RF_RDPORT_SPILL_n261, DataPath_RF_RDPORT_SPILL_n260, 
      DataPath_RF_RDPORT_SPILL_n259, DataPath_RF_RDPORT_SPILL_n258, 
      DataPath_RF_RDPORT_SPILL_n257, DataPath_RF_RDPORT_SPILL_n256, 
      DataPath_RF_RDPORT_SPILL_n255, DataPath_RF_RDPORT_SPILL_n254, 
      DataPath_RF_RDPORT_SPILL_n253, DataPath_RF_RDPORT_SPILL_n252, 
      DataPath_RF_RDPORT_SPILL_n251, DataPath_RF_RDPORT_SPILL_n250, 
      DataPath_RF_RDPORT_SPILL_n249, DataPath_RF_RDPORT_SPILL_n248, 
      DataPath_RF_RDPORT_SPILL_n247, DataPath_RF_RDPORT_SPILL_n246, 
      DataPath_RF_RDPORT_SPILL_n245, DataPath_RF_RDPORT_SPILL_n244, 
      DataPath_RF_RDPORT_SPILL_n243, DataPath_RF_RDPORT_SPILL_n242, 
      DataPath_RF_RDPORT_SPILL_n241, DataPath_RF_RDPORT_SPILL_n240, 
      DataPath_RF_RDPORT_SPILL_n239, DataPath_RF_RDPORT_SPILL_n238, 
      DataPath_RF_RDPORT_SPILL_n237, DataPath_RF_RDPORT_SPILL_n236, 
      DataPath_RF_RDPORT_SPILL_n235, DataPath_RF_RDPORT_SPILL_n234, 
      DataPath_RF_RDPORT_SPILL_n233, DataPath_RF_RDPORT_SPILL_n232, 
      DataPath_RF_RDPORT_SPILL_n231, DataPath_RF_RDPORT_SPILL_n230, 
      DataPath_RF_RDPORT_SPILL_n229, DataPath_RF_RDPORT_SPILL_n228, 
      DataPath_RF_RDPORT_SPILL_n227, DataPath_RF_RDPORT_SPILL_n226, 
      DataPath_RF_RDPORT_SPILL_n225, DataPath_RF_RDPORT_SPILL_n224, 
      DataPath_RF_RDPORT_SPILL_n223, DataPath_RF_RDPORT_SPILL_n222, 
      DataPath_RF_RDPORT_SPILL_n221, DataPath_RF_RDPORT_SPILL_n220, 
      DataPath_RF_RDPORT_SPILL_n219, DataPath_RF_RDPORT_SPILL_n218, 
      DataPath_RF_RDPORT_SPILL_n217, DataPath_RF_RDPORT_SPILL_n216, 
      DataPath_RF_RDPORT_SPILL_n215, DataPath_RF_RDPORT_SPILL_n214, 
      DataPath_RF_RDPORT_SPILL_n213, DataPath_RF_RDPORT_SPILL_n212, 
      DataPath_RF_RDPORT_SPILL_n211, DataPath_RF_RDPORT_SPILL_n210, 
      DataPath_RF_RDPORT_SPILL_n209, DataPath_RF_RDPORT_SPILL_n208, 
      DataPath_RF_RDPORT_SPILL_n207, DataPath_RF_RDPORT_SPILL_n206, 
      DataPath_RF_RDPORT_SPILL_n205, DataPath_RF_RDPORT_SPILL_n204, 
      DataPath_RF_RDPORT_SPILL_n203, DataPath_RF_RDPORT_SPILL_n202, 
      DataPath_RF_RDPORT_SPILL_n201, DataPath_RF_RDPORT_SPILL_n200, 
      DataPath_RF_RDPORT_SPILL_n199, DataPath_RF_RDPORT_SPILL_n198, 
      DataPath_RF_RDPORT_SPILL_n197, DataPath_RF_RDPORT_SPILL_n196, 
      DataPath_RF_RDPORT_SPILL_n195, DataPath_RF_RDPORT_SPILL_n194, 
      DataPath_RF_RDPORT_SPILL_n193, DataPath_RF_RDPORT_SPILL_n192, 
      DataPath_RF_RDPORT_SPILL_n191, DataPath_RF_RDPORT_SPILL_n190, 
      DataPath_RF_RDPORT_SPILL_n189, DataPath_RF_RDPORT_SPILL_n188, 
      DataPath_RF_RDPORT_SPILL_n187, DataPath_RF_RDPORT_SPILL_n186, 
      DataPath_RF_RDPORT_SPILL_n185, DataPath_RF_RDPORT_SPILL_n184, 
      DataPath_RF_RDPORT_SPILL_n183, DataPath_RF_RDPORT_SPILL_n182, 
      DataPath_RF_RDPORT_SPILL_n181, DataPath_RF_RDPORT_SPILL_n180, 
      DataPath_RF_RDPORT_SPILL_n179, DataPath_RF_RDPORT_SPILL_n178, 
      DataPath_RF_RDPORT_SPILL_n177, DataPath_RF_RDPORT_SPILL_n176, 
      DataPath_RF_RDPORT_SPILL_n175, DataPath_RF_RDPORT_SPILL_n174, 
      DataPath_RF_RDPORT_SPILL_n173, DataPath_RF_RDPORT_SPILL_n172, 
      DataPath_RF_RDPORT_SPILL_n171, DataPath_RF_RDPORT_SPILL_n170, 
      DataPath_RF_RDPORT_SPILL_n169, DataPath_RF_RDPORT_SPILL_n168, 
      DataPath_RF_RDPORT_SPILL_n167, DataPath_RF_RDPORT_SPILL_n166, 
      DataPath_RF_RDPORT_SPILL_n165, DataPath_RF_RDPORT_SPILL_n164, 
      DataPath_RF_RDPORT_SPILL_n163, DataPath_RF_RDPORT_SPILL_n162, 
      DataPath_RF_RDPORT_SPILL_n161, DataPath_RF_RDPORT_SPILL_n160, 
      DataPath_RF_RDPORT_SPILL_n159, DataPath_RF_RDPORT_SPILL_n158, 
      DataPath_RF_RDPORT_SPILL_n157, DataPath_RF_RDPORT_SPILL_n156, 
      DataPath_RF_RDPORT_SPILL_n155, DataPath_RF_RDPORT_SPILL_n154, 
      DataPath_RF_RDPORT_SPILL_n153, DataPath_RF_RDPORT_SPILL_n152, 
      DataPath_RF_RDPORT_SPILL_n151, DataPath_RF_RDPORT_SPILL_n150, 
      DataPath_RF_RDPORT_SPILL_n149, DataPath_RF_RDPORT_SPILL_n148, 
      DataPath_RF_RDPORT_SPILL_n147, DataPath_RF_RDPORT_SPILL_n146, 
      DataPath_RF_RDPORT_SPILL_n145, DataPath_RF_RDPORT_SPILL_n144, 
      DataPath_RF_RDPORT_SPILL_n143, DataPath_RF_RDPORT_SPILL_n142, 
      DataPath_RF_RDPORT_SPILL_n141, DataPath_RF_RDPORT_SPILL_n140, 
      DataPath_RF_RDPORT_SPILL_n139, DataPath_RF_RDPORT_SPILL_n138, 
      DataPath_RF_RDPORT_SPILL_n137, DataPath_RF_RDPORT_SPILL_n136, 
      DataPath_RF_RDPORT_SPILL_n135, DataPath_RF_RDPORT_SPILL_n134, 
      DataPath_RF_RDPORT_SPILL_n133, DataPath_RF_RDPORT_SPILL_n132, 
      DataPath_RF_RDPORT_SPILL_n131, DataPath_RF_RDPORT_SPILL_n130, 
      DataPath_RF_RDPORT_SPILL_n129, DataPath_RF_RDPORT_SPILL_n128, 
      DataPath_RF_RDPORT_SPILL_n127, DataPath_RF_RDPORT_SPILL_n126, 
      DataPath_RF_RDPORT_SPILL_n125, DataPath_RF_RDPORT_SPILL_n124, 
      DataPath_RF_RDPORT_SPILL_n123, DataPath_RF_RDPORT_SPILL_n122, 
      DataPath_RF_RDPORT_SPILL_n121, DataPath_RF_RDPORT_SPILL_n120, 
      DataPath_RF_RDPORT_SPILL_n119, DataPath_RF_RDPORT_SPILL_n118, 
      DataPath_RF_RDPORT_SPILL_n117, DataPath_RF_RDPORT_SPILL_n116, 
      DataPath_RF_RDPORT_SPILL_n115, DataPath_RF_RDPORT_SPILL_n114, 
      DataPath_RF_RDPORT_SPILL_n113, DataPath_RF_RDPORT_SPILL_n112, 
      DataPath_RF_RDPORT_SPILL_n111, DataPath_RF_RDPORT_SPILL_n110, 
      DataPath_RF_RDPORT_SPILL_n109, DataPath_RF_RDPORT_SPILL_n108, 
      DataPath_RF_RDPORT_SPILL_n107, DataPath_RF_RDPORT_SPILL_n106, 
      DataPath_RF_RDPORT_SPILL_n105, DataPath_RF_RDPORT_SPILL_n104, 
      DataPath_RF_RDPORT_SPILL_n103, DataPath_RF_RDPORT_SPILL_n102, 
      DataPath_RF_RDPORT_SPILL_n101, DataPath_RF_RDPORT_SPILL_n100, 
      DataPath_RF_RDPORT_SPILL_n99, DataPath_RF_RDPORT_SPILL_n98, 
      DataPath_RF_RDPORT_SPILL_n97, DataPath_RF_RDPORT_SPILL_n96, 
      DataPath_RF_RDPORT_SPILL_n95, DataPath_RF_RDPORT_SPILL_n94, 
      DataPath_RF_RDPORT_SPILL_n93, DataPath_RF_RDPORT_SPILL_n92, 
      DataPath_RF_RDPORT_SPILL_n91, DataPath_RF_RDPORT_SPILL_n90, 
      DataPath_RF_RDPORT_SPILL_n89, DataPath_RF_RDPORT_SPILL_n88, 
      DataPath_RF_RDPORT_SPILL_n87, DataPath_RF_RDPORT_SPILL_n86, 
      DataPath_RF_RDPORT_SPILL_n85, DataPath_RF_RDPORT_SPILL_n84, 
      DataPath_RF_RDPORT_SPILL_n83, DataPath_RF_RDPORT_SPILL_n82, 
      DataPath_RF_RDPORT_SPILL_n81, DataPath_RF_RDPORT_SPILL_n80, 
      DataPath_RF_RDPORT_SPILL_n79, DataPath_RF_RDPORT_SPILL_n78, 
      DataPath_RF_RDPORT_SPILL_n77, DataPath_RF_RDPORT_SPILL_n76, 
      DataPath_RF_RDPORT_SPILL_n75, DataPath_RF_RDPORT_SPILL_n74, 
      DataPath_RF_RDPORT_SPILL_n73, DataPath_RF_RDPORT_SPILL_n72, 
      DataPath_RF_RDPORT_SPILL_n71, DataPath_RF_RDPORT_SPILL_n70, 
      DataPath_RF_RDPORT_SPILL_n69, DataPath_RF_RDPORT_SPILL_n68, 
      DataPath_RF_RDPORT_SPILL_n67, DataPath_RF_RDPORT_SPILL_n66, 
      DataPath_RF_RDPORT_SPILL_n65, DataPath_RF_RDPORT_SPILL_n64, 
      DataPath_RF_RDPORT_SPILL_n63, DataPath_RF_RDPORT_SPILL_n62, 
      DataPath_RF_RDPORT_SPILL_n61, DataPath_RF_RDPORT_SPILL_n60, 
      DataPath_RF_RDPORT_SPILL_n59, DataPath_RF_RDPORT_SPILL_n58, 
      DataPath_RF_RDPORT_SPILL_n57, DataPath_RF_RDPORT_SPILL_n56, 
      DataPath_RF_RDPORT_SPILL_n55, DataPath_RF_RDPORT_SPILL_n54, 
      DataPath_RF_RDPORT_SPILL_n53, DataPath_RF_RDPORT_SPILL_n52, 
      DataPath_RF_RDPORT_SPILL_n51, DataPath_RF_RDPORT_SPILL_n50, 
      DataPath_RF_RDPORT_SPILL_n49, DataPath_RF_RDPORT_SPILL_n48, 
      DataPath_RF_RDPORT_SPILL_n47, DataPath_RF_RDPORT_SPILL_n46, 
      DataPath_RF_RDPORT_SPILL_n45, DataPath_RF_RDPORT_SPILL_n44, 
      DataPath_RF_RDPORT_SPILL_n43, DataPath_RF_RDPORT_SPILL_n42, 
      DataPath_RF_RDPORT_SPILL_n41, DataPath_RF_RDPORT_SPILL_n40, 
      DataPath_RF_RDPORT_SPILL_n39, DataPath_RF_RDPORT_SPILL_n38, 
      DataPath_RF_RDPORT_SPILL_n37, DataPath_RF_RDPORT_SPILL_n36, 
      DataPath_RF_RDPORT_SPILL_n35, DataPath_RF_RDPORT_SPILL_n34, 
      DataPath_RF_RDPORT_SPILL_n33, DataPath_RF_RDPORT_SPILL_n32, 
      DataPath_RF_RDPORT_SPILL_n31, DataPath_RF_RDPORT_SPILL_n30, 
      DataPath_RF_RDPORT_SPILL_n29, DataPath_RF_RDPORT_SPILL_n28, 
      DataPath_RF_RDPORT_SPILL_n27, DataPath_RF_RDPORT_SPILL_n26, 
      DataPath_RF_RDPORT_SPILL_n25, DataPath_RF_RDPORT_SPILL_n24, 
      DataPath_RF_RDPORT_SPILL_n23, DataPath_RF_RDPORT_SPILL_n22, 
      DataPath_RF_RDPORT_SPILL_n21, DataPath_RF_RDPORT_SPILL_n20, 
      DataPath_RF_RDPORT_SPILL_n19, DataPath_RF_RDPORT_SPILL_n18, 
      DataPath_RF_RDPORT_SPILL_n17, DataPath_RF_RDPORT_SPILL_n16, 
      DataPath_RF_RDPORT_SPILL_n15, DataPath_RF_RDPORT_SPILL_n14, 
      DataPath_RF_RDPORT_SPILL_n13, DataPath_RF_RDPORT_SPILL_n12, 
      DataPath_RF_RDPORT_SPILL_n11, DataPath_RF_RDPORT_SPILL_n10, 
      DataPath_RF_RDPORT_SPILL_n9, DataPath_RF_RDPORT_SPILL_n8, 
      DataPath_RF_RDPORT_SPILL_n7, DataPath_RF_RDPORT_SPILL_n6, 
      DataPath_RF_RDPORT_SPILL_n5, DataPath_RF_RDPORT_SPILL_n4, 
      DataPath_ALUhw_MUXOUT_n69, DataPath_ALUhw_MUXOUT_n68, 
      DataPath_ALUhw_MUXOUT_n67, DataPath_ALUhw_MUXOUT_n66, 
      DataPath_ALUhw_MUXOUT_n65, DataPath_ALUhw_MUXOUT_n64, 
      DataPath_ALUhw_MUXOUT_n63, DataPath_ALUhw_MUXOUT_n62, 
      DataPath_ALUhw_MUXOUT_n61, DataPath_ALUhw_MUXOUT_n60, 
      DataPath_ALUhw_MUXOUT_n59, DataPath_ALUhw_MUXOUT_n58, 
      DataPath_ALUhw_MUXOUT_n57, DataPath_ALUhw_MUXOUT_n56, 
      DataPath_ALUhw_MUXOUT_n55, DataPath_ALUhw_MUXOUT_n54, 
      DataPath_ALUhw_MUXOUT_n47, DataPath_ALUhw_MUXOUT_n46, 
      DataPath_ALUhw_MUXOUT_n25, DataPath_ALUhw_MUXOUT_n24, 
      DataPath_ALUhw_MUXOUT_n19, DataPath_ALUhw_MUXOUT_n18, 
      DataPath_ALUhw_MUXOUT_n17, DataPath_ALUhw_MUXOUT_n16, 
      DataPath_ALUhw_MUXOUT_n15, DataPath_ALUhw_MUXOUT_n14, 
      DataPath_ALUhw_MUXOUT_n13, DataPath_ALUhw_MUXOUT_n12, 
      DataPath_ALUhw_MUXOUT_n11, DataPath_ALUhw_MUXOUT_n10, 
      DataPath_ALUhw_MUXOUT_n9, DataPath_ALUhw_MUXOUT_n8, 
      DataPath_ALUhw_MUXOUT_n3, DataPath_ALUhw_MUXOUT_n2, 
      DataPath_ALUhw_BWISE_n137, DataPath_ALUhw_BWISE_n136, 
      DataPath_ALUhw_BWISE_n135, DataPath_ALUhw_BWISE_n72, 
      DataPath_ALUhw_BWISE_n71, DataPath_ALUhw_BWISE_n70, 
      DataPath_ALUhw_SHIFTER_HW_n641, DataPath_ALUhw_SHIFTER_HW_n639, 
      DataPath_ALUhw_SHIFTER_HW_n636, DataPath_ALUhw_SHIFTER_HW_n635, 
      DataPath_ALUhw_SHIFTER_HW_n626, DataPath_ALUhw_SHIFTER_HW_n625, 
      DataPath_ALUhw_SHIFTER_HW_n622, DataPath_ALUhw_SHIFTER_HW_n621, 
      DataPath_ALUhw_SHIFTER_HW_n606, DataPath_ALUhw_SHIFTER_HW_n603, 
      DataPath_ALUhw_SHIFTER_HW_n600, DataPath_ALUhw_SHIFTER_HW_n598, 
      DataPath_ALUhw_SHIFTER_HW_n597, DataPath_ALUhw_SHIFTER_HW_n588, 
      DataPath_ALUhw_SHIFTER_HW_n587, DataPath_ALUhw_SHIFTER_HW_n586, 
      DataPath_ALUhw_SHIFTER_HW_n585, DataPath_ALUhw_SHIFTER_HW_n584, 
      DataPath_ALUhw_SHIFTER_HW_n583, DataPath_ALUhw_SHIFTER_HW_n582, 
      DataPath_ALUhw_SHIFTER_HW_n576, DataPath_ALUhw_SHIFTER_HW_n552, 
      DataPath_ALUhw_SHIFTER_HW_n551, DataPath_ALUhw_SHIFTER_HW_n549, 
      DataPath_ALUhw_SHIFTER_HW_n548, DataPath_ALUhw_SHIFTER_HW_n540, 
      DataPath_ALUhw_SHIFTER_HW_n539, DataPath_ALUhw_SHIFTER_HW_n538, 
      DataPath_ALUhw_SHIFTER_HW_n537, DataPath_ALUhw_SHIFTER_HW_n536, 
      DataPath_ALUhw_SHIFTER_HW_n535, DataPath_ALUhw_SHIFTER_HW_n533, 
      DataPath_ALUhw_SHIFTER_HW_n529, DataPath_ALUhw_SHIFTER_HW_n526, 
      DataPath_ALUhw_SHIFTER_HW_n525, DataPath_ALUhw_SHIFTER_HW_n524, 
      DataPath_ALUhw_SHIFTER_HW_n523, DataPath_ALUhw_SHIFTER_HW_n522, 
      DataPath_ALUhw_SHIFTER_HW_n520, DataPath_ALUhw_SHIFTER_HW_n513, 
      DataPath_ALUhw_SHIFTER_HW_n512, DataPath_ALUhw_SHIFTER_HW_n511, 
      DataPath_ALUhw_SHIFTER_HW_n510, DataPath_ALUhw_SHIFTER_HW_n509, 
      DataPath_ALUhw_SHIFTER_HW_n508, DataPath_ALUhw_SHIFTER_HW_n507, 
      DataPath_ALUhw_SHIFTER_HW_n500, DataPath_ALUhw_SHIFTER_HW_n499, 
      DataPath_ALUhw_SHIFTER_HW_n498, DataPath_ALUhw_SHIFTER_HW_n497, 
      DataPath_ALUhw_SHIFTER_HW_n496, DataPath_ALUhw_SHIFTER_HW_n495, 
      DataPath_ALUhw_SHIFTER_HW_n494, DataPath_ALUhw_SHIFTER_HW_n487, 
      DataPath_ALUhw_SHIFTER_HW_n486, DataPath_ALUhw_SHIFTER_HW_n485, 
      DataPath_ALUhw_SHIFTER_HW_n484, DataPath_ALUhw_SHIFTER_HW_n483, 
      DataPath_ALUhw_SHIFTER_HW_n482, DataPath_ALUhw_SHIFTER_HW_n481, 
      DataPath_ALUhw_SHIFTER_HW_n478, DataPath_ALUhw_SHIFTER_HW_n472, 
      DataPath_ALUhw_SHIFTER_HW_n471, DataPath_ALUhw_SHIFTER_HW_n470, 
      DataPath_ALUhw_SHIFTER_HW_n469, DataPath_ALUhw_SHIFTER_HW_n468, 
      DataPath_ALUhw_SHIFTER_HW_n467, DataPath_ALUhw_SHIFTER_HW_n466, 
      DataPath_ALUhw_SHIFTER_HW_n460, DataPath_ALUhw_SHIFTER_HW_n459, 
      DataPath_ALUhw_SHIFTER_HW_n458, DataPath_ALUhw_SHIFTER_HW_n457, 
      DataPath_ALUhw_SHIFTER_HW_n456, DataPath_ALUhw_SHIFTER_HW_n455, 
      DataPath_ALUhw_SHIFTER_HW_n453, DataPath_ALUhw_SHIFTER_HW_n450, 
      DataPath_ALUhw_SHIFTER_HW_n445, DataPath_ALUhw_SHIFTER_HW_n443, 
      DataPath_ALUhw_SHIFTER_HW_n437, DataPath_ALUhw_SHIFTER_HW_n432, 
      DataPath_ALUhw_SHIFTER_HW_n430, DataPath_ALUhw_SHIFTER_HW_n424, 
      DataPath_ALUhw_SHIFTER_HW_n419, DataPath_ALUhw_SHIFTER_HW_n418, 
      DataPath_ALUhw_SHIFTER_HW_n417, DataPath_ALUhw_SHIFTER_HW_n411, 
      DataPath_ALUhw_SHIFTER_HW_n410, DataPath_ALUhw_SHIFTER_HW_n409, 
      DataPath_ALUhw_SHIFTER_HW_n408, DataPath_ALUhw_SHIFTER_HW_n407, 
      DataPath_ALUhw_SHIFTER_HW_n406, DataPath_ALUhw_SHIFTER_HW_n405, 
      DataPath_ALUhw_SHIFTER_HW_n403, DataPath_ALUhw_SHIFTER_HW_n397, 
      DataPath_ALUhw_SHIFTER_HW_n392, DataPath_ALUhw_SHIFTER_HW_n390, 
      DataPath_ALUhw_SHIFTER_HW_n385, DataPath_ALUhw_SHIFTER_HW_n380, 
      DataPath_ALUhw_SHIFTER_HW_n378, DataPath_ALUhw_SHIFTER_HW_n373, 
      DataPath_ALUhw_SHIFTER_HW_n367, DataPath_ALUhw_SHIFTER_HW_n360, 
      DataPath_ALUhw_SHIFTER_HW_n354, DataPath_ALUhw_SHIFTER_HW_n349, 
      DataPath_ALUhw_SHIFTER_HW_n345, DataPath_ALUhw_SHIFTER_HW_n344, 
      DataPath_ALUhw_SHIFTER_HW_n338, DataPath_ALUhw_SHIFTER_HW_n331, 
      DataPath_ALUhw_SHIFTER_HW_n324, DataPath_ALUhw_SHIFTER_HW_n317, 
      DataPath_ALUhw_SHIFTER_HW_n310, DataPath_ALUhw_SHIFTER_HW_n303, 
      DataPath_ALUhw_SHIFTER_HW_n296, DataPath_ALUhw_SHIFTER_HW_n289, 
      DataPath_ALUhw_SHIFTER_HW_n282, DataPath_ALUhw_SHIFTER_HW_n275, 
      DataPath_ALUhw_SHIFTER_HW_n269, DataPath_ALUhw_SHIFTER_HW_n268, 
      DataPath_ALUhw_SHIFTER_HW_n267, DataPath_ALUhw_SHIFTER_HW_n266, 
      DataPath_ALUhw_SHIFTER_HW_n265, DataPath_ALUhw_SHIFTER_HW_n264, 
      DataPath_ALUhw_SHIFTER_HW_n263, DataPath_ALUhw_SHIFTER_HW_n262, 
      DataPath_ALUhw_SHIFTER_HW_n260, DataPath_ALUhw_SHIFTER_HW_n250, 
      DataPath_ALUhw_SHIFTER_HW_n219, DataPath_ALUhw_SHIFTER_HW_n217, 
      DataPath_ALUhw_SHIFTER_HW_n216, DataPath_ALUhw_SHIFTER_HW_n215, 
      DataPath_ALUhw_SHIFTER_HW_n214, DataPath_ALUhw_SHIFTER_HW_n213, 
      DataPath_ALUhw_SHIFTER_HW_n212, DataPath_ALUhw_SHIFTER_HW_n211, 
      DataPath_ALUhw_SHIFTER_HW_n207, DataPath_ALUhw_SHIFTER_HW_n206, 
      DataPath_ALUhw_SHIFTER_HW_n205, DataPath_ALUhw_SHIFTER_HW_n204, 
      DataPath_ALUhw_SHIFTER_HW_n203, DataPath_ALUhw_SHIFTER_HW_n202, 
      DataPath_ALUhw_SHIFTER_HW_n201, DataPath_ALUhw_SHIFTER_HW_n200, 
      DataPath_ALUhw_SHIFTER_HW_n199, DataPath_ALUhw_SHIFTER_HW_n198, 
      DataPath_ALUhw_SHIFTER_HW_n197, DataPath_ALUhw_SHIFTER_HW_n196, 
      DataPath_ALUhw_SHIFTER_HW_n195, DataPath_ALUhw_SHIFTER_HW_n194, 
      DataPath_ALUhw_SHIFTER_HW_n193, DataPath_ALUhw_SHIFTER_HW_n192, 
      DataPath_ALUhw_SHIFTER_HW_n191, DataPath_ALUhw_SHIFTER_HW_n190, 
      DataPath_ALUhw_SHIFTER_HW_n189, DataPath_ALUhw_SHIFTER_HW_n188, 
      DataPath_ALUhw_SHIFTER_HW_n187, DataPath_ALUhw_SHIFTER_HW_n186, 
      DataPath_ALUhw_SHIFTER_HW_n185, DataPath_ALUhw_SHIFTER_HW_n184, 
      DataPath_ALUhw_SHIFTER_HW_n183, DataPath_ALUhw_SHIFTER_HW_n182, 
      DataPath_ALUhw_SHIFTER_HW_n181, DataPath_ALUhw_SHIFTER_HW_n180, 
      DataPath_ALUhw_SHIFTER_HW_n179, DataPath_ALUhw_SHIFTER_HW_n178, 
      DataPath_ALUhw_SHIFTER_HW_n177, DataPath_ALUhw_SHIFTER_HW_n176, 
      DataPath_ALUhw_SHIFTER_HW_n175, DataPath_ALUhw_SHIFTER_HW_n174, 
      DataPath_ALUhw_SHIFTER_HW_n173, DataPath_ALUhw_SHIFTER_HW_n172, 
      DataPath_ALUhw_SHIFTER_HW_n171, DataPath_ALUhw_SHIFTER_HW_n170, 
      DataPath_ALUhw_SHIFTER_HW_n169, DataPath_ALUhw_SHIFTER_HW_n168, 
      DataPath_ALUhw_SHIFTER_HW_n167, DataPath_ALUhw_SHIFTER_HW_n166, 
      DataPath_ALUhw_SHIFTER_HW_n165, DataPath_ALUhw_SHIFTER_HW_n164, 
      DataPath_ALUhw_SHIFTER_HW_n161, DataPath_ALUhw_SHIFTER_HW_n157, 
      DataPath_ALUhw_SHIFTER_HW_n156, DataPath_ALUhw_SHIFTER_HW_n155, 
      DataPath_ALUhw_SHIFTER_HW_n153, DataPath_ALUhw_SHIFTER_HW_n152, 
      DataPath_ALUhw_SHIFTER_HW_n151, DataPath_ALUhw_SHIFTER_HW_n150, 
      DataPath_ALUhw_SHIFTER_HW_n148, DataPath_ALUhw_SHIFTER_HW_n147, 
      DataPath_ALUhw_SHIFTER_HW_n146, DataPath_ALUhw_SHIFTER_HW_n145, 
      DataPath_ALUhw_SHIFTER_HW_n144, DataPath_ALUhw_SHIFTER_HW_n143, 
      DataPath_ALUhw_SHIFTER_HW_n142, DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n15, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n14, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n13, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n12, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n11, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n10, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n9, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n8, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n6, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n3, 
      DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n2, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_4_28_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_3_16_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_3_24_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_8_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_12_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_16_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_20_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_24_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_28_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_6_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_10_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_14_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_18_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_22_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_26_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_28_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_25_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_26_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_27_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_26_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_27_port, 
      DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_28_port, 
      DataPath_RF_POP_ADDRGEN_N61, DataPath_RF_POP_ADDRGEN_N60, 
      DataPath_RF_POP_ADDRGEN_N59, DataPath_RF_POP_ADDRGEN_N58, 
      DataPath_RF_POP_ADDRGEN_N57, DataPath_RF_POP_ADDRGEN_N56, 
      DataPath_RF_POP_ADDRGEN_N55, DataPath_RF_POP_ADDRGEN_N54, 
      DataPath_RF_POP_ADDRGEN_N53, DataPath_RF_POP_ADDRGEN_N52, 
      DataPath_RF_POP_ADDRGEN_N51, DataPath_RF_POP_ADDRGEN_N50, 
      DataPath_RF_POP_ADDRGEN_N49, DataPath_RF_POP_ADDRGEN_N48, 
      DataPath_RF_POP_ADDRGEN_N47, DataPath_RF_POP_ADDRGEN_N46, 
      DataPath_RF_POP_ADDRGEN_curr_state_0_port, 
      DataPath_RF_POP_ADDRGEN_curr_state_1_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_0_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_1_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_2_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_3_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_4_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_5_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_6_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_7_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_8_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_9_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_10_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_11_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_12_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_13_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_14_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_15_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_3_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_3_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_3_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_3_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_3_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_3_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_3_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_1_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_2_port, 
      DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_3_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_3_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_4_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_5_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_6_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_7_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_8_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_9_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_10_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_11_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_12_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_13_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_14_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_15_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_16_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_17_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_18_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_19_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_20_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_21_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_22_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_23_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_24_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_25_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_26_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_27_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_28_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_29_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_30_port, 
      DataPath_WRF_CUhw_sub_85_aco_carry_31_port, WS1_4_port, n200, n201, n202,
      n203, n204, n205, n207, n208, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
      n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
      n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n554, n555, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, 
      n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, 
      n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n692, n693, n694, n695, n696, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n950, n951, n952, n953, n954, n955, n956, 
      n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
      n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, 
      n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, 
      n993, n994, n995, n996, n997, n998, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
      n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
      n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, 
      n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, 
      n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, 
      n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, 
      n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, 
      n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
      n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
      n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, 
      n1136, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, 
      n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, 
      n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, 
      n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, 
      n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, 
      n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, 
      n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, 
      n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
      n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
      n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, 
      n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, 
      n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, 
      n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, 
      n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, 
      n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, 
      n1437, n1438, n1439, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1777, n1778, n1780, 
      n1781, n1782, n1783, n1785, n1786, n1787, n1788, n1789, n1790, n1791, 
      n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
      n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, 
      n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, 
      n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, 
      n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, 
      n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, 
      n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, 
      n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, 
      n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, 
      n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, 
      n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, 
      n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, 
      n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, 
      n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, 
      n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, 
      n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, 
      n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, 
      n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, 
      n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, 
      n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, 
      n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, 
      n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, 
      n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, 
      n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, 
      n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, 
      n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, 
      n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, 
      n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, 
      n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, 
      n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, 
      n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, 
      n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, 
      n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, 
      n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, 
      n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, 
      n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, 
      n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, 
      n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, 
      n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, 
      n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, 
      n2192, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, 
      n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, 
      n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, 
      n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, 
      n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, 
      n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
      n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, 
      n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, 
      n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, 
      n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, 
      n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, 
      n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, 
      n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, 
      n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
      n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, 
      n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, 
      n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, 
      n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, 
      n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, 
      n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, 
      n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, 
      n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, 
      n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, 
      n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, 
      n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, 
      n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, 
      n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
      n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, 
      n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, 
      n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, 
      n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, 
      n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
      n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, 
      n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, 
      n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, 
      n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, 
      n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, 
      n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, 
      n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, 
      n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, 
      n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, 
      n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, 
      n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, 
      n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, 
      n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, 
      n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
      n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
      n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
      n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
      n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
      n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
      n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
      n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
      n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
      n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, 
      n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, 
      n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
      n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
      n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, 
      n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
      n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
      n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
      n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
      n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
      n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
      n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
      n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
      n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
      n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
      n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
      n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
      n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
      n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
      n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
      n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
      n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, 
      n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
      n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, 
      n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
      n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
      n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, 
      n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, 
      n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
      n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
      n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
      n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
      n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
      n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, 
      n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
      n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, 
      n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, 
      n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, 
      n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, 
      n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, 
      n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, 
      n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, 
      n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, 
      n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, 
      n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, 
      n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, 
      n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, 
      n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, 
      n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, 
      n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, 
      n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, 
      n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, 
      n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, 
      n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, 
      n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, 
      n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, 
      n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, 
      n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
      n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, 
      n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
      n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, 
      n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
      n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
      n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
      n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, 
      n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, 
      n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, 
      n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, 
      n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, 
      n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, 
      n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, 
      n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, 
      n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, 
      n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, 
      n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, 
      n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, 
      n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, 
      n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, 
      n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, 
      n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, 
      n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, 
      n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, 
      n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, 
      n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, 
      n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, 
      n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, 
      n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, 
      n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, 
      n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, 
      n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, 
      n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, 
      n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, 
      n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, 
      n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, 
      n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, 
      n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
      n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, 
      n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, 
      n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, 
      n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, 
      n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
      n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, 
      n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, 
      n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4142, n4143, n4144, 
      n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, 
      n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, 
      n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, 
      n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, 
      n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, 
      n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, 
      n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, 
      n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, 
      n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
      n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, 
      n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, 
      n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, 
      n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
      n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, 
      n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, 
      n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, 
      n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, 
      n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, 
      n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, 
      n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, 
      n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, 
      n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, 
      n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, 
      n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, 
      n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
      n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, 
      n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, 
      n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, 
      n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, 
      n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, 
      n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, 
      n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, 
      n4465, n4466, n4467, n4468, n4470, n4471, n4472, n4474, n4475, n4476, 
      n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, 
      n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, 
      n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, 
      n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, 
      n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, 
      n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, 
      n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
      n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, 
      n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, 
      n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, 
      n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, 
      n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, 
      n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, 
      n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, 
      n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, 
      n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, 
      n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, 
      n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, 
      n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, 
      n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, 
      n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, 
      n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, 
      n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, 
      n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, 
      n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, 
      n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, 
      n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, 
      n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, 
      n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, 
      n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, 
      n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, 
      n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, 
      n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, 
      n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, 
      n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, 
      n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, 
      n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, 
      n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, 
      n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, 
      n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, 
      n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, 
      n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, 
      n4898, n4899, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, 
      n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, 
      n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, 
      n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, 
      n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, 
      n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, 
      n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, 
      n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, 
      n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, 
      n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, 
      n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, 
      n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, 
      n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, 
      n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, 
      n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, 
      n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, 
      n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, 
      n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, 
      n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, 
      n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, 
      n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, 
      n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, 
      n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, 
      n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, 
      n5139, n5140, n5141, n5142, n5143, n5145, n5146, n5147, n5148, n5149, 
      n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, 
      n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, 
      n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, 
      n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, 
      n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, 
      n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, 
      n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, 
      n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, 
      n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, 
      n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, 
      n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, 
      n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, 
      n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, 
      n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, 
      n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, 
      n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
      n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, 
      n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, 
      n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
      n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, 
      n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, 
      n5360, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, 
      n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, 
      n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, 
      n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, 
      n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, 
      n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, 
      n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, 
      n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, 
      n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, 
      n5451, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, 
      n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
      n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, 
      n5482, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, 
      n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, 
      n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, 
      n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, 
      n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, 
      n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, 
      n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, 
      n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, 
      n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, 
      n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, 
      n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, 
      n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, 
      n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, 
      n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, 
      n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, 
      n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, 
      n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, 
      n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, 
      n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
      n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, 
      n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, 
      n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, 
      n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
      n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, 
      n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, 
      n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
      n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5877, n5878, n5879, n5880, n5881, n5882, n5883, 
      n5884, n5885, n5886, n5887, n5889, n5890, n5891, n5892, n5893, n5894, 
      n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, 
      n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, 
      n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, 
      n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, 
      n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, 
      n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, 
      n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, 
      n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, 
      n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, 
      n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, 
      n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, 
      n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, 
      n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, 
      n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, 
      n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, 
      n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, 
      n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, 
      n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, 
      n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, 
      n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, 
      n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, 
      n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, 
      n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, 
      n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, 
      n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, 
      n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, 
      n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, 
      n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, 
      n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, 
      n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, 
      n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, 
      n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, 
      n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, 
      n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, 
      n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6244, n6245, 
      n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, 
      n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, 
      n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, 
      n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, 
      n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, 
      n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, 
      n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, 
      n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
      n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, 
      n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, 
      n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, 
      n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, 
      n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, 
      n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6384, n6385, n6386, 
      n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, 
      n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, 
      n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, 
      n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, 
      n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, 
      n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, 
      n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, 
      n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, 
      n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, 
      n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6486, n6487, 
      n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, 
      n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, 
      n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, 
      n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, 
      n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, 
      n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, 
      n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, 
      n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, 
      n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, 
      n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, 
      n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, 
      n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, 
      n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, 
      n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, 
      n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, 
      n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, 
      n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, 
      n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, 
      n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, 
      n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, 
      n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, 
      n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, 
      n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, 
      n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, 
      n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, 
      n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, 
      n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, 
      n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, 
      n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, 
      n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6786, n6787, n6788, 
      n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, 
      n6799, n6800, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, 
      n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, 
      n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, 
      n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, 
      n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, 
      n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, 
      n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, 
      n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, 
      n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, 
      n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, 
      n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, 
      n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, 
      n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, 
      n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, 
      n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, 
      n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, 
      n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, 
      n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, 
      n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, 
      n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, 
      n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, 
      n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, 
      n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, 
      n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, 
      n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, 
      n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, 
      n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7069, n7070, 
      n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, 
      n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, 
      n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, 
      n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, 
      n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, 
      n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, 
      n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, 
      n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, 
      n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, 
      n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, 
      n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, 
      n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, 
      n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, 
      n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, 
      n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, 
      n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7229, n7230, n7231, 
      n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, 
      n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, 
      n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, 
      n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, 
      n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, 
      n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, 
      n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, 
      n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, 
      n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, 
      n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, 
      n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, 
      n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, 
      n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, 
      n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, 
      n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7382, 
      n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, 
      n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, 
      n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, 
      n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, 
      n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, 
      n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, 
      n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, 
      n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, 
      n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, 
      n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, 
      n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, 
      n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, 
      n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, 
      n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, 
      n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, 
      n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, 
      n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, 
      n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, 
      n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, 
      n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, 
      n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, 
      n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, 
      n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, 
      n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, 
      n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, 
      n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, 
      n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, 
      n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, 
      n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, 
      n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, 
      n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, 
      n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, 
      n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, 
      n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, 
      n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, 
      n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, 
      n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, 
      n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, 
      n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, 
      n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, 
      n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, 
      n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, 
      n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, 
      n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, 
      n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, 
      n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, 
      n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, 
      n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, 
      n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, 
      n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, 
      n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, 
      n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, 
      n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, 
      n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, 
      n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, 
      n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, 
      n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, 
      n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, 
      n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, 
      n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, 
      n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, 
      n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, 
      n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, 
      n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, 
      n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, 
      n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, 
      n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, 
      n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, 
      n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, 
      n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, 
      n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, 
      n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, 
      n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, 
      n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, 
      n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, 
      n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, 
      n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, 
      n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, 
      n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, 
      n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, 
      n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, 
      n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, 
      n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, 
      n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, 
      n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, 
      n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, 
      n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, 
      n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, 
      n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, 
      n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, 
      n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, 
      n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, 
      n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, 
      n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, 
      n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, 
      n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, 
      n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, 
      n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, 
      n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, 
      n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, 
      n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, 
      n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, 
      n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, 
      n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, 
      n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, 
      n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, 
      n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, 
      n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, 
      n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, 
      n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, 
      n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, 
      n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, 
      n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, 
      n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, 
      n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, 
      n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, 
      n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, 
      n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, 
      n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, 
      n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, 
      n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, 
      n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, 
      n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, 
      n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, 
      n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, 
      n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, 
      n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, 
      n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, 
      n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, 
      n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, 
      n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, 
      n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, 
      n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, 
      n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, 
      n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, 
      n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, 
      n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, 
      n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, 
      n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, 
      n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, 
      n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, 
      n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, 
      n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, 
      n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, 
      n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, 
      n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, 
      n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, 
      n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, 
      n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, 
      n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, 
      n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, 
      n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, 
      n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, 
      n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, 
      n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, 
      n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, 
      n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, 
      n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, 
      n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, 
      n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, 
      n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, 
      n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, 
      n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, 
      n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, 
      n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, 
      n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, 
      n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, 
      n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, 
      n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, 
      n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, 
      n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, 
      n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, 
      n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, 
      n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, 
      n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, 
      n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, 
      n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, 
      n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, 
      n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, 
      n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, 
      n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, 
      n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, 
      n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, 
      n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, 
      n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, 
      n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, 
      n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, 
      n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, 
      n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, 
      n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, 
      n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, 
      n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, 
      n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, 
      n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, 
      n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, 
      n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, 
      n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, 
      n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, 
      n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, 
      n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, 
      n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, 
      n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, 
      n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, 
      n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, 
      n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, 
      n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, 
      n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, 
      n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, 
      n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, 
      n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, 
      n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, 
      n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, 
      n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, 
      n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, 
      n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, 
      n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, 
      n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, 
      n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, 
      n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, 
      n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, 
      n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, 
      n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, 
      n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, 
      n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, 
      n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, 
      n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, 
      n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, 
      n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, 
      n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, 
      n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, 
      n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, 
      n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, 
      n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, 
      n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, 
      n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, 
      n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, 
      n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, 
      n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, 
      n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, 
      n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, 
      n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, 
      n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, 
      n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, 
      n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, 
      n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, 
      n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, 
      n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, 
      n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, 
      n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, 
      n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, 
      n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, 
      n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, 
      n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, 
      n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, 
      n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, 
      n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, 
      n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, 
      n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, 
      n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, 
      n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, 
      n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, 
      n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, 
      n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, 
      n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, 
      n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, 
      n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, 
      n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, 
      n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, 
      n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, 
      n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, 
      n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, 
      n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, 
      n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, 
      n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, 
      n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, 
      n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, 
      n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, 
      n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, 
      n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, 
      n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, 
      n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, 
      n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, 
      n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, 
      n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, 
      n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, 
      n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, 
      n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, 
      n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, 
      n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, 
      n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, 
      n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, 
      n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, 
      n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, 
      n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, 
      n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, 
      n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, 
      n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, 
      n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, 
      n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, 
      n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, 
      n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, 
      n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, 
      n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, 
      n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, 
      n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, 
      n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, 
      n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, 
      n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, 
      n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, 
      n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, 
      n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, 
      n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, 
      n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, 
      n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, 
      n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, 
      n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, 
      n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, 
      n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, 
      n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, 
      n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, 
      n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, 
      n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, 
      n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, 
      n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, 
      n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, 
      n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, 
      n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, 
      n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, 
      n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, 
      n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, 
      n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, 
      n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, 
      n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, 
      n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, 
      n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, 
      n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, 
      n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, 
      n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, 
      n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, 
      n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, 
      n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, 
      n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, 
      n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, 
      n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, 
      n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, 
      n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, 
      n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, 
      n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, 
      n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, 
      n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, 
      n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, 
      n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, 
      n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, 
      n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, 
      n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, 
      n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, 
      n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, 
      n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, 
      n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, 
      n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, 
      n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, 
      n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, 
      n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, 
      n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, 
      n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, 
      n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, 
      n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, 
      n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, 
      n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, 
      n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, 
      n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, 
      n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, 
      n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, 
      n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, 
      n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, 
      n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, 
      n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, 
      n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, 
      n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, 
      n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, 
      n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, 
      n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, 
      n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, 
      n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, 
      n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, 
      n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, 
      n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, 
      n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, 
      n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, 
      n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, 
      n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, 
      n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, 
      n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, 
      n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, 
      n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, 
      n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, 
      n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, 
      n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, 
      n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, 
      n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, 
      n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, 
      n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, 
      n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, 
      n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, 
      n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, 
      n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, 
      n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, 
      n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, 
      n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, 
      n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, 
      n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, 
      n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, 
      n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, 
      n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, 
      n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, 
      n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, 
      n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, 
      n11398, n11399, n11400, n11431, n11432, n11433, n11434, n11435, n11436, 
      n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, 
      n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, 
      n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, 
      n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, 
      n11473, n11474, n11475, n11476, n11477, n11478, n11480, n11481, n11482, 
      n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, 
      n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, 
      n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, 
      n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, 
      n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, 
      n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, 
      n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, 
      n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, 
      n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, 
      n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, 
      n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, 
      DRAM_ADDRESS_1_port, n11582, DRAM_READNOTWRITE_port, n11584, n11585, 
      n11586, n11587, n11590, n11591, n11592, n11593, n11594, n11595, n11596, 
      n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, 
      n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, 
      n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, 
      n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, 
      n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, 
      n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, 
      n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, 
      n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, 
      n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, 
      n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, 
      n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, 
      n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, 
      n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, 
      n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, 
      n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, 
      n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, 
      n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, 
      n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, 
      n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, 
      n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, 
      n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, 
      n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, 
      n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, 
      n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, 
      n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, 
      n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, 
      n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, 
      n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, 
      n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, 
      n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, 
      n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, 
      n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, 
      n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, 
      n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, 
      n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, 
      n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, 
      n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, 
      n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, 
      n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, 
      n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, 
      n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, 
      n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, 
      n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, 
      n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, 
      n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, 
      n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, 
      n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, 
      n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, 
      n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, 
      n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, 
      n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, 
      n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, 
      n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, 
      n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, 
      n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, 
      n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, 
      n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, 
      n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, 
      n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, 
      n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, 
      n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, 
      n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, 
      n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, 
      n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, 
      n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, 
      n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, 
      n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, 
      n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, 
      n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, 
      n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, 
      n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, 
      n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, 
      n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, 
      n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, 
      n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, 
      n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, 
      n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, 
      n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, 
      n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, 
      n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, 
      n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, 
      n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, 
      n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, 
      n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, 
      n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, 
      n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, 
      n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, 
      n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, 
      n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, 
      n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, 
      n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, 
      n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, 
      n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, 
      n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, 
      n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, 
      n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, 
      n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, 
      n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, 
      n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, 
      n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, 
      n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, 
      n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, 
      n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, 
      n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, 
      n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, 
      n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, 
      n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, 
      n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, 
      n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, 
      n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, 
      n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, 
      n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, 
      n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, 
      n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, 
      n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, 
      n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, 
      n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, 
      n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, 
      n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, 
      n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, 
      n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, 
      n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, 
      n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, 
      n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, 
      n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, 
      n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, 
      n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, 
      n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, 
      n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, 
      n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, 
      n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, 
      n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, 
      n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, 
      n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, 
      n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, 
      n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, 
      n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, 
      n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, 
      n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, 
      n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, 
      n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, 
      n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, 
      n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, 
      n12884, n12885, n12886, n12887, RS2_4_port, n12889, n12890, n12891, 
      n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, 
      n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, 
      n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, 
      n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, 
      n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, 
      n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, 
      n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, 
      n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, 
      n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, 
      n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, 
      n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, 
      n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, 
      n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, 
      n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, 
      n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, 
      n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, 
      n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, 
      n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, 
      n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, 
      n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, 
      n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, 
      n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, 
      n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, 
      n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, 
      n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, 
      n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, 
      n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, 
      n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, 
      n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, 
      n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, 
      n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, 
      n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, 
      n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, 
      n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, 
      n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, 
      n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, 
      n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, 
      n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, 
      n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, 
      n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, 
      n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, 
      n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, 
      n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, 
      n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, 
      n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, 
      n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, 
      n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, 
      n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, 
      n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, 
      n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, 
      n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, 
      n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, 
      n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, 
      n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, 
      n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, 
      n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, 
      n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, 
      n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, 
      n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, 
      n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, 
      n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, 
      n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, 
      n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, 
      n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, 
      n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, 
      n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, 
      n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, 
      n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, 
      n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, 
      n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, 
      n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, 
      n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, 
      n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, 
      n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, 
      n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, 
      n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, 
      n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, 
      n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, 
      n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, 
      n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, 
      n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, 
      n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, 
      n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, 
      n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, 
      n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, 
      n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, 
      n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, 
      n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, 
      n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, 
      n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, 
      n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, 
      n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, 
      n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, 
      n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, 
      n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, 
      n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, 
      n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, 
      n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, 
      n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, 
      n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, 
      n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, 
      n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, 
      n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, 
      n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, 
      n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, 
      n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, 
      n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, 
      n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, 
      n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, 
      n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, 
      n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, 
      n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, 
      n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, 
      n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, 
      n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, 
      n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, 
      n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, 
      n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, 
      n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, 
      n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, 
      n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, 
      n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, 
      n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, 
      n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, 
      n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, 
      n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, 
      n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, 
      n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, 
      n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, 
      n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, 
      n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, 
      n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, 
      n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, 
      n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, 
      n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, 
      n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, 
      n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, 
      n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, 
      n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, 
      n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, 
      n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, 
      n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, 
      n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, 
      n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, 
      n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, 
      n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, 
      n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, 
      n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, 
      n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, 
      n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, 
      n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, 
      n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, 
      n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, 
      n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, 
      n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, 
      n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, 
      n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, 
      n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, 
      n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, 
      n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, 
      n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, 
      n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, 
      n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, 
      n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, 
      n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, 
      n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, 
      n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, 
      n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, 
      n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, 
      n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, 
      n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, 
      n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, 
      n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, 
      n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, 
      n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, 
      n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, 
      n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, 
      n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, 
      n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, 
      n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, 
      n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, 
      n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, 
      n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, 
      n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, 
      n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, 
      n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, 
      n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, 
      n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, 
      n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, 
      n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, 
      n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, 
      n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, 
      n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, 
      n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, 
      n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, 
      n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, 
      n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, 
      n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, 
      n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, 
      n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, 
      n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, 
      n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, 
      n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, 
      n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, 
      n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, 
      n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, 
      n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, 
      n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, 
      n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, 
      n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, 
      n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, 
      n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, 
      n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, 
      n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, 
      n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, 
      n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, 
      n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, 
      n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, 
      n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, 
      n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, 
      n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, 
      n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, 
      n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, 
      n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, 
      n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, 
      n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, 
      n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, 
      n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, 
      n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, 
      n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, 
      n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, 
      n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, 
      n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, 
      n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, 
      n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, 
      n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, 
      n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, 
      n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, 
      n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, 
      n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, 
      n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, 
      n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, 
      n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, 
      n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, 
      n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, 
      n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, 
      n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, 
      n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, 
      n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, 
      n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, 
      n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, 
      n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, 
      n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, 
      n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, 
      n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, 
      n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, 
      n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, 
      n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, 
      n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, 
      n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, 
      n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, 
      n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, 
      n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, 
      n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, 
      n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, 
      n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, 
      n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, 
      n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, 
      n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, 
      n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, 
      n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, 
      n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, 
      n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, 
      n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, 
      n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, 
      n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, 
      n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, 
      n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, 
      n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, 
      n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, 
      n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, 
      n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, 
      n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, 
      n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, 
      n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, 
      n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, 
      n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, 
      n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, 
      n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, 
      n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, 
      n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, 
      n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, 
      n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, 
      n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, 
      n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, 
      n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, 
      n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, 
      n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, 
      n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, 
      n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, 
      n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, 
      n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, 
      n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, 
      n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, 
      n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, 
      n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, 
      n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, 
      n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, 
      n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, 
      n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, 
      n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, 
      n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, 
      n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, 
      n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, 
      n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, 
      n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, 
      n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, 
      n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, 
      n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, 
      n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, 
      n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, 
      n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, 
      n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, 
      n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, 
      n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, 
      n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, 
      n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, 
      n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, 
      n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, 
      n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, 
      n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, 
      n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, 
      n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, 
      n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, 
      n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, 
      n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, 
      n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, 
      n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, 
      n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, 
      n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, 
      n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, 
      n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, 
      n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, 
      n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, 
      n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, 
      n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, 
      n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, 
      n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, 
      n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, 
      n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, 
      n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, 
      n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, 
      n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, 
      n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, 
      n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, 
      n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, 
      n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, 
      n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, 
      n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, 
      n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, 
      n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, 
      n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, 
      n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, 
      n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, 
      n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, 
      n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, 
      n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, 
      n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, 
      n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, 
      n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, 
      n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, 
      n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, 
      n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, 
      n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, 
      n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, 
      n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, 
      n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, 
      n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, 
      n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, 
      n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, 
      n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, 
      n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, 
      n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, 
      n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, 
      n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, 
      n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, 
      n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, 
      n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, 
      n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, 
      n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, 
      n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, 
      n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, 
      n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, 
      n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, 
      n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, 
      n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, 
      n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, 
      n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, 
      n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, 
      n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, 
      n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, 
      n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, 
      n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, 
      n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, 
      n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, 
      n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, 
      n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, 
      n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, 
      n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, 
      n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, 
      n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, 
      n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, 
      n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, 
      n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, 
      n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, 
      n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, 
      n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, 
      n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, 
      n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, 
      n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, 
      n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, 
      n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, 
      n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, 
      n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, 
      n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, 
      n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, 
      n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, 
      n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, 
      n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, 
      n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, 
      n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, 
      n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, 
      n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, 
      n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, 
      n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, 
      n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, 
      n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, 
      n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, 
      n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, 
      n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, 
      n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, 
      n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, 
      n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, 
      n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, 
      n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, 
      n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, 
      n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, 
      n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, 
      n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, 
      n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, 
      n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, 
      n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, 
      n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, 
      n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, 
      n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, 
      n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, 
      n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, 
      n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, 
      n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, 
      n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, 
      n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, 
      n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, 
      n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, 
      n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, 
      n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, 
      n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, 
      n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, 
      n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, 
      n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, 
      n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, 
      n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, 
      n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, 
      n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17148, n17149, 
      n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, 
      n17159, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, 
      n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, 
      n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, 
      n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, 
      n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, 
      n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, 
      n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, 
      n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, 
      n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, 
      n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, 
      n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, 
      n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, 
      n17268, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, 
      n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, 
      n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, 
      n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, 
      n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, 
      n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, 
      n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, 
      n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, 
      n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, 
      n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, 
      n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, 
      n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, 
      n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, 
      n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, 
      n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, 
      n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, 
      n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, 
      n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, 
      n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, 
      n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, 
      n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, 
      n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, 
      n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, 
      n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, 
      n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, 
      n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, 
      n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, 
      n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, 
      n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, 
      n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, 
      n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, 
      n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, 
      n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, 
      n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, 
      n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, 
      n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, 
      n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, 
      n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, 
      n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, 
      n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, 
      n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, 
      n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, 
      n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, 
      n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, 
      n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, 
      n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, 
      n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, 
      n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, 
      n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, 
      n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, 
      n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, 
      n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, 
      n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, 
      n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, 
      n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, 
      n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, 
      n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, 
      n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, 
      n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, 
      n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, 
      n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, 
      n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, 
      n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, 
      n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, 
      n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, 
      n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, 
      n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, 
      n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, 
      n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, 
      n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, 
      n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, 
      n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, 
      n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, 
      n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, 
      n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, 
      n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, 
      n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, 
      n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, 
      n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, 
      n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, 
      n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, 
      n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, 
      n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, 
      n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, 
      n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, 
      n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, 
      n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, 
      n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, 
      n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, 
      n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, 
      n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, 
      n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, 
      n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, 
      n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, 
      n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, 
      n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, 
      n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, 
      n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, 
      n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, 
      n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, 
      n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, 
      n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, 
      n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, 
      n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, 
      n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, 
      n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, 
      n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, 
      n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, 
      n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, 
      n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, 
      n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, 
      n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, 
      n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, 
      n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, 
      n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, 
      n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, 
      n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, 
      n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, 
      n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, 
      n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, 
      n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, 
      n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, 
      n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, 
      n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, 
      n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, 
      n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, 
      n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, 
      n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, 
      n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, 
      n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, 
      n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, 
      n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, 
      n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, 
      n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, 
      n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, 
      n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, 
      n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, 
      n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, 
      n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, 
      n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, 
      n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, 
      n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, 
      n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, 
      n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, 
      n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, 
      n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, 
      n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, 
      n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, 
      n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, 
      n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, 
      n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, 
      n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, 
      n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, 
      n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, 
      n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, 
      n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, 
      n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, 
      n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, 
      n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, 
      n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, 
      n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, 
      n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, 
      n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, 
      n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, 
      n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, 
      n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, 
      n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, 
      n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, 
      n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, 
      n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, 
      n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, 
      n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, 
      n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, 
      n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, 
      n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, 
      n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, 
      n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, 
      n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, 
      n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, 
      n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, 
      n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, 
      n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, 
      n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, 
      n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, 
      n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, 
      n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, 
      n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, 
      n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, 
      n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, 
      n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, 
      n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, 
      n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, 
      n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, 
      n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, 
      n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, 
      n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, 
      n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, 
      n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, 
      n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, 
      n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, 
      n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, 
      n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, 
      n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, 
      n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, 
      n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, 
      n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, 
      n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, 
      n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, 
      n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, 
      n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, 
      n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, 
      n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, 
      n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, 
      n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, 
      n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, 
      n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, 
      n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, 
      n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, 
      n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, 
      n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, 
      n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, 
      n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, 
      n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, 
      n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, 
      n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, 
      n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, 
      n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, 
      n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, 
      n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, 
      n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, 
      n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, 
      n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, 
      n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, 
      n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, 
      n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, 
      n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, 
      n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, 
      n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, 
      n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, 
      n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, 
      n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, 
      n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, 
      n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, 
      n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, 
      n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, 
      n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, 
      n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, 
      n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, 
      n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, 
      n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, 
      n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, 
      n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, 
      n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, 
      n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, 
      n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, 
      n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, 
      n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, 
      n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, 
      n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, 
      n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, 
      n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, 
      n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, 
      n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, 
      n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, 
      n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, 
      n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, 
      n_3780, n_3781, n_3782 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, DRAM_ADDRESS_0_port );
   DRAM_ISSUE <= DRAM_ISSUE_port;
   DRAM_READNOTWRITE <= DRAM_READNOTWRITE_port;
   DRAM_DATA_OUT <= ( DRAM_DATA_OUT_31_port, DRAM_DATA_OUT_30_port, 
      DRAM_DATA_OUT_29_port, DRAM_DATA_OUT_28_port, DRAM_DATA_OUT_27_port, 
      DRAM_DATA_OUT_26_port, DRAM_DATA_OUT_25_port, DRAM_DATA_OUT_24_port, 
      DRAM_DATA_OUT_23_port, DRAM_DATA_OUT_22_port, DRAM_DATA_OUT_21_port, 
      DRAM_DATA_OUT_20_port, DRAM_DATA_OUT_19_port, DRAM_DATA_OUT_18_port, 
      DRAM_DATA_OUT_17_port, DRAM_DATA_OUT_16_port, DRAM_DATA_OUT_15_port, 
      DRAM_DATA_OUT_14_port, DRAM_DATA_OUT_13_port, DRAM_DATA_OUT_12_port, 
      DRAM_DATA_OUT_11_port, DRAM_DATA_OUT_10_port, DRAM_DATA_OUT_9_port, 
      DRAM_DATA_OUT_8_port, DRAM_DATA_OUT_7_port, DRAM_DATA_OUT_6_port, 
      DRAM_DATA_OUT_5_port, DRAM_DATA_OUT_4_port, DRAM_DATA_OUT_3_port, 
      DRAM_DATA_OUT_2_port, DRAM_DATA_OUT_1_port, DRAM_DATA_OUT_0_port );
   DATA_SIZE <= ( DATA_SIZE_1_port, DATA_SIZE_0_port );
   DRAMRF_READNOTWRITE <= DRAMRF_READNOTWRITE_port;
   DATA_SIZE_RF <= ( X_Logic0_port, X_Logic0_port );
   OPCODE <= ( OPCODE_5_port, OPCODE_4_port, OPCODE_3_port, OPCODE_2_port, 
      OPCODE_1_port, OPCODE_0_port );
   RS2 <= ( RS2_4_port, RS2_4_port, RS2_4_port, RS2_4_port, RS2_4_port );
   WS1 <= ( WS1_4_port, WS1_4_port, WS1_4_port, WS1_4_port, WS1_4_port );
   IRO <= ( OPCODE_5_port, OPCODE_4_port, OPCODE_3_port, OPCODE_2_port, 
      OPCODE_1_port, OPCODE_0_port, IRO_25_port, IRO_24_port, IRO_23_port, 
      IRO_22_port, IRO_21_port, IRO_20_port, IRO_19_port, IRO_18_port, 
      IRO_17_port, IRO_16_port, IRO_15_port, IRO_14_port, IRO_13_port, 
      IRO_12_port, IRO_11_port, IRO_10_port, IRO_9_port, IRO_8_port, IRO_7_port
      , IRO_6_port, IRO_5_port, IRO_4_port, IRO_3_port, IRO_2_port, IRO_1_port,
      IRO_0_port );
   PCO <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   
   IRAM_ISSUE <= '1';
   X_Logic0_port <= '0';
   DIR_EN <= '0';
   DataPath_REG_A_Q_reg_3_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_3_port, QN => n_1000);
   DataPath_REG_A_Q_reg_5_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_5_port, QN => n_1001);
   DataPath_REG_A_Q_reg_11_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_11_port, QN => n_1002);
   DataPath_SETCMP_U11 : NAND3_X1 port map( A1 => n11483, A2 => n11484, A3 => 
                           i_SEL_LGET_1_port, ZN => DataPath_SETCMP_n4);
   DataPath_SETCMP_U10 : OAI33_X1 port map( A1 => n11484, A2 => 
                           i_SEL_LGET_1_port, A3 => i_SEL_LGET_0_port, B1 => 
                           n11483, B2 => i_SEL_LGET_1_port, B3 => n11591, ZN =>
                           DataPath_SETCMP_n7);
   DataPath_SETCMP_U9 : NAND3_X1 port map( A1 => DataPath_i_LGET_0_port, A2 => 
                           n11484, A3 => i_SEL_LGET_0_port, ZN => 
                           DataPath_SETCMP_n9);
   DataPath_LDSTR_U119 : NAND3_X1 port map( A1 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_1_port, A2 =>
                           n11578, A3 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_0_port, ZN =>
                           DataPath_LDSTR_n86);
   DataPath_LDSTR_U118 : NAND3_X1 port map( A1 => DRAM_DATA_OUT_7_port, A2 => 
                           n11480, A3 => n11578, ZN => DataPath_LDSTR_n62);
   DataPath_LDSTR_U117 : NAND3_X1 port map( A1 => DataPath_LDSTR_n61, A2 => 
                           DataPath_LDSTR_n62, A3 => DataPath_LDSTR_n63, ZN => 
                           DRAM_DATA_OUT_23_port);
   DataPath_LDSTR_U69 : NOR4_X2 port map( A1 => DataPath_LDSTR_n69, A2 => 
                           DataPath_LDSTR_n80, A3 => DataPath_LDSTR_n83, A4 => 
                           DataPath_LDSTR_n84, ZN => DataPath_LDSTR_n68);
   DataPath_WRB1_Q_reg_0_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB1_0_port, QN => n_1003);
   DataPath_WRB1_Q_reg_1_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB1_1_port, QN => n_1004);
   DataPath_WRB1_Q_reg_2_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB1_2_port, QN => n_1005);
   DataPath_WRB1_Q_reg_3_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB1_3_port, QN => n_1006);
   DataPath_WRB1_Q_reg_4_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB1_4_port, QN => n_1007);
   DataPath_RF_DEC_U49 : NAND3_X1 port map( A1 => i_ADD_WB_1_port, A2 => 
                           i_ADD_WB_0_port, A3 => i_ADD_WB_2_port, ZN => 
                           DataPath_RF_DEC_n14);
   DataPath_RF_DEC_U48 : NAND3_X1 port map( A1 => i_ADD_WB_1_port, A2 => n11598
                           , A3 => i_ADD_WB_2_port, ZN => DataPath_RF_DEC_n13);
   DataPath_RF_DEC_U47 : NAND3_X1 port map( A1 => i_ADD_WB_0_port, A2 => n11599
                           , A3 => i_ADD_WB_2_port, ZN => DataPath_RF_DEC_n12);
   DataPath_RF_DEC_U46 : NAND3_X1 port map( A1 => n11598, A2 => n11599, A3 => 
                           i_ADD_WB_2_port, ZN => DataPath_RF_DEC_n11);
   DataPath_RF_DEC_U45 : NAND3_X1 port map( A1 => i_ADD_WB_0_port, A2 => n11600
                           , A3 => i_ADD_WB_1_port, ZN => DataPath_RF_DEC_n10);
   DataPath_RF_DEC_U44 : NAND3_X1 port map( A1 => n11598, A2 => n11600, A3 => 
                           i_ADD_WB_1_port, ZN => DataPath_RF_DEC_n9);
   DataPath_RF_DEC_U43 : NAND3_X1 port map( A1 => n11599, A2 => n11600, A3 => 
                           i_ADD_WB_0_port, ZN => DataPath_RF_DEC_n8);
   DataPath_RF_DEC_U42 : NAND3_X1 port map( A1 => n11599, A2 => n11600, A3 => 
                           n11598, ZN => DataPath_RF_DEC_n7);
   DataPath_RF_SPILLADDR_ENC_U40 : NAND3_X1 port map( A1 => n11437, A2 => 
                           n11438, A3 => DataPath_RF_SPILLADDR_ENC_n25, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n24);
   DataPath_RF_SPILLADDR_ENC_U39 : NAND3_X1 port map( A1 => n11439, A2 => 
                           n11440, A3 => n11442, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n15);
   DataPath_ALUhw_BWISE_U101 : OAI22_X2 port map( A1 => i_ALU_OP_4_port, A2 => 
                           n4129, B1 => n11540, B2 => n11500, ZN => 
                           DataPath_ALUhw_BWISE_n72);
   DataPath_ALUhw_BWISE_U96 : OAI21_X2 port map( B1 => i_ALU_OP_4_port, B2 => 
                           n4133, A => n11500, ZN => DataPath_ALUhw_BWISE_n71);
   DataPath_RF_BLOCKi_87_Q_reg_0_inst : DFF_X1 port map( D => n11347, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2528_port, QN => 
                           n_1008);
   DataPath_RF_BLOCKi_87_Q_reg_1_inst : DFF_X1 port map( D => n11346, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2529_port, QN => 
                           n_1009);
   DataPath_RF_BLOCKi_87_Q_reg_2_inst : DFF_X1 port map( D => n11345, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2530_port, QN => 
                           n_1010);
   DataPath_RF_BLOCKi_87_Q_reg_3_inst : DFF_X1 port map( D => n11344, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2531_port, QN => 
                           n_1011);
   DataPath_RF_BLOCKi_87_Q_reg_4_inst : DFF_X1 port map( D => n11343, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2532_port, QN => 
                           n_1012);
   DataPath_RF_BLOCKi_87_Q_reg_5_inst : DFF_X1 port map( D => n11342, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2533_port, QN => 
                           n_1013);
   DataPath_RF_BLOCKi_87_Q_reg_6_inst : DFF_X1 port map( D => n11341, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2534_port, QN => 
                           n_1014);
   DataPath_RF_BLOCKi_87_Q_reg_7_inst : DFF_X1 port map( D => n11340, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2535_port, QN => 
                           n_1015);
   DataPath_RF_BLOCKi_87_Q_reg_8_inst : DFF_X1 port map( D => n11339, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2536_port, QN => 
                           n_1016);
   DataPath_RF_BLOCKi_87_Q_reg_9_inst : DFF_X1 port map( D => n11338, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2537_port, QN => 
                           n_1017);
   DataPath_RF_BLOCKi_87_Q_reg_10_inst : DFF_X1 port map( D => n11337, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2538_port, QN 
                           => n_1018);
   DataPath_RF_BLOCKi_87_Q_reg_11_inst : DFF_X1 port map( D => n11336, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2539_port, QN 
                           => n_1019);
   DataPath_RF_BLOCKi_87_Q_reg_12_inst : DFF_X1 port map( D => n11335, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2540_port, QN 
                           => n_1020);
   DataPath_RF_BLOCKi_87_Q_reg_13_inst : DFF_X1 port map( D => n11334, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2541_port, QN 
                           => n_1021);
   DataPath_RF_BLOCKi_87_Q_reg_14_inst : DFF_X1 port map( D => n11333, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2542_port, QN 
                           => n_1022);
   DataPath_RF_BLOCKi_87_Q_reg_15_inst : DFF_X1 port map( D => n11332, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2543_port, QN 
                           => n_1023);
   DataPath_RF_BLOCKi_87_Q_reg_16_inst : DFF_X1 port map( D => n11331, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2544_port, QN 
                           => n_1024);
   DataPath_RF_BLOCKi_87_Q_reg_17_inst : DFF_X1 port map( D => n11330, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2545_port, QN 
                           => n_1025);
   DataPath_RF_BLOCKi_87_Q_reg_18_inst : DFF_X1 port map( D => n11329, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2546_port, QN 
                           => n_1026);
   DataPath_RF_BLOCKi_87_Q_reg_19_inst : DFF_X1 port map( D => n11328, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2547_port, QN 
                           => n_1027);
   DataPath_RF_BLOCKi_87_Q_reg_20_inst : DFF_X1 port map( D => n11327, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2548_port, QN 
                           => n_1028);
   DataPath_RF_BLOCKi_87_Q_reg_21_inst : DFF_X1 port map( D => n11326, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2549_port, QN 
                           => n_1029);
   DataPath_RF_BLOCKi_87_Q_reg_22_inst : DFF_X1 port map( D => n11325, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2550_port, QN 
                           => n_1030);
   DataPath_RF_BLOCKi_87_Q_reg_23_inst : DFF_X1 port map( D => n11324, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2551_port, QN 
                           => n_1031);
   DataPath_RF_BLOCKi_87_Q_reg_24_inst : DFF_X1 port map( D => n11323, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2552_port, QN 
                           => n_1032);
   DataPath_RF_BLOCKi_87_Q_reg_25_inst : DFF_X1 port map( D => n11322, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2553_port, QN 
                           => n_1033);
   DataPath_RF_BLOCKi_87_Q_reg_26_inst : DFF_X1 port map( D => n11321, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2554_port, QN 
                           => n_1034);
   DataPath_RF_BLOCKi_87_Q_reg_27_inst : DFF_X1 port map( D => n11320, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2555_port, QN 
                           => n_1035);
   DataPath_RF_BLOCKi_87_Q_reg_28_inst : DFF_X1 port map( D => n11319, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2556_port, QN 
                           => n_1036);
   DataPath_RF_BLOCKi_87_Q_reg_29_inst : DFF_X1 port map( D => n11318, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2557_port, QN 
                           => n_1037);
   DataPath_RF_BLOCKi_87_Q_reg_30_inst : DFF_X1 port map( D => n11317, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2558_port, QN 
                           => n_1038);
   DataPath_RF_BLOCKi_87_Q_reg_31_inst : DFF_X1 port map( D => n11316, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2559_port, QN 
                           => n_1039);
   DataPath_RF_BLOCKi_86_Q_reg_0_inst : DFF_X1 port map( D => n11315, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2496_port, QN => 
                           n_1040);
   DataPath_RF_BLOCKi_86_Q_reg_1_inst : DFF_X1 port map( D => n11314, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2497_port, QN => 
                           n_1041);
   DataPath_RF_BLOCKi_86_Q_reg_2_inst : DFF_X1 port map( D => n11313, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2498_port, QN => 
                           n_1042);
   DataPath_RF_BLOCKi_86_Q_reg_3_inst : DFF_X1 port map( D => n11312, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2499_port, QN => 
                           n_1043);
   DataPath_RF_BLOCKi_86_Q_reg_4_inst : DFF_X1 port map( D => n11311, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2500_port, QN => 
                           n_1044);
   DataPath_RF_BLOCKi_86_Q_reg_5_inst : DFF_X1 port map( D => n11310, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2501_port, QN => 
                           n_1045);
   DataPath_RF_BLOCKi_86_Q_reg_6_inst : DFF_X1 port map( D => n11309, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2502_port, QN => 
                           n_1046);
   DataPath_RF_BLOCKi_86_Q_reg_7_inst : DFF_X1 port map( D => n11308, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2503_port, QN => 
                           n_1047);
   DataPath_RF_BLOCKi_86_Q_reg_8_inst : DFF_X1 port map( D => n11307, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2504_port, QN => 
                           n_1048);
   DataPath_RF_BLOCKi_86_Q_reg_9_inst : DFF_X1 port map( D => n11306, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2505_port, QN => 
                           n_1049);
   DataPath_RF_BLOCKi_86_Q_reg_10_inst : DFF_X1 port map( D => n11305, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2506_port, QN 
                           => n_1050);
   DataPath_RF_BLOCKi_86_Q_reg_11_inst : DFF_X1 port map( D => n11304, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2507_port, QN 
                           => n_1051);
   DataPath_RF_BLOCKi_86_Q_reg_12_inst : DFF_X1 port map( D => n11303, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2508_port, QN 
                           => n_1052);
   DataPath_RF_BLOCKi_86_Q_reg_13_inst : DFF_X1 port map( D => n11302, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2509_port, QN 
                           => n_1053);
   DataPath_RF_BLOCKi_86_Q_reg_14_inst : DFF_X1 port map( D => n11301, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2510_port, QN 
                           => n_1054);
   DataPath_RF_BLOCKi_86_Q_reg_15_inst : DFF_X1 port map( D => n11300, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2511_port, QN 
                           => n_1055);
   DataPath_RF_BLOCKi_86_Q_reg_16_inst : DFF_X1 port map( D => n11299, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2512_port, QN 
                           => n_1056);
   DataPath_RF_BLOCKi_86_Q_reg_17_inst : DFF_X1 port map( D => n11298, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2513_port, QN 
                           => n_1057);
   DataPath_RF_BLOCKi_86_Q_reg_18_inst : DFF_X1 port map( D => n11297, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2514_port, QN 
                           => n_1058);
   DataPath_RF_BLOCKi_86_Q_reg_19_inst : DFF_X1 port map( D => n11296, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2515_port, QN 
                           => n_1059);
   DataPath_RF_BLOCKi_86_Q_reg_20_inst : DFF_X1 port map( D => n11295, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2516_port, QN 
                           => n_1060);
   DataPath_RF_BLOCKi_86_Q_reg_21_inst : DFF_X1 port map( D => n11294, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2517_port, QN 
                           => n_1061);
   DataPath_RF_BLOCKi_86_Q_reg_22_inst : DFF_X1 port map( D => n11293, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2518_port, QN 
                           => n_1062);
   DataPath_RF_BLOCKi_86_Q_reg_23_inst : DFF_X1 port map( D => n11292, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2519_port, QN 
                           => n_1063);
   DataPath_RF_BLOCKi_86_Q_reg_24_inst : DFF_X1 port map( D => n11291, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2520_port, QN 
                           => n_1064);
   DataPath_RF_BLOCKi_86_Q_reg_25_inst : DFF_X1 port map( D => n11290, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2521_port, QN 
                           => n_1065);
   DataPath_RF_BLOCKi_86_Q_reg_26_inst : DFF_X1 port map( D => n11289, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2522_port, QN 
                           => n_1066);
   DataPath_RF_BLOCKi_86_Q_reg_27_inst : DFF_X1 port map( D => n11288, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2523_port, QN 
                           => n_1067);
   DataPath_RF_BLOCKi_86_Q_reg_28_inst : DFF_X1 port map( D => n11287, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2524_port, QN 
                           => n_1068);
   DataPath_RF_BLOCKi_86_Q_reg_29_inst : DFF_X1 port map( D => n11286, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2525_port, QN 
                           => n_1069);
   DataPath_RF_BLOCKi_86_Q_reg_30_inst : DFF_X1 port map( D => n11285, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2526_port, QN 
                           => n_1070);
   DataPath_RF_BLOCKi_86_Q_reg_31_inst : DFF_X1 port map( D => n11284, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2527_port, QN 
                           => n_1071);
   DataPath_RF_BLOCKi_85_Q_reg_0_inst : DFF_X1 port map( D => n11283, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2464_port, QN => 
                           n_1072);
   DataPath_RF_BLOCKi_85_Q_reg_1_inst : DFF_X1 port map( D => n11282, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2465_port, QN => 
                           n_1073);
   DataPath_RF_BLOCKi_85_Q_reg_2_inst : DFF_X1 port map( D => n11281, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2466_port, QN => 
                           n_1074);
   DataPath_RF_BLOCKi_85_Q_reg_3_inst : DFF_X1 port map( D => n11280, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2467_port, QN => 
                           n_1075);
   DataPath_RF_BLOCKi_85_Q_reg_4_inst : DFF_X1 port map( D => n11279, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2468_port, QN => 
                           n_1076);
   DataPath_RF_BLOCKi_85_Q_reg_5_inst : DFF_X1 port map( D => n11278, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2469_port, QN => 
                           n_1077);
   DataPath_RF_BLOCKi_85_Q_reg_6_inst : DFF_X1 port map( D => n11277, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2470_port, QN => 
                           n_1078);
   DataPath_RF_BLOCKi_85_Q_reg_7_inst : DFF_X1 port map( D => n11276, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2471_port, QN => 
                           n_1079);
   DataPath_RF_BLOCKi_85_Q_reg_8_inst : DFF_X1 port map( D => n11275, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2472_port, QN => 
                           n_1080);
   DataPath_RF_BLOCKi_85_Q_reg_9_inst : DFF_X1 port map( D => n11274, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2473_port, QN => 
                           n_1081);
   DataPath_RF_BLOCKi_85_Q_reg_10_inst : DFF_X1 port map( D => n11273, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2474_port, QN 
                           => n_1082);
   DataPath_RF_BLOCKi_85_Q_reg_11_inst : DFF_X1 port map( D => n11272, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2475_port, QN 
                           => n_1083);
   DataPath_RF_BLOCKi_85_Q_reg_12_inst : DFF_X1 port map( D => n11271, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2476_port, QN 
                           => n_1084);
   DataPath_RF_BLOCKi_85_Q_reg_13_inst : DFF_X1 port map( D => n11270, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2477_port, QN 
                           => n_1085);
   DataPath_RF_BLOCKi_85_Q_reg_14_inst : DFF_X1 port map( D => n11269, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2478_port, QN 
                           => n_1086);
   DataPath_RF_BLOCKi_85_Q_reg_15_inst : DFF_X1 port map( D => n11268, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2479_port, QN 
                           => n_1087);
   DataPath_RF_BLOCKi_85_Q_reg_16_inst : DFF_X1 port map( D => n11267, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2480_port, QN 
                           => n_1088);
   DataPath_RF_BLOCKi_85_Q_reg_17_inst : DFF_X1 port map( D => n11266, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2481_port, QN 
                           => n_1089);
   DataPath_RF_BLOCKi_85_Q_reg_18_inst : DFF_X1 port map( D => n11265, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2482_port, QN 
                           => n_1090);
   DataPath_RF_BLOCKi_85_Q_reg_19_inst : DFF_X1 port map( D => n11264, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2483_port, QN 
                           => n_1091);
   DataPath_RF_BLOCKi_85_Q_reg_20_inst : DFF_X1 port map( D => n11263, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2484_port, QN 
                           => n_1092);
   DataPath_RF_BLOCKi_85_Q_reg_21_inst : DFF_X1 port map( D => n11262, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2485_port, QN 
                           => n_1093);
   DataPath_RF_BLOCKi_85_Q_reg_22_inst : DFF_X1 port map( D => n11261, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2486_port, QN 
                           => n_1094);
   DataPath_RF_BLOCKi_85_Q_reg_23_inst : DFF_X1 port map( D => n11260, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2487_port, QN 
                           => n_1095);
   DataPath_RF_BLOCKi_85_Q_reg_24_inst : DFF_X1 port map( D => n11259, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2488_port, QN 
                           => n_1096);
   DataPath_RF_BLOCKi_85_Q_reg_25_inst : DFF_X1 port map( D => n11258, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2489_port, QN 
                           => n_1097);
   DataPath_RF_BLOCKi_85_Q_reg_26_inst : DFF_X1 port map( D => n11257, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2490_port, QN 
                           => n_1098);
   DataPath_RF_BLOCKi_85_Q_reg_27_inst : DFF_X1 port map( D => n11256, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2491_port, QN 
                           => n_1099);
   DataPath_RF_BLOCKi_85_Q_reg_28_inst : DFF_X1 port map( D => n11255, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2492_port, QN 
                           => n_1100);
   DataPath_RF_BLOCKi_85_Q_reg_29_inst : DFF_X1 port map( D => n11254, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2493_port, QN 
                           => n_1101);
   DataPath_RF_BLOCKi_85_Q_reg_30_inst : DFF_X1 port map( D => n11253, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2494_port, QN 
                           => n_1102);
   DataPath_RF_BLOCKi_85_Q_reg_31_inst : DFF_X1 port map( D => n11252, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2495_port, QN 
                           => n_1103);
   DataPath_RF_BLOCKi_84_Q_reg_0_inst : DFF_X1 port map( D => n11251, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2432_port, QN => 
                           n_1104);
   DataPath_RF_BLOCKi_84_Q_reg_1_inst : DFF_X1 port map( D => n11250, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2433_port, QN => 
                           n_1105);
   DataPath_RF_BLOCKi_84_Q_reg_2_inst : DFF_X1 port map( D => n11249, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2434_port, QN => 
                           n_1106);
   DataPath_RF_BLOCKi_84_Q_reg_3_inst : DFF_X1 port map( D => n11248, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2435_port, QN => 
                           n_1107);
   DataPath_RF_BLOCKi_84_Q_reg_4_inst : DFF_X1 port map( D => n11247, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2436_port, QN => 
                           n_1108);
   DataPath_RF_BLOCKi_84_Q_reg_5_inst : DFF_X1 port map( D => n11246, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2437_port, QN => 
                           n_1109);
   DataPath_RF_BLOCKi_84_Q_reg_6_inst : DFF_X1 port map( D => n11245, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2438_port, QN => 
                           n_1110);
   DataPath_RF_BLOCKi_84_Q_reg_7_inst : DFF_X1 port map( D => n11244, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2439_port, QN => 
                           n_1111);
   DataPath_RF_BLOCKi_84_Q_reg_8_inst : DFF_X1 port map( D => n11243, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2440_port, QN => 
                           n_1112);
   DataPath_RF_BLOCKi_84_Q_reg_9_inst : DFF_X1 port map( D => n11242, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2441_port, QN => 
                           n_1113);
   DataPath_RF_BLOCKi_84_Q_reg_10_inst : DFF_X1 port map( D => n11241, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2442_port, QN 
                           => n_1114);
   DataPath_RF_BLOCKi_84_Q_reg_11_inst : DFF_X1 port map( D => n11240, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2443_port, QN 
                           => n_1115);
   DataPath_RF_BLOCKi_84_Q_reg_12_inst : DFF_X1 port map( D => n11239, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2444_port, QN 
                           => n_1116);
   DataPath_RF_BLOCKi_84_Q_reg_13_inst : DFF_X1 port map( D => n11238, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2445_port, QN 
                           => n_1117);
   DataPath_RF_BLOCKi_84_Q_reg_14_inst : DFF_X1 port map( D => n11237, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2446_port, QN 
                           => n_1118);
   DataPath_RF_BLOCKi_84_Q_reg_15_inst : DFF_X1 port map( D => n11236, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2447_port, QN 
                           => n_1119);
   DataPath_RF_BLOCKi_84_Q_reg_16_inst : DFF_X1 port map( D => n11235, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2448_port, QN 
                           => n_1120);
   DataPath_RF_BLOCKi_84_Q_reg_17_inst : DFF_X1 port map( D => n11234, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2449_port, QN 
                           => n_1121);
   DataPath_RF_BLOCKi_84_Q_reg_18_inst : DFF_X1 port map( D => n11233, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2450_port, QN 
                           => n_1122);
   DataPath_RF_BLOCKi_84_Q_reg_19_inst : DFF_X1 port map( D => n11232, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2451_port, QN 
                           => n_1123);
   DataPath_RF_BLOCKi_84_Q_reg_20_inst : DFF_X1 port map( D => n11231, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2452_port, QN 
                           => n_1124);
   DataPath_RF_BLOCKi_84_Q_reg_21_inst : DFF_X1 port map( D => n11230, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2453_port, QN 
                           => n_1125);
   DataPath_RF_BLOCKi_84_Q_reg_22_inst : DFF_X1 port map( D => n11229, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2454_port, QN 
                           => n_1126);
   DataPath_RF_BLOCKi_84_Q_reg_23_inst : DFF_X1 port map( D => n11228, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2455_port, QN 
                           => n_1127);
   DataPath_RF_BLOCKi_84_Q_reg_24_inst : DFF_X1 port map( D => n11227, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2456_port, QN 
                           => n_1128);
   DataPath_RF_BLOCKi_84_Q_reg_25_inst : DFF_X1 port map( D => n11226, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2457_port, QN 
                           => n_1129);
   DataPath_RF_BLOCKi_84_Q_reg_26_inst : DFF_X1 port map( D => n11225, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2458_port, QN 
                           => n_1130);
   DataPath_RF_BLOCKi_84_Q_reg_27_inst : DFF_X1 port map( D => n11224, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2459_port, QN 
                           => n_1131);
   DataPath_RF_BLOCKi_84_Q_reg_28_inst : DFF_X1 port map( D => n11223, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2460_port, QN 
                           => n_1132);
   DataPath_RF_BLOCKi_84_Q_reg_29_inst : DFF_X1 port map( D => n11222, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2461_port, QN 
                           => n_1133);
   DataPath_RF_BLOCKi_84_Q_reg_30_inst : DFF_X1 port map( D => n11221, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2462_port, QN 
                           => n_1134);
   DataPath_RF_BLOCKi_84_Q_reg_31_inst : DFF_X1 port map( D => n11220, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2463_port, QN 
                           => n_1135);
   DataPath_RF_BLOCKi_83_Q_reg_0_inst : DFF_X1 port map( D => n11219, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2400_port, QN => 
                           n_1136);
   DataPath_RF_BLOCKi_83_Q_reg_1_inst : DFF_X1 port map( D => n11218, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2401_port, QN => 
                           n_1137);
   DataPath_RF_BLOCKi_83_Q_reg_2_inst : DFF_X1 port map( D => n11217, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2402_port, QN => 
                           n_1138);
   DataPath_RF_BLOCKi_83_Q_reg_3_inst : DFF_X1 port map( D => n11216, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2403_port, QN => 
                           n_1139);
   DataPath_RF_BLOCKi_83_Q_reg_4_inst : DFF_X1 port map( D => n11215, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2404_port, QN => 
                           n_1140);
   DataPath_RF_BLOCKi_83_Q_reg_5_inst : DFF_X1 port map( D => n11214, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2405_port, QN => 
                           n_1141);
   DataPath_RF_BLOCKi_83_Q_reg_6_inst : DFF_X1 port map( D => n11213, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2406_port, QN => 
                           n_1142);
   DataPath_RF_BLOCKi_83_Q_reg_7_inst : DFF_X1 port map( D => n11212, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2407_port, QN => 
                           n_1143);
   DataPath_RF_BLOCKi_83_Q_reg_8_inst : DFF_X1 port map( D => n11211, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2408_port, QN => 
                           n_1144);
   DataPath_RF_BLOCKi_83_Q_reg_9_inst : DFF_X1 port map( D => n11210, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2409_port, QN => 
                           n_1145);
   DataPath_RF_BLOCKi_83_Q_reg_10_inst : DFF_X1 port map( D => n11209, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2410_port, QN 
                           => n_1146);
   DataPath_RF_BLOCKi_83_Q_reg_11_inst : DFF_X1 port map( D => n11208, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2411_port, QN 
                           => n_1147);
   DataPath_RF_BLOCKi_83_Q_reg_12_inst : DFF_X1 port map( D => n11207, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2412_port, QN 
                           => n_1148);
   DataPath_RF_BLOCKi_83_Q_reg_13_inst : DFF_X1 port map( D => n11206, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2413_port, QN 
                           => n_1149);
   DataPath_RF_BLOCKi_83_Q_reg_14_inst : DFF_X1 port map( D => n11205, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2414_port, QN 
                           => n_1150);
   DataPath_RF_BLOCKi_83_Q_reg_15_inst : DFF_X1 port map( D => n11204, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2415_port, QN 
                           => n_1151);
   DataPath_RF_BLOCKi_83_Q_reg_16_inst : DFF_X1 port map( D => n11203, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2416_port, QN 
                           => n_1152);
   DataPath_RF_BLOCKi_83_Q_reg_17_inst : DFF_X1 port map( D => n11202, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2417_port, QN 
                           => n_1153);
   DataPath_RF_BLOCKi_83_Q_reg_18_inst : DFF_X1 port map( D => n11201, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2418_port, QN 
                           => n_1154);
   DataPath_RF_BLOCKi_83_Q_reg_19_inst : DFF_X1 port map( D => n11200, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2419_port, QN 
                           => n_1155);
   DataPath_RF_BLOCKi_83_Q_reg_20_inst : DFF_X1 port map( D => n11199, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2420_port, QN 
                           => n_1156);
   DataPath_RF_BLOCKi_83_Q_reg_21_inst : DFF_X1 port map( D => n11198, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2421_port, QN 
                           => n_1157);
   DataPath_RF_BLOCKi_83_Q_reg_22_inst : DFF_X1 port map( D => n11197, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2422_port, QN 
                           => n_1158);
   DataPath_RF_BLOCKi_83_Q_reg_23_inst : DFF_X1 port map( D => n11196, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2423_port, QN 
                           => n_1159);
   DataPath_RF_BLOCKi_83_Q_reg_24_inst : DFF_X1 port map( D => n11195, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2424_port, QN 
                           => n_1160);
   DataPath_RF_BLOCKi_83_Q_reg_25_inst : DFF_X1 port map( D => n11194, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2425_port, QN 
                           => n_1161);
   DataPath_RF_BLOCKi_83_Q_reg_26_inst : DFF_X1 port map( D => n11193, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2426_port, QN 
                           => n_1162);
   DataPath_RF_BLOCKi_83_Q_reg_27_inst : DFF_X1 port map( D => n11192, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2427_port, QN 
                           => n_1163);
   DataPath_RF_BLOCKi_83_Q_reg_28_inst : DFF_X1 port map( D => n11191, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2428_port, QN 
                           => n_1164);
   DataPath_RF_BLOCKi_83_Q_reg_29_inst : DFF_X1 port map( D => n11190, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2429_port, QN 
                           => n_1165);
   DataPath_RF_BLOCKi_83_Q_reg_30_inst : DFF_X1 port map( D => n11189, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2430_port, QN 
                           => n_1166);
   DataPath_RF_BLOCKi_83_Q_reg_31_inst : DFF_X1 port map( D => n11188, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2431_port, QN 
                           => n_1167);
   DataPath_RF_BLOCKi_82_Q_reg_0_inst : DFF_X1 port map( D => n11187, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2368_port, QN => 
                           n_1168);
   DataPath_RF_BLOCKi_82_Q_reg_1_inst : DFF_X1 port map( D => n11186, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2369_port, QN => 
                           n_1169);
   DataPath_RF_BLOCKi_82_Q_reg_2_inst : DFF_X1 port map( D => n11185, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2370_port, QN => 
                           n_1170);
   DataPath_RF_BLOCKi_82_Q_reg_3_inst : DFF_X1 port map( D => n11184, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2371_port, QN => 
                           n_1171);
   DataPath_RF_BLOCKi_82_Q_reg_4_inst : DFF_X1 port map( D => n11183, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2372_port, QN => 
                           n_1172);
   DataPath_RF_BLOCKi_82_Q_reg_5_inst : DFF_X1 port map( D => n11182, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2373_port, QN => 
                           n_1173);
   DataPath_RF_BLOCKi_82_Q_reg_6_inst : DFF_X1 port map( D => n11181, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2374_port, QN => 
                           n_1174);
   DataPath_RF_BLOCKi_82_Q_reg_7_inst : DFF_X1 port map( D => n11180, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2375_port, QN => 
                           n_1175);
   DataPath_RF_BLOCKi_82_Q_reg_8_inst : DFF_X1 port map( D => n11179, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2376_port, QN => 
                           n_1176);
   DataPath_RF_BLOCKi_82_Q_reg_9_inst : DFF_X1 port map( D => n11178, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2377_port, QN => 
                           n_1177);
   DataPath_RF_BLOCKi_82_Q_reg_10_inst : DFF_X1 port map( D => n11177, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2378_port, QN 
                           => n_1178);
   DataPath_RF_BLOCKi_82_Q_reg_11_inst : DFF_X1 port map( D => n11176, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2379_port, QN 
                           => n_1179);
   DataPath_RF_BLOCKi_82_Q_reg_12_inst : DFF_X1 port map( D => n11175, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2380_port, QN 
                           => n_1180);
   DataPath_RF_BLOCKi_82_Q_reg_13_inst : DFF_X1 port map( D => n11174, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2381_port, QN 
                           => n_1181);
   DataPath_RF_BLOCKi_82_Q_reg_14_inst : DFF_X1 port map( D => n11173, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2382_port, QN 
                           => n_1182);
   DataPath_RF_BLOCKi_82_Q_reg_15_inst : DFF_X1 port map( D => n11172, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2383_port, QN 
                           => n_1183);
   DataPath_RF_BLOCKi_82_Q_reg_16_inst : DFF_X1 port map( D => n11171, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2384_port, QN 
                           => n_1184);
   DataPath_RF_BLOCKi_82_Q_reg_17_inst : DFF_X1 port map( D => n11170, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2385_port, QN 
                           => n_1185);
   DataPath_RF_BLOCKi_82_Q_reg_18_inst : DFF_X1 port map( D => n11169, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2386_port, QN 
                           => n_1186);
   DataPath_RF_BLOCKi_82_Q_reg_19_inst : DFF_X1 port map( D => n11168, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2387_port, QN 
                           => n_1187);
   DataPath_RF_BLOCKi_82_Q_reg_20_inst : DFF_X1 port map( D => n11167, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2388_port, QN 
                           => n_1188);
   DataPath_RF_BLOCKi_82_Q_reg_21_inst : DFF_X1 port map( D => n11166, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2389_port, QN 
                           => n_1189);
   DataPath_RF_BLOCKi_82_Q_reg_22_inst : DFF_X1 port map( D => n11165, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2390_port, QN 
                           => n_1190);
   DataPath_RF_BLOCKi_82_Q_reg_23_inst : DFF_X1 port map( D => n11164, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2391_port, QN 
                           => n_1191);
   DataPath_RF_BLOCKi_82_Q_reg_24_inst : DFF_X1 port map( D => n11163, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2392_port, QN 
                           => n_1192);
   DataPath_RF_BLOCKi_82_Q_reg_25_inst : DFF_X1 port map( D => n11162, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2393_port, QN 
                           => n_1193);
   DataPath_RF_BLOCKi_82_Q_reg_26_inst : DFF_X1 port map( D => n11161, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2394_port, QN 
                           => n_1194);
   DataPath_RF_BLOCKi_82_Q_reg_27_inst : DFF_X1 port map( D => n11160, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2395_port, QN 
                           => n_1195);
   DataPath_RF_BLOCKi_82_Q_reg_28_inst : DFF_X1 port map( D => n11159, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2396_port, QN 
                           => n_1196);
   DataPath_RF_BLOCKi_82_Q_reg_29_inst : DFF_X1 port map( D => n11158, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2397_port, QN 
                           => n_1197);
   DataPath_RF_BLOCKi_82_Q_reg_30_inst : DFF_X1 port map( D => n11157, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2398_port, QN 
                           => n_1198);
   DataPath_RF_BLOCKi_82_Q_reg_31_inst : DFF_X1 port map( D => n11156, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2399_port, QN 
                           => n_1199);
   DataPath_RF_BLOCKi_81_Q_reg_0_inst : DFF_X1 port map( D => n11155, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2336_port, QN => 
                           n_1200);
   DataPath_RF_BLOCKi_81_Q_reg_1_inst : DFF_X1 port map( D => n11154, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2337_port, QN => 
                           n_1201);
   DataPath_RF_BLOCKi_81_Q_reg_2_inst : DFF_X1 port map( D => n11153, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2338_port, QN => 
                           n_1202);
   DataPath_RF_BLOCKi_81_Q_reg_3_inst : DFF_X1 port map( D => n11152, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2339_port, QN => 
                           n_1203);
   DataPath_RF_BLOCKi_81_Q_reg_4_inst : DFF_X1 port map( D => n11151, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2340_port, QN => 
                           n_1204);
   DataPath_RF_BLOCKi_81_Q_reg_5_inst : DFF_X1 port map( D => n11150, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2341_port, QN => 
                           n_1205);
   DataPath_RF_BLOCKi_81_Q_reg_6_inst : DFF_X1 port map( D => n11149, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2342_port, QN => 
                           n_1206);
   DataPath_RF_BLOCKi_81_Q_reg_7_inst : DFF_X1 port map( D => n11148, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2343_port, QN => 
                           n_1207);
   DataPath_RF_BLOCKi_81_Q_reg_8_inst : DFF_X1 port map( D => n11147, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2344_port, QN => 
                           n_1208);
   DataPath_RF_BLOCKi_81_Q_reg_9_inst : DFF_X1 port map( D => n11146, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2345_port, QN => 
                           n_1209);
   DataPath_RF_BLOCKi_81_Q_reg_10_inst : DFF_X1 port map( D => n11145, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2346_port, QN 
                           => n_1210);
   DataPath_RF_BLOCKi_81_Q_reg_11_inst : DFF_X1 port map( D => n11144, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2347_port, QN 
                           => n_1211);
   DataPath_RF_BLOCKi_81_Q_reg_12_inst : DFF_X1 port map( D => n11143, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2348_port, QN 
                           => n_1212);
   DataPath_RF_BLOCKi_81_Q_reg_13_inst : DFF_X1 port map( D => n11142, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2349_port, QN 
                           => n_1213);
   DataPath_RF_BLOCKi_81_Q_reg_14_inst : DFF_X1 port map( D => n11141, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2350_port, QN 
                           => n_1214);
   DataPath_RF_BLOCKi_81_Q_reg_15_inst : DFF_X1 port map( D => n11140, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2351_port, QN 
                           => n_1215);
   DataPath_RF_BLOCKi_81_Q_reg_16_inst : DFF_X1 port map( D => n11139, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2352_port, QN 
                           => n_1216);
   DataPath_RF_BLOCKi_81_Q_reg_17_inst : DFF_X1 port map( D => n11138, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2353_port, QN 
                           => n_1217);
   DataPath_RF_BLOCKi_81_Q_reg_18_inst : DFF_X1 port map( D => n11137, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2354_port, QN 
                           => n_1218);
   DataPath_RF_BLOCKi_81_Q_reg_19_inst : DFF_X1 port map( D => n11136, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2355_port, QN 
                           => n_1219);
   DataPath_RF_BLOCKi_81_Q_reg_20_inst : DFF_X1 port map( D => n11135, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2356_port, QN 
                           => n_1220);
   DataPath_RF_BLOCKi_81_Q_reg_21_inst : DFF_X1 port map( D => n11134, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2357_port, QN 
                           => n_1221);
   DataPath_RF_BLOCKi_81_Q_reg_22_inst : DFF_X1 port map( D => n11133, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2358_port, QN 
                           => n_1222);
   DataPath_RF_BLOCKi_81_Q_reg_23_inst : DFF_X1 port map( D => n11132, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2359_port, QN 
                           => n_1223);
   DataPath_RF_BLOCKi_81_Q_reg_24_inst : DFF_X1 port map( D => n11131, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2360_port, QN 
                           => n_1224);
   DataPath_RF_BLOCKi_81_Q_reg_25_inst : DFF_X1 port map( D => n11130, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2361_port, QN 
                           => n_1225);
   DataPath_RF_BLOCKi_81_Q_reg_26_inst : DFF_X1 port map( D => n11129, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2362_port, QN 
                           => n_1226);
   DataPath_RF_BLOCKi_81_Q_reg_27_inst : DFF_X1 port map( D => n11128, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2363_port, QN 
                           => n_1227);
   DataPath_RF_BLOCKi_81_Q_reg_28_inst : DFF_X1 port map( D => n11127, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2364_port, QN 
                           => n_1228);
   DataPath_RF_BLOCKi_81_Q_reg_29_inst : DFF_X1 port map( D => n11126, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2365_port, QN 
                           => n_1229);
   DataPath_RF_BLOCKi_81_Q_reg_30_inst : DFF_X1 port map( D => n11125, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2366_port, QN 
                           => n_1230);
   DataPath_RF_BLOCKi_81_Q_reg_31_inst : DFF_X1 port map( D => n11124, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2367_port, QN 
                           => n_1231);
   DataPath_RF_BLOCKi_80_Q_reg_0_inst : DFF_X1 port map( D => n11123, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2304_port, QN => 
                           n_1232);
   DataPath_RF_BLOCKi_80_Q_reg_1_inst : DFF_X1 port map( D => n11122, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2305_port, QN => 
                           n_1233);
   DataPath_RF_BLOCKi_80_Q_reg_2_inst : DFF_X1 port map( D => n11121, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2306_port, QN => 
                           n_1234);
   DataPath_RF_BLOCKi_80_Q_reg_3_inst : DFF_X1 port map( D => n11120, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2307_port, QN => 
                           n_1235);
   DataPath_RF_BLOCKi_80_Q_reg_4_inst : DFF_X1 port map( D => n11119, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2308_port, QN => 
                           n_1236);
   DataPath_RF_BLOCKi_80_Q_reg_5_inst : DFF_X1 port map( D => n11118, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2309_port, QN => 
                           n_1237);
   DataPath_RF_BLOCKi_80_Q_reg_6_inst : DFF_X1 port map( D => n11117, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2310_port, QN => 
                           n_1238);
   DataPath_RF_BLOCKi_80_Q_reg_7_inst : DFF_X1 port map( D => n11116, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2311_port, QN => 
                           n_1239);
   DataPath_RF_BLOCKi_80_Q_reg_8_inst : DFF_X1 port map( D => n11115, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2312_port, QN => 
                           n_1240);
   DataPath_RF_BLOCKi_80_Q_reg_9_inst : DFF_X1 port map( D => n11114, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2313_port, QN => 
                           n_1241);
   DataPath_RF_BLOCKi_80_Q_reg_10_inst : DFF_X1 port map( D => n11113, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2314_port, QN 
                           => n_1242);
   DataPath_RF_BLOCKi_80_Q_reg_11_inst : DFF_X1 port map( D => n11112, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2315_port, QN 
                           => n_1243);
   DataPath_RF_BLOCKi_80_Q_reg_12_inst : DFF_X1 port map( D => n11111, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2316_port, QN 
                           => n_1244);
   DataPath_RF_BLOCKi_80_Q_reg_13_inst : DFF_X1 port map( D => n11110, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2317_port, QN 
                           => n_1245);
   DataPath_RF_BLOCKi_80_Q_reg_14_inst : DFF_X1 port map( D => n11109, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2318_port, QN 
                           => n_1246);
   DataPath_RF_BLOCKi_80_Q_reg_15_inst : DFF_X1 port map( D => n11108, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2319_port, QN 
                           => n_1247);
   DataPath_RF_BLOCKi_80_Q_reg_16_inst : DFF_X1 port map( D => n11107, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2320_port, QN 
                           => n_1248);
   DataPath_RF_BLOCKi_80_Q_reg_17_inst : DFF_X1 port map( D => n11106, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2321_port, QN 
                           => n_1249);
   DataPath_RF_BLOCKi_80_Q_reg_18_inst : DFF_X1 port map( D => n11105, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2322_port, QN 
                           => n_1250);
   DataPath_RF_BLOCKi_80_Q_reg_19_inst : DFF_X1 port map( D => n11104, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2323_port, QN 
                           => n_1251);
   DataPath_RF_BLOCKi_80_Q_reg_20_inst : DFF_X1 port map( D => n11103, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2324_port, QN 
                           => n_1252);
   DataPath_RF_BLOCKi_80_Q_reg_21_inst : DFF_X1 port map( D => n11102, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2325_port, QN 
                           => n_1253);
   DataPath_RF_BLOCKi_80_Q_reg_22_inst : DFF_X1 port map( D => n11101, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2326_port, QN 
                           => n_1254);
   DataPath_RF_BLOCKi_80_Q_reg_23_inst : DFF_X1 port map( D => n11100, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2327_port, QN 
                           => n_1255);
   DataPath_RF_BLOCKi_80_Q_reg_24_inst : DFF_X1 port map( D => n11099, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2328_port, QN 
                           => n_1256);
   DataPath_RF_BLOCKi_80_Q_reg_25_inst : DFF_X1 port map( D => n11098, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2329_port, QN 
                           => n_1257);
   DataPath_RF_BLOCKi_80_Q_reg_26_inst : DFF_X1 port map( D => n11097, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2330_port, QN 
                           => n_1258);
   DataPath_RF_BLOCKi_80_Q_reg_27_inst : DFF_X1 port map( D => n11096, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2331_port, QN 
                           => n_1259);
   DataPath_RF_BLOCKi_80_Q_reg_28_inst : DFF_X1 port map( D => n11095, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2332_port, QN 
                           => n_1260);
   DataPath_RF_BLOCKi_80_Q_reg_29_inst : DFF_X1 port map( D => n11094, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2333_port, QN 
                           => n_1261);
   DataPath_RF_BLOCKi_80_Q_reg_30_inst : DFF_X1 port map( D => n11093, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2334_port, QN 
                           => n_1262);
   DataPath_RF_BLOCKi_80_Q_reg_31_inst : DFF_X1 port map( D => n11092, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2335_port, QN 
                           => n_1263);
   DataPath_RF_BLOCKi_79_Q_reg_0_inst : DFF_X1 port map( D => n11091, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2272_port, QN => 
                           n_1264);
   DataPath_RF_BLOCKi_79_Q_reg_1_inst : DFF_X1 port map( D => n11090, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2273_port, QN => 
                           n_1265);
   DataPath_RF_BLOCKi_79_Q_reg_2_inst : DFF_X1 port map( D => n11089, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2274_port, QN => 
                           n_1266);
   DataPath_RF_BLOCKi_79_Q_reg_3_inst : DFF_X1 port map( D => n11088, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2275_port, QN => 
                           n_1267);
   DataPath_RF_BLOCKi_79_Q_reg_4_inst : DFF_X1 port map( D => n11087, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2276_port, QN => 
                           n_1268);
   DataPath_RF_BLOCKi_79_Q_reg_5_inst : DFF_X1 port map( D => n11086, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2277_port, QN => 
                           n_1269);
   DataPath_RF_BLOCKi_79_Q_reg_6_inst : DFF_X1 port map( D => n11085, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2278_port, QN => 
                           n_1270);
   DataPath_RF_BLOCKi_79_Q_reg_7_inst : DFF_X1 port map( D => n11084, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2279_port, QN => 
                           n_1271);
   DataPath_RF_BLOCKi_79_Q_reg_8_inst : DFF_X1 port map( D => n11083, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2280_port, QN => 
                           n_1272);
   DataPath_RF_BLOCKi_79_Q_reg_9_inst : DFF_X1 port map( D => n11082, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2281_port, QN => 
                           n_1273);
   DataPath_RF_BLOCKi_79_Q_reg_10_inst : DFF_X1 port map( D => n11081, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2282_port, QN 
                           => n_1274);
   DataPath_RF_BLOCKi_79_Q_reg_11_inst : DFF_X1 port map( D => n11080, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2283_port, QN 
                           => n_1275);
   DataPath_RF_BLOCKi_79_Q_reg_12_inst : DFF_X1 port map( D => n11079, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2284_port, QN 
                           => n_1276);
   DataPath_RF_BLOCKi_79_Q_reg_13_inst : DFF_X1 port map( D => n11078, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2285_port, QN 
                           => n_1277);
   DataPath_RF_BLOCKi_79_Q_reg_14_inst : DFF_X1 port map( D => n11077, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2286_port, QN 
                           => n_1278);
   DataPath_RF_BLOCKi_79_Q_reg_15_inst : DFF_X1 port map( D => n11076, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2287_port, QN 
                           => n_1279);
   DataPath_RF_BLOCKi_79_Q_reg_16_inst : DFF_X1 port map( D => n11075, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2288_port, QN 
                           => n_1280);
   DataPath_RF_BLOCKi_79_Q_reg_17_inst : DFF_X1 port map( D => n11074, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2289_port, QN 
                           => n_1281);
   DataPath_RF_BLOCKi_79_Q_reg_18_inst : DFF_X1 port map( D => n11073, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2290_port, QN 
                           => n_1282);
   DataPath_RF_BLOCKi_79_Q_reg_19_inst : DFF_X1 port map( D => n11072, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2291_port, QN 
                           => n_1283);
   DataPath_RF_BLOCKi_79_Q_reg_20_inst : DFF_X1 port map( D => n11071, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2292_port, QN 
                           => n_1284);
   DataPath_RF_BLOCKi_79_Q_reg_21_inst : DFF_X1 port map( D => n11070, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2293_port, QN 
                           => n_1285);
   DataPath_RF_BLOCKi_79_Q_reg_22_inst : DFF_X1 port map( D => n11069, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2294_port, QN 
                           => n_1286);
   DataPath_RF_BLOCKi_79_Q_reg_23_inst : DFF_X1 port map( D => n11068, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2295_port, QN 
                           => n_1287);
   DataPath_RF_BLOCKi_79_Q_reg_24_inst : DFF_X1 port map( D => n11067, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2296_port, QN 
                           => n_1288);
   DataPath_RF_BLOCKi_79_Q_reg_25_inst : DFF_X1 port map( D => n11066, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2297_port, QN 
                           => n_1289);
   DataPath_RF_BLOCKi_79_Q_reg_26_inst : DFF_X1 port map( D => n11065, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2298_port, QN 
                           => n_1290);
   DataPath_RF_BLOCKi_79_Q_reg_27_inst : DFF_X1 port map( D => n11064, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2299_port, QN 
                           => n_1291);
   DataPath_RF_BLOCKi_79_Q_reg_28_inst : DFF_X1 port map( D => n11063, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2300_port, QN 
                           => n_1292);
   DataPath_RF_BLOCKi_79_Q_reg_29_inst : DFF_X1 port map( D => n11062, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2301_port, QN 
                           => n_1293);
   DataPath_RF_BLOCKi_79_Q_reg_30_inst : DFF_X1 port map( D => n11061, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2302_port, QN 
                           => n_1294);
   DataPath_RF_BLOCKi_79_Q_reg_31_inst : DFF_X1 port map( D => n11060, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2303_port, QN 
                           => n_1295);
   DataPath_RF_BLOCKi_78_Q_reg_0_inst : DFF_X1 port map( D => n11059, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2240_port, QN => 
                           n_1296);
   DataPath_RF_BLOCKi_78_Q_reg_1_inst : DFF_X1 port map( D => n11058, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2241_port, QN => 
                           n_1297);
   DataPath_RF_BLOCKi_78_Q_reg_2_inst : DFF_X1 port map( D => n11057, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2242_port, QN => 
                           n_1298);
   DataPath_RF_BLOCKi_78_Q_reg_3_inst : DFF_X1 port map( D => n11056, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2243_port, QN => 
                           n_1299);
   DataPath_RF_BLOCKi_78_Q_reg_4_inst : DFF_X1 port map( D => n11055, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2244_port, QN => 
                           n_1300);
   DataPath_RF_BLOCKi_78_Q_reg_5_inst : DFF_X1 port map( D => n11054, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2245_port, QN => 
                           n_1301);
   DataPath_RF_BLOCKi_78_Q_reg_6_inst : DFF_X1 port map( D => n11053, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2246_port, QN => 
                           n_1302);
   DataPath_RF_BLOCKi_78_Q_reg_7_inst : DFF_X1 port map( D => n11052, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2247_port, QN => 
                           n_1303);
   DataPath_RF_BLOCKi_78_Q_reg_8_inst : DFF_X1 port map( D => n11051, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2248_port, QN => 
                           n_1304);
   DataPath_RF_BLOCKi_78_Q_reg_9_inst : DFF_X1 port map( D => n11050, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2249_port, QN => 
                           n_1305);
   DataPath_RF_BLOCKi_78_Q_reg_10_inst : DFF_X1 port map( D => n11049, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2250_port, QN 
                           => n_1306);
   DataPath_RF_BLOCKi_78_Q_reg_11_inst : DFF_X1 port map( D => n11048, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2251_port, QN 
                           => n_1307);
   DataPath_RF_BLOCKi_78_Q_reg_12_inst : DFF_X1 port map( D => n11047, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2252_port, QN 
                           => n_1308);
   DataPath_RF_BLOCKi_78_Q_reg_13_inst : DFF_X1 port map( D => n11046, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2253_port, QN 
                           => n_1309);
   DataPath_RF_BLOCKi_78_Q_reg_14_inst : DFF_X1 port map( D => n11045, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2254_port, QN 
                           => n_1310);
   DataPath_RF_BLOCKi_78_Q_reg_15_inst : DFF_X1 port map( D => n11044, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2255_port, QN 
                           => n_1311);
   DataPath_RF_BLOCKi_78_Q_reg_16_inst : DFF_X1 port map( D => n11043, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2256_port, QN 
                           => n_1312);
   DataPath_RF_BLOCKi_78_Q_reg_17_inst : DFF_X1 port map( D => n11042, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2257_port, QN 
                           => n_1313);
   DataPath_RF_BLOCKi_78_Q_reg_18_inst : DFF_X1 port map( D => n11041, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2258_port, QN 
                           => n_1314);
   DataPath_RF_BLOCKi_78_Q_reg_19_inst : DFF_X1 port map( D => n11040, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2259_port, QN 
                           => n_1315);
   DataPath_RF_BLOCKi_78_Q_reg_20_inst : DFF_X1 port map( D => n11039, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2260_port, QN 
                           => n_1316);
   DataPath_RF_BLOCKi_78_Q_reg_21_inst : DFF_X1 port map( D => n11038, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2261_port, QN 
                           => n_1317);
   DataPath_RF_BLOCKi_78_Q_reg_22_inst : DFF_X1 port map( D => n11037, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2262_port, QN 
                           => n_1318);
   DataPath_RF_BLOCKi_78_Q_reg_23_inst : DFF_X1 port map( D => n11036, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2263_port, QN 
                           => n_1319);
   DataPath_RF_BLOCKi_78_Q_reg_24_inst : DFF_X1 port map( D => n11035, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2264_port, QN 
                           => n_1320);
   DataPath_RF_BLOCKi_78_Q_reg_25_inst : DFF_X1 port map( D => n11034, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2265_port, QN 
                           => n_1321);
   DataPath_RF_BLOCKi_78_Q_reg_26_inst : DFF_X1 port map( D => n11033, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2266_port, QN 
                           => n_1322);
   DataPath_RF_BLOCKi_78_Q_reg_27_inst : DFF_X1 port map( D => n11032, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2267_port, QN 
                           => n_1323);
   DataPath_RF_BLOCKi_78_Q_reg_28_inst : DFF_X1 port map( D => n11031, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2268_port, QN 
                           => n_1324);
   DataPath_RF_BLOCKi_78_Q_reg_29_inst : DFF_X1 port map( D => n11030, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2269_port, QN 
                           => n_1325);
   DataPath_RF_BLOCKi_78_Q_reg_30_inst : DFF_X1 port map( D => n11029, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2270_port, QN 
                           => n_1326);
   DataPath_RF_BLOCKi_78_Q_reg_31_inst : DFF_X1 port map( D => n11028, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2271_port, QN 
                           => n_1327);
   DataPath_RF_BLOCKi_77_Q_reg_0_inst : DFF_X1 port map( D => n11027, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2208_port, QN => 
                           n_1328);
   DataPath_RF_BLOCKi_77_Q_reg_1_inst : DFF_X1 port map( D => n11026, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2209_port, QN => 
                           n_1329);
   DataPath_RF_BLOCKi_77_Q_reg_2_inst : DFF_X1 port map( D => n11025, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2210_port, QN => 
                           n_1330);
   DataPath_RF_BLOCKi_77_Q_reg_3_inst : DFF_X1 port map( D => n11024, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2211_port, QN => 
                           n_1331);
   DataPath_RF_BLOCKi_77_Q_reg_4_inst : DFF_X1 port map( D => n11023, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2212_port, QN => 
                           n_1332);
   DataPath_RF_BLOCKi_77_Q_reg_5_inst : DFF_X1 port map( D => n11022, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2213_port, QN => 
                           n_1333);
   DataPath_RF_BLOCKi_77_Q_reg_6_inst : DFF_X1 port map( D => n11021, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2214_port, QN => 
                           n_1334);
   DataPath_RF_BLOCKi_77_Q_reg_7_inst : DFF_X1 port map( D => n11020, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2215_port, QN => 
                           n_1335);
   DataPath_RF_BLOCKi_77_Q_reg_8_inst : DFF_X1 port map( D => n11019, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2216_port, QN => 
                           n_1336);
   DataPath_RF_BLOCKi_77_Q_reg_9_inst : DFF_X1 port map( D => n11018, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2217_port, QN => 
                           n_1337);
   DataPath_RF_BLOCKi_77_Q_reg_10_inst : DFF_X1 port map( D => n11017, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2218_port, QN 
                           => n_1338);
   DataPath_RF_BLOCKi_77_Q_reg_11_inst : DFF_X1 port map( D => n11016, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2219_port, QN 
                           => n_1339);
   DataPath_RF_BLOCKi_77_Q_reg_12_inst : DFF_X1 port map( D => n11015, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2220_port, QN 
                           => n_1340);
   DataPath_RF_BLOCKi_77_Q_reg_13_inst : DFF_X1 port map( D => n11014, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2221_port, QN 
                           => n_1341);
   DataPath_RF_BLOCKi_77_Q_reg_14_inst : DFF_X1 port map( D => n11013, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2222_port, QN 
                           => n_1342);
   DataPath_RF_BLOCKi_77_Q_reg_15_inst : DFF_X1 port map( D => n11012, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2223_port, QN 
                           => n_1343);
   DataPath_RF_BLOCKi_77_Q_reg_16_inst : DFF_X1 port map( D => n11011, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2224_port, QN 
                           => n_1344);
   DataPath_RF_BLOCKi_77_Q_reg_17_inst : DFF_X1 port map( D => n11010, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2225_port, QN 
                           => n_1345);
   DataPath_RF_BLOCKi_77_Q_reg_18_inst : DFF_X1 port map( D => n11009, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2226_port, QN 
                           => n_1346);
   DataPath_RF_BLOCKi_77_Q_reg_19_inst : DFF_X1 port map( D => n11008, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2227_port, QN 
                           => n_1347);
   DataPath_RF_BLOCKi_77_Q_reg_20_inst : DFF_X1 port map( D => n11007, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2228_port, QN 
                           => n_1348);
   DataPath_RF_BLOCKi_77_Q_reg_21_inst : DFF_X1 port map( D => n11006, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2229_port, QN 
                           => n_1349);
   DataPath_RF_BLOCKi_77_Q_reg_22_inst : DFF_X1 port map( D => n11005, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2230_port, QN 
                           => n_1350);
   DataPath_RF_BLOCKi_77_Q_reg_23_inst : DFF_X1 port map( D => n11004, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2231_port, QN 
                           => n_1351);
   DataPath_RF_BLOCKi_77_Q_reg_24_inst : DFF_X1 port map( D => n11003, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2232_port, QN 
                           => n_1352);
   DataPath_RF_BLOCKi_77_Q_reg_25_inst : DFF_X1 port map( D => n11002, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2233_port, QN 
                           => n_1353);
   DataPath_RF_BLOCKi_77_Q_reg_26_inst : DFF_X1 port map( D => n11001, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2234_port, QN 
                           => n_1354);
   DataPath_RF_BLOCKi_77_Q_reg_27_inst : DFF_X1 port map( D => n11000, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2235_port, QN 
                           => n_1355);
   DataPath_RF_BLOCKi_77_Q_reg_28_inst : DFF_X1 port map( D => n10999, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2236_port, QN 
                           => n_1356);
   DataPath_RF_BLOCKi_77_Q_reg_29_inst : DFF_X1 port map( D => n10998, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2237_port, QN 
                           => n_1357);
   DataPath_RF_BLOCKi_77_Q_reg_30_inst : DFF_X1 port map( D => n10997, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2238_port, QN 
                           => n_1358);
   DataPath_RF_BLOCKi_77_Q_reg_31_inst : DFF_X1 port map( D => n10996, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2239_port, QN 
                           => n_1359);
   DataPath_RF_BLOCKi_76_Q_reg_0_inst : DFF_X1 port map( D => n10995, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2176_port, QN => 
                           n_1360);
   DataPath_RF_BLOCKi_76_Q_reg_1_inst : DFF_X1 port map( D => n10994, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2177_port, QN => 
                           n_1361);
   DataPath_RF_BLOCKi_76_Q_reg_2_inst : DFF_X1 port map( D => n10993, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2178_port, QN => 
                           n_1362);
   DataPath_RF_BLOCKi_76_Q_reg_3_inst : DFF_X1 port map( D => n10992, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2179_port, QN => 
                           n_1363);
   DataPath_RF_BLOCKi_76_Q_reg_4_inst : DFF_X1 port map( D => n10991, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2180_port, QN => 
                           n_1364);
   DataPath_RF_BLOCKi_76_Q_reg_5_inst : DFF_X1 port map( D => n10990, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2181_port, QN => 
                           n_1365);
   DataPath_RF_BLOCKi_76_Q_reg_6_inst : DFF_X1 port map( D => n10989, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2182_port, QN => 
                           n_1366);
   DataPath_RF_BLOCKi_76_Q_reg_7_inst : DFF_X1 port map( D => n10988, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2183_port, QN => 
                           n_1367);
   DataPath_RF_BLOCKi_76_Q_reg_8_inst : DFF_X1 port map( D => n10987, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2184_port, QN => 
                           n_1368);
   DataPath_RF_BLOCKi_76_Q_reg_9_inst : DFF_X1 port map( D => n10986, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2185_port, QN => 
                           n_1369);
   DataPath_RF_BLOCKi_76_Q_reg_10_inst : DFF_X1 port map( D => n10985, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2186_port, QN 
                           => n_1370);
   DataPath_RF_BLOCKi_76_Q_reg_11_inst : DFF_X1 port map( D => n10984, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2187_port, QN 
                           => n_1371);
   DataPath_RF_BLOCKi_76_Q_reg_12_inst : DFF_X1 port map( D => n10983, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2188_port, QN 
                           => n_1372);
   DataPath_RF_BLOCKi_76_Q_reg_13_inst : DFF_X1 port map( D => n10982, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2189_port, QN 
                           => n_1373);
   DataPath_RF_BLOCKi_76_Q_reg_14_inst : DFF_X1 port map( D => n10981, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2190_port, QN 
                           => n_1374);
   DataPath_RF_BLOCKi_76_Q_reg_15_inst : DFF_X1 port map( D => n10980, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2191_port, QN 
                           => n_1375);
   DataPath_RF_BLOCKi_76_Q_reg_16_inst : DFF_X1 port map( D => n10979, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2192_port, QN 
                           => n_1376);
   DataPath_RF_BLOCKi_76_Q_reg_17_inst : DFF_X1 port map( D => n10978, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2193_port, QN 
                           => n_1377);
   DataPath_RF_BLOCKi_76_Q_reg_18_inst : DFF_X1 port map( D => n10977, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2194_port, QN 
                           => n_1378);
   DataPath_RF_BLOCKi_76_Q_reg_19_inst : DFF_X1 port map( D => n10976, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2195_port, QN 
                           => n_1379);
   DataPath_RF_BLOCKi_76_Q_reg_20_inst : DFF_X1 port map( D => n10975, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2196_port, QN 
                           => n_1380);
   DataPath_RF_BLOCKi_76_Q_reg_21_inst : DFF_X1 port map( D => n10974, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2197_port, QN 
                           => n_1381);
   DataPath_RF_BLOCKi_76_Q_reg_22_inst : DFF_X1 port map( D => n10973, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2198_port, QN 
                           => n_1382);
   DataPath_RF_BLOCKi_76_Q_reg_23_inst : DFF_X1 port map( D => n10972, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2199_port, QN 
                           => n_1383);
   DataPath_RF_BLOCKi_76_Q_reg_24_inst : DFF_X1 port map( D => n10971, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2200_port, QN 
                           => n_1384);
   DataPath_RF_BLOCKi_76_Q_reg_25_inst : DFF_X1 port map( D => n10970, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2201_port, QN 
                           => n_1385);
   DataPath_RF_BLOCKi_76_Q_reg_26_inst : DFF_X1 port map( D => n10969, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2202_port, QN 
                           => n_1386);
   DataPath_RF_BLOCKi_76_Q_reg_27_inst : DFF_X1 port map( D => n10968, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2203_port, QN 
                           => n_1387);
   DataPath_RF_BLOCKi_76_Q_reg_28_inst : DFF_X1 port map( D => n10967, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2204_port, QN 
                           => n_1388);
   DataPath_RF_BLOCKi_76_Q_reg_29_inst : DFF_X1 port map( D => n10966, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2205_port, QN 
                           => n_1389);
   DataPath_RF_BLOCKi_76_Q_reg_30_inst : DFF_X1 port map( D => n10965, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2206_port, QN 
                           => n_1390);
   DataPath_RF_BLOCKi_76_Q_reg_31_inst : DFF_X1 port map( D => n10964, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2207_port, QN 
                           => n_1391);
   DataPath_RF_BLOCKi_75_Q_reg_0_inst : DFF_X1 port map( D => n10963, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2144_port, QN => 
                           n_1392);
   DataPath_RF_BLOCKi_75_Q_reg_1_inst : DFF_X1 port map( D => n10962, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2145_port, QN => 
                           n_1393);
   DataPath_RF_BLOCKi_75_Q_reg_2_inst : DFF_X1 port map( D => n10961, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2146_port, QN => 
                           n_1394);
   DataPath_RF_BLOCKi_75_Q_reg_3_inst : DFF_X1 port map( D => n10960, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2147_port, QN => 
                           n_1395);
   DataPath_RF_BLOCKi_75_Q_reg_4_inst : DFF_X1 port map( D => n10959, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2148_port, QN => 
                           n_1396);
   DataPath_RF_BLOCKi_75_Q_reg_5_inst : DFF_X1 port map( D => n10958, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2149_port, QN => 
                           n_1397);
   DataPath_RF_BLOCKi_75_Q_reg_6_inst : DFF_X1 port map( D => n10957, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2150_port, QN => 
                           n_1398);
   DataPath_RF_BLOCKi_75_Q_reg_7_inst : DFF_X1 port map( D => n10956, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2151_port, QN => 
                           n_1399);
   DataPath_RF_BLOCKi_75_Q_reg_8_inst : DFF_X1 port map( D => n10955, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2152_port, QN => 
                           n_1400);
   DataPath_RF_BLOCKi_75_Q_reg_9_inst : DFF_X1 port map( D => n10954, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2153_port, QN => 
                           n_1401);
   DataPath_RF_BLOCKi_75_Q_reg_10_inst : DFF_X1 port map( D => n10953, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2154_port, QN 
                           => n_1402);
   DataPath_RF_BLOCKi_75_Q_reg_11_inst : DFF_X1 port map( D => n10952, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2155_port, QN 
                           => n_1403);
   DataPath_RF_BLOCKi_75_Q_reg_12_inst : DFF_X1 port map( D => n10951, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2156_port, QN 
                           => n_1404);
   DataPath_RF_BLOCKi_75_Q_reg_13_inst : DFF_X1 port map( D => n10950, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2157_port, QN 
                           => n_1405);
   DataPath_RF_BLOCKi_75_Q_reg_14_inst : DFF_X1 port map( D => n10949, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2158_port, QN 
                           => n_1406);
   DataPath_RF_BLOCKi_75_Q_reg_15_inst : DFF_X1 port map( D => n10948, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2159_port, QN 
                           => n_1407);
   DataPath_RF_BLOCKi_75_Q_reg_16_inst : DFF_X1 port map( D => n10947, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2160_port, QN 
                           => n_1408);
   DataPath_RF_BLOCKi_75_Q_reg_17_inst : DFF_X1 port map( D => n10946, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2161_port, QN 
                           => n_1409);
   DataPath_RF_BLOCKi_75_Q_reg_18_inst : DFF_X1 port map( D => n10945, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2162_port, QN 
                           => n_1410);
   DataPath_RF_BLOCKi_75_Q_reg_19_inst : DFF_X1 port map( D => n10944, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2163_port, QN 
                           => n_1411);
   DataPath_RF_BLOCKi_75_Q_reg_20_inst : DFF_X1 port map( D => n10943, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2164_port, QN 
                           => n_1412);
   DataPath_RF_BLOCKi_75_Q_reg_21_inst : DFF_X1 port map( D => n10942, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2165_port, QN 
                           => n_1413);
   DataPath_RF_BLOCKi_75_Q_reg_22_inst : DFF_X1 port map( D => n10941, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2166_port, QN 
                           => n_1414);
   DataPath_RF_BLOCKi_75_Q_reg_23_inst : DFF_X1 port map( D => n10940, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2167_port, QN 
                           => n_1415);
   DataPath_RF_BLOCKi_75_Q_reg_24_inst : DFF_X1 port map( D => n10939, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2168_port, QN 
                           => n_1416);
   DataPath_RF_BLOCKi_75_Q_reg_25_inst : DFF_X1 port map( D => n10938, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2169_port, QN 
                           => n_1417);
   DataPath_RF_BLOCKi_75_Q_reg_26_inst : DFF_X1 port map( D => n10937, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2170_port, QN 
                           => n_1418);
   DataPath_RF_BLOCKi_75_Q_reg_27_inst : DFF_X1 port map( D => n10936, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2171_port, QN 
                           => n_1419);
   DataPath_RF_BLOCKi_75_Q_reg_28_inst : DFF_X1 port map( D => n10935, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2172_port, QN 
                           => n_1420);
   DataPath_RF_BLOCKi_75_Q_reg_29_inst : DFF_X1 port map( D => n10934, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2173_port, QN 
                           => n_1421);
   DataPath_RF_BLOCKi_75_Q_reg_30_inst : DFF_X1 port map( D => n10933, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2174_port, QN 
                           => n_1422);
   DataPath_RF_BLOCKi_75_Q_reg_31_inst : DFF_X1 port map( D => n10932, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2175_port, QN 
                           => n_1423);
   DataPath_RF_BLOCKi_74_Q_reg_0_inst : DFF_X1 port map( D => n10931, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2112_port, QN => 
                           n_1424);
   DataPath_RF_BLOCKi_74_Q_reg_1_inst : DFF_X1 port map( D => n10930, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2113_port, QN => 
                           n_1425);
   DataPath_RF_BLOCKi_74_Q_reg_2_inst : DFF_X1 port map( D => n10929, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2114_port, QN => 
                           n_1426);
   DataPath_RF_BLOCKi_74_Q_reg_3_inst : DFF_X1 port map( D => n10928, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2115_port, QN => 
                           n_1427);
   DataPath_RF_BLOCKi_74_Q_reg_4_inst : DFF_X1 port map( D => n10927, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2116_port, QN => 
                           n_1428);
   DataPath_RF_BLOCKi_74_Q_reg_5_inst : DFF_X1 port map( D => n10926, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2117_port, QN => 
                           n_1429);
   DataPath_RF_BLOCKi_74_Q_reg_6_inst : DFF_X1 port map( D => n10925, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2118_port, QN => 
                           n_1430);
   DataPath_RF_BLOCKi_74_Q_reg_7_inst : DFF_X1 port map( D => n10924, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2119_port, QN => 
                           n_1431);
   DataPath_RF_BLOCKi_74_Q_reg_8_inst : DFF_X1 port map( D => n10923, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2120_port, QN => 
                           n_1432);
   DataPath_RF_BLOCKi_74_Q_reg_9_inst : DFF_X1 port map( D => n10922, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2121_port, QN => 
                           n_1433);
   DataPath_RF_BLOCKi_74_Q_reg_10_inst : DFF_X1 port map( D => n10921, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2122_port, QN 
                           => n_1434);
   DataPath_RF_BLOCKi_74_Q_reg_11_inst : DFF_X1 port map( D => n10920, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2123_port, QN 
                           => n_1435);
   DataPath_RF_BLOCKi_74_Q_reg_12_inst : DFF_X1 port map( D => n10919, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2124_port, QN 
                           => n_1436);
   DataPath_RF_BLOCKi_74_Q_reg_13_inst : DFF_X1 port map( D => n10918, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2125_port, QN 
                           => n_1437);
   DataPath_RF_BLOCKi_74_Q_reg_14_inst : DFF_X1 port map( D => n10917, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2126_port, QN 
                           => n_1438);
   DataPath_RF_BLOCKi_74_Q_reg_15_inst : DFF_X1 port map( D => n10916, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2127_port, QN 
                           => n_1439);
   DataPath_RF_BLOCKi_74_Q_reg_16_inst : DFF_X1 port map( D => n10915, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2128_port, QN 
                           => n_1440);
   DataPath_RF_BLOCKi_74_Q_reg_17_inst : DFF_X1 port map( D => n10914, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2129_port, QN 
                           => n_1441);
   DataPath_RF_BLOCKi_74_Q_reg_18_inst : DFF_X1 port map( D => n10913, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2130_port, QN 
                           => n_1442);
   DataPath_RF_BLOCKi_74_Q_reg_19_inst : DFF_X1 port map( D => n10912, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2131_port, QN 
                           => n_1443);
   DataPath_RF_BLOCKi_74_Q_reg_20_inst : DFF_X1 port map( D => n10911, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2132_port, QN 
                           => n_1444);
   DataPath_RF_BLOCKi_74_Q_reg_21_inst : DFF_X1 port map( D => n10910, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2133_port, QN 
                           => n_1445);
   DataPath_RF_BLOCKi_74_Q_reg_22_inst : DFF_X1 port map( D => n10909, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2134_port, QN 
                           => n_1446);
   DataPath_RF_BLOCKi_74_Q_reg_23_inst : DFF_X1 port map( D => n10908, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2135_port, QN 
                           => n_1447);
   DataPath_RF_BLOCKi_74_Q_reg_24_inst : DFF_X1 port map( D => n10907, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2136_port, QN 
                           => n_1448);
   DataPath_RF_BLOCKi_74_Q_reg_25_inst : DFF_X1 port map( D => n10906, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2137_port, QN 
                           => n_1449);
   DataPath_RF_BLOCKi_74_Q_reg_26_inst : DFF_X1 port map( D => n10905, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2138_port, QN 
                           => n_1450);
   DataPath_RF_BLOCKi_74_Q_reg_27_inst : DFF_X1 port map( D => n10904, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2139_port, QN 
                           => n_1451);
   DataPath_RF_BLOCKi_74_Q_reg_28_inst : DFF_X1 port map( D => n10903, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2140_port, QN 
                           => n_1452);
   DataPath_RF_BLOCKi_74_Q_reg_29_inst : DFF_X1 port map( D => n10902, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2141_port, QN 
                           => n_1453);
   DataPath_RF_BLOCKi_74_Q_reg_30_inst : DFF_X1 port map( D => n10901, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2142_port, QN 
                           => n_1454);
   DataPath_RF_BLOCKi_74_Q_reg_31_inst : DFF_X1 port map( D => n10900, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2143_port, QN 
                           => n_1455);
   DataPath_RF_BLOCKi_73_Q_reg_0_inst : DFF_X1 port map( D => n10899, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2080_port, QN => 
                           n_1456);
   DataPath_RF_BLOCKi_73_Q_reg_1_inst : DFF_X1 port map( D => n10898, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2081_port, QN => 
                           n_1457);
   DataPath_RF_BLOCKi_73_Q_reg_2_inst : DFF_X1 port map( D => n10897, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2082_port, QN => 
                           n_1458);
   DataPath_RF_BLOCKi_73_Q_reg_3_inst : DFF_X1 port map( D => n10896, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2083_port, QN => 
                           n_1459);
   DataPath_RF_BLOCKi_73_Q_reg_4_inst : DFF_X1 port map( D => n10895, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2084_port, QN => 
                           n_1460);
   DataPath_RF_BLOCKi_73_Q_reg_5_inst : DFF_X1 port map( D => n10894, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2085_port, QN => 
                           n_1461);
   DataPath_RF_BLOCKi_73_Q_reg_6_inst : DFF_X1 port map( D => n10893, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2086_port, QN => 
                           n_1462);
   DataPath_RF_BLOCKi_73_Q_reg_7_inst : DFF_X1 port map( D => n10892, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2087_port, QN => 
                           n_1463);
   DataPath_RF_BLOCKi_73_Q_reg_8_inst : DFF_X1 port map( D => n10891, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2088_port, QN => 
                           n_1464);
   DataPath_RF_BLOCKi_73_Q_reg_9_inst : DFF_X1 port map( D => n10890, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2089_port, QN => 
                           n_1465);
   DataPath_RF_BLOCKi_73_Q_reg_10_inst : DFF_X1 port map( D => n10889, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2090_port, QN 
                           => n_1466);
   DataPath_RF_BLOCKi_73_Q_reg_11_inst : DFF_X1 port map( D => n10888, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2091_port, QN 
                           => n_1467);
   DataPath_RF_BLOCKi_73_Q_reg_12_inst : DFF_X1 port map( D => n10887, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2092_port, QN 
                           => n_1468);
   DataPath_RF_BLOCKi_73_Q_reg_13_inst : DFF_X1 port map( D => n10886, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2093_port, QN 
                           => n_1469);
   DataPath_RF_BLOCKi_73_Q_reg_14_inst : DFF_X1 port map( D => n10885, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2094_port, QN 
                           => n_1470);
   DataPath_RF_BLOCKi_73_Q_reg_15_inst : DFF_X1 port map( D => n10884, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2095_port, QN 
                           => n_1471);
   DataPath_RF_BLOCKi_73_Q_reg_16_inst : DFF_X1 port map( D => n10883, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2096_port, QN 
                           => n_1472);
   DataPath_RF_BLOCKi_73_Q_reg_17_inst : DFF_X1 port map( D => n10882, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2097_port, QN 
                           => n_1473);
   DataPath_RF_BLOCKi_73_Q_reg_18_inst : DFF_X1 port map( D => n10881, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2098_port, QN 
                           => n_1474);
   DataPath_RF_BLOCKi_73_Q_reg_19_inst : DFF_X1 port map( D => n10880, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2099_port, QN 
                           => n_1475);
   DataPath_RF_BLOCKi_73_Q_reg_20_inst : DFF_X1 port map( D => n10879, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2100_port, QN 
                           => n_1476);
   DataPath_RF_BLOCKi_73_Q_reg_21_inst : DFF_X1 port map( D => n10878, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2101_port, QN 
                           => n_1477);
   DataPath_RF_BLOCKi_73_Q_reg_22_inst : DFF_X1 port map( D => n10877, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2102_port, QN 
                           => n_1478);
   DataPath_RF_BLOCKi_73_Q_reg_23_inst : DFF_X1 port map( D => n10876, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2103_port, QN 
                           => n_1479);
   DataPath_RF_BLOCKi_73_Q_reg_24_inst : DFF_X1 port map( D => n10875, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2104_port, QN 
                           => n_1480);
   DataPath_RF_BLOCKi_73_Q_reg_25_inst : DFF_X1 port map( D => n10874, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2105_port, QN 
                           => n_1481);
   DataPath_RF_BLOCKi_73_Q_reg_26_inst : DFF_X1 port map( D => n10873, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2106_port, QN 
                           => n_1482);
   DataPath_RF_BLOCKi_73_Q_reg_27_inst : DFF_X1 port map( D => n10872, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2107_port, QN 
                           => n_1483);
   DataPath_RF_BLOCKi_73_Q_reg_28_inst : DFF_X1 port map( D => n10871, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2108_port, QN 
                           => n_1484);
   DataPath_RF_BLOCKi_73_Q_reg_29_inst : DFF_X1 port map( D => n10870, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2109_port, QN 
                           => n_1485);
   DataPath_RF_BLOCKi_73_Q_reg_30_inst : DFF_X1 port map( D => n10869, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2110_port, QN 
                           => n_1486);
   DataPath_RF_BLOCKi_73_Q_reg_31_inst : DFF_X1 port map( D => n10868, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2111_port, QN 
                           => n_1487);
   DataPath_RF_BLOCKi_72_Q_reg_0_inst : DFF_X1 port map( D => n10867, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2048_port, QN => 
                           n_1488);
   DataPath_RF_BLOCKi_72_Q_reg_1_inst : DFF_X1 port map( D => n10866, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2049_port, QN => 
                           n_1489);
   DataPath_RF_BLOCKi_72_Q_reg_2_inst : DFF_X1 port map( D => n10865, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2050_port, QN => 
                           n_1490);
   DataPath_RF_BLOCKi_72_Q_reg_3_inst : DFF_X1 port map( D => n10864, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2051_port, QN => 
                           n_1491);
   DataPath_RF_BLOCKi_72_Q_reg_4_inst : DFF_X1 port map( D => n10863, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2052_port, QN => 
                           n_1492);
   DataPath_RF_BLOCKi_72_Q_reg_5_inst : DFF_X1 port map( D => n10862, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2053_port, QN => 
                           n_1493);
   DataPath_RF_BLOCKi_72_Q_reg_6_inst : DFF_X1 port map( D => n10861, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2054_port, QN => 
                           n_1494);
   DataPath_RF_BLOCKi_72_Q_reg_7_inst : DFF_X1 port map( D => n10860, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2055_port, QN => 
                           n_1495);
   DataPath_RF_BLOCKi_72_Q_reg_8_inst : DFF_X1 port map( D => n10859, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2056_port, QN => 
                           n_1496);
   DataPath_RF_BLOCKi_72_Q_reg_9_inst : DFF_X1 port map( D => n10858, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2057_port, QN => 
                           n_1497);
   DataPath_RF_BLOCKi_72_Q_reg_10_inst : DFF_X1 port map( D => n10857, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2058_port, QN 
                           => n_1498);
   DataPath_RF_BLOCKi_72_Q_reg_11_inst : DFF_X1 port map( D => n10856, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2059_port, QN 
                           => n_1499);
   DataPath_RF_BLOCKi_72_Q_reg_12_inst : DFF_X1 port map( D => n10855, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2060_port, QN 
                           => n_1500);
   DataPath_RF_BLOCKi_72_Q_reg_13_inst : DFF_X1 port map( D => n10854, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2061_port, QN 
                           => n_1501);
   DataPath_RF_BLOCKi_72_Q_reg_14_inst : DFF_X1 port map( D => n10853, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2062_port, QN 
                           => n_1502);
   DataPath_RF_BLOCKi_72_Q_reg_15_inst : DFF_X1 port map( D => n10852, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2063_port, QN 
                           => n_1503);
   DataPath_RF_BLOCKi_72_Q_reg_16_inst : DFF_X1 port map( D => n10851, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2064_port, QN 
                           => n_1504);
   DataPath_RF_BLOCKi_72_Q_reg_17_inst : DFF_X1 port map( D => n10850, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2065_port, QN 
                           => n_1505);
   DataPath_RF_BLOCKi_72_Q_reg_18_inst : DFF_X1 port map( D => n10849, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2066_port, QN 
                           => n_1506);
   DataPath_RF_BLOCKi_72_Q_reg_19_inst : DFF_X1 port map( D => n10848, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2067_port, QN 
                           => n_1507);
   DataPath_RF_BLOCKi_72_Q_reg_20_inst : DFF_X1 port map( D => n10847, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2068_port, QN 
                           => n_1508);
   DataPath_RF_BLOCKi_72_Q_reg_21_inst : DFF_X1 port map( D => n10846, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2069_port, QN 
                           => n_1509);
   DataPath_RF_BLOCKi_72_Q_reg_22_inst : DFF_X1 port map( D => n10845, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2070_port, QN 
                           => n_1510);
   DataPath_RF_BLOCKi_72_Q_reg_23_inst : DFF_X1 port map( D => n10844, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2071_port, QN 
                           => n_1511);
   DataPath_RF_BLOCKi_72_Q_reg_24_inst : DFF_X1 port map( D => n10843, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2072_port, QN 
                           => n_1512);
   DataPath_RF_BLOCKi_72_Q_reg_25_inst : DFF_X1 port map( D => n10842, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2073_port, QN 
                           => n_1513);
   DataPath_RF_BLOCKi_72_Q_reg_26_inst : DFF_X1 port map( D => n10841, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2074_port, QN 
                           => n_1514);
   DataPath_RF_BLOCKi_72_Q_reg_27_inst : DFF_X1 port map( D => n10840, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2075_port, QN 
                           => n_1515);
   DataPath_RF_BLOCKi_72_Q_reg_28_inst : DFF_X1 port map( D => n10839, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2076_port, QN 
                           => n_1516);
   DataPath_RF_BLOCKi_72_Q_reg_29_inst : DFF_X1 port map( D => n10838, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2077_port, QN 
                           => n_1517);
   DataPath_RF_BLOCKi_72_Q_reg_30_inst : DFF_X1 port map( D => n10837, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2078_port, QN 
                           => n_1518);
   DataPath_RF_BLOCKi_72_Q_reg_31_inst : DFF_X1 port map( D => n10836, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2079_port, QN 
                           => n_1519);
   DataPath_RF_BLOCKi_71_Q_reg_0_inst : DFF_X1 port map( D => n10835, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2016_port, QN => 
                           n_1520);
   DataPath_RF_BLOCKi_71_Q_reg_1_inst : DFF_X1 port map( D => n10834, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2017_port, QN => 
                           n_1521);
   DataPath_RF_BLOCKi_71_Q_reg_2_inst : DFF_X1 port map( D => n10833, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2018_port, QN => 
                           n_1522);
   DataPath_RF_BLOCKi_71_Q_reg_3_inst : DFF_X1 port map( D => n10832, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2019_port, QN => 
                           n_1523);
   DataPath_RF_BLOCKi_71_Q_reg_4_inst : DFF_X1 port map( D => n10831, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2020_port, QN => 
                           n_1524);
   DataPath_RF_BLOCKi_71_Q_reg_5_inst : DFF_X1 port map( D => n10830, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2021_port, QN => 
                           n_1525);
   DataPath_RF_BLOCKi_71_Q_reg_6_inst : DFF_X1 port map( D => n10829, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2022_port, QN => 
                           n_1526);
   DataPath_RF_BLOCKi_71_Q_reg_7_inst : DFF_X1 port map( D => n10828, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2023_port, QN => 
                           n_1527);
   DataPath_RF_BLOCKi_71_Q_reg_8_inst : DFF_X1 port map( D => n10827, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2024_port, QN => 
                           n_1528);
   DataPath_RF_BLOCKi_71_Q_reg_9_inst : DFF_X1 port map( D => n10826, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_2025_port, QN => 
                           n_1529);
   DataPath_RF_BLOCKi_71_Q_reg_10_inst : DFF_X1 port map( D => n10825, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2026_port, QN 
                           => n_1530);
   DataPath_RF_BLOCKi_71_Q_reg_11_inst : DFF_X1 port map( D => n10824, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2027_port, QN 
                           => n_1531);
   DataPath_RF_BLOCKi_71_Q_reg_12_inst : DFF_X1 port map( D => n10823, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2028_port, QN 
                           => n_1532);
   DataPath_RF_BLOCKi_71_Q_reg_13_inst : DFF_X1 port map( D => n10822, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2029_port, QN 
                           => n_1533);
   DataPath_RF_BLOCKi_71_Q_reg_14_inst : DFF_X1 port map( D => n10821, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2030_port, QN 
                           => n_1534);
   DataPath_RF_BLOCKi_71_Q_reg_15_inst : DFF_X1 port map( D => n10820, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2031_port, QN 
                           => n_1535);
   DataPath_RF_BLOCKi_71_Q_reg_16_inst : DFF_X1 port map( D => n10819, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2032_port, QN 
                           => n_1536);
   DataPath_RF_BLOCKi_71_Q_reg_17_inst : DFF_X1 port map( D => n10818, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2033_port, QN 
                           => n_1537);
   DataPath_RF_BLOCKi_71_Q_reg_18_inst : DFF_X1 port map( D => n10817, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2034_port, QN 
                           => n_1538);
   DataPath_RF_BLOCKi_71_Q_reg_19_inst : DFF_X1 port map( D => n10816, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2035_port, QN 
                           => n_1539);
   DataPath_RF_BLOCKi_71_Q_reg_20_inst : DFF_X1 port map( D => n10815, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2036_port, QN 
                           => n_1540);
   DataPath_RF_BLOCKi_71_Q_reg_21_inst : DFF_X1 port map( D => n10814, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2037_port, QN 
                           => n_1541);
   DataPath_RF_BLOCKi_71_Q_reg_22_inst : DFF_X1 port map( D => n10813, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2038_port, QN 
                           => n_1542);
   DataPath_RF_BLOCKi_71_Q_reg_23_inst : DFF_X1 port map( D => n10812, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2039_port, QN 
                           => n_1543);
   DataPath_RF_BLOCKi_71_Q_reg_24_inst : DFF_X1 port map( D => n10811, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2040_port, QN 
                           => n_1544);
   DataPath_RF_BLOCKi_71_Q_reg_25_inst : DFF_X1 port map( D => n10810, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2041_port, QN 
                           => n_1545);
   DataPath_RF_BLOCKi_71_Q_reg_26_inst : DFF_X1 port map( D => n10809, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2042_port, QN 
                           => n_1546);
   DataPath_RF_BLOCKi_71_Q_reg_27_inst : DFF_X1 port map( D => n10808, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2043_port, QN 
                           => n_1547);
   DataPath_RF_BLOCKi_71_Q_reg_28_inst : DFF_X1 port map( D => n10807, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2044_port, QN 
                           => n_1548);
   DataPath_RF_BLOCKi_71_Q_reg_29_inst : DFF_X1 port map( D => n10806, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2045_port, QN 
                           => n_1549);
   DataPath_RF_BLOCKi_71_Q_reg_30_inst : DFF_X1 port map( D => n10805, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2046_port, QN 
                           => n_1550);
   DataPath_RF_BLOCKi_71_Q_reg_31_inst : DFF_X1 port map( D => n10804, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2047_port, QN 
                           => n_1551);
   DataPath_RF_BLOCKi_70_Q_reg_0_inst : DFF_X1 port map( D => n10803, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1984_port, QN => 
                           n_1552);
   DataPath_RF_BLOCKi_70_Q_reg_1_inst : DFF_X1 port map( D => n10802, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1985_port, QN => 
                           n_1553);
   DataPath_RF_BLOCKi_70_Q_reg_2_inst : DFF_X1 port map( D => n10801, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1986_port, QN => 
                           n_1554);
   DataPath_RF_BLOCKi_70_Q_reg_3_inst : DFF_X1 port map( D => n10800, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1987_port, QN => 
                           n_1555);
   DataPath_RF_BLOCKi_70_Q_reg_4_inst : DFF_X1 port map( D => n10799, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1988_port, QN => 
                           n_1556);
   DataPath_RF_BLOCKi_70_Q_reg_5_inst : DFF_X1 port map( D => n10798, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1989_port, QN => 
                           n_1557);
   DataPath_RF_BLOCKi_70_Q_reg_6_inst : DFF_X1 port map( D => n10797, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1990_port, QN => 
                           n_1558);
   DataPath_RF_BLOCKi_70_Q_reg_7_inst : DFF_X1 port map( D => n10796, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1991_port, QN => 
                           n_1559);
   DataPath_RF_BLOCKi_70_Q_reg_8_inst : DFF_X1 port map( D => n10795, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1992_port, QN => 
                           n_1560);
   DataPath_RF_BLOCKi_70_Q_reg_9_inst : DFF_X1 port map( D => n10794, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1993_port, QN => 
                           n_1561);
   DataPath_RF_BLOCKi_70_Q_reg_10_inst : DFF_X1 port map( D => n10793, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1994_port, QN 
                           => n_1562);
   DataPath_RF_BLOCKi_70_Q_reg_11_inst : DFF_X1 port map( D => n10792, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1995_port, QN 
                           => n_1563);
   DataPath_RF_BLOCKi_70_Q_reg_12_inst : DFF_X1 port map( D => n10791, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1996_port, QN 
                           => n_1564);
   DataPath_RF_BLOCKi_70_Q_reg_13_inst : DFF_X1 port map( D => n10790, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1997_port, QN 
                           => n_1565);
   DataPath_RF_BLOCKi_70_Q_reg_14_inst : DFF_X1 port map( D => n10789, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1998_port, QN 
                           => n_1566);
   DataPath_RF_BLOCKi_70_Q_reg_15_inst : DFF_X1 port map( D => n10788, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1999_port, QN 
                           => n_1567);
   DataPath_RF_BLOCKi_70_Q_reg_16_inst : DFF_X1 port map( D => n10787, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2000_port, QN 
                           => n_1568);
   DataPath_RF_BLOCKi_70_Q_reg_17_inst : DFF_X1 port map( D => n10786, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2001_port, QN 
                           => n_1569);
   DataPath_RF_BLOCKi_70_Q_reg_18_inst : DFF_X1 port map( D => n10785, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2002_port, QN 
                           => n_1570);
   DataPath_RF_BLOCKi_70_Q_reg_19_inst : DFF_X1 port map( D => n10784, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2003_port, QN 
                           => n_1571);
   DataPath_RF_BLOCKi_70_Q_reg_20_inst : DFF_X1 port map( D => n10783, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2004_port, QN 
                           => n_1572);
   DataPath_RF_BLOCKi_70_Q_reg_21_inst : DFF_X1 port map( D => n10782, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2005_port, QN 
                           => n_1573);
   DataPath_RF_BLOCKi_70_Q_reg_22_inst : DFF_X1 port map( D => n10781, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2006_port, QN 
                           => n_1574);
   DataPath_RF_BLOCKi_70_Q_reg_23_inst : DFF_X1 port map( D => n10780, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2007_port, QN 
                           => n_1575);
   DataPath_RF_BLOCKi_70_Q_reg_24_inst : DFF_X1 port map( D => n10779, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2008_port, QN 
                           => n_1576);
   DataPath_RF_BLOCKi_70_Q_reg_25_inst : DFF_X1 port map( D => n10778, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2009_port, QN 
                           => n_1577);
   DataPath_RF_BLOCKi_70_Q_reg_26_inst : DFF_X1 port map( D => n10777, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2010_port, QN 
                           => n_1578);
   DataPath_RF_BLOCKi_70_Q_reg_27_inst : DFF_X1 port map( D => n10776, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2011_port, QN 
                           => n_1579);
   DataPath_RF_BLOCKi_70_Q_reg_28_inst : DFF_X1 port map( D => n10775, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2012_port, QN 
                           => n_1580);
   DataPath_RF_BLOCKi_70_Q_reg_29_inst : DFF_X1 port map( D => n10774, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2013_port, QN 
                           => n_1581);
   DataPath_RF_BLOCKi_70_Q_reg_30_inst : DFF_X1 port map( D => n10773, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2014_port, QN 
                           => n_1582);
   DataPath_RF_BLOCKi_70_Q_reg_31_inst : DFF_X1 port map( D => n10772, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_2015_port, QN 
                           => n_1583);
   DataPath_RF_BLOCKi_69_Q_reg_0_inst : DFF_X1 port map( D => n10771, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1952_port, QN => 
                           n_1584);
   DataPath_RF_BLOCKi_69_Q_reg_1_inst : DFF_X1 port map( D => n10770, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1953_port, QN => 
                           n_1585);
   DataPath_RF_BLOCKi_69_Q_reg_2_inst : DFF_X1 port map( D => n10769, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1954_port, QN => 
                           n_1586);
   DataPath_RF_BLOCKi_69_Q_reg_3_inst : DFF_X1 port map( D => n10768, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1955_port, QN => 
                           n_1587);
   DataPath_RF_BLOCKi_69_Q_reg_4_inst : DFF_X1 port map( D => n10767, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1956_port, QN => 
                           n_1588);
   DataPath_RF_BLOCKi_69_Q_reg_5_inst : DFF_X1 port map( D => n10766, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1957_port, QN => 
                           n_1589);
   DataPath_RF_BLOCKi_69_Q_reg_6_inst : DFF_X1 port map( D => n10765, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1958_port, QN => 
                           n_1590);
   DataPath_RF_BLOCKi_69_Q_reg_7_inst : DFF_X1 port map( D => n10764, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1959_port, QN => 
                           n_1591);
   DataPath_RF_BLOCKi_69_Q_reg_8_inst : DFF_X1 port map( D => n10763, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1960_port, QN => 
                           n_1592);
   DataPath_RF_BLOCKi_69_Q_reg_9_inst : DFF_X1 port map( D => n10762, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1961_port, QN => 
                           n_1593);
   DataPath_RF_BLOCKi_69_Q_reg_10_inst : DFF_X1 port map( D => n10761, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1962_port, QN 
                           => n_1594);
   DataPath_RF_BLOCKi_69_Q_reg_11_inst : DFF_X1 port map( D => n10760, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1963_port, QN 
                           => n_1595);
   DataPath_RF_BLOCKi_69_Q_reg_12_inst : DFF_X1 port map( D => n10759, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1964_port, QN 
                           => n_1596);
   DataPath_RF_BLOCKi_69_Q_reg_13_inst : DFF_X1 port map( D => n10758, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1965_port, QN 
                           => n_1597);
   DataPath_RF_BLOCKi_69_Q_reg_14_inst : DFF_X1 port map( D => n10757, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1966_port, QN 
                           => n_1598);
   DataPath_RF_BLOCKi_69_Q_reg_15_inst : DFF_X1 port map( D => n10756, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1967_port, QN 
                           => n_1599);
   DataPath_RF_BLOCKi_69_Q_reg_16_inst : DFF_X1 port map( D => n10755, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1968_port, QN 
                           => n_1600);
   DataPath_RF_BLOCKi_69_Q_reg_17_inst : DFF_X1 port map( D => n10754, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1969_port, QN 
                           => n_1601);
   DataPath_RF_BLOCKi_69_Q_reg_18_inst : DFF_X1 port map( D => n10753, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1970_port, QN 
                           => n_1602);
   DataPath_RF_BLOCKi_69_Q_reg_19_inst : DFF_X1 port map( D => n10752, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1971_port, QN 
                           => n_1603);
   DataPath_RF_BLOCKi_69_Q_reg_20_inst : DFF_X1 port map( D => n10751, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1972_port, QN 
                           => n_1604);
   DataPath_RF_BLOCKi_69_Q_reg_21_inst : DFF_X1 port map( D => n10750, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1973_port, QN 
                           => n_1605);
   DataPath_RF_BLOCKi_69_Q_reg_22_inst : DFF_X1 port map( D => n10749, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1974_port, QN 
                           => n_1606);
   DataPath_RF_BLOCKi_69_Q_reg_23_inst : DFF_X1 port map( D => n10748, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1975_port, QN 
                           => n_1607);
   DataPath_RF_BLOCKi_69_Q_reg_24_inst : DFF_X1 port map( D => n10747, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1976_port, QN 
                           => n_1608);
   DataPath_RF_BLOCKi_69_Q_reg_25_inst : DFF_X1 port map( D => n10746, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1977_port, QN 
                           => n_1609);
   DataPath_RF_BLOCKi_69_Q_reg_26_inst : DFF_X1 port map( D => n10745, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1978_port, QN 
                           => n_1610);
   DataPath_RF_BLOCKi_69_Q_reg_27_inst : DFF_X1 port map( D => n10744, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1979_port, QN 
                           => n_1611);
   DataPath_RF_BLOCKi_69_Q_reg_28_inst : DFF_X1 port map( D => n10743, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1980_port, QN 
                           => n_1612);
   DataPath_RF_BLOCKi_69_Q_reg_29_inst : DFF_X1 port map( D => n10742, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1981_port, QN 
                           => n_1613);
   DataPath_RF_BLOCKi_69_Q_reg_30_inst : DFF_X1 port map( D => n10741, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1982_port, QN 
                           => n_1614);
   DataPath_RF_BLOCKi_69_Q_reg_31_inst : DFF_X1 port map( D => n10740, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1983_port, QN 
                           => n_1615);
   DataPath_RF_BLOCKi_68_Q_reg_0_inst : DFF_X1 port map( D => n10739, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1920_port, QN => 
                           n_1616);
   DataPath_RF_BLOCKi_68_Q_reg_1_inst : DFF_X1 port map( D => n10738, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1921_port, QN => 
                           n_1617);
   DataPath_RF_BLOCKi_68_Q_reg_2_inst : DFF_X1 port map( D => n10737, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1922_port, QN => 
                           n_1618);
   DataPath_RF_BLOCKi_68_Q_reg_3_inst : DFF_X1 port map( D => n10736, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1923_port, QN => 
                           n_1619);
   DataPath_RF_BLOCKi_68_Q_reg_4_inst : DFF_X1 port map( D => n10735, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1924_port, QN => 
                           n_1620);
   DataPath_RF_BLOCKi_68_Q_reg_5_inst : DFF_X1 port map( D => n10734, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1925_port, QN => 
                           n_1621);
   DataPath_RF_BLOCKi_68_Q_reg_6_inst : DFF_X1 port map( D => n10733, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1926_port, QN => 
                           n_1622);
   DataPath_RF_BLOCKi_68_Q_reg_7_inst : DFF_X1 port map( D => n10732, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1927_port, QN => 
                           n_1623);
   DataPath_RF_BLOCKi_68_Q_reg_8_inst : DFF_X1 port map( D => n10731, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1928_port, QN => 
                           n_1624);
   DataPath_RF_BLOCKi_68_Q_reg_9_inst : DFF_X1 port map( D => n10730, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1929_port, QN => 
                           n_1625);
   DataPath_RF_BLOCKi_68_Q_reg_10_inst : DFF_X1 port map( D => n10729, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1930_port, QN 
                           => n_1626);
   DataPath_RF_BLOCKi_68_Q_reg_11_inst : DFF_X1 port map( D => n10728, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1931_port, QN 
                           => n_1627);
   DataPath_RF_BLOCKi_68_Q_reg_12_inst : DFF_X1 port map( D => n10727, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1932_port, QN 
                           => n_1628);
   DataPath_RF_BLOCKi_68_Q_reg_13_inst : DFF_X1 port map( D => n10726, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1933_port, QN 
                           => n_1629);
   DataPath_RF_BLOCKi_68_Q_reg_14_inst : DFF_X1 port map( D => n10725, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1934_port, QN 
                           => n_1630);
   DataPath_RF_BLOCKi_68_Q_reg_15_inst : DFF_X1 port map( D => n10724, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1935_port, QN 
                           => n_1631);
   DataPath_RF_BLOCKi_68_Q_reg_16_inst : DFF_X1 port map( D => n10723, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1936_port, QN 
                           => n_1632);
   DataPath_RF_BLOCKi_68_Q_reg_17_inst : DFF_X1 port map( D => n10722, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1937_port, QN 
                           => n_1633);
   DataPath_RF_BLOCKi_68_Q_reg_18_inst : DFF_X1 port map( D => n10721, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1938_port, QN 
                           => n_1634);
   DataPath_RF_BLOCKi_68_Q_reg_19_inst : DFF_X1 port map( D => n10720, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1939_port, QN 
                           => n_1635);
   DataPath_RF_BLOCKi_68_Q_reg_20_inst : DFF_X1 port map( D => n10719, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1940_port, QN 
                           => n_1636);
   DataPath_RF_BLOCKi_68_Q_reg_21_inst : DFF_X1 port map( D => n10718, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1941_port, QN 
                           => n_1637);
   DataPath_RF_BLOCKi_68_Q_reg_22_inst : DFF_X1 port map( D => n10717, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1942_port, QN 
                           => n_1638);
   DataPath_RF_BLOCKi_68_Q_reg_23_inst : DFF_X1 port map( D => n10716, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1943_port, QN 
                           => n_1639);
   DataPath_RF_BLOCKi_68_Q_reg_24_inst : DFF_X1 port map( D => n10715, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1944_port, QN 
                           => n_1640);
   DataPath_RF_BLOCKi_68_Q_reg_25_inst : DFF_X1 port map( D => n10714, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1945_port, QN 
                           => n_1641);
   DataPath_RF_BLOCKi_68_Q_reg_26_inst : DFF_X1 port map( D => n10713, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1946_port, QN 
                           => n_1642);
   DataPath_RF_BLOCKi_68_Q_reg_27_inst : DFF_X1 port map( D => n10712, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1947_port, QN 
                           => n_1643);
   DataPath_RF_BLOCKi_68_Q_reg_28_inst : DFF_X1 port map( D => n10711, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1948_port, QN 
                           => n_1644);
   DataPath_RF_BLOCKi_68_Q_reg_29_inst : DFF_X1 port map( D => n10710, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1949_port, QN 
                           => n_1645);
   DataPath_RF_BLOCKi_68_Q_reg_30_inst : DFF_X1 port map( D => n10709, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1950_port, QN 
                           => n_1646);
   DataPath_RF_BLOCKi_68_Q_reg_31_inst : DFF_X1 port map( D => n10708, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1951_port, QN 
                           => n_1647);
   DataPath_RF_BLOCKi_67_Q_reg_0_inst : DFF_X1 port map( D => n10707, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1888_port, QN => 
                           n_1648);
   DataPath_RF_BLOCKi_67_Q_reg_1_inst : DFF_X1 port map( D => n10706, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1889_port, QN => 
                           n_1649);
   DataPath_RF_BLOCKi_67_Q_reg_2_inst : DFF_X1 port map( D => n10705, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1890_port, QN => 
                           n_1650);
   DataPath_RF_BLOCKi_67_Q_reg_3_inst : DFF_X1 port map( D => n10704, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1891_port, QN => 
                           n_1651);
   DataPath_RF_BLOCKi_67_Q_reg_4_inst : DFF_X1 port map( D => n10703, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1892_port, QN => 
                           n_1652);
   DataPath_RF_BLOCKi_67_Q_reg_5_inst : DFF_X1 port map( D => n10702, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1893_port, QN => 
                           n_1653);
   DataPath_RF_BLOCKi_67_Q_reg_6_inst : DFF_X1 port map( D => n10701, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1894_port, QN => 
                           n_1654);
   DataPath_RF_BLOCKi_67_Q_reg_7_inst : DFF_X1 port map( D => n10700, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1895_port, QN => 
                           n_1655);
   DataPath_RF_BLOCKi_67_Q_reg_8_inst : DFF_X1 port map( D => n10699, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1896_port, QN => 
                           n_1656);
   DataPath_RF_BLOCKi_67_Q_reg_9_inst : DFF_X1 port map( D => n10698, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1897_port, QN => 
                           n_1657);
   DataPath_RF_BLOCKi_67_Q_reg_10_inst : DFF_X1 port map( D => n10697, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1898_port, QN 
                           => n_1658);
   DataPath_RF_BLOCKi_67_Q_reg_11_inst : DFF_X1 port map( D => n10696, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1899_port, QN 
                           => n_1659);
   DataPath_RF_BLOCKi_67_Q_reg_12_inst : DFF_X1 port map( D => n10695, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1900_port, QN 
                           => n_1660);
   DataPath_RF_BLOCKi_67_Q_reg_13_inst : DFF_X1 port map( D => n10694, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1901_port, QN 
                           => n_1661);
   DataPath_RF_BLOCKi_67_Q_reg_14_inst : DFF_X1 port map( D => n10693, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1902_port, QN 
                           => n_1662);
   DataPath_RF_BLOCKi_67_Q_reg_15_inst : DFF_X1 port map( D => n10692, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1903_port, QN 
                           => n_1663);
   DataPath_RF_BLOCKi_67_Q_reg_16_inst : DFF_X1 port map( D => n10691, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1904_port, QN 
                           => n_1664);
   DataPath_RF_BLOCKi_67_Q_reg_17_inst : DFF_X1 port map( D => n10690, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1905_port, QN 
                           => n_1665);
   DataPath_RF_BLOCKi_67_Q_reg_18_inst : DFF_X1 port map( D => n10689, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1906_port, QN 
                           => n_1666);
   DataPath_RF_BLOCKi_67_Q_reg_19_inst : DFF_X1 port map( D => n10688, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1907_port, QN 
                           => n_1667);
   DataPath_RF_BLOCKi_67_Q_reg_20_inst : DFF_X1 port map( D => n10687, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1908_port, QN 
                           => n_1668);
   DataPath_RF_BLOCKi_67_Q_reg_21_inst : DFF_X1 port map( D => n10686, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1909_port, QN 
                           => n_1669);
   DataPath_RF_BLOCKi_67_Q_reg_22_inst : DFF_X1 port map( D => n10685, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1910_port, QN 
                           => n_1670);
   DataPath_RF_BLOCKi_67_Q_reg_23_inst : DFF_X1 port map( D => n10684, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1911_port, QN 
                           => n_1671);
   DataPath_RF_BLOCKi_67_Q_reg_24_inst : DFF_X1 port map( D => n10683, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1912_port, QN 
                           => n_1672);
   DataPath_RF_BLOCKi_67_Q_reg_25_inst : DFF_X1 port map( D => n10682, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1913_port, QN 
                           => n_1673);
   DataPath_RF_BLOCKi_67_Q_reg_26_inst : DFF_X1 port map( D => n10681, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1914_port, QN 
                           => n_1674);
   DataPath_RF_BLOCKi_67_Q_reg_27_inst : DFF_X1 port map( D => n10680, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1915_port, QN 
                           => n_1675);
   DataPath_RF_BLOCKi_67_Q_reg_28_inst : DFF_X1 port map( D => n10679, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1916_port, QN 
                           => n_1676);
   DataPath_RF_BLOCKi_67_Q_reg_29_inst : DFF_X1 port map( D => n10678, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1917_port, QN 
                           => n_1677);
   DataPath_RF_BLOCKi_67_Q_reg_30_inst : DFF_X1 port map( D => n10677, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1918_port, QN 
                           => n_1678);
   DataPath_RF_BLOCKi_67_Q_reg_31_inst : DFF_X1 port map( D => n10676, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1919_port, QN 
                           => n_1679);
   DataPath_RF_BLOCKi_66_Q_reg_0_inst : DFF_X1 port map( D => n10675, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1856_port, QN => 
                           n_1680);
   DataPath_RF_BLOCKi_66_Q_reg_1_inst : DFF_X1 port map( D => n10674, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1857_port, QN => 
                           n_1681);
   DataPath_RF_BLOCKi_66_Q_reg_2_inst : DFF_X1 port map( D => n10673, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1858_port, QN => 
                           n_1682);
   DataPath_RF_BLOCKi_66_Q_reg_3_inst : DFF_X1 port map( D => n10672, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1859_port, QN => 
                           n_1683);
   DataPath_RF_BLOCKi_66_Q_reg_4_inst : DFF_X1 port map( D => n10671, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1860_port, QN => 
                           n_1684);
   DataPath_RF_BLOCKi_66_Q_reg_5_inst : DFF_X1 port map( D => n10670, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1861_port, QN => 
                           n_1685);
   DataPath_RF_BLOCKi_66_Q_reg_6_inst : DFF_X1 port map( D => n10669, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1862_port, QN => 
                           n_1686);
   DataPath_RF_BLOCKi_66_Q_reg_7_inst : DFF_X1 port map( D => n10668, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1863_port, QN => 
                           n_1687);
   DataPath_RF_BLOCKi_66_Q_reg_8_inst : DFF_X1 port map( D => n10667, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1864_port, QN => 
                           n_1688);
   DataPath_RF_BLOCKi_66_Q_reg_9_inst : DFF_X1 port map( D => n10666, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1865_port, QN => 
                           n_1689);
   DataPath_RF_BLOCKi_66_Q_reg_10_inst : DFF_X1 port map( D => n10665, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1866_port, QN 
                           => n_1690);
   DataPath_RF_BLOCKi_66_Q_reg_11_inst : DFF_X1 port map( D => n10664, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1867_port, QN 
                           => n_1691);
   DataPath_RF_BLOCKi_66_Q_reg_12_inst : DFF_X1 port map( D => n10663, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1868_port, QN 
                           => n_1692);
   DataPath_RF_BLOCKi_66_Q_reg_13_inst : DFF_X1 port map( D => n10662, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1869_port, QN 
                           => n_1693);
   DataPath_RF_BLOCKi_66_Q_reg_14_inst : DFF_X1 port map( D => n10661, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1870_port, QN 
                           => n_1694);
   DataPath_RF_BLOCKi_66_Q_reg_15_inst : DFF_X1 port map( D => n10660, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1871_port, QN 
                           => n_1695);
   DataPath_RF_BLOCKi_66_Q_reg_16_inst : DFF_X1 port map( D => n10659, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1872_port, QN 
                           => n_1696);
   DataPath_RF_BLOCKi_66_Q_reg_17_inst : DFF_X1 port map( D => n10658, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1873_port, QN 
                           => n_1697);
   DataPath_RF_BLOCKi_66_Q_reg_18_inst : DFF_X1 port map( D => n10657, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1874_port, QN 
                           => n_1698);
   DataPath_RF_BLOCKi_66_Q_reg_19_inst : DFF_X1 port map( D => n10656, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1875_port, QN 
                           => n_1699);
   DataPath_RF_BLOCKi_66_Q_reg_20_inst : DFF_X1 port map( D => n10655, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1876_port, QN 
                           => n_1700);
   DataPath_RF_BLOCKi_66_Q_reg_21_inst : DFF_X1 port map( D => n10654, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1877_port, QN 
                           => n_1701);
   DataPath_RF_BLOCKi_66_Q_reg_22_inst : DFF_X1 port map( D => n10653, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1878_port, QN 
                           => n_1702);
   DataPath_RF_BLOCKi_66_Q_reg_23_inst : DFF_X1 port map( D => n10652, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1879_port, QN 
                           => n_1703);
   DataPath_RF_BLOCKi_66_Q_reg_24_inst : DFF_X1 port map( D => n10651, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1880_port, QN 
                           => n_1704);
   DataPath_RF_BLOCKi_66_Q_reg_25_inst : DFF_X1 port map( D => n10650, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1881_port, QN 
                           => n_1705);
   DataPath_RF_BLOCKi_66_Q_reg_26_inst : DFF_X1 port map( D => n10649, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1882_port, QN 
                           => n_1706);
   DataPath_RF_BLOCKi_66_Q_reg_27_inst : DFF_X1 port map( D => n10648, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1883_port, QN 
                           => n_1707);
   DataPath_RF_BLOCKi_66_Q_reg_28_inst : DFF_X1 port map( D => n10647, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1884_port, QN 
                           => n_1708);
   DataPath_RF_BLOCKi_66_Q_reg_29_inst : DFF_X1 port map( D => n10646, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1885_port, QN 
                           => n_1709);
   DataPath_RF_BLOCKi_66_Q_reg_30_inst : DFF_X1 port map( D => n10645, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1886_port, QN 
                           => n_1710);
   DataPath_RF_BLOCKi_66_Q_reg_31_inst : DFF_X1 port map( D => n10644, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1887_port, QN 
                           => n_1711);
   DataPath_RF_BLOCKi_65_Q_reg_0_inst : DFF_X1 port map( D => n10643, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1824_port, QN => 
                           n_1712);
   DataPath_RF_BLOCKi_65_Q_reg_1_inst : DFF_X1 port map( D => n10642, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1825_port, QN => 
                           n_1713);
   DataPath_RF_BLOCKi_65_Q_reg_2_inst : DFF_X1 port map( D => n10641, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1826_port, QN => 
                           n_1714);
   DataPath_RF_BLOCKi_65_Q_reg_3_inst : DFF_X1 port map( D => n10640, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1827_port, QN => 
                           n_1715);
   DataPath_RF_BLOCKi_65_Q_reg_4_inst : DFF_X1 port map( D => n10639, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1828_port, QN => 
                           n_1716);
   DataPath_RF_BLOCKi_65_Q_reg_5_inst : DFF_X1 port map( D => n10638, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1829_port, QN => 
                           n_1717);
   DataPath_RF_BLOCKi_65_Q_reg_6_inst : DFF_X1 port map( D => n10637, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1830_port, QN => 
                           n_1718);
   DataPath_RF_BLOCKi_65_Q_reg_7_inst : DFF_X1 port map( D => n10636, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1831_port, QN => 
                           n_1719);
   DataPath_RF_BLOCKi_65_Q_reg_8_inst : DFF_X1 port map( D => n10635, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1832_port, QN => 
                           n_1720);
   DataPath_RF_BLOCKi_65_Q_reg_9_inst : DFF_X1 port map( D => n10634, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1833_port, QN => 
                           n_1721);
   DataPath_RF_BLOCKi_65_Q_reg_10_inst : DFF_X1 port map( D => n10633, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1834_port, QN 
                           => n_1722);
   DataPath_RF_BLOCKi_65_Q_reg_11_inst : DFF_X1 port map( D => n10632, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1835_port, QN 
                           => n_1723);
   DataPath_RF_BLOCKi_65_Q_reg_12_inst : DFF_X1 port map( D => n10631, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1836_port, QN 
                           => n_1724);
   DataPath_RF_BLOCKi_65_Q_reg_13_inst : DFF_X1 port map( D => n10630, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1837_port, QN 
                           => n_1725);
   DataPath_RF_BLOCKi_65_Q_reg_14_inst : DFF_X1 port map( D => n10629, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1838_port, QN 
                           => n_1726);
   DataPath_RF_BLOCKi_65_Q_reg_15_inst : DFF_X1 port map( D => n10628, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1839_port, QN 
                           => n_1727);
   DataPath_RF_BLOCKi_65_Q_reg_16_inst : DFF_X1 port map( D => n10627, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1840_port, QN 
                           => n_1728);
   DataPath_RF_BLOCKi_65_Q_reg_17_inst : DFF_X1 port map( D => n10626, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1841_port, QN 
                           => n_1729);
   DataPath_RF_BLOCKi_65_Q_reg_18_inst : DFF_X1 port map( D => n10625, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1842_port, QN 
                           => n_1730);
   DataPath_RF_BLOCKi_65_Q_reg_19_inst : DFF_X1 port map( D => n10624, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1843_port, QN 
                           => n_1731);
   DataPath_RF_BLOCKi_65_Q_reg_20_inst : DFF_X1 port map( D => n10623, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1844_port, QN 
                           => n_1732);
   DataPath_RF_BLOCKi_65_Q_reg_21_inst : DFF_X1 port map( D => n10622, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1845_port, QN 
                           => n_1733);
   DataPath_RF_BLOCKi_65_Q_reg_22_inst : DFF_X1 port map( D => n10621, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1846_port, QN 
                           => n_1734);
   DataPath_RF_BLOCKi_65_Q_reg_23_inst : DFF_X1 port map( D => n10620, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1847_port, QN 
                           => n_1735);
   DataPath_RF_BLOCKi_65_Q_reg_24_inst : DFF_X1 port map( D => n10619, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1848_port, QN 
                           => n_1736);
   DataPath_RF_BLOCKi_65_Q_reg_25_inst : DFF_X1 port map( D => n10618, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1849_port, QN 
                           => n_1737);
   DataPath_RF_BLOCKi_65_Q_reg_26_inst : DFF_X1 port map( D => n10617, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1850_port, QN 
                           => n_1738);
   DataPath_RF_BLOCKi_65_Q_reg_27_inst : DFF_X1 port map( D => n10616, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1851_port, QN 
                           => n_1739);
   DataPath_RF_BLOCKi_65_Q_reg_28_inst : DFF_X1 port map( D => n10615, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1852_port, QN 
                           => n_1740);
   DataPath_RF_BLOCKi_65_Q_reg_29_inst : DFF_X1 port map( D => n10614, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1853_port, QN 
                           => n_1741);
   DataPath_RF_BLOCKi_65_Q_reg_30_inst : DFF_X1 port map( D => n10613, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1854_port, QN 
                           => n_1742);
   DataPath_RF_BLOCKi_65_Q_reg_31_inst : DFF_X1 port map( D => n10612, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1855_port, QN 
                           => n_1743);
   DataPath_RF_BLOCKi_64_Q_reg_0_inst : DFF_X1 port map( D => n10611, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1792_port, QN => 
                           n_1744);
   DataPath_RF_BLOCKi_64_Q_reg_1_inst : DFF_X1 port map( D => n10610, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1793_port, QN => 
                           n_1745);
   DataPath_RF_BLOCKi_64_Q_reg_2_inst : DFF_X1 port map( D => n10609, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1794_port, QN => 
                           n_1746);
   DataPath_RF_BLOCKi_64_Q_reg_3_inst : DFF_X1 port map( D => n10608, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1795_port, QN => 
                           n_1747);
   DataPath_RF_BLOCKi_64_Q_reg_4_inst : DFF_X1 port map( D => n10607, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1796_port, QN => 
                           n_1748);
   DataPath_RF_BLOCKi_64_Q_reg_5_inst : DFF_X1 port map( D => n10606, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1797_port, QN => 
                           n_1749);
   DataPath_RF_BLOCKi_64_Q_reg_6_inst : DFF_X1 port map( D => n10605, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1798_port, QN => 
                           n_1750);
   DataPath_RF_BLOCKi_64_Q_reg_7_inst : DFF_X1 port map( D => n10604, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1799_port, QN => 
                           n_1751);
   DataPath_RF_BLOCKi_64_Q_reg_8_inst : DFF_X1 port map( D => n10603, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1800_port, QN => 
                           n_1752);
   DataPath_RF_BLOCKi_64_Q_reg_9_inst : DFF_X1 port map( D => n10602, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1801_port, QN => 
                           n_1753);
   DataPath_RF_BLOCKi_64_Q_reg_10_inst : DFF_X1 port map( D => n10601, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1802_port, QN 
                           => n_1754);
   DataPath_RF_BLOCKi_64_Q_reg_11_inst : DFF_X1 port map( D => n10600, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1803_port, QN 
                           => n_1755);
   DataPath_RF_BLOCKi_64_Q_reg_12_inst : DFF_X1 port map( D => n10599, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1804_port, QN 
                           => n_1756);
   DataPath_RF_BLOCKi_64_Q_reg_13_inst : DFF_X1 port map( D => n10598, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1805_port, QN 
                           => n_1757);
   DataPath_RF_BLOCKi_64_Q_reg_14_inst : DFF_X1 port map( D => n10597, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1806_port, QN 
                           => n_1758);
   DataPath_RF_BLOCKi_64_Q_reg_15_inst : DFF_X1 port map( D => n10596, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1807_port, QN 
                           => n_1759);
   DataPath_RF_BLOCKi_64_Q_reg_16_inst : DFF_X1 port map( D => n10595, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1808_port, QN 
                           => n_1760);
   DataPath_RF_BLOCKi_64_Q_reg_17_inst : DFF_X1 port map( D => n10594, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1809_port, QN 
                           => n_1761);
   DataPath_RF_BLOCKi_64_Q_reg_18_inst : DFF_X1 port map( D => n10593, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1810_port, QN 
                           => n_1762);
   DataPath_RF_BLOCKi_64_Q_reg_19_inst : DFF_X1 port map( D => n10592, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1811_port, QN 
                           => n_1763);
   DataPath_RF_BLOCKi_64_Q_reg_20_inst : DFF_X1 port map( D => n10591, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1812_port, QN 
                           => n_1764);
   DataPath_RF_BLOCKi_64_Q_reg_21_inst : DFF_X1 port map( D => n10590, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1813_port, QN 
                           => n_1765);
   DataPath_RF_BLOCKi_64_Q_reg_22_inst : DFF_X1 port map( D => n10589, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1814_port, QN 
                           => n_1766);
   DataPath_RF_BLOCKi_64_Q_reg_23_inst : DFF_X1 port map( D => n10588, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1815_port, QN 
                           => n_1767);
   DataPath_RF_BLOCKi_64_Q_reg_24_inst : DFF_X1 port map( D => n10587, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1816_port, QN 
                           => n_1768);
   DataPath_RF_BLOCKi_64_Q_reg_25_inst : DFF_X1 port map( D => n10586, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1817_port, QN 
                           => n_1769);
   DataPath_RF_BLOCKi_64_Q_reg_26_inst : DFF_X1 port map( D => n10585, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1818_port, QN 
                           => n_1770);
   DataPath_RF_BLOCKi_64_Q_reg_27_inst : DFF_X1 port map( D => n10584, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1819_port, QN 
                           => n_1771);
   DataPath_RF_BLOCKi_64_Q_reg_28_inst : DFF_X1 port map( D => n10583, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1820_port, QN 
                           => n_1772);
   DataPath_RF_BLOCKi_64_Q_reg_29_inst : DFF_X1 port map( D => n10582, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1821_port, QN 
                           => n_1773);
   DataPath_RF_BLOCKi_64_Q_reg_30_inst : DFF_X1 port map( D => n10581, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1822_port, QN 
                           => n_1774);
   DataPath_RF_BLOCKi_64_Q_reg_31_inst : DFF_X1 port map( D => n10580, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1823_port, QN 
                           => n_1775);
   DataPath_RF_BLOCKi_63_Q_reg_0_inst : DFF_X1 port map( D => n10579, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1760_port, QN => 
                           n_1776);
   DataPath_RF_BLOCKi_63_Q_reg_1_inst : DFF_X1 port map( D => n10578, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1761_port, QN => 
                           n_1777);
   DataPath_RF_BLOCKi_63_Q_reg_2_inst : DFF_X1 port map( D => n10577, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1762_port, QN => 
                           n_1778);
   DataPath_RF_BLOCKi_63_Q_reg_3_inst : DFF_X1 port map( D => n10576, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1763_port, QN => 
                           n_1779);
   DataPath_RF_BLOCKi_63_Q_reg_4_inst : DFF_X1 port map( D => n10575, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1764_port, QN => 
                           n_1780);
   DataPath_RF_BLOCKi_63_Q_reg_5_inst : DFF_X1 port map( D => n10574, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1765_port, QN => 
                           n_1781);
   DataPath_RF_BLOCKi_63_Q_reg_6_inst : DFF_X1 port map( D => n10573, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1766_port, QN => 
                           n_1782);
   DataPath_RF_BLOCKi_63_Q_reg_7_inst : DFF_X1 port map( D => n10572, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1767_port, QN => 
                           n_1783);
   DataPath_RF_BLOCKi_63_Q_reg_8_inst : DFF_X1 port map( D => n10571, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1768_port, QN => 
                           n_1784);
   DataPath_RF_BLOCKi_63_Q_reg_9_inst : DFF_X1 port map( D => n10570, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1769_port, QN => 
                           n_1785);
   DataPath_RF_BLOCKi_63_Q_reg_10_inst : DFF_X1 port map( D => n10569, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1770_port, QN 
                           => n_1786);
   DataPath_RF_BLOCKi_63_Q_reg_11_inst : DFF_X1 port map( D => n10568, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1771_port, QN 
                           => n_1787);
   DataPath_RF_BLOCKi_63_Q_reg_12_inst : DFF_X1 port map( D => n10567, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1772_port, QN 
                           => n_1788);
   DataPath_RF_BLOCKi_63_Q_reg_13_inst : DFF_X1 port map( D => n10566, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1773_port, QN 
                           => n_1789);
   DataPath_RF_BLOCKi_63_Q_reg_14_inst : DFF_X1 port map( D => n10565, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1774_port, QN 
                           => n_1790);
   DataPath_RF_BLOCKi_63_Q_reg_15_inst : DFF_X1 port map( D => n10564, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1775_port, QN 
                           => n_1791);
   DataPath_RF_BLOCKi_63_Q_reg_16_inst : DFF_X1 port map( D => n10563, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1776_port, QN 
                           => n_1792);
   DataPath_RF_BLOCKi_63_Q_reg_17_inst : DFF_X1 port map( D => n10562, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1777_port, QN 
                           => n_1793);
   DataPath_RF_BLOCKi_63_Q_reg_18_inst : DFF_X1 port map( D => n10561, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1778_port, QN 
                           => n_1794);
   DataPath_RF_BLOCKi_63_Q_reg_19_inst : DFF_X1 port map( D => n10560, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1779_port, QN 
                           => n_1795);
   DataPath_RF_BLOCKi_63_Q_reg_20_inst : DFF_X1 port map( D => n10559, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1780_port, QN 
                           => n_1796);
   DataPath_RF_BLOCKi_63_Q_reg_21_inst : DFF_X1 port map( D => n10558, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1781_port, QN 
                           => n_1797);
   DataPath_RF_BLOCKi_63_Q_reg_22_inst : DFF_X1 port map( D => n10557, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1782_port, QN 
                           => n_1798);
   DataPath_RF_BLOCKi_63_Q_reg_23_inst : DFF_X1 port map( D => n10556, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1783_port, QN 
                           => n_1799);
   DataPath_RF_BLOCKi_63_Q_reg_24_inst : DFF_X1 port map( D => n10555, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1784_port, QN 
                           => n_1800);
   DataPath_RF_BLOCKi_63_Q_reg_25_inst : DFF_X1 port map( D => n10554, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1785_port, QN 
                           => n_1801);
   DataPath_RF_BLOCKi_63_Q_reg_26_inst : DFF_X1 port map( D => n10553, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1786_port, QN 
                           => n_1802);
   DataPath_RF_BLOCKi_63_Q_reg_27_inst : DFF_X1 port map( D => n10552, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1787_port, QN 
                           => n_1803);
   DataPath_RF_BLOCKi_63_Q_reg_28_inst : DFF_X1 port map( D => n10551, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1788_port, QN 
                           => n_1804);
   DataPath_RF_BLOCKi_63_Q_reg_29_inst : DFF_X1 port map( D => n10550, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1789_port, QN 
                           => n_1805);
   DataPath_RF_BLOCKi_63_Q_reg_30_inst : DFF_X1 port map( D => n10549, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1790_port, QN 
                           => n_1806);
   DataPath_RF_BLOCKi_63_Q_reg_31_inst : DFF_X1 port map( D => n10548, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1791_port, QN 
                           => n_1807);
   DataPath_RF_BLOCKi_62_Q_reg_0_inst : DFF_X1 port map( D => n10547, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1728_port, QN => 
                           n_1808);
   DataPath_RF_BLOCKi_62_Q_reg_1_inst : DFF_X1 port map( D => n10546, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1729_port, QN => 
                           n_1809);
   DataPath_RF_BLOCKi_62_Q_reg_2_inst : DFF_X1 port map( D => n10545, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1730_port, QN => 
                           n_1810);
   DataPath_RF_BLOCKi_62_Q_reg_3_inst : DFF_X1 port map( D => n10544, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1731_port, QN => 
                           n_1811);
   DataPath_RF_BLOCKi_62_Q_reg_4_inst : DFF_X1 port map( D => n10543, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1732_port, QN => 
                           n_1812);
   DataPath_RF_BLOCKi_62_Q_reg_5_inst : DFF_X1 port map( D => n10542, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1733_port, QN => 
                           n_1813);
   DataPath_RF_BLOCKi_62_Q_reg_6_inst : DFF_X1 port map( D => n10541, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1734_port, QN => 
                           n_1814);
   DataPath_RF_BLOCKi_62_Q_reg_7_inst : DFF_X1 port map( D => n10540, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1735_port, QN => 
                           n_1815);
   DataPath_RF_BLOCKi_62_Q_reg_8_inst : DFF_X1 port map( D => n10539, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1736_port, QN => 
                           n_1816);
   DataPath_RF_BLOCKi_62_Q_reg_9_inst : DFF_X1 port map( D => n10538, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1737_port, QN => 
                           n_1817);
   DataPath_RF_BLOCKi_62_Q_reg_10_inst : DFF_X1 port map( D => n10537, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1738_port, QN 
                           => n_1818);
   DataPath_RF_BLOCKi_62_Q_reg_11_inst : DFF_X1 port map( D => n10536, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1739_port, QN 
                           => n_1819);
   DataPath_RF_BLOCKi_62_Q_reg_12_inst : DFF_X1 port map( D => n10535, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1740_port, QN 
                           => n_1820);
   DataPath_RF_BLOCKi_62_Q_reg_13_inst : DFF_X1 port map( D => n10534, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1741_port, QN 
                           => n_1821);
   DataPath_RF_BLOCKi_62_Q_reg_14_inst : DFF_X1 port map( D => n10533, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1742_port, QN 
                           => n_1822);
   DataPath_RF_BLOCKi_62_Q_reg_15_inst : DFF_X1 port map( D => n10532, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1743_port, QN 
                           => n_1823);
   DataPath_RF_BLOCKi_62_Q_reg_16_inst : DFF_X1 port map( D => n10531, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1744_port, QN 
                           => n_1824);
   DataPath_RF_BLOCKi_62_Q_reg_17_inst : DFF_X1 port map( D => n10530, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1745_port, QN 
                           => n_1825);
   DataPath_RF_BLOCKi_62_Q_reg_18_inst : DFF_X1 port map( D => n10529, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1746_port, QN 
                           => n_1826);
   DataPath_RF_BLOCKi_62_Q_reg_19_inst : DFF_X1 port map( D => n10528, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1747_port, QN 
                           => n_1827);
   DataPath_RF_BLOCKi_62_Q_reg_20_inst : DFF_X1 port map( D => n10527, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1748_port, QN 
                           => n_1828);
   DataPath_RF_BLOCKi_62_Q_reg_21_inst : DFF_X1 port map( D => n10526, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1749_port, QN 
                           => n_1829);
   DataPath_RF_BLOCKi_62_Q_reg_22_inst : DFF_X1 port map( D => n10525, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1750_port, QN 
                           => n_1830);
   DataPath_RF_BLOCKi_62_Q_reg_23_inst : DFF_X1 port map( D => n10524, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1751_port, QN 
                           => n_1831);
   DataPath_RF_BLOCKi_62_Q_reg_24_inst : DFF_X1 port map( D => n10523, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1752_port, QN 
                           => n_1832);
   DataPath_RF_BLOCKi_62_Q_reg_25_inst : DFF_X1 port map( D => n10522, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1753_port, QN 
                           => n_1833);
   DataPath_RF_BLOCKi_62_Q_reg_26_inst : DFF_X1 port map( D => n10521, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1754_port, QN 
                           => n_1834);
   DataPath_RF_BLOCKi_62_Q_reg_27_inst : DFF_X1 port map( D => n10520, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1755_port, QN 
                           => n_1835);
   DataPath_RF_BLOCKi_62_Q_reg_28_inst : DFF_X1 port map( D => n10519, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1756_port, QN 
                           => n_1836);
   DataPath_RF_BLOCKi_62_Q_reg_29_inst : DFF_X1 port map( D => n10518, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1757_port, QN 
                           => n_1837);
   DataPath_RF_BLOCKi_62_Q_reg_30_inst : DFF_X1 port map( D => n10517, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1758_port, QN 
                           => n_1838);
   DataPath_RF_BLOCKi_62_Q_reg_31_inst : DFF_X1 port map( D => n10516, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1759_port, QN 
                           => n_1839);
   DataPath_RF_BLOCKi_61_Q_reg_0_inst : DFF_X1 port map( D => n10515, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1696_port, QN => 
                           n_1840);
   DataPath_RF_BLOCKi_61_Q_reg_1_inst : DFF_X1 port map( D => n10514, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1697_port, QN => 
                           n_1841);
   DataPath_RF_BLOCKi_61_Q_reg_2_inst : DFF_X1 port map( D => n10513, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1698_port, QN => 
                           n_1842);
   DataPath_RF_BLOCKi_61_Q_reg_3_inst : DFF_X1 port map( D => n10512, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1699_port, QN => 
                           n_1843);
   DataPath_RF_BLOCKi_61_Q_reg_4_inst : DFF_X1 port map( D => n10511, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1700_port, QN => 
                           n_1844);
   DataPath_RF_BLOCKi_61_Q_reg_5_inst : DFF_X1 port map( D => n10510, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1701_port, QN => 
                           n_1845);
   DataPath_RF_BLOCKi_61_Q_reg_6_inst : DFF_X1 port map( D => n10509, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1702_port, QN => 
                           n_1846);
   DataPath_RF_BLOCKi_61_Q_reg_7_inst : DFF_X1 port map( D => n10508, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1703_port, QN => 
                           n_1847);
   DataPath_RF_BLOCKi_61_Q_reg_8_inst : DFF_X1 port map( D => n10507, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1704_port, QN => 
                           n_1848);
   DataPath_RF_BLOCKi_61_Q_reg_9_inst : DFF_X1 port map( D => n10506, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1705_port, QN => 
                           n_1849);
   DataPath_RF_BLOCKi_61_Q_reg_10_inst : DFF_X1 port map( D => n10505, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1706_port, QN 
                           => n_1850);
   DataPath_RF_BLOCKi_61_Q_reg_11_inst : DFF_X1 port map( D => n10504, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1707_port, QN 
                           => n_1851);
   DataPath_RF_BLOCKi_61_Q_reg_12_inst : DFF_X1 port map( D => n10503, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1708_port, QN 
                           => n_1852);
   DataPath_RF_BLOCKi_61_Q_reg_13_inst : DFF_X1 port map( D => n10502, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1709_port, QN 
                           => n_1853);
   DataPath_RF_BLOCKi_61_Q_reg_14_inst : DFF_X1 port map( D => n10501, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1710_port, QN 
                           => n_1854);
   DataPath_RF_BLOCKi_61_Q_reg_15_inst : DFF_X1 port map( D => n10500, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1711_port, QN 
                           => n_1855);
   DataPath_RF_BLOCKi_61_Q_reg_16_inst : DFF_X1 port map( D => n10499, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1712_port, QN 
                           => n_1856);
   DataPath_RF_BLOCKi_61_Q_reg_17_inst : DFF_X1 port map( D => n10498, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1713_port, QN 
                           => n_1857);
   DataPath_RF_BLOCKi_61_Q_reg_18_inst : DFF_X1 port map( D => n10497, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1714_port, QN 
                           => n_1858);
   DataPath_RF_BLOCKi_61_Q_reg_19_inst : DFF_X1 port map( D => n10496, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1715_port, QN 
                           => n_1859);
   DataPath_RF_BLOCKi_61_Q_reg_20_inst : DFF_X1 port map( D => n10495, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1716_port, QN 
                           => n_1860);
   DataPath_RF_BLOCKi_61_Q_reg_21_inst : DFF_X1 port map( D => n10494, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1717_port, QN 
                           => n_1861);
   DataPath_RF_BLOCKi_61_Q_reg_22_inst : DFF_X1 port map( D => n10493, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1718_port, QN 
                           => n_1862);
   DataPath_RF_BLOCKi_61_Q_reg_23_inst : DFF_X1 port map( D => n10492, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1719_port, QN 
                           => n_1863);
   DataPath_RF_BLOCKi_61_Q_reg_24_inst : DFF_X1 port map( D => n10491, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1720_port, QN 
                           => n_1864);
   DataPath_RF_BLOCKi_61_Q_reg_25_inst : DFF_X1 port map( D => n10490, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1721_port, QN 
                           => n_1865);
   DataPath_RF_BLOCKi_61_Q_reg_26_inst : DFF_X1 port map( D => n10489, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1722_port, QN 
                           => n_1866);
   DataPath_RF_BLOCKi_61_Q_reg_27_inst : DFF_X1 port map( D => n10488, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1723_port, QN 
                           => n_1867);
   DataPath_RF_BLOCKi_61_Q_reg_28_inst : DFF_X1 port map( D => n10487, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1724_port, QN 
                           => n_1868);
   DataPath_RF_BLOCKi_61_Q_reg_29_inst : DFF_X1 port map( D => n10486, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1725_port, QN 
                           => n_1869);
   DataPath_RF_BLOCKi_61_Q_reg_30_inst : DFF_X1 port map( D => n10485, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1726_port, QN 
                           => n_1870);
   DataPath_RF_BLOCKi_61_Q_reg_31_inst : DFF_X1 port map( D => n10484, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1727_port, QN 
                           => n_1871);
   DataPath_RF_BLOCKi_60_Q_reg_0_inst : DFF_X1 port map( D => n10483, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1664_port, QN => 
                           n_1872);
   DataPath_RF_BLOCKi_60_Q_reg_1_inst : DFF_X1 port map( D => n10482, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1665_port, QN => 
                           n_1873);
   DataPath_RF_BLOCKi_60_Q_reg_2_inst : DFF_X1 port map( D => n10481, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1666_port, QN => 
                           n_1874);
   DataPath_RF_BLOCKi_60_Q_reg_3_inst : DFF_X1 port map( D => n10480, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1667_port, QN => 
                           n_1875);
   DataPath_RF_BLOCKi_60_Q_reg_4_inst : DFF_X1 port map( D => n10479, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1668_port, QN => 
                           n_1876);
   DataPath_RF_BLOCKi_60_Q_reg_5_inst : DFF_X1 port map( D => n10478, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1669_port, QN => 
                           n_1877);
   DataPath_RF_BLOCKi_60_Q_reg_6_inst : DFF_X1 port map( D => n10477, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1670_port, QN => 
                           n_1878);
   DataPath_RF_BLOCKi_60_Q_reg_7_inst : DFF_X1 port map( D => n10476, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1671_port, QN => 
                           n_1879);
   DataPath_RF_BLOCKi_60_Q_reg_8_inst : DFF_X1 port map( D => n10475, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1672_port, QN => 
                           n_1880);
   DataPath_RF_BLOCKi_60_Q_reg_9_inst : DFF_X1 port map( D => n10474, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1673_port, QN => 
                           n_1881);
   DataPath_RF_BLOCKi_60_Q_reg_10_inst : DFF_X1 port map( D => n10473, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1674_port, QN 
                           => n_1882);
   DataPath_RF_BLOCKi_60_Q_reg_11_inst : DFF_X1 port map( D => n10472, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1675_port, QN 
                           => n_1883);
   DataPath_RF_BLOCKi_60_Q_reg_12_inst : DFF_X1 port map( D => n10471, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1676_port, QN 
                           => n_1884);
   DataPath_RF_BLOCKi_60_Q_reg_13_inst : DFF_X1 port map( D => n10470, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1677_port, QN 
                           => n_1885);
   DataPath_RF_BLOCKi_60_Q_reg_14_inst : DFF_X1 port map( D => n10469, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1678_port, QN 
                           => n_1886);
   DataPath_RF_BLOCKi_60_Q_reg_15_inst : DFF_X1 port map( D => n10468, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1679_port, QN 
                           => n_1887);
   DataPath_RF_BLOCKi_60_Q_reg_16_inst : DFF_X1 port map( D => n10467, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1680_port, QN 
                           => n_1888);
   DataPath_RF_BLOCKi_60_Q_reg_17_inst : DFF_X1 port map( D => n10466, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1681_port, QN 
                           => n_1889);
   DataPath_RF_BLOCKi_60_Q_reg_18_inst : DFF_X1 port map( D => n10465, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1682_port, QN 
                           => n_1890);
   DataPath_RF_BLOCKi_60_Q_reg_19_inst : DFF_X1 port map( D => n10464, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1683_port, QN 
                           => n_1891);
   DataPath_RF_BLOCKi_60_Q_reg_20_inst : DFF_X1 port map( D => n10463, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1684_port, QN 
                           => n_1892);
   DataPath_RF_BLOCKi_60_Q_reg_21_inst : DFF_X1 port map( D => n10462, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1685_port, QN 
                           => n_1893);
   DataPath_RF_BLOCKi_60_Q_reg_22_inst : DFF_X1 port map( D => n10461, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1686_port, QN 
                           => n_1894);
   DataPath_RF_BLOCKi_60_Q_reg_23_inst : DFF_X1 port map( D => n10460, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1687_port, QN 
                           => n_1895);
   DataPath_RF_BLOCKi_60_Q_reg_24_inst : DFF_X1 port map( D => n10459, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1688_port, QN 
                           => n_1896);
   DataPath_RF_BLOCKi_60_Q_reg_25_inst : DFF_X1 port map( D => n10458, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1689_port, QN 
                           => n_1897);
   DataPath_RF_BLOCKi_60_Q_reg_26_inst : DFF_X1 port map( D => n10457, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1690_port, QN 
                           => n_1898);
   DataPath_RF_BLOCKi_60_Q_reg_27_inst : DFF_X1 port map( D => n10456, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1691_port, QN 
                           => n_1899);
   DataPath_RF_BLOCKi_60_Q_reg_28_inst : DFF_X1 port map( D => n10455, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1692_port, QN 
                           => n_1900);
   DataPath_RF_BLOCKi_60_Q_reg_29_inst : DFF_X1 port map( D => n10454, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1693_port, QN 
                           => n_1901);
   DataPath_RF_BLOCKi_60_Q_reg_30_inst : DFF_X1 port map( D => n10453, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1694_port, QN 
                           => n_1902);
   DataPath_RF_BLOCKi_60_Q_reg_31_inst : DFF_X1 port map( D => n10452, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1695_port, QN 
                           => n_1903);
   DataPath_RF_BLOCKi_59_Q_reg_0_inst : DFF_X1 port map( D => n10451, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1632_port, QN => 
                           n_1904);
   DataPath_RF_BLOCKi_59_Q_reg_1_inst : DFF_X1 port map( D => n10450, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1633_port, QN => 
                           n_1905);
   DataPath_RF_BLOCKi_59_Q_reg_2_inst : DFF_X1 port map( D => n10449, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1634_port, QN => 
                           n_1906);
   DataPath_RF_BLOCKi_59_Q_reg_3_inst : DFF_X1 port map( D => n10448, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1635_port, QN => 
                           n_1907);
   DataPath_RF_BLOCKi_59_Q_reg_4_inst : DFF_X1 port map( D => n10447, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1636_port, QN => 
                           n_1908);
   DataPath_RF_BLOCKi_59_Q_reg_5_inst : DFF_X1 port map( D => n10446, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1637_port, QN => 
                           n_1909);
   DataPath_RF_BLOCKi_59_Q_reg_6_inst : DFF_X1 port map( D => n10445, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1638_port, QN => 
                           n_1910);
   DataPath_RF_BLOCKi_59_Q_reg_7_inst : DFF_X1 port map( D => n10444, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1639_port, QN => 
                           n_1911);
   DataPath_RF_BLOCKi_59_Q_reg_8_inst : DFF_X1 port map( D => n10443, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1640_port, QN => 
                           n_1912);
   DataPath_RF_BLOCKi_59_Q_reg_9_inst : DFF_X1 port map( D => n10442, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1641_port, QN => 
                           n_1913);
   DataPath_RF_BLOCKi_59_Q_reg_10_inst : DFF_X1 port map( D => n10441, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1642_port, QN 
                           => n_1914);
   DataPath_RF_BLOCKi_59_Q_reg_11_inst : DFF_X1 port map( D => n10440, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1643_port, QN 
                           => n_1915);
   DataPath_RF_BLOCKi_59_Q_reg_12_inst : DFF_X1 port map( D => n10439, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1644_port, QN 
                           => n_1916);
   DataPath_RF_BLOCKi_59_Q_reg_13_inst : DFF_X1 port map( D => n10438, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1645_port, QN 
                           => n_1917);
   DataPath_RF_BLOCKi_59_Q_reg_14_inst : DFF_X1 port map( D => n10437, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1646_port, QN 
                           => n_1918);
   DataPath_RF_BLOCKi_59_Q_reg_15_inst : DFF_X1 port map( D => n10436, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1647_port, QN 
                           => n_1919);
   DataPath_RF_BLOCKi_59_Q_reg_16_inst : DFF_X1 port map( D => n10435, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1648_port, QN 
                           => n_1920);
   DataPath_RF_BLOCKi_59_Q_reg_17_inst : DFF_X1 port map( D => n10434, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1649_port, QN 
                           => n_1921);
   DataPath_RF_BLOCKi_59_Q_reg_18_inst : DFF_X1 port map( D => n10433, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1650_port, QN 
                           => n_1922);
   DataPath_RF_BLOCKi_59_Q_reg_19_inst : DFF_X1 port map( D => n10432, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1651_port, QN 
                           => n_1923);
   DataPath_RF_BLOCKi_59_Q_reg_20_inst : DFF_X1 port map( D => n10431, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1652_port, QN 
                           => n_1924);
   DataPath_RF_BLOCKi_59_Q_reg_21_inst : DFF_X1 port map( D => n10430, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1653_port, QN 
                           => n_1925);
   DataPath_RF_BLOCKi_59_Q_reg_22_inst : DFF_X1 port map( D => n10429, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1654_port, QN 
                           => n_1926);
   DataPath_RF_BLOCKi_59_Q_reg_23_inst : DFF_X1 port map( D => n10428, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1655_port, QN 
                           => n_1927);
   DataPath_RF_BLOCKi_59_Q_reg_24_inst : DFF_X1 port map( D => n10427, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1656_port, QN 
                           => n_1928);
   DataPath_RF_BLOCKi_59_Q_reg_25_inst : DFF_X1 port map( D => n10426, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1657_port, QN 
                           => n_1929);
   DataPath_RF_BLOCKi_59_Q_reg_26_inst : DFF_X1 port map( D => n10425, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1658_port, QN 
                           => n_1930);
   DataPath_RF_BLOCKi_59_Q_reg_27_inst : DFF_X1 port map( D => n10424, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1659_port, QN 
                           => n_1931);
   DataPath_RF_BLOCKi_59_Q_reg_28_inst : DFF_X1 port map( D => n10423, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1660_port, QN 
                           => n_1932);
   DataPath_RF_BLOCKi_59_Q_reg_29_inst : DFF_X1 port map( D => n10422, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1661_port, QN 
                           => n_1933);
   DataPath_RF_BLOCKi_59_Q_reg_30_inst : DFF_X1 port map( D => n10421, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1662_port, QN 
                           => n_1934);
   DataPath_RF_BLOCKi_59_Q_reg_31_inst : DFF_X1 port map( D => n10420, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1663_port, QN 
                           => n_1935);
   DataPath_RF_BLOCKi_58_Q_reg_0_inst : DFF_X1 port map( D => n10419, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1600_port, QN => 
                           n_1936);
   DataPath_RF_BLOCKi_58_Q_reg_1_inst : DFF_X1 port map( D => n10418, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1601_port, QN => 
                           n_1937);
   DataPath_RF_BLOCKi_58_Q_reg_2_inst : DFF_X1 port map( D => n10417, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1602_port, QN => 
                           n_1938);
   DataPath_RF_BLOCKi_58_Q_reg_3_inst : DFF_X1 port map( D => n10416, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1603_port, QN => 
                           n_1939);
   DataPath_RF_BLOCKi_58_Q_reg_4_inst : DFF_X1 port map( D => n10415, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1604_port, QN => 
                           n_1940);
   DataPath_RF_BLOCKi_58_Q_reg_5_inst : DFF_X1 port map( D => n10414, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1605_port, QN => 
                           n_1941);
   DataPath_RF_BLOCKi_58_Q_reg_6_inst : DFF_X1 port map( D => n10413, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1606_port, QN => 
                           n_1942);
   DataPath_RF_BLOCKi_58_Q_reg_7_inst : DFF_X1 port map( D => n10412, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1607_port, QN => 
                           n_1943);
   DataPath_RF_BLOCKi_58_Q_reg_8_inst : DFF_X1 port map( D => n10411, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1608_port, QN => 
                           n_1944);
   DataPath_RF_BLOCKi_58_Q_reg_9_inst : DFF_X1 port map( D => n10410, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1609_port, QN => 
                           n_1945);
   DataPath_RF_BLOCKi_58_Q_reg_10_inst : DFF_X1 port map( D => n10409, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1610_port, QN 
                           => n_1946);
   DataPath_RF_BLOCKi_58_Q_reg_11_inst : DFF_X1 port map( D => n10408, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1611_port, QN 
                           => n_1947);
   DataPath_RF_BLOCKi_58_Q_reg_12_inst : DFF_X1 port map( D => n10407, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1612_port, QN 
                           => n_1948);
   DataPath_RF_BLOCKi_58_Q_reg_13_inst : DFF_X1 port map( D => n10406, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1613_port, QN 
                           => n_1949);
   DataPath_RF_BLOCKi_58_Q_reg_14_inst : DFF_X1 port map( D => n10405, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1614_port, QN 
                           => n_1950);
   DataPath_RF_BLOCKi_58_Q_reg_15_inst : DFF_X1 port map( D => n10404, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1615_port, QN 
                           => n_1951);
   DataPath_RF_BLOCKi_58_Q_reg_16_inst : DFF_X1 port map( D => n10403, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1616_port, QN 
                           => n_1952);
   DataPath_RF_BLOCKi_58_Q_reg_17_inst : DFF_X1 port map( D => n10402, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1617_port, QN 
                           => n_1953);
   DataPath_RF_BLOCKi_58_Q_reg_18_inst : DFF_X1 port map( D => n10401, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1618_port, QN 
                           => n_1954);
   DataPath_RF_BLOCKi_58_Q_reg_19_inst : DFF_X1 port map( D => n10400, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1619_port, QN 
                           => n_1955);
   DataPath_RF_BLOCKi_58_Q_reg_20_inst : DFF_X1 port map( D => n10399, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1620_port, QN 
                           => n_1956);
   DataPath_RF_BLOCKi_58_Q_reg_21_inst : DFF_X1 port map( D => n10398, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1621_port, QN 
                           => n_1957);
   DataPath_RF_BLOCKi_58_Q_reg_22_inst : DFF_X1 port map( D => n10397, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1622_port, QN 
                           => n_1958);
   DataPath_RF_BLOCKi_58_Q_reg_23_inst : DFF_X1 port map( D => n10396, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1623_port, QN 
                           => n_1959);
   DataPath_RF_BLOCKi_58_Q_reg_24_inst : DFF_X1 port map( D => n10395, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1624_port, QN 
                           => n_1960);
   DataPath_RF_BLOCKi_58_Q_reg_25_inst : DFF_X1 port map( D => n10394, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1625_port, QN 
                           => n_1961);
   DataPath_RF_BLOCKi_58_Q_reg_26_inst : DFF_X1 port map( D => n10393, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1626_port, QN 
                           => n_1962);
   DataPath_RF_BLOCKi_58_Q_reg_27_inst : DFF_X1 port map( D => n10392, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1627_port, QN 
                           => n_1963);
   DataPath_RF_BLOCKi_58_Q_reg_28_inst : DFF_X1 port map( D => n10391, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1628_port, QN 
                           => n_1964);
   DataPath_RF_BLOCKi_58_Q_reg_29_inst : DFF_X1 port map( D => n10390, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1629_port, QN 
                           => n_1965);
   DataPath_RF_BLOCKi_58_Q_reg_30_inst : DFF_X1 port map( D => n10389, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1630_port, QN 
                           => n_1966);
   DataPath_RF_BLOCKi_58_Q_reg_31_inst : DFF_X1 port map( D => n10388, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1631_port, QN 
                           => n_1967);
   DataPath_RF_BLOCKi_57_Q_reg_0_inst : DFF_X1 port map( D => n10387, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1568_port, QN => 
                           n_1968);
   DataPath_RF_BLOCKi_57_Q_reg_1_inst : DFF_X1 port map( D => n10386, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1569_port, QN => 
                           n_1969);
   DataPath_RF_BLOCKi_57_Q_reg_2_inst : DFF_X1 port map( D => n10385, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1570_port, QN => 
                           n_1970);
   DataPath_RF_BLOCKi_57_Q_reg_3_inst : DFF_X1 port map( D => n10384, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1571_port, QN => 
                           n_1971);
   DataPath_RF_BLOCKi_57_Q_reg_4_inst : DFF_X1 port map( D => n10383, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1572_port, QN => 
                           n_1972);
   DataPath_RF_BLOCKi_57_Q_reg_5_inst : DFF_X1 port map( D => n10382, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1573_port, QN => 
                           n_1973);
   DataPath_RF_BLOCKi_57_Q_reg_6_inst : DFF_X1 port map( D => n10381, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1574_port, QN => 
                           n_1974);
   DataPath_RF_BLOCKi_57_Q_reg_7_inst : DFF_X1 port map( D => n10380, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1575_port, QN => 
                           n_1975);
   DataPath_RF_BLOCKi_57_Q_reg_8_inst : DFF_X1 port map( D => n10379, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1576_port, QN => 
                           n_1976);
   DataPath_RF_BLOCKi_57_Q_reg_9_inst : DFF_X1 port map( D => n10378, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1577_port, QN => 
                           n_1977);
   DataPath_RF_BLOCKi_57_Q_reg_10_inst : DFF_X1 port map( D => n10377, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1578_port, QN 
                           => n_1978);
   DataPath_RF_BLOCKi_57_Q_reg_11_inst : DFF_X1 port map( D => n10376, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1579_port, QN 
                           => n_1979);
   DataPath_RF_BLOCKi_57_Q_reg_12_inst : DFF_X1 port map( D => n10375, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1580_port, QN 
                           => n_1980);
   DataPath_RF_BLOCKi_57_Q_reg_13_inst : DFF_X1 port map( D => n10374, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1581_port, QN 
                           => n_1981);
   DataPath_RF_BLOCKi_57_Q_reg_14_inst : DFF_X1 port map( D => n10373, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1582_port, QN 
                           => n_1982);
   DataPath_RF_BLOCKi_57_Q_reg_15_inst : DFF_X1 port map( D => n10372, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1583_port, QN 
                           => n_1983);
   DataPath_RF_BLOCKi_57_Q_reg_16_inst : DFF_X1 port map( D => n10371, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1584_port, QN 
                           => n_1984);
   DataPath_RF_BLOCKi_57_Q_reg_17_inst : DFF_X1 port map( D => n10370, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1585_port, QN 
                           => n_1985);
   DataPath_RF_BLOCKi_57_Q_reg_18_inst : DFF_X1 port map( D => n10369, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1586_port, QN 
                           => n_1986);
   DataPath_RF_BLOCKi_57_Q_reg_19_inst : DFF_X1 port map( D => n10368, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1587_port, QN 
                           => n_1987);
   DataPath_RF_BLOCKi_57_Q_reg_20_inst : DFF_X1 port map( D => n10367, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1588_port, QN 
                           => n_1988);
   DataPath_RF_BLOCKi_57_Q_reg_21_inst : DFF_X1 port map( D => n10366, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1589_port, QN 
                           => n_1989);
   DataPath_RF_BLOCKi_57_Q_reg_22_inst : DFF_X1 port map( D => n10365, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1590_port, QN 
                           => n_1990);
   DataPath_RF_BLOCKi_57_Q_reg_23_inst : DFF_X1 port map( D => n10364, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1591_port, QN 
                           => n_1991);
   DataPath_RF_BLOCKi_57_Q_reg_24_inst : DFF_X1 port map( D => n10363, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1592_port, QN 
                           => n_1992);
   DataPath_RF_BLOCKi_57_Q_reg_25_inst : DFF_X1 port map( D => n10362, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1593_port, QN 
                           => n_1993);
   DataPath_RF_BLOCKi_57_Q_reg_26_inst : DFF_X1 port map( D => n10361, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1594_port, QN 
                           => n_1994);
   DataPath_RF_BLOCKi_57_Q_reg_27_inst : DFF_X1 port map( D => n10360, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1595_port, QN 
                           => n_1995);
   DataPath_RF_BLOCKi_57_Q_reg_28_inst : DFF_X1 port map( D => n10359, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1596_port, QN 
                           => n_1996);
   DataPath_RF_BLOCKi_57_Q_reg_29_inst : DFF_X1 port map( D => n10358, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1597_port, QN 
                           => n_1997);
   DataPath_RF_BLOCKi_57_Q_reg_30_inst : DFF_X1 port map( D => n10357, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1598_port, QN 
                           => n_1998);
   DataPath_RF_BLOCKi_57_Q_reg_31_inst : DFF_X1 port map( D => n10356, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1599_port, QN 
                           => n_1999);
   DataPath_RF_BLOCKi_56_Q_reg_0_inst : DFF_X1 port map( D => n10355, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1536_port, QN => 
                           n_2000);
   DataPath_RF_BLOCKi_56_Q_reg_1_inst : DFF_X1 port map( D => n10354, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1537_port, QN => 
                           n_2001);
   DataPath_RF_BLOCKi_56_Q_reg_2_inst : DFF_X1 port map( D => n10353, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1538_port, QN => 
                           n_2002);
   DataPath_RF_BLOCKi_56_Q_reg_3_inst : DFF_X1 port map( D => n10352, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1539_port, QN => 
                           n_2003);
   DataPath_RF_BLOCKi_56_Q_reg_4_inst : DFF_X1 port map( D => n10351, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1540_port, QN => 
                           n_2004);
   DataPath_RF_BLOCKi_56_Q_reg_5_inst : DFF_X1 port map( D => n10350, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1541_port, QN => 
                           n_2005);
   DataPath_RF_BLOCKi_56_Q_reg_6_inst : DFF_X1 port map( D => n10349, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1542_port, QN => 
                           n_2006);
   DataPath_RF_BLOCKi_56_Q_reg_7_inst : DFF_X1 port map( D => n10348, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1543_port, QN => 
                           n_2007);
   DataPath_RF_BLOCKi_56_Q_reg_8_inst : DFF_X1 port map( D => n10347, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1544_port, QN => 
                           n_2008);
   DataPath_RF_BLOCKi_56_Q_reg_9_inst : DFF_X1 port map( D => n10346, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1545_port, QN => 
                           n_2009);
   DataPath_RF_BLOCKi_56_Q_reg_10_inst : DFF_X1 port map( D => n10345, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1546_port, QN 
                           => n_2010);
   DataPath_RF_BLOCKi_56_Q_reg_11_inst : DFF_X1 port map( D => n10344, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1547_port, QN 
                           => n_2011);
   DataPath_RF_BLOCKi_56_Q_reg_12_inst : DFF_X1 port map( D => n10343, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1548_port, QN 
                           => n_2012);
   DataPath_RF_BLOCKi_56_Q_reg_13_inst : DFF_X1 port map( D => n10342, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1549_port, QN 
                           => n_2013);
   DataPath_RF_BLOCKi_56_Q_reg_14_inst : DFF_X1 port map( D => n10341, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1550_port, QN 
                           => n_2014);
   DataPath_RF_BLOCKi_56_Q_reg_15_inst : DFF_X1 port map( D => n10340, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1551_port, QN 
                           => n_2015);
   DataPath_RF_BLOCKi_56_Q_reg_16_inst : DFF_X1 port map( D => n10339, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1552_port, QN 
                           => n_2016);
   DataPath_RF_BLOCKi_56_Q_reg_17_inst : DFF_X1 port map( D => n10338, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1553_port, QN 
                           => n_2017);
   DataPath_RF_BLOCKi_56_Q_reg_18_inst : DFF_X1 port map( D => n10337, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1554_port, QN 
                           => n_2018);
   DataPath_RF_BLOCKi_56_Q_reg_19_inst : DFF_X1 port map( D => n10336, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1555_port, QN 
                           => n_2019);
   DataPath_RF_BLOCKi_56_Q_reg_20_inst : DFF_X1 port map( D => n10335, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1556_port, QN 
                           => n_2020);
   DataPath_RF_BLOCKi_56_Q_reg_21_inst : DFF_X1 port map( D => n10334, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1557_port, QN 
                           => n_2021);
   DataPath_RF_BLOCKi_56_Q_reg_22_inst : DFF_X1 port map( D => n10333, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1558_port, QN 
                           => n_2022);
   DataPath_RF_BLOCKi_56_Q_reg_23_inst : DFF_X1 port map( D => n10332, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1559_port, QN 
                           => n_2023);
   DataPath_RF_BLOCKi_56_Q_reg_24_inst : DFF_X1 port map( D => n10331, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1560_port, QN 
                           => n_2024);
   DataPath_RF_BLOCKi_56_Q_reg_25_inst : DFF_X1 port map( D => n10330, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1561_port, QN 
                           => n_2025);
   DataPath_RF_BLOCKi_56_Q_reg_26_inst : DFF_X1 port map( D => n10329, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1562_port, QN 
                           => n_2026);
   DataPath_RF_BLOCKi_56_Q_reg_27_inst : DFF_X1 port map( D => n10328, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1563_port, QN 
                           => n_2027);
   DataPath_RF_BLOCKi_56_Q_reg_28_inst : DFF_X1 port map( D => n10327, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1564_port, QN 
                           => n_2028);
   DataPath_RF_BLOCKi_56_Q_reg_29_inst : DFF_X1 port map( D => n10326, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1565_port, QN 
                           => n_2029);
   DataPath_RF_BLOCKi_56_Q_reg_30_inst : DFF_X1 port map( D => n10325, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1566_port, QN 
                           => n_2030);
   DataPath_RF_BLOCKi_56_Q_reg_31_inst : DFF_X1 port map( D => n10324, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1567_port, QN 
                           => n_2031);
   DataPath_RF_BLOCKi_55_Q_reg_0_inst : DFF_X1 port map( D => n10323, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1504_port, QN => 
                           n_2032);
   DataPath_RF_BLOCKi_55_Q_reg_1_inst : DFF_X1 port map( D => n10322, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1505_port, QN => 
                           n_2033);
   DataPath_RF_BLOCKi_55_Q_reg_2_inst : DFF_X1 port map( D => n10321, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1506_port, QN => 
                           n_2034);
   DataPath_RF_BLOCKi_55_Q_reg_3_inst : DFF_X1 port map( D => n10320, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1507_port, QN => 
                           n_2035);
   DataPath_RF_BLOCKi_55_Q_reg_4_inst : DFF_X1 port map( D => n10319, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1508_port, QN => 
                           n_2036);
   DataPath_RF_BLOCKi_55_Q_reg_5_inst : DFF_X1 port map( D => n10318, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1509_port, QN => 
                           n_2037);
   DataPath_RF_BLOCKi_55_Q_reg_6_inst : DFF_X1 port map( D => n10317, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1510_port, QN => 
                           n_2038);
   DataPath_RF_BLOCKi_55_Q_reg_7_inst : DFF_X1 port map( D => n10316, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1511_port, QN => 
                           n_2039);
   DataPath_RF_BLOCKi_55_Q_reg_8_inst : DFF_X1 port map( D => n10315, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1512_port, QN => 
                           n_2040);
   DataPath_RF_BLOCKi_55_Q_reg_9_inst : DFF_X1 port map( D => n10314, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1513_port, QN => 
                           n_2041);
   DataPath_RF_BLOCKi_55_Q_reg_10_inst : DFF_X1 port map( D => n10313, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1514_port, QN 
                           => n_2042);
   DataPath_RF_BLOCKi_55_Q_reg_11_inst : DFF_X1 port map( D => n10312, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1515_port, QN 
                           => n_2043);
   DataPath_RF_BLOCKi_55_Q_reg_12_inst : DFF_X1 port map( D => n10311, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1516_port, QN 
                           => n_2044);
   DataPath_RF_BLOCKi_55_Q_reg_13_inst : DFF_X1 port map( D => n10310, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1517_port, QN 
                           => n_2045);
   DataPath_RF_BLOCKi_55_Q_reg_14_inst : DFF_X1 port map( D => n10309, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1518_port, QN 
                           => n_2046);
   DataPath_RF_BLOCKi_55_Q_reg_15_inst : DFF_X1 port map( D => n10308, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1519_port, QN 
                           => n_2047);
   DataPath_RF_BLOCKi_55_Q_reg_16_inst : DFF_X1 port map( D => n10307, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1520_port, QN 
                           => n_2048);
   DataPath_RF_BLOCKi_55_Q_reg_17_inst : DFF_X1 port map( D => n10306, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1521_port, QN 
                           => n_2049);
   DataPath_RF_BLOCKi_55_Q_reg_18_inst : DFF_X1 port map( D => n10305, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1522_port, QN 
                           => n_2050);
   DataPath_RF_BLOCKi_55_Q_reg_19_inst : DFF_X1 port map( D => n10304, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1523_port, QN 
                           => n_2051);
   DataPath_RF_BLOCKi_55_Q_reg_20_inst : DFF_X1 port map( D => n10303, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1524_port, QN 
                           => n_2052);
   DataPath_RF_BLOCKi_55_Q_reg_21_inst : DFF_X1 port map( D => n10302, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1525_port, QN 
                           => n_2053);
   DataPath_RF_BLOCKi_55_Q_reg_22_inst : DFF_X1 port map( D => n10301, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1526_port, QN 
                           => n_2054);
   DataPath_RF_BLOCKi_55_Q_reg_23_inst : DFF_X1 port map( D => n10300, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1527_port, QN 
                           => n_2055);
   DataPath_RF_BLOCKi_55_Q_reg_24_inst : DFF_X1 port map( D => n10299, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1528_port, QN 
                           => n_2056);
   DataPath_RF_BLOCKi_55_Q_reg_25_inst : DFF_X1 port map( D => n10298, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1529_port, QN 
                           => n_2057);
   DataPath_RF_BLOCKi_55_Q_reg_26_inst : DFF_X1 port map( D => n10297, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1530_port, QN 
                           => n_2058);
   DataPath_RF_BLOCKi_55_Q_reg_27_inst : DFF_X1 port map( D => n10296, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1531_port, QN 
                           => n_2059);
   DataPath_RF_BLOCKi_55_Q_reg_28_inst : DFF_X1 port map( D => n10295, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1532_port, QN 
                           => n_2060);
   DataPath_RF_BLOCKi_55_Q_reg_29_inst : DFF_X1 port map( D => n10294, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1533_port, QN 
                           => n_2061);
   DataPath_RF_BLOCKi_55_Q_reg_30_inst : DFF_X1 port map( D => n10293, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1534_port, QN 
                           => n_2062);
   DataPath_RF_BLOCKi_55_Q_reg_31_inst : DFF_X1 port map( D => n10292, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1535_port, QN 
                           => n_2063);
   DataPath_RF_BLOCKi_54_Q_reg_0_inst : DFF_X1 port map( D => n10291, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1472_port, QN => 
                           n_2064);
   DataPath_RF_BLOCKi_54_Q_reg_1_inst : DFF_X1 port map( D => n10290, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1473_port, QN => 
                           n_2065);
   DataPath_RF_BLOCKi_54_Q_reg_2_inst : DFF_X1 port map( D => n10289, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1474_port, QN => 
                           n_2066);
   DataPath_RF_BLOCKi_54_Q_reg_3_inst : DFF_X1 port map( D => n10288, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1475_port, QN => 
                           n_2067);
   DataPath_RF_BLOCKi_54_Q_reg_4_inst : DFF_X1 port map( D => n10287, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1476_port, QN => 
                           n_2068);
   DataPath_RF_BLOCKi_54_Q_reg_5_inst : DFF_X1 port map( D => n10286, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1477_port, QN => 
                           n_2069);
   DataPath_RF_BLOCKi_54_Q_reg_6_inst : DFF_X1 port map( D => n10285, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1478_port, QN => 
                           n_2070);
   DataPath_RF_BLOCKi_54_Q_reg_7_inst : DFF_X1 port map( D => n10284, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1479_port, QN => 
                           n_2071);
   DataPath_RF_BLOCKi_54_Q_reg_8_inst : DFF_X1 port map( D => n10283, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1480_port, QN => 
                           n_2072);
   DataPath_RF_BLOCKi_54_Q_reg_9_inst : DFF_X1 port map( D => n10282, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1481_port, QN => 
                           n_2073);
   DataPath_RF_BLOCKi_54_Q_reg_10_inst : DFF_X1 port map( D => n10281, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1482_port, QN 
                           => n_2074);
   DataPath_RF_BLOCKi_54_Q_reg_11_inst : DFF_X1 port map( D => n10280, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1483_port, QN 
                           => n_2075);
   DataPath_RF_BLOCKi_54_Q_reg_12_inst : DFF_X1 port map( D => n10279, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1484_port, QN 
                           => n_2076);
   DataPath_RF_BLOCKi_54_Q_reg_13_inst : DFF_X1 port map( D => n10278, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1485_port, QN 
                           => n_2077);
   DataPath_RF_BLOCKi_54_Q_reg_14_inst : DFF_X1 port map( D => n10277, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1486_port, QN 
                           => n_2078);
   DataPath_RF_BLOCKi_54_Q_reg_15_inst : DFF_X1 port map( D => n10276, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1487_port, QN 
                           => n_2079);
   DataPath_RF_BLOCKi_54_Q_reg_16_inst : DFF_X1 port map( D => n10275, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1488_port, QN 
                           => n_2080);
   DataPath_RF_BLOCKi_54_Q_reg_17_inst : DFF_X1 port map( D => n10274, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1489_port, QN 
                           => n_2081);
   DataPath_RF_BLOCKi_54_Q_reg_18_inst : DFF_X1 port map( D => n10273, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1490_port, QN 
                           => n_2082);
   DataPath_RF_BLOCKi_54_Q_reg_19_inst : DFF_X1 port map( D => n10272, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1491_port, QN 
                           => n_2083);
   DataPath_RF_BLOCKi_54_Q_reg_20_inst : DFF_X1 port map( D => n10271, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1492_port, QN 
                           => n_2084);
   DataPath_RF_BLOCKi_54_Q_reg_21_inst : DFF_X1 port map( D => n10270, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1493_port, QN 
                           => n_2085);
   DataPath_RF_BLOCKi_54_Q_reg_22_inst : DFF_X1 port map( D => n10269, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1494_port, QN 
                           => n_2086);
   DataPath_RF_BLOCKi_54_Q_reg_23_inst : DFF_X1 port map( D => n10268, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1495_port, QN 
                           => n_2087);
   DataPath_RF_BLOCKi_54_Q_reg_24_inst : DFF_X1 port map( D => n10267, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1496_port, QN 
                           => n_2088);
   DataPath_RF_BLOCKi_54_Q_reg_25_inst : DFF_X1 port map( D => n10266, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1497_port, QN 
                           => n_2089);
   DataPath_RF_BLOCKi_54_Q_reg_26_inst : DFF_X1 port map( D => n10265, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1498_port, QN 
                           => n_2090);
   DataPath_RF_BLOCKi_54_Q_reg_27_inst : DFF_X1 port map( D => n10264, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1499_port, QN 
                           => n_2091);
   DataPath_RF_BLOCKi_54_Q_reg_28_inst : DFF_X1 port map( D => n10263, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1500_port, QN 
                           => n_2092);
   DataPath_RF_BLOCKi_54_Q_reg_29_inst : DFF_X1 port map( D => n10262, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1501_port, QN 
                           => n_2093);
   DataPath_RF_BLOCKi_54_Q_reg_30_inst : DFF_X1 port map( D => n10261, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1502_port, QN 
                           => n_2094);
   DataPath_RF_BLOCKi_54_Q_reg_31_inst : DFF_X1 port map( D => n10260, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1503_port, QN 
                           => n_2095);
   DataPath_RF_BLOCKi_53_Q_reg_0_inst : DFF_X1 port map( D => n10259, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1440_port, QN => 
                           n_2096);
   DataPath_RF_BLOCKi_53_Q_reg_1_inst : DFF_X1 port map( D => n10258, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1441_port, QN => 
                           n_2097);
   DataPath_RF_BLOCKi_53_Q_reg_2_inst : DFF_X1 port map( D => n10257, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1442_port, QN => 
                           n_2098);
   DataPath_RF_BLOCKi_53_Q_reg_3_inst : DFF_X1 port map( D => n10256, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1443_port, QN => 
                           n_2099);
   DataPath_RF_BLOCKi_53_Q_reg_4_inst : DFF_X1 port map( D => n10255, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1444_port, QN => 
                           n_2100);
   DataPath_RF_BLOCKi_53_Q_reg_5_inst : DFF_X1 port map( D => n10254, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1445_port, QN => 
                           n_2101);
   DataPath_RF_BLOCKi_53_Q_reg_6_inst : DFF_X1 port map( D => n10253, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1446_port, QN => 
                           n_2102);
   DataPath_RF_BLOCKi_53_Q_reg_7_inst : DFF_X1 port map( D => n10252, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1447_port, QN => 
                           n_2103);
   DataPath_RF_BLOCKi_53_Q_reg_8_inst : DFF_X1 port map( D => n10251, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1448_port, QN => 
                           n_2104);
   DataPath_RF_BLOCKi_53_Q_reg_9_inst : DFF_X1 port map( D => n10250, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1449_port, QN => 
                           n_2105);
   DataPath_RF_BLOCKi_53_Q_reg_10_inst : DFF_X1 port map( D => n10249, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1450_port, QN 
                           => n_2106);
   DataPath_RF_BLOCKi_53_Q_reg_11_inst : DFF_X1 port map( D => n10248, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1451_port, QN 
                           => n_2107);
   DataPath_RF_BLOCKi_53_Q_reg_12_inst : DFF_X1 port map( D => n10247, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1452_port, QN 
                           => n_2108);
   DataPath_RF_BLOCKi_53_Q_reg_13_inst : DFF_X1 port map( D => n10246, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1453_port, QN 
                           => n_2109);
   DataPath_RF_BLOCKi_53_Q_reg_14_inst : DFF_X1 port map( D => n10245, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1454_port, QN 
                           => n_2110);
   DataPath_RF_BLOCKi_53_Q_reg_15_inst : DFF_X1 port map( D => n10244, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1455_port, QN 
                           => n_2111);
   DataPath_RF_BLOCKi_53_Q_reg_16_inst : DFF_X1 port map( D => n10243, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1456_port, QN 
                           => n_2112);
   DataPath_RF_BLOCKi_53_Q_reg_17_inst : DFF_X1 port map( D => n10242, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1457_port, QN 
                           => n_2113);
   DataPath_RF_BLOCKi_53_Q_reg_18_inst : DFF_X1 port map( D => n10241, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1458_port, QN 
                           => n_2114);
   DataPath_RF_BLOCKi_53_Q_reg_19_inst : DFF_X1 port map( D => n10240, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1459_port, QN 
                           => n_2115);
   DataPath_RF_BLOCKi_53_Q_reg_20_inst : DFF_X1 port map( D => n10239, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1460_port, QN 
                           => n_2116);
   DataPath_RF_BLOCKi_53_Q_reg_21_inst : DFF_X1 port map( D => n10238, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1461_port, QN 
                           => n_2117);
   DataPath_RF_BLOCKi_53_Q_reg_22_inst : DFF_X1 port map( D => n10237, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1462_port, QN 
                           => n_2118);
   DataPath_RF_BLOCKi_53_Q_reg_23_inst : DFF_X1 port map( D => n10236, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1463_port, QN 
                           => n_2119);
   DataPath_RF_BLOCKi_53_Q_reg_24_inst : DFF_X1 port map( D => n10235, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1464_port, QN 
                           => n_2120);
   DataPath_RF_BLOCKi_53_Q_reg_25_inst : DFF_X1 port map( D => n10234, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1465_port, QN 
                           => n_2121);
   DataPath_RF_BLOCKi_53_Q_reg_26_inst : DFF_X1 port map( D => n10233, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1466_port, QN 
                           => n_2122);
   DataPath_RF_BLOCKi_53_Q_reg_27_inst : DFF_X1 port map( D => n10232, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1467_port, QN 
                           => n_2123);
   DataPath_RF_BLOCKi_53_Q_reg_28_inst : DFF_X1 port map( D => n10231, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1468_port, QN 
                           => n_2124);
   DataPath_RF_BLOCKi_53_Q_reg_29_inst : DFF_X1 port map( D => n10230, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1469_port, QN 
                           => n_2125);
   DataPath_RF_BLOCKi_53_Q_reg_30_inst : DFF_X1 port map( D => n10229, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1470_port, QN 
                           => n_2126);
   DataPath_RF_BLOCKi_53_Q_reg_31_inst : DFF_X1 port map( D => n10228, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1471_port, QN 
                           => n_2127);
   DataPath_RF_BLOCKi_52_Q_reg_0_inst : DFF_X1 port map( D => n10227, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1408_port, QN => 
                           n_2128);
   DataPath_RF_BLOCKi_52_Q_reg_1_inst : DFF_X1 port map( D => n10226, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1409_port, QN => 
                           n_2129);
   DataPath_RF_BLOCKi_52_Q_reg_2_inst : DFF_X1 port map( D => n10225, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1410_port, QN => 
                           n_2130);
   DataPath_RF_BLOCKi_52_Q_reg_3_inst : DFF_X1 port map( D => n10224, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1411_port, QN => 
                           n_2131);
   DataPath_RF_BLOCKi_52_Q_reg_4_inst : DFF_X1 port map( D => n10223, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1412_port, QN => 
                           n_2132);
   DataPath_RF_BLOCKi_52_Q_reg_5_inst : DFF_X1 port map( D => n10222, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1413_port, QN => 
                           n_2133);
   DataPath_RF_BLOCKi_52_Q_reg_6_inst : DFF_X1 port map( D => n10221, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1414_port, QN => 
                           n_2134);
   DataPath_RF_BLOCKi_52_Q_reg_7_inst : DFF_X1 port map( D => n10220, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1415_port, QN => 
                           n_2135);
   DataPath_RF_BLOCKi_52_Q_reg_8_inst : DFF_X1 port map( D => n10219, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1416_port, QN => 
                           n_2136);
   DataPath_RF_BLOCKi_52_Q_reg_9_inst : DFF_X1 port map( D => n10218, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1417_port, QN => 
                           n_2137);
   DataPath_RF_BLOCKi_52_Q_reg_10_inst : DFF_X1 port map( D => n10217, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1418_port, QN 
                           => n_2138);
   DataPath_RF_BLOCKi_52_Q_reg_11_inst : DFF_X1 port map( D => n10216, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1419_port, QN 
                           => n_2139);
   DataPath_RF_BLOCKi_52_Q_reg_12_inst : DFF_X1 port map( D => n10215, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1420_port, QN 
                           => n_2140);
   DataPath_RF_BLOCKi_52_Q_reg_13_inst : DFF_X1 port map( D => n10214, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1421_port, QN 
                           => n_2141);
   DataPath_RF_BLOCKi_52_Q_reg_14_inst : DFF_X1 port map( D => n10213, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1422_port, QN 
                           => n_2142);
   DataPath_RF_BLOCKi_52_Q_reg_15_inst : DFF_X1 port map( D => n10212, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1423_port, QN 
                           => n_2143);
   DataPath_RF_BLOCKi_52_Q_reg_16_inst : DFF_X1 port map( D => n10211, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1424_port, QN 
                           => n_2144);
   DataPath_RF_BLOCKi_52_Q_reg_17_inst : DFF_X1 port map( D => n10210, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1425_port, QN 
                           => n_2145);
   DataPath_RF_BLOCKi_52_Q_reg_18_inst : DFF_X1 port map( D => n10209, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1426_port, QN 
                           => n_2146);
   DataPath_RF_BLOCKi_52_Q_reg_19_inst : DFF_X1 port map( D => n10208, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1427_port, QN 
                           => n_2147);
   DataPath_RF_BLOCKi_52_Q_reg_20_inst : DFF_X1 port map( D => n10207, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1428_port, QN 
                           => n_2148);
   DataPath_RF_BLOCKi_52_Q_reg_21_inst : DFF_X1 port map( D => n10206, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1429_port, QN 
                           => n_2149);
   DataPath_RF_BLOCKi_52_Q_reg_22_inst : DFF_X1 port map( D => n10205, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1430_port, QN 
                           => n_2150);
   DataPath_RF_BLOCKi_52_Q_reg_23_inst : DFF_X1 port map( D => n10204, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1431_port, QN 
                           => n_2151);
   DataPath_RF_BLOCKi_52_Q_reg_24_inst : DFF_X1 port map( D => n10203, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1432_port, QN 
                           => n_2152);
   DataPath_RF_BLOCKi_52_Q_reg_25_inst : DFF_X1 port map( D => n10202, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1433_port, QN 
                           => n_2153);
   DataPath_RF_BLOCKi_52_Q_reg_26_inst : DFF_X1 port map( D => n10201, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1434_port, QN 
                           => n_2154);
   DataPath_RF_BLOCKi_52_Q_reg_27_inst : DFF_X1 port map( D => n10200, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1435_port, QN 
                           => n_2155);
   DataPath_RF_BLOCKi_52_Q_reg_28_inst : DFF_X1 port map( D => n10199, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1436_port, QN 
                           => n_2156);
   DataPath_RF_BLOCKi_52_Q_reg_29_inst : DFF_X1 port map( D => n10198, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1437_port, QN 
                           => n_2157);
   DataPath_RF_BLOCKi_52_Q_reg_30_inst : DFF_X1 port map( D => n10197, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1438_port, QN 
                           => n_2158);
   DataPath_RF_BLOCKi_52_Q_reg_31_inst : DFF_X1 port map( D => n10196, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1439_port, QN 
                           => n_2159);
   DataPath_RF_BLOCKi_51_Q_reg_0_inst : DFF_X1 port map( D => n10195, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1376_port, QN => 
                           n_2160);
   DataPath_RF_BLOCKi_51_Q_reg_1_inst : DFF_X1 port map( D => n10194, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1377_port, QN => 
                           n_2161);
   DataPath_RF_BLOCKi_51_Q_reg_2_inst : DFF_X1 port map( D => n10193, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1378_port, QN => 
                           n_2162);
   DataPath_RF_BLOCKi_51_Q_reg_3_inst : DFF_X1 port map( D => n10192, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1379_port, QN => 
                           n_2163);
   DataPath_RF_BLOCKi_51_Q_reg_4_inst : DFF_X1 port map( D => n10191, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1380_port, QN => 
                           n_2164);
   DataPath_RF_BLOCKi_51_Q_reg_5_inst : DFF_X1 port map( D => n10190, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1381_port, QN => 
                           n_2165);
   DataPath_RF_BLOCKi_51_Q_reg_6_inst : DFF_X1 port map( D => n10189, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1382_port, QN => 
                           n_2166);
   DataPath_RF_BLOCKi_51_Q_reg_7_inst : DFF_X1 port map( D => n10188, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1383_port, QN => 
                           n_2167);
   DataPath_RF_BLOCKi_51_Q_reg_8_inst : DFF_X1 port map( D => n10187, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1384_port, QN => 
                           n_2168);
   DataPath_RF_BLOCKi_51_Q_reg_9_inst : DFF_X1 port map( D => n10186, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1385_port, QN => 
                           n_2169);
   DataPath_RF_BLOCKi_51_Q_reg_10_inst : DFF_X1 port map( D => n10185, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1386_port, QN 
                           => n_2170);
   DataPath_RF_BLOCKi_51_Q_reg_11_inst : DFF_X1 port map( D => n10184, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1387_port, QN 
                           => n_2171);
   DataPath_RF_BLOCKi_51_Q_reg_12_inst : DFF_X1 port map( D => n10183, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1388_port, QN 
                           => n_2172);
   DataPath_RF_BLOCKi_51_Q_reg_13_inst : DFF_X1 port map( D => n10182, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1389_port, QN 
                           => n_2173);
   DataPath_RF_BLOCKi_51_Q_reg_14_inst : DFF_X1 port map( D => n10181, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1390_port, QN 
                           => n_2174);
   DataPath_RF_BLOCKi_51_Q_reg_15_inst : DFF_X1 port map( D => n10180, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1391_port, QN 
                           => n_2175);
   DataPath_RF_BLOCKi_51_Q_reg_16_inst : DFF_X1 port map( D => n10179, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1392_port, QN 
                           => n_2176);
   DataPath_RF_BLOCKi_51_Q_reg_17_inst : DFF_X1 port map( D => n10178, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1393_port, QN 
                           => n_2177);
   DataPath_RF_BLOCKi_51_Q_reg_18_inst : DFF_X1 port map( D => n10177, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1394_port, QN 
                           => n_2178);
   DataPath_RF_BLOCKi_51_Q_reg_19_inst : DFF_X1 port map( D => n10176, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1395_port, QN 
                           => n_2179);
   DataPath_RF_BLOCKi_51_Q_reg_20_inst : DFF_X1 port map( D => n10175, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1396_port, QN 
                           => n_2180);
   DataPath_RF_BLOCKi_51_Q_reg_21_inst : DFF_X1 port map( D => n10174, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1397_port, QN 
                           => n_2181);
   DataPath_RF_BLOCKi_51_Q_reg_22_inst : DFF_X1 port map( D => n10173, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1398_port, QN 
                           => n_2182);
   DataPath_RF_BLOCKi_51_Q_reg_23_inst : DFF_X1 port map( D => n10172, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1399_port, QN 
                           => n_2183);
   DataPath_RF_BLOCKi_51_Q_reg_24_inst : DFF_X1 port map( D => n10171, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1400_port, QN 
                           => n_2184);
   DataPath_RF_BLOCKi_51_Q_reg_25_inst : DFF_X1 port map( D => n10170, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1401_port, QN 
                           => n_2185);
   DataPath_RF_BLOCKi_51_Q_reg_26_inst : DFF_X1 port map( D => n10169, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1402_port, QN 
                           => n_2186);
   DataPath_RF_BLOCKi_51_Q_reg_27_inst : DFF_X1 port map( D => n10168, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1403_port, QN 
                           => n_2187);
   DataPath_RF_BLOCKi_51_Q_reg_28_inst : DFF_X1 port map( D => n10167, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1404_port, QN 
                           => n_2188);
   DataPath_RF_BLOCKi_51_Q_reg_29_inst : DFF_X1 port map( D => n10166, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1405_port, QN 
                           => n_2189);
   DataPath_RF_BLOCKi_51_Q_reg_30_inst : DFF_X1 port map( D => n10165, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1406_port, QN 
                           => n_2190);
   DataPath_RF_BLOCKi_51_Q_reg_31_inst : DFF_X1 port map( D => n10164, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1407_port, QN 
                           => n_2191);
   DataPath_RF_BLOCKi_50_Q_reg_0_inst : DFF_X1 port map( D => n10163, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1344_port, QN => 
                           n_2192);
   DataPath_RF_BLOCKi_50_Q_reg_1_inst : DFF_X1 port map( D => n10162, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1345_port, QN => 
                           n_2193);
   DataPath_RF_BLOCKi_50_Q_reg_2_inst : DFF_X1 port map( D => n10161, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1346_port, QN => 
                           n_2194);
   DataPath_RF_BLOCKi_50_Q_reg_3_inst : DFF_X1 port map( D => n10160, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1347_port, QN => 
                           n_2195);
   DataPath_RF_BLOCKi_50_Q_reg_4_inst : DFF_X1 port map( D => n10159, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1348_port, QN => 
                           n_2196);
   DataPath_RF_BLOCKi_50_Q_reg_5_inst : DFF_X1 port map( D => n10158, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1349_port, QN => 
                           n_2197);
   DataPath_RF_BLOCKi_50_Q_reg_6_inst : DFF_X1 port map( D => n10157, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1350_port, QN => 
                           n_2198);
   DataPath_RF_BLOCKi_50_Q_reg_7_inst : DFF_X1 port map( D => n10156, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1351_port, QN => 
                           n_2199);
   DataPath_RF_BLOCKi_50_Q_reg_8_inst : DFF_X1 port map( D => n10155, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1352_port, QN => 
                           n_2200);
   DataPath_RF_BLOCKi_50_Q_reg_9_inst : DFF_X1 port map( D => n10154, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1353_port, QN => 
                           n_2201);
   DataPath_RF_BLOCKi_50_Q_reg_10_inst : DFF_X1 port map( D => n10153, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1354_port, QN 
                           => n_2202);
   DataPath_RF_BLOCKi_50_Q_reg_11_inst : DFF_X1 port map( D => n10152, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1355_port, QN 
                           => n_2203);
   DataPath_RF_BLOCKi_50_Q_reg_12_inst : DFF_X1 port map( D => n10151, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1356_port, QN 
                           => n_2204);
   DataPath_RF_BLOCKi_50_Q_reg_13_inst : DFF_X1 port map( D => n10150, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1357_port, QN 
                           => n_2205);
   DataPath_RF_BLOCKi_50_Q_reg_14_inst : DFF_X1 port map( D => n10149, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1358_port, QN 
                           => n_2206);
   DataPath_RF_BLOCKi_50_Q_reg_15_inst : DFF_X1 port map( D => n10148, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1359_port, QN 
                           => n_2207);
   DataPath_RF_BLOCKi_50_Q_reg_16_inst : DFF_X1 port map( D => n10147, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1360_port, QN 
                           => n_2208);
   DataPath_RF_BLOCKi_50_Q_reg_17_inst : DFF_X1 port map( D => n10146, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1361_port, QN 
                           => n_2209);
   DataPath_RF_BLOCKi_50_Q_reg_18_inst : DFF_X1 port map( D => n10145, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1362_port, QN 
                           => n_2210);
   DataPath_RF_BLOCKi_50_Q_reg_19_inst : DFF_X1 port map( D => n10144, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1363_port, QN 
                           => n_2211);
   DataPath_RF_BLOCKi_50_Q_reg_20_inst : DFF_X1 port map( D => n10143, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1364_port, QN 
                           => n_2212);
   DataPath_RF_BLOCKi_50_Q_reg_21_inst : DFF_X1 port map( D => n10142, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1365_port, QN 
                           => n_2213);
   DataPath_RF_BLOCKi_50_Q_reg_22_inst : DFF_X1 port map( D => n10141, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1366_port, QN 
                           => n_2214);
   DataPath_RF_BLOCKi_50_Q_reg_23_inst : DFF_X1 port map( D => n10140, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1367_port, QN 
                           => n_2215);
   DataPath_RF_BLOCKi_50_Q_reg_24_inst : DFF_X1 port map( D => n10139, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1368_port, QN 
                           => n_2216);
   DataPath_RF_BLOCKi_50_Q_reg_25_inst : DFF_X1 port map( D => n10138, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1369_port, QN 
                           => n_2217);
   DataPath_RF_BLOCKi_50_Q_reg_26_inst : DFF_X1 port map( D => n10137, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1370_port, QN 
                           => n_2218);
   DataPath_RF_BLOCKi_50_Q_reg_27_inst : DFF_X1 port map( D => n10136, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1371_port, QN 
                           => n_2219);
   DataPath_RF_BLOCKi_50_Q_reg_28_inst : DFF_X1 port map( D => n10135, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1372_port, QN 
                           => n_2220);
   DataPath_RF_BLOCKi_50_Q_reg_29_inst : DFF_X1 port map( D => n10134, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1373_port, QN 
                           => n_2221);
   DataPath_RF_BLOCKi_50_Q_reg_30_inst : DFF_X1 port map( D => n10133, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1374_port, QN 
                           => n_2222);
   DataPath_RF_BLOCKi_50_Q_reg_31_inst : DFF_X1 port map( D => n10132, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1375_port, QN 
                           => n_2223);
   DataPath_RF_BLOCKi_49_Q_reg_0_inst : DFF_X1 port map( D => n10131, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1312_port, QN => 
                           n_2224);
   DataPath_RF_BLOCKi_49_Q_reg_1_inst : DFF_X1 port map( D => n10130, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1313_port, QN => 
                           n_2225);
   DataPath_RF_BLOCKi_49_Q_reg_2_inst : DFF_X1 port map( D => n10129, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1314_port, QN => 
                           n_2226);
   DataPath_RF_BLOCKi_49_Q_reg_3_inst : DFF_X1 port map( D => n10128, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1315_port, QN => 
                           n_2227);
   DataPath_RF_BLOCKi_49_Q_reg_4_inst : DFF_X1 port map( D => n10127, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1316_port, QN => 
                           n_2228);
   DataPath_RF_BLOCKi_49_Q_reg_5_inst : DFF_X1 port map( D => n10126, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1317_port, QN => 
                           n_2229);
   DataPath_RF_BLOCKi_49_Q_reg_6_inst : DFF_X1 port map( D => n10125, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1318_port, QN => 
                           n_2230);
   DataPath_RF_BLOCKi_49_Q_reg_7_inst : DFF_X1 port map( D => n10124, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1319_port, QN => 
                           n_2231);
   DataPath_RF_BLOCKi_49_Q_reg_8_inst : DFF_X1 port map( D => n10123, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1320_port, QN => 
                           n_2232);
   DataPath_RF_BLOCKi_49_Q_reg_9_inst : DFF_X1 port map( D => n10122, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1321_port, QN => 
                           n_2233);
   DataPath_RF_BLOCKi_49_Q_reg_10_inst : DFF_X1 port map( D => n10121, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1322_port, QN 
                           => n_2234);
   DataPath_RF_BLOCKi_49_Q_reg_11_inst : DFF_X1 port map( D => n10120, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1323_port, QN 
                           => n_2235);
   DataPath_RF_BLOCKi_49_Q_reg_12_inst : DFF_X1 port map( D => n10119, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1324_port, QN 
                           => n_2236);
   DataPath_RF_BLOCKi_49_Q_reg_13_inst : DFF_X1 port map( D => n10118, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1325_port, QN 
                           => n_2237);
   DataPath_RF_BLOCKi_49_Q_reg_14_inst : DFF_X1 port map( D => n10117, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1326_port, QN 
                           => n_2238);
   DataPath_RF_BLOCKi_49_Q_reg_15_inst : DFF_X1 port map( D => n10116, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1327_port, QN 
                           => n_2239);
   DataPath_RF_BLOCKi_49_Q_reg_16_inst : DFF_X1 port map( D => n10115, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1328_port, QN 
                           => n_2240);
   DataPath_RF_BLOCKi_49_Q_reg_17_inst : DFF_X1 port map( D => n10114, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1329_port, QN 
                           => n_2241);
   DataPath_RF_BLOCKi_49_Q_reg_18_inst : DFF_X1 port map( D => n10113, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1330_port, QN 
                           => n_2242);
   DataPath_RF_BLOCKi_49_Q_reg_19_inst : DFF_X1 port map( D => n10112, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1331_port, QN 
                           => n_2243);
   DataPath_RF_BLOCKi_49_Q_reg_20_inst : DFF_X1 port map( D => n10111, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1332_port, QN 
                           => n_2244);
   DataPath_RF_BLOCKi_49_Q_reg_21_inst : DFF_X1 port map( D => n10110, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1333_port, QN 
                           => n_2245);
   DataPath_RF_BLOCKi_49_Q_reg_22_inst : DFF_X1 port map( D => n10109, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1334_port, QN 
                           => n_2246);
   DataPath_RF_BLOCKi_49_Q_reg_23_inst : DFF_X1 port map( D => n10108, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1335_port, QN 
                           => n_2247);
   DataPath_RF_BLOCKi_49_Q_reg_24_inst : DFF_X1 port map( D => n10107, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1336_port, QN 
                           => n_2248);
   DataPath_RF_BLOCKi_49_Q_reg_25_inst : DFF_X1 port map( D => n10106, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1337_port, QN 
                           => n_2249);
   DataPath_RF_BLOCKi_49_Q_reg_26_inst : DFF_X1 port map( D => n10105, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1338_port, QN 
                           => n_2250);
   DataPath_RF_BLOCKi_49_Q_reg_27_inst : DFF_X1 port map( D => n10104, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1339_port, QN 
                           => n_2251);
   DataPath_RF_BLOCKi_49_Q_reg_28_inst : DFF_X1 port map( D => n10103, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1340_port, QN 
                           => n_2252);
   DataPath_RF_BLOCKi_49_Q_reg_29_inst : DFF_X1 port map( D => n10102, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1341_port, QN 
                           => n_2253);
   DataPath_RF_BLOCKi_49_Q_reg_30_inst : DFF_X1 port map( D => n10101, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1342_port, QN 
                           => n_2254);
   DataPath_RF_BLOCKi_49_Q_reg_31_inst : DFF_X1 port map( D => n10100, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1343_port, QN 
                           => n_2255);
   DataPath_RF_BLOCKi_48_Q_reg_0_inst : DFF_X1 port map( D => n10099, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1280_port, QN => 
                           n_2256);
   DataPath_RF_BLOCKi_48_Q_reg_1_inst : DFF_X1 port map( D => n10098, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1281_port, QN => 
                           n_2257);
   DataPath_RF_BLOCKi_48_Q_reg_2_inst : DFF_X1 port map( D => n10097, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1282_port, QN => 
                           n_2258);
   DataPath_RF_BLOCKi_48_Q_reg_3_inst : DFF_X1 port map( D => n10096, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1283_port, QN => 
                           n_2259);
   DataPath_RF_BLOCKi_48_Q_reg_4_inst : DFF_X1 port map( D => n10095, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1284_port, QN => 
                           n_2260);
   DataPath_RF_BLOCKi_48_Q_reg_5_inst : DFF_X1 port map( D => n10094, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1285_port, QN => 
                           n_2261);
   DataPath_RF_BLOCKi_48_Q_reg_6_inst : DFF_X1 port map( D => n10093, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1286_port, QN => 
                           n_2262);
   DataPath_RF_BLOCKi_48_Q_reg_7_inst : DFF_X1 port map( D => n10092, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1287_port, QN => 
                           n_2263);
   DataPath_RF_BLOCKi_48_Q_reg_8_inst : DFF_X1 port map( D => n10091, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1288_port, QN => 
                           n_2264);
   DataPath_RF_BLOCKi_48_Q_reg_9_inst : DFF_X1 port map( D => n10090, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1289_port, QN => 
                           n_2265);
   DataPath_RF_BLOCKi_48_Q_reg_10_inst : DFF_X1 port map( D => n10089, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1290_port, QN 
                           => n_2266);
   DataPath_RF_BLOCKi_48_Q_reg_11_inst : DFF_X1 port map( D => n10088, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1291_port, QN 
                           => n_2267);
   DataPath_RF_BLOCKi_48_Q_reg_12_inst : DFF_X1 port map( D => n10087, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1292_port, QN 
                           => n_2268);
   DataPath_RF_BLOCKi_48_Q_reg_13_inst : DFF_X1 port map( D => n10086, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1293_port, QN 
                           => n_2269);
   DataPath_RF_BLOCKi_48_Q_reg_14_inst : DFF_X1 port map( D => n10085, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1294_port, QN 
                           => n_2270);
   DataPath_RF_BLOCKi_48_Q_reg_15_inst : DFF_X1 port map( D => n10084, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1295_port, QN 
                           => n_2271);
   DataPath_RF_BLOCKi_48_Q_reg_16_inst : DFF_X1 port map( D => n10083, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1296_port, QN 
                           => n_2272);
   DataPath_RF_BLOCKi_48_Q_reg_17_inst : DFF_X1 port map( D => n10082, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1297_port, QN 
                           => n_2273);
   DataPath_RF_BLOCKi_48_Q_reg_18_inst : DFF_X1 port map( D => n10081, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1298_port, QN 
                           => n_2274);
   DataPath_RF_BLOCKi_48_Q_reg_19_inst : DFF_X1 port map( D => n10080, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1299_port, QN 
                           => n_2275);
   DataPath_RF_BLOCKi_48_Q_reg_20_inst : DFF_X1 port map( D => n10079, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1300_port, QN 
                           => n_2276);
   DataPath_RF_BLOCKi_48_Q_reg_21_inst : DFF_X1 port map( D => n10078, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1301_port, QN 
                           => n_2277);
   DataPath_RF_BLOCKi_48_Q_reg_22_inst : DFF_X1 port map( D => n10077, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1302_port, QN 
                           => n_2278);
   DataPath_RF_BLOCKi_48_Q_reg_23_inst : DFF_X1 port map( D => n10076, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1303_port, QN 
                           => n_2279);
   DataPath_RF_BLOCKi_48_Q_reg_24_inst : DFF_X1 port map( D => n10075, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1304_port, QN 
                           => n_2280);
   DataPath_RF_BLOCKi_48_Q_reg_25_inst : DFF_X1 port map( D => n10074, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1305_port, QN 
                           => n_2281);
   DataPath_RF_BLOCKi_48_Q_reg_26_inst : DFF_X1 port map( D => n10073, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1306_port, QN 
                           => n_2282);
   DataPath_RF_BLOCKi_48_Q_reg_27_inst : DFF_X1 port map( D => n10072, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1307_port, QN 
                           => n_2283);
   DataPath_RF_BLOCKi_48_Q_reg_28_inst : DFF_X1 port map( D => n10071, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1308_port, QN 
                           => n_2284);
   DataPath_RF_BLOCKi_48_Q_reg_29_inst : DFF_X1 port map( D => n10070, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1309_port, QN 
                           => n_2285);
   DataPath_RF_BLOCKi_48_Q_reg_30_inst : DFF_X1 port map( D => n10069, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1310_port, QN 
                           => n_2286);
   DataPath_RF_BLOCKi_48_Q_reg_31_inst : DFF_X1 port map( D => n10068, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1311_port, QN 
                           => n_2287);
   DataPath_RF_BLOCKi_47_Q_reg_0_inst : DFF_X1 port map( D => n10067, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1248_port, QN => 
                           n_2288);
   DataPath_RF_BLOCKi_47_Q_reg_1_inst : DFF_X1 port map( D => n10066, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1249_port, QN => 
                           n_2289);
   DataPath_RF_BLOCKi_47_Q_reg_2_inst : DFF_X1 port map( D => n10065, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1250_port, QN => 
                           n_2290);
   DataPath_RF_BLOCKi_47_Q_reg_3_inst : DFF_X1 port map( D => n10064, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1251_port, QN => 
                           n_2291);
   DataPath_RF_BLOCKi_47_Q_reg_4_inst : DFF_X1 port map( D => n10063, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1252_port, QN => 
                           n_2292);
   DataPath_RF_BLOCKi_47_Q_reg_5_inst : DFF_X1 port map( D => n10062, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1253_port, QN => 
                           n_2293);
   DataPath_RF_BLOCKi_47_Q_reg_6_inst : DFF_X1 port map( D => n10061, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1254_port, QN => 
                           n_2294);
   DataPath_RF_BLOCKi_47_Q_reg_7_inst : DFF_X1 port map( D => n10060, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1255_port, QN => 
                           n_2295);
   DataPath_RF_BLOCKi_47_Q_reg_8_inst : DFF_X1 port map( D => n10059, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1256_port, QN => 
                           n_2296);
   DataPath_RF_BLOCKi_47_Q_reg_9_inst : DFF_X1 port map( D => n10058, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1257_port, QN => 
                           n_2297);
   DataPath_RF_BLOCKi_47_Q_reg_10_inst : DFF_X1 port map( D => n10057, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1258_port, QN 
                           => n_2298);
   DataPath_RF_BLOCKi_47_Q_reg_11_inst : DFF_X1 port map( D => n10056, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1259_port, QN 
                           => n_2299);
   DataPath_RF_BLOCKi_47_Q_reg_12_inst : DFF_X1 port map( D => n10055, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1260_port, QN 
                           => n_2300);
   DataPath_RF_BLOCKi_47_Q_reg_13_inst : DFF_X1 port map( D => n10054, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1261_port, QN 
                           => n_2301);
   DataPath_RF_BLOCKi_47_Q_reg_14_inst : DFF_X1 port map( D => n10053, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1262_port, QN 
                           => n_2302);
   DataPath_RF_BLOCKi_47_Q_reg_15_inst : DFF_X1 port map( D => n10052, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1263_port, QN 
                           => n_2303);
   DataPath_RF_BLOCKi_47_Q_reg_16_inst : DFF_X1 port map( D => n10051, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1264_port, QN 
                           => n_2304);
   DataPath_RF_BLOCKi_47_Q_reg_17_inst : DFF_X1 port map( D => n10050, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1265_port, QN 
                           => n_2305);
   DataPath_RF_BLOCKi_47_Q_reg_18_inst : DFF_X1 port map( D => n10049, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1266_port, QN 
                           => n_2306);
   DataPath_RF_BLOCKi_47_Q_reg_19_inst : DFF_X1 port map( D => n10048, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1267_port, QN 
                           => n_2307);
   DataPath_RF_BLOCKi_47_Q_reg_20_inst : DFF_X1 port map( D => n10047, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1268_port, QN 
                           => n_2308);
   DataPath_RF_BLOCKi_47_Q_reg_21_inst : DFF_X1 port map( D => n10046, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1269_port, QN 
                           => n_2309);
   DataPath_RF_BLOCKi_47_Q_reg_22_inst : DFF_X1 port map( D => n10045, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1270_port, QN 
                           => n_2310);
   DataPath_RF_BLOCKi_47_Q_reg_23_inst : DFF_X1 port map( D => n10044, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1271_port, QN 
                           => n_2311);
   DataPath_RF_BLOCKi_47_Q_reg_24_inst : DFF_X1 port map( D => n10043, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1272_port, QN 
                           => n_2312);
   DataPath_RF_BLOCKi_47_Q_reg_25_inst : DFF_X1 port map( D => n10042, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1273_port, QN 
                           => n_2313);
   DataPath_RF_BLOCKi_47_Q_reg_26_inst : DFF_X1 port map( D => n10041, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1274_port, QN 
                           => n_2314);
   DataPath_RF_BLOCKi_47_Q_reg_27_inst : DFF_X1 port map( D => n10040, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1275_port, QN 
                           => n_2315);
   DataPath_RF_BLOCKi_47_Q_reg_28_inst : DFF_X1 port map( D => n10039, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1276_port, QN 
                           => n_2316);
   DataPath_RF_BLOCKi_47_Q_reg_29_inst : DFF_X1 port map( D => n10038, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1277_port, QN 
                           => n_2317);
   DataPath_RF_BLOCKi_47_Q_reg_30_inst : DFF_X1 port map( D => n10037, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1278_port, QN 
                           => n_2318);
   DataPath_RF_BLOCKi_47_Q_reg_31_inst : DFF_X1 port map( D => n10036, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1279_port, QN 
                           => n_2319);
   DataPath_RF_BLOCKi_46_Q_reg_0_inst : DFF_X1 port map( D => n10035, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1216_port, QN => 
                           n_2320);
   DataPath_RF_BLOCKi_46_Q_reg_1_inst : DFF_X1 port map( D => n10034, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1217_port, QN => 
                           n_2321);
   DataPath_RF_BLOCKi_46_Q_reg_2_inst : DFF_X1 port map( D => n10033, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1218_port, QN => 
                           n_2322);
   DataPath_RF_BLOCKi_46_Q_reg_3_inst : DFF_X1 port map( D => n10032, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1219_port, QN => 
                           n_2323);
   DataPath_RF_BLOCKi_46_Q_reg_4_inst : DFF_X1 port map( D => n10031, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1220_port, QN => 
                           n_2324);
   DataPath_RF_BLOCKi_46_Q_reg_5_inst : DFF_X1 port map( D => n10030, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1221_port, QN => 
                           n_2325);
   DataPath_RF_BLOCKi_46_Q_reg_6_inst : DFF_X1 port map( D => n10029, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1222_port, QN => 
                           n_2326);
   DataPath_RF_BLOCKi_46_Q_reg_7_inst : DFF_X1 port map( D => n10028, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1223_port, QN => 
                           n_2327);
   DataPath_RF_BLOCKi_46_Q_reg_8_inst : DFF_X1 port map( D => n10027, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1224_port, QN => 
                           n_2328);
   DataPath_RF_BLOCKi_46_Q_reg_9_inst : DFF_X1 port map( D => n10026, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1225_port, QN => 
                           n_2329);
   DataPath_RF_BLOCKi_46_Q_reg_10_inst : DFF_X1 port map( D => n10025, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1226_port, QN 
                           => n_2330);
   DataPath_RF_BLOCKi_46_Q_reg_11_inst : DFF_X1 port map( D => n10024, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1227_port, QN 
                           => n_2331);
   DataPath_RF_BLOCKi_46_Q_reg_12_inst : DFF_X1 port map( D => n10023, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1228_port, QN 
                           => n_2332);
   DataPath_RF_BLOCKi_46_Q_reg_13_inst : DFF_X1 port map( D => n10022, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1229_port, QN 
                           => n_2333);
   DataPath_RF_BLOCKi_46_Q_reg_14_inst : DFF_X1 port map( D => n10021, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1230_port, QN 
                           => n_2334);
   DataPath_RF_BLOCKi_46_Q_reg_15_inst : DFF_X1 port map( D => n10020, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1231_port, QN 
                           => n_2335);
   DataPath_RF_BLOCKi_46_Q_reg_16_inst : DFF_X1 port map( D => n10019, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1232_port, QN 
                           => n_2336);
   DataPath_RF_BLOCKi_46_Q_reg_17_inst : DFF_X1 port map( D => n10018, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1233_port, QN 
                           => n_2337);
   DataPath_RF_BLOCKi_46_Q_reg_18_inst : DFF_X1 port map( D => n10017, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1234_port, QN 
                           => n_2338);
   DataPath_RF_BLOCKi_46_Q_reg_19_inst : DFF_X1 port map( D => n10016, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1235_port, QN 
                           => n_2339);
   DataPath_RF_BLOCKi_46_Q_reg_20_inst : DFF_X1 port map( D => n10015, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1236_port, QN 
                           => n_2340);
   DataPath_RF_BLOCKi_46_Q_reg_21_inst : DFF_X1 port map( D => n10014, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1237_port, QN 
                           => n_2341);
   DataPath_RF_BLOCKi_46_Q_reg_22_inst : DFF_X1 port map( D => n10013, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1238_port, QN 
                           => n_2342);
   DataPath_RF_BLOCKi_46_Q_reg_23_inst : DFF_X1 port map( D => n10012, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1239_port, QN 
                           => n_2343);
   DataPath_RF_BLOCKi_46_Q_reg_24_inst : DFF_X1 port map( D => n10011, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1240_port, QN 
                           => n_2344);
   DataPath_RF_BLOCKi_46_Q_reg_25_inst : DFF_X1 port map( D => n10010, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1241_port, QN 
                           => n_2345);
   DataPath_RF_BLOCKi_46_Q_reg_26_inst : DFF_X1 port map( D => n10009, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1242_port, QN 
                           => n_2346);
   DataPath_RF_BLOCKi_46_Q_reg_27_inst : DFF_X1 port map( D => n10008, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1243_port, QN 
                           => n_2347);
   DataPath_RF_BLOCKi_46_Q_reg_28_inst : DFF_X1 port map( D => n10007, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1244_port, QN 
                           => n_2348);
   DataPath_RF_BLOCKi_46_Q_reg_29_inst : DFF_X1 port map( D => n10006, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1245_port, QN 
                           => n_2349);
   DataPath_RF_BLOCKi_46_Q_reg_30_inst : DFF_X1 port map( D => n10005, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1246_port, QN 
                           => n_2350);
   DataPath_RF_BLOCKi_46_Q_reg_31_inst : DFF_X1 port map( D => n10004, CK => 
                           CLK, Q => DataPath_RF_bus_reg_dataout_1247_port, QN 
                           => n_2351);
   DataPath_RF_BLOCKi_45_Q_reg_0_inst : DFF_X1 port map( D => n10003, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1184_port, QN => 
                           n_2352);
   DataPath_RF_BLOCKi_45_Q_reg_1_inst : DFF_X1 port map( D => n10002, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1185_port, QN => 
                           n_2353);
   DataPath_RF_BLOCKi_45_Q_reg_2_inst : DFF_X1 port map( D => n10001, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1186_port, QN => 
                           n_2354);
   DataPath_RF_BLOCKi_45_Q_reg_3_inst : DFF_X1 port map( D => n10000, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1187_port, QN => 
                           n_2355);
   DataPath_RF_BLOCKi_45_Q_reg_4_inst : DFF_X1 port map( D => n9999, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1188_port, QN => 
                           n_2356);
   DataPath_RF_BLOCKi_45_Q_reg_5_inst : DFF_X1 port map( D => n9998, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1189_port, QN => 
                           n_2357);
   DataPath_RF_BLOCKi_45_Q_reg_6_inst : DFF_X1 port map( D => n9997, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1190_port, QN => 
                           n_2358);
   DataPath_RF_BLOCKi_45_Q_reg_7_inst : DFF_X1 port map( D => n9996, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1191_port, QN => 
                           n_2359);
   DataPath_RF_BLOCKi_45_Q_reg_8_inst : DFF_X1 port map( D => n9995, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1192_port, QN => 
                           n_2360);
   DataPath_RF_BLOCKi_45_Q_reg_9_inst : DFF_X1 port map( D => n9994, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1193_port, QN => 
                           n_2361);
   DataPath_RF_BLOCKi_45_Q_reg_10_inst : DFF_X1 port map( D => n9993, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1194_port, QN => 
                           n_2362);
   DataPath_RF_BLOCKi_45_Q_reg_11_inst : DFF_X1 port map( D => n9992, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1195_port, QN => 
                           n_2363);
   DataPath_RF_BLOCKi_45_Q_reg_12_inst : DFF_X1 port map( D => n9991, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1196_port, QN => 
                           n_2364);
   DataPath_RF_BLOCKi_45_Q_reg_13_inst : DFF_X1 port map( D => n9990, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1197_port, QN => 
                           n_2365);
   DataPath_RF_BLOCKi_45_Q_reg_14_inst : DFF_X1 port map( D => n9989, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1198_port, QN => 
                           n_2366);
   DataPath_RF_BLOCKi_45_Q_reg_15_inst : DFF_X1 port map( D => n9988, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1199_port, QN => 
                           n_2367);
   DataPath_RF_BLOCKi_45_Q_reg_16_inst : DFF_X1 port map( D => n9987, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1200_port, QN => 
                           n_2368);
   DataPath_RF_BLOCKi_45_Q_reg_17_inst : DFF_X1 port map( D => n9986, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1201_port, QN => 
                           n_2369);
   DataPath_RF_BLOCKi_45_Q_reg_18_inst : DFF_X1 port map( D => n9985, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1202_port, QN => 
                           n_2370);
   DataPath_RF_BLOCKi_45_Q_reg_19_inst : DFF_X1 port map( D => n9984, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1203_port, QN => 
                           n_2371);
   DataPath_RF_BLOCKi_45_Q_reg_20_inst : DFF_X1 port map( D => n9983, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1204_port, QN => 
                           n_2372);
   DataPath_RF_BLOCKi_45_Q_reg_21_inst : DFF_X1 port map( D => n9982, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1205_port, QN => 
                           n_2373);
   DataPath_RF_BLOCKi_45_Q_reg_22_inst : DFF_X1 port map( D => n9981, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1206_port, QN => 
                           n_2374);
   DataPath_RF_BLOCKi_45_Q_reg_23_inst : DFF_X1 port map( D => n9980, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1207_port, QN => 
                           n_2375);
   DataPath_RF_BLOCKi_45_Q_reg_24_inst : DFF_X1 port map( D => n9979, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1208_port, QN => 
                           n_2376);
   DataPath_RF_BLOCKi_45_Q_reg_25_inst : DFF_X1 port map( D => n9978, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1209_port, QN => 
                           n_2377);
   DataPath_RF_BLOCKi_45_Q_reg_26_inst : DFF_X1 port map( D => n9977, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1210_port, QN => 
                           n_2378);
   DataPath_RF_BLOCKi_45_Q_reg_27_inst : DFF_X1 port map( D => n9976, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1211_port, QN => 
                           n_2379);
   DataPath_RF_BLOCKi_45_Q_reg_28_inst : DFF_X1 port map( D => n9975, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1212_port, QN => 
                           n_2380);
   DataPath_RF_BLOCKi_45_Q_reg_29_inst : DFF_X1 port map( D => n9974, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1213_port, QN => 
                           n_2381);
   DataPath_RF_BLOCKi_45_Q_reg_30_inst : DFF_X1 port map( D => n9973, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1214_port, QN => 
                           n_2382);
   DataPath_RF_BLOCKi_45_Q_reg_31_inst : DFF_X1 port map( D => n9972, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1215_port, QN => 
                           n_2383);
   DataPath_RF_BLOCKi_44_Q_reg_0_inst : DFF_X1 port map( D => n9971, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1152_port, QN => 
                           n_2384);
   DataPath_RF_BLOCKi_44_Q_reg_1_inst : DFF_X1 port map( D => n9970, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1153_port, QN => 
                           n_2385);
   DataPath_RF_BLOCKi_44_Q_reg_2_inst : DFF_X1 port map( D => n9969, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1154_port, QN => 
                           n_2386);
   DataPath_RF_BLOCKi_44_Q_reg_3_inst : DFF_X1 port map( D => n9968, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1155_port, QN => 
                           n_2387);
   DataPath_RF_BLOCKi_44_Q_reg_4_inst : DFF_X1 port map( D => n9967, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1156_port, QN => 
                           n_2388);
   DataPath_RF_BLOCKi_44_Q_reg_5_inst : DFF_X1 port map( D => n9966, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1157_port, QN => 
                           n_2389);
   DataPath_RF_BLOCKi_44_Q_reg_6_inst : DFF_X1 port map( D => n9965, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1158_port, QN => 
                           n_2390);
   DataPath_RF_BLOCKi_44_Q_reg_7_inst : DFF_X1 port map( D => n9964, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1159_port, QN => 
                           n_2391);
   DataPath_RF_BLOCKi_44_Q_reg_8_inst : DFF_X1 port map( D => n9963, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1160_port, QN => 
                           n_2392);
   DataPath_RF_BLOCKi_44_Q_reg_9_inst : DFF_X1 port map( D => n9962, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1161_port, QN => 
                           n_2393);
   DataPath_RF_BLOCKi_44_Q_reg_10_inst : DFF_X1 port map( D => n9961, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1162_port, QN => 
                           n_2394);
   DataPath_RF_BLOCKi_44_Q_reg_11_inst : DFF_X1 port map( D => n9960, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1163_port, QN => 
                           n_2395);
   DataPath_RF_BLOCKi_44_Q_reg_12_inst : DFF_X1 port map( D => n9959, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1164_port, QN => 
                           n_2396);
   DataPath_RF_BLOCKi_44_Q_reg_13_inst : DFF_X1 port map( D => n9958, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1165_port, QN => 
                           n_2397);
   DataPath_RF_BLOCKi_44_Q_reg_14_inst : DFF_X1 port map( D => n9957, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1166_port, QN => 
                           n_2398);
   DataPath_RF_BLOCKi_44_Q_reg_15_inst : DFF_X1 port map( D => n9956, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1167_port, QN => 
                           n_2399);
   DataPath_RF_BLOCKi_44_Q_reg_16_inst : DFF_X1 port map( D => n9955, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1168_port, QN => 
                           n_2400);
   DataPath_RF_BLOCKi_44_Q_reg_17_inst : DFF_X1 port map( D => n9954, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1169_port, QN => 
                           n_2401);
   DataPath_RF_BLOCKi_44_Q_reg_18_inst : DFF_X1 port map( D => n9953, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1170_port, QN => 
                           n_2402);
   DataPath_RF_BLOCKi_44_Q_reg_19_inst : DFF_X1 port map( D => n9952, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1171_port, QN => 
                           n_2403);
   DataPath_RF_BLOCKi_44_Q_reg_20_inst : DFF_X1 port map( D => n9951, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1172_port, QN => 
                           n_2404);
   DataPath_RF_BLOCKi_44_Q_reg_21_inst : DFF_X1 port map( D => n9950, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1173_port, QN => 
                           n_2405);
   DataPath_RF_BLOCKi_44_Q_reg_22_inst : DFF_X1 port map( D => n9949, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1174_port, QN => 
                           n_2406);
   DataPath_RF_BLOCKi_44_Q_reg_23_inst : DFF_X1 port map( D => n9948, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1175_port, QN => 
                           n_2407);
   DataPath_RF_BLOCKi_44_Q_reg_24_inst : DFF_X1 port map( D => n9947, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1176_port, QN => 
                           n_2408);
   DataPath_RF_BLOCKi_44_Q_reg_25_inst : DFF_X1 port map( D => n9946, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1177_port, QN => 
                           n_2409);
   DataPath_RF_BLOCKi_44_Q_reg_26_inst : DFF_X1 port map( D => n9945, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1178_port, QN => 
                           n_2410);
   DataPath_RF_BLOCKi_44_Q_reg_27_inst : DFF_X1 port map( D => n9944, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1179_port, QN => 
                           n_2411);
   DataPath_RF_BLOCKi_44_Q_reg_28_inst : DFF_X1 port map( D => n9943, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1180_port, QN => 
                           n_2412);
   DataPath_RF_BLOCKi_44_Q_reg_29_inst : DFF_X1 port map( D => n9942, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1181_port, QN => 
                           n_2413);
   DataPath_RF_BLOCKi_44_Q_reg_30_inst : DFF_X1 port map( D => n9941, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1182_port, QN => 
                           n_2414);
   DataPath_RF_BLOCKi_44_Q_reg_31_inst : DFF_X1 port map( D => n9940, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1183_port, QN => 
                           n_2415);
   DataPath_RF_BLOCKi_43_Q_reg_0_inst : DFF_X1 port map( D => n9939, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1120_port, QN => 
                           n_2416);
   DataPath_RF_BLOCKi_43_Q_reg_1_inst : DFF_X1 port map( D => n9938, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1121_port, QN => 
                           n_2417);
   DataPath_RF_BLOCKi_43_Q_reg_2_inst : DFF_X1 port map( D => n9937, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1122_port, QN => 
                           n_2418);
   DataPath_RF_BLOCKi_43_Q_reg_3_inst : DFF_X1 port map( D => n9936, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1123_port, QN => 
                           n_2419);
   DataPath_RF_BLOCKi_43_Q_reg_4_inst : DFF_X1 port map( D => n9935, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1124_port, QN => 
                           n_2420);
   DataPath_RF_BLOCKi_43_Q_reg_5_inst : DFF_X1 port map( D => n9934, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1125_port, QN => 
                           n_2421);
   DataPath_RF_BLOCKi_43_Q_reg_6_inst : DFF_X1 port map( D => n9933, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1126_port, QN => 
                           n_2422);
   DataPath_RF_BLOCKi_43_Q_reg_7_inst : DFF_X1 port map( D => n9932, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1127_port, QN => 
                           n_2423);
   DataPath_RF_BLOCKi_43_Q_reg_8_inst : DFF_X1 port map( D => n9931, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1128_port, QN => 
                           n_2424);
   DataPath_RF_BLOCKi_43_Q_reg_9_inst : DFF_X1 port map( D => n9930, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1129_port, QN => 
                           n_2425);
   DataPath_RF_BLOCKi_43_Q_reg_10_inst : DFF_X1 port map( D => n9929, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1130_port, QN => 
                           n_2426);
   DataPath_RF_BLOCKi_43_Q_reg_11_inst : DFF_X1 port map( D => n9928, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1131_port, QN => 
                           n_2427);
   DataPath_RF_BLOCKi_43_Q_reg_12_inst : DFF_X1 port map( D => n9927, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1132_port, QN => 
                           n_2428);
   DataPath_RF_BLOCKi_43_Q_reg_13_inst : DFF_X1 port map( D => n9926, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1133_port, QN => 
                           n_2429);
   DataPath_RF_BLOCKi_43_Q_reg_14_inst : DFF_X1 port map( D => n9925, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1134_port, QN => 
                           n_2430);
   DataPath_RF_BLOCKi_43_Q_reg_15_inst : DFF_X1 port map( D => n9924, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1135_port, QN => 
                           n_2431);
   DataPath_RF_BLOCKi_43_Q_reg_16_inst : DFF_X1 port map( D => n9923, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1136_port, QN => 
                           n_2432);
   DataPath_RF_BLOCKi_43_Q_reg_17_inst : DFF_X1 port map( D => n9922, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1137_port, QN => 
                           n_2433);
   DataPath_RF_BLOCKi_43_Q_reg_18_inst : DFF_X1 port map( D => n9921, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1138_port, QN => 
                           n_2434);
   DataPath_RF_BLOCKi_43_Q_reg_19_inst : DFF_X1 port map( D => n9920, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1139_port, QN => 
                           n_2435);
   DataPath_RF_BLOCKi_43_Q_reg_20_inst : DFF_X1 port map( D => n9919, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1140_port, QN => 
                           n_2436);
   DataPath_RF_BLOCKi_43_Q_reg_21_inst : DFF_X1 port map( D => n9918, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1141_port, QN => 
                           n_2437);
   DataPath_RF_BLOCKi_43_Q_reg_22_inst : DFF_X1 port map( D => n9917, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1142_port, QN => 
                           n_2438);
   DataPath_RF_BLOCKi_43_Q_reg_23_inst : DFF_X1 port map( D => n9916, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1143_port, QN => 
                           n_2439);
   DataPath_RF_BLOCKi_43_Q_reg_24_inst : DFF_X1 port map( D => n9915, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1144_port, QN => 
                           n_2440);
   DataPath_RF_BLOCKi_43_Q_reg_25_inst : DFF_X1 port map( D => n9914, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1145_port, QN => 
                           n_2441);
   DataPath_RF_BLOCKi_43_Q_reg_26_inst : DFF_X1 port map( D => n9913, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1146_port, QN => 
                           n_2442);
   DataPath_RF_BLOCKi_43_Q_reg_27_inst : DFF_X1 port map( D => n9912, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1147_port, QN => 
                           n_2443);
   DataPath_RF_BLOCKi_43_Q_reg_28_inst : DFF_X1 port map( D => n9911, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1148_port, QN => 
                           n_2444);
   DataPath_RF_BLOCKi_43_Q_reg_29_inst : DFF_X1 port map( D => n9910, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1149_port, QN => 
                           n_2445);
   DataPath_RF_BLOCKi_43_Q_reg_30_inst : DFF_X1 port map( D => n9909, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1150_port, QN => 
                           n_2446);
   DataPath_RF_BLOCKi_43_Q_reg_31_inst : DFF_X1 port map( D => n9908, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1151_port, QN => 
                           n_2447);
   DataPath_RF_BLOCKi_42_Q_reg_0_inst : DFF_X1 port map( D => n9907, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1088_port, QN => 
                           n_2448);
   DataPath_RF_BLOCKi_42_Q_reg_1_inst : DFF_X1 port map( D => n9906, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1089_port, QN => 
                           n_2449);
   DataPath_RF_BLOCKi_42_Q_reg_2_inst : DFF_X1 port map( D => n9905, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1090_port, QN => 
                           n_2450);
   DataPath_RF_BLOCKi_42_Q_reg_3_inst : DFF_X1 port map( D => n9904, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1091_port, QN => 
                           n_2451);
   DataPath_RF_BLOCKi_42_Q_reg_4_inst : DFF_X1 port map( D => n9903, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1092_port, QN => 
                           n_2452);
   DataPath_RF_BLOCKi_42_Q_reg_5_inst : DFF_X1 port map( D => n9902, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1093_port, QN => 
                           n_2453);
   DataPath_RF_BLOCKi_42_Q_reg_6_inst : DFF_X1 port map( D => n9901, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1094_port, QN => 
                           n_2454);
   DataPath_RF_BLOCKi_42_Q_reg_7_inst : DFF_X1 port map( D => n9900, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1095_port, QN => 
                           n_2455);
   DataPath_RF_BLOCKi_42_Q_reg_8_inst : DFF_X1 port map( D => n9899, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1096_port, QN => 
                           n_2456);
   DataPath_RF_BLOCKi_42_Q_reg_9_inst : DFF_X1 port map( D => n9898, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1097_port, QN => 
                           n_2457);
   DataPath_RF_BLOCKi_42_Q_reg_10_inst : DFF_X1 port map( D => n9897, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1098_port, QN => 
                           n_2458);
   DataPath_RF_BLOCKi_42_Q_reg_11_inst : DFF_X1 port map( D => n9896, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1099_port, QN => 
                           n_2459);
   DataPath_RF_BLOCKi_42_Q_reg_12_inst : DFF_X1 port map( D => n9895, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1100_port, QN => 
                           n_2460);
   DataPath_RF_BLOCKi_42_Q_reg_13_inst : DFF_X1 port map( D => n9894, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1101_port, QN => 
                           n_2461);
   DataPath_RF_BLOCKi_42_Q_reg_14_inst : DFF_X1 port map( D => n9893, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1102_port, QN => 
                           n_2462);
   DataPath_RF_BLOCKi_42_Q_reg_15_inst : DFF_X1 port map( D => n9892, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1103_port, QN => 
                           n_2463);
   DataPath_RF_BLOCKi_42_Q_reg_16_inst : DFF_X1 port map( D => n9891, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1104_port, QN => 
                           n_2464);
   DataPath_RF_BLOCKi_42_Q_reg_17_inst : DFF_X1 port map( D => n9890, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1105_port, QN => 
                           n_2465);
   DataPath_RF_BLOCKi_42_Q_reg_18_inst : DFF_X1 port map( D => n9889, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1106_port, QN => 
                           n_2466);
   DataPath_RF_BLOCKi_42_Q_reg_19_inst : DFF_X1 port map( D => n9888, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1107_port, QN => 
                           n_2467);
   DataPath_RF_BLOCKi_42_Q_reg_20_inst : DFF_X1 port map( D => n9887, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1108_port, QN => 
                           n_2468);
   DataPath_RF_BLOCKi_42_Q_reg_21_inst : DFF_X1 port map( D => n9886, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1109_port, QN => 
                           n_2469);
   DataPath_RF_BLOCKi_42_Q_reg_22_inst : DFF_X1 port map( D => n9885, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1110_port, QN => 
                           n_2470);
   DataPath_RF_BLOCKi_42_Q_reg_23_inst : DFF_X1 port map( D => n9884, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1111_port, QN => 
                           n_2471);
   DataPath_RF_BLOCKi_42_Q_reg_24_inst : DFF_X1 port map( D => n9883, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1112_port, QN => 
                           n_2472);
   DataPath_RF_BLOCKi_42_Q_reg_25_inst : DFF_X1 port map( D => n9882, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1113_port, QN => 
                           n_2473);
   DataPath_RF_BLOCKi_42_Q_reg_26_inst : DFF_X1 port map( D => n9881, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1114_port, QN => 
                           n_2474);
   DataPath_RF_BLOCKi_42_Q_reg_27_inst : DFF_X1 port map( D => n9880, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1115_port, QN => 
                           n_2475);
   DataPath_RF_BLOCKi_42_Q_reg_28_inst : DFF_X1 port map( D => n9879, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1116_port, QN => 
                           n_2476);
   DataPath_RF_BLOCKi_42_Q_reg_29_inst : DFF_X1 port map( D => n9878, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1117_port, QN => 
                           n_2477);
   DataPath_RF_BLOCKi_42_Q_reg_30_inst : DFF_X1 port map( D => n9877, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1118_port, QN => 
                           n_2478);
   DataPath_RF_BLOCKi_42_Q_reg_31_inst : DFF_X1 port map( D => n9876, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1119_port, QN => 
                           n_2479);
   DataPath_RF_BLOCKi_41_Q_reg_0_inst : DFF_X1 port map( D => n9875, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1056_port, QN => 
                           n_2480);
   DataPath_RF_BLOCKi_41_Q_reg_1_inst : DFF_X1 port map( D => n9874, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1057_port, QN => 
                           n_2481);
   DataPath_RF_BLOCKi_41_Q_reg_2_inst : DFF_X1 port map( D => n9873, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1058_port, QN => 
                           n_2482);
   DataPath_RF_BLOCKi_41_Q_reg_3_inst : DFF_X1 port map( D => n9872, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1059_port, QN => 
                           n_2483);
   DataPath_RF_BLOCKi_41_Q_reg_4_inst : DFF_X1 port map( D => n9871, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1060_port, QN => 
                           n_2484);
   DataPath_RF_BLOCKi_41_Q_reg_5_inst : DFF_X1 port map( D => n9870, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1061_port, QN => 
                           n_2485);
   DataPath_RF_BLOCKi_41_Q_reg_6_inst : DFF_X1 port map( D => n9869, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1062_port, QN => 
                           n_2486);
   DataPath_RF_BLOCKi_41_Q_reg_7_inst : DFF_X1 port map( D => n9868, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1063_port, QN => 
                           n_2487);
   DataPath_RF_BLOCKi_41_Q_reg_8_inst : DFF_X1 port map( D => n9867, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1064_port, QN => 
                           n_2488);
   DataPath_RF_BLOCKi_41_Q_reg_9_inst : DFF_X1 port map( D => n9866, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1065_port, QN => 
                           n_2489);
   DataPath_RF_BLOCKi_41_Q_reg_10_inst : DFF_X1 port map( D => n9865, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1066_port, QN => 
                           n_2490);
   DataPath_RF_BLOCKi_41_Q_reg_11_inst : DFF_X1 port map( D => n9864, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1067_port, QN => 
                           n_2491);
   DataPath_RF_BLOCKi_41_Q_reg_12_inst : DFF_X1 port map( D => n9863, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1068_port, QN => 
                           n_2492);
   DataPath_RF_BLOCKi_41_Q_reg_13_inst : DFF_X1 port map( D => n9862, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1069_port, QN => 
                           n_2493);
   DataPath_RF_BLOCKi_41_Q_reg_14_inst : DFF_X1 port map( D => n9861, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1070_port, QN => 
                           n_2494);
   DataPath_RF_BLOCKi_41_Q_reg_15_inst : DFF_X1 port map( D => n9860, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1071_port, QN => 
                           n_2495);
   DataPath_RF_BLOCKi_41_Q_reg_16_inst : DFF_X1 port map( D => n9859, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1072_port, QN => 
                           n_2496);
   DataPath_RF_BLOCKi_41_Q_reg_17_inst : DFF_X1 port map( D => n9858, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1073_port, QN => 
                           n_2497);
   DataPath_RF_BLOCKi_41_Q_reg_18_inst : DFF_X1 port map( D => n9857, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1074_port, QN => 
                           n_2498);
   DataPath_RF_BLOCKi_41_Q_reg_19_inst : DFF_X1 port map( D => n9856, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1075_port, QN => 
                           n_2499);
   DataPath_RF_BLOCKi_41_Q_reg_20_inst : DFF_X1 port map( D => n9855, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1076_port, QN => 
                           n_2500);
   DataPath_RF_BLOCKi_41_Q_reg_21_inst : DFF_X1 port map( D => n9854, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1077_port, QN => 
                           n_2501);
   DataPath_RF_BLOCKi_41_Q_reg_22_inst : DFF_X1 port map( D => n9853, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1078_port, QN => 
                           n_2502);
   DataPath_RF_BLOCKi_41_Q_reg_23_inst : DFF_X1 port map( D => n9852, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1079_port, QN => 
                           n_2503);
   DataPath_RF_BLOCKi_41_Q_reg_24_inst : DFF_X1 port map( D => n9851, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1080_port, QN => 
                           n_2504);
   DataPath_RF_BLOCKi_41_Q_reg_25_inst : DFF_X1 port map( D => n9850, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1081_port, QN => 
                           n_2505);
   DataPath_RF_BLOCKi_41_Q_reg_26_inst : DFF_X1 port map( D => n9849, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1082_port, QN => 
                           n_2506);
   DataPath_RF_BLOCKi_41_Q_reg_27_inst : DFF_X1 port map( D => n9848, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1083_port, QN => 
                           n_2507);
   DataPath_RF_BLOCKi_41_Q_reg_28_inst : DFF_X1 port map( D => n9847, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1084_port, QN => 
                           n_2508);
   DataPath_RF_BLOCKi_41_Q_reg_29_inst : DFF_X1 port map( D => n9846, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1085_port, QN => 
                           n_2509);
   DataPath_RF_BLOCKi_41_Q_reg_30_inst : DFF_X1 port map( D => n9845, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1086_port, QN => 
                           n_2510);
   DataPath_RF_BLOCKi_41_Q_reg_31_inst : DFF_X1 port map( D => n9844, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1087_port, QN => 
                           n_2511);
   DataPath_RF_BLOCKi_40_Q_reg_0_inst : DFF_X1 port map( D => n9843, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1024_port, QN => 
                           n_2512);
   DataPath_RF_BLOCKi_40_Q_reg_1_inst : DFF_X1 port map( D => n9842, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1025_port, QN => 
                           n_2513);
   DataPath_RF_BLOCKi_40_Q_reg_2_inst : DFF_X1 port map( D => n9841, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1026_port, QN => 
                           n_2514);
   DataPath_RF_BLOCKi_40_Q_reg_3_inst : DFF_X1 port map( D => n9840, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1027_port, QN => 
                           n_2515);
   DataPath_RF_BLOCKi_40_Q_reg_4_inst : DFF_X1 port map( D => n9839, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1028_port, QN => 
                           n_2516);
   DataPath_RF_BLOCKi_40_Q_reg_5_inst : DFF_X1 port map( D => n9838, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1029_port, QN => 
                           n_2517);
   DataPath_RF_BLOCKi_40_Q_reg_6_inst : DFF_X1 port map( D => n9837, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1030_port, QN => 
                           n_2518);
   DataPath_RF_BLOCKi_40_Q_reg_7_inst : DFF_X1 port map( D => n9836, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1031_port, QN => 
                           n_2519);
   DataPath_RF_BLOCKi_40_Q_reg_8_inst : DFF_X1 port map( D => n9835, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1032_port, QN => 
                           n_2520);
   DataPath_RF_BLOCKi_40_Q_reg_9_inst : DFF_X1 port map( D => n9834, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1033_port, QN => 
                           n_2521);
   DataPath_RF_BLOCKi_40_Q_reg_10_inst : DFF_X1 port map( D => n9833, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1034_port, QN => 
                           n_2522);
   DataPath_RF_BLOCKi_40_Q_reg_11_inst : DFF_X1 port map( D => n9832, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1035_port, QN => 
                           n_2523);
   DataPath_RF_BLOCKi_40_Q_reg_12_inst : DFF_X1 port map( D => n9831, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1036_port, QN => 
                           n_2524);
   DataPath_RF_BLOCKi_40_Q_reg_13_inst : DFF_X1 port map( D => n9830, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1037_port, QN => 
                           n_2525);
   DataPath_RF_BLOCKi_40_Q_reg_14_inst : DFF_X1 port map( D => n9829, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1038_port, QN => 
                           n_2526);
   DataPath_RF_BLOCKi_40_Q_reg_15_inst : DFF_X1 port map( D => n9828, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1039_port, QN => 
                           n_2527);
   DataPath_RF_BLOCKi_40_Q_reg_16_inst : DFF_X1 port map( D => n9827, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1040_port, QN => 
                           n_2528);
   DataPath_RF_BLOCKi_40_Q_reg_17_inst : DFF_X1 port map( D => n9826, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1041_port, QN => 
                           n_2529);
   DataPath_RF_BLOCKi_40_Q_reg_18_inst : DFF_X1 port map( D => n9825, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1042_port, QN => 
                           n_2530);
   DataPath_RF_BLOCKi_40_Q_reg_19_inst : DFF_X1 port map( D => n9824, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1043_port, QN => 
                           n_2531);
   DataPath_RF_BLOCKi_40_Q_reg_20_inst : DFF_X1 port map( D => n9823, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1044_port, QN => 
                           n_2532);
   DataPath_RF_BLOCKi_40_Q_reg_21_inst : DFF_X1 port map( D => n9822, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1045_port, QN => 
                           n_2533);
   DataPath_RF_BLOCKi_40_Q_reg_22_inst : DFF_X1 port map( D => n9821, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1046_port, QN => 
                           n_2534);
   DataPath_RF_BLOCKi_40_Q_reg_23_inst : DFF_X1 port map( D => n9820, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1047_port, QN => 
                           n_2535);
   DataPath_RF_BLOCKi_40_Q_reg_24_inst : DFF_X1 port map( D => n9819, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1048_port, QN => 
                           n_2536);
   DataPath_RF_BLOCKi_40_Q_reg_25_inst : DFF_X1 port map( D => n9818, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1049_port, QN => 
                           n_2537);
   DataPath_RF_BLOCKi_40_Q_reg_26_inst : DFF_X1 port map( D => n9817, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1050_port, QN => 
                           n_2538);
   DataPath_RF_BLOCKi_40_Q_reg_27_inst : DFF_X1 port map( D => n9816, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1051_port, QN => 
                           n_2539);
   DataPath_RF_BLOCKi_40_Q_reg_28_inst : DFF_X1 port map( D => n9815, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1052_port, QN => 
                           n_2540);
   DataPath_RF_BLOCKi_40_Q_reg_29_inst : DFF_X1 port map( D => n9814, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1053_port, QN => 
                           n_2541);
   DataPath_RF_BLOCKi_40_Q_reg_30_inst : DFF_X1 port map( D => n9813, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1054_port, QN => 
                           n_2542);
   DataPath_RF_BLOCKi_40_Q_reg_31_inst : DFF_X1 port map( D => n9812, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1055_port, QN => 
                           n_2543);
   DataPath_RF_BLOCKi_39_Q_reg_0_inst : DFF_X1 port map( D => n9811, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_992_port, QN => 
                           n_2544);
   DataPath_RF_BLOCKi_39_Q_reg_1_inst : DFF_X1 port map( D => n9810, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_993_port, QN => 
                           n_2545);
   DataPath_RF_BLOCKi_39_Q_reg_2_inst : DFF_X1 port map( D => n9809, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_994_port, QN => 
                           n_2546);
   DataPath_RF_BLOCKi_39_Q_reg_3_inst : DFF_X1 port map( D => n9808, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_995_port, QN => 
                           n_2547);
   DataPath_RF_BLOCKi_39_Q_reg_4_inst : DFF_X1 port map( D => n9807, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_996_port, QN => 
                           n_2548);
   DataPath_RF_BLOCKi_39_Q_reg_5_inst : DFF_X1 port map( D => n9806, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_997_port, QN => 
                           n_2549);
   DataPath_RF_BLOCKi_39_Q_reg_6_inst : DFF_X1 port map( D => n9805, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_998_port, QN => 
                           n_2550);
   DataPath_RF_BLOCKi_39_Q_reg_7_inst : DFF_X1 port map( D => n9804, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_999_port, QN => 
                           n_2551);
   DataPath_RF_BLOCKi_39_Q_reg_8_inst : DFF_X1 port map( D => n9803, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1000_port, QN => 
                           n_2552);
   DataPath_RF_BLOCKi_39_Q_reg_9_inst : DFF_X1 port map( D => n9802, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_1001_port, QN => 
                           n_2553);
   DataPath_RF_BLOCKi_39_Q_reg_10_inst : DFF_X1 port map( D => n9801, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1002_port, QN => 
                           n_2554);
   DataPath_RF_BLOCKi_39_Q_reg_11_inst : DFF_X1 port map( D => n9800, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1003_port, QN => 
                           n_2555);
   DataPath_RF_BLOCKi_39_Q_reg_12_inst : DFF_X1 port map( D => n9799, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1004_port, QN => 
                           n_2556);
   DataPath_RF_BLOCKi_39_Q_reg_13_inst : DFF_X1 port map( D => n9798, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1005_port, QN => 
                           n_2557);
   DataPath_RF_BLOCKi_39_Q_reg_14_inst : DFF_X1 port map( D => n9797, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1006_port, QN => 
                           n_2558);
   DataPath_RF_BLOCKi_39_Q_reg_15_inst : DFF_X1 port map( D => n9796, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1007_port, QN => 
                           n_2559);
   DataPath_RF_BLOCKi_39_Q_reg_16_inst : DFF_X1 port map( D => n9795, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1008_port, QN => 
                           n_2560);
   DataPath_RF_BLOCKi_39_Q_reg_17_inst : DFF_X1 port map( D => n9794, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1009_port, QN => 
                           n_2561);
   DataPath_RF_BLOCKi_39_Q_reg_18_inst : DFF_X1 port map( D => n9793, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1010_port, QN => 
                           n_2562);
   DataPath_RF_BLOCKi_39_Q_reg_19_inst : DFF_X1 port map( D => n9792, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1011_port, QN => 
                           n_2563);
   DataPath_RF_BLOCKi_39_Q_reg_20_inst : DFF_X1 port map( D => n9791, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1012_port, QN => 
                           n_2564);
   DataPath_RF_BLOCKi_39_Q_reg_21_inst : DFF_X1 port map( D => n9790, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1013_port, QN => 
                           n_2565);
   DataPath_RF_BLOCKi_39_Q_reg_22_inst : DFF_X1 port map( D => n9789, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1014_port, QN => 
                           n_2566);
   DataPath_RF_BLOCKi_39_Q_reg_23_inst : DFF_X1 port map( D => n9788, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1015_port, QN => 
                           n_2567);
   DataPath_RF_BLOCKi_39_Q_reg_24_inst : DFF_X1 port map( D => n9787, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1016_port, QN => 
                           n_2568);
   DataPath_RF_BLOCKi_39_Q_reg_25_inst : DFF_X1 port map( D => n9786, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1017_port, QN => 
                           n_2569);
   DataPath_RF_BLOCKi_39_Q_reg_26_inst : DFF_X1 port map( D => n9785, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1018_port, QN => 
                           n_2570);
   DataPath_RF_BLOCKi_39_Q_reg_27_inst : DFF_X1 port map( D => n9784, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1019_port, QN => 
                           n_2571);
   DataPath_RF_BLOCKi_39_Q_reg_28_inst : DFF_X1 port map( D => n9783, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1020_port, QN => 
                           n_2572);
   DataPath_RF_BLOCKi_39_Q_reg_29_inst : DFF_X1 port map( D => n9782, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1021_port, QN => 
                           n_2573);
   DataPath_RF_BLOCKi_39_Q_reg_30_inst : DFF_X1 port map( D => n9781, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1022_port, QN => 
                           n_2574);
   DataPath_RF_BLOCKi_39_Q_reg_31_inst : DFF_X1 port map( D => n9780, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_1023_port, QN => 
                           n_2575);
   DataPath_RF_BLOCKi_38_Q_reg_0_inst : DFF_X1 port map( D => n9779, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_960_port, QN => 
                           n_2576);
   DataPath_RF_BLOCKi_38_Q_reg_1_inst : DFF_X1 port map( D => n9778, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_961_port, QN => 
                           n_2577);
   DataPath_RF_BLOCKi_38_Q_reg_2_inst : DFF_X1 port map( D => n9777, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_962_port, QN => 
                           n_2578);
   DataPath_RF_BLOCKi_38_Q_reg_3_inst : DFF_X1 port map( D => n9776, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_963_port, QN => 
                           n_2579);
   DataPath_RF_BLOCKi_38_Q_reg_4_inst : DFF_X1 port map( D => n9775, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_964_port, QN => 
                           n_2580);
   DataPath_RF_BLOCKi_38_Q_reg_5_inst : DFF_X1 port map( D => n9774, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_965_port, QN => 
                           n_2581);
   DataPath_RF_BLOCKi_38_Q_reg_6_inst : DFF_X1 port map( D => n9773, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_966_port, QN => 
                           n_2582);
   DataPath_RF_BLOCKi_38_Q_reg_7_inst : DFF_X1 port map( D => n9772, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_967_port, QN => 
                           n_2583);
   DataPath_RF_BLOCKi_38_Q_reg_8_inst : DFF_X1 port map( D => n9771, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_968_port, QN => 
                           n_2584);
   DataPath_RF_BLOCKi_38_Q_reg_9_inst : DFF_X1 port map( D => n9770, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_969_port, QN => 
                           n_2585);
   DataPath_RF_BLOCKi_38_Q_reg_10_inst : DFF_X1 port map( D => n9769, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_970_port, QN => 
                           n_2586);
   DataPath_RF_BLOCKi_38_Q_reg_11_inst : DFF_X1 port map( D => n9768, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_971_port, QN => 
                           n_2587);
   DataPath_RF_BLOCKi_38_Q_reg_12_inst : DFF_X1 port map( D => n9767, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_972_port, QN => 
                           n_2588);
   DataPath_RF_BLOCKi_38_Q_reg_13_inst : DFF_X1 port map( D => n9766, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_973_port, QN => 
                           n_2589);
   DataPath_RF_BLOCKi_38_Q_reg_14_inst : DFF_X1 port map( D => n9765, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_974_port, QN => 
                           n_2590);
   DataPath_RF_BLOCKi_38_Q_reg_15_inst : DFF_X1 port map( D => n9764, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_975_port, QN => 
                           n_2591);
   DataPath_RF_BLOCKi_38_Q_reg_16_inst : DFF_X1 port map( D => n9763, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_976_port, QN => 
                           n_2592);
   DataPath_RF_BLOCKi_38_Q_reg_17_inst : DFF_X1 port map( D => n9762, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_977_port, QN => 
                           n_2593);
   DataPath_RF_BLOCKi_38_Q_reg_18_inst : DFF_X1 port map( D => n9761, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_978_port, QN => 
                           n_2594);
   DataPath_RF_BLOCKi_38_Q_reg_19_inst : DFF_X1 port map( D => n9760, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_979_port, QN => 
                           n_2595);
   DataPath_RF_BLOCKi_38_Q_reg_20_inst : DFF_X1 port map( D => n9759, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_980_port, QN => 
                           n_2596);
   DataPath_RF_BLOCKi_38_Q_reg_21_inst : DFF_X1 port map( D => n9758, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_981_port, QN => 
                           n_2597);
   DataPath_RF_BLOCKi_38_Q_reg_22_inst : DFF_X1 port map( D => n9757, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_982_port, QN => 
                           n_2598);
   DataPath_RF_BLOCKi_38_Q_reg_23_inst : DFF_X1 port map( D => n9756, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_983_port, QN => 
                           n_2599);
   DataPath_RF_BLOCKi_38_Q_reg_24_inst : DFF_X1 port map( D => n9755, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_984_port, QN => 
                           n_2600);
   DataPath_RF_BLOCKi_38_Q_reg_25_inst : DFF_X1 port map( D => n9754, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_985_port, QN => 
                           n_2601);
   DataPath_RF_BLOCKi_38_Q_reg_26_inst : DFF_X1 port map( D => n9753, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_986_port, QN => 
                           n_2602);
   DataPath_RF_BLOCKi_38_Q_reg_27_inst : DFF_X1 port map( D => n9752, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_987_port, QN => 
                           n_2603);
   DataPath_RF_BLOCKi_38_Q_reg_28_inst : DFF_X1 port map( D => n9751, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_988_port, QN => 
                           n_2604);
   DataPath_RF_BLOCKi_38_Q_reg_29_inst : DFF_X1 port map( D => n9750, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_989_port, QN => 
                           n_2605);
   DataPath_RF_BLOCKi_38_Q_reg_30_inst : DFF_X1 port map( D => n9749, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_990_port, QN => 
                           n_2606);
   DataPath_RF_BLOCKi_38_Q_reg_31_inst : DFF_X1 port map( D => n9748, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_991_port, QN => 
                           n_2607);
   DataPath_RF_BLOCKi_37_Q_reg_0_inst : DFF_X1 port map( D => n9747, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_928_port, QN => 
                           n_2608);
   DataPath_RF_BLOCKi_37_Q_reg_1_inst : DFF_X1 port map( D => n9746, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_929_port, QN => 
                           n_2609);
   DataPath_RF_BLOCKi_37_Q_reg_2_inst : DFF_X1 port map( D => n9745, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_930_port, QN => 
                           n_2610);
   DataPath_RF_BLOCKi_37_Q_reg_3_inst : DFF_X1 port map( D => n9744, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_931_port, QN => 
                           n_2611);
   DataPath_RF_BLOCKi_37_Q_reg_4_inst : DFF_X1 port map( D => n9743, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_932_port, QN => 
                           n_2612);
   DataPath_RF_BLOCKi_37_Q_reg_5_inst : DFF_X1 port map( D => n9742, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_933_port, QN => 
                           n_2613);
   DataPath_RF_BLOCKi_37_Q_reg_6_inst : DFF_X1 port map( D => n9741, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_934_port, QN => 
                           n_2614);
   DataPath_RF_BLOCKi_37_Q_reg_7_inst : DFF_X1 port map( D => n9740, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_935_port, QN => 
                           n_2615);
   DataPath_RF_BLOCKi_37_Q_reg_8_inst : DFF_X1 port map( D => n9739, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_936_port, QN => 
                           n_2616);
   DataPath_RF_BLOCKi_37_Q_reg_9_inst : DFF_X1 port map( D => n9738, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_937_port, QN => 
                           n_2617);
   DataPath_RF_BLOCKi_37_Q_reg_10_inst : DFF_X1 port map( D => n9737, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_938_port, QN => 
                           n_2618);
   DataPath_RF_BLOCKi_37_Q_reg_11_inst : DFF_X1 port map( D => n9736, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_939_port, QN => 
                           n_2619);
   DataPath_RF_BLOCKi_37_Q_reg_12_inst : DFF_X1 port map( D => n9735, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_940_port, QN => 
                           n_2620);
   DataPath_RF_BLOCKi_37_Q_reg_13_inst : DFF_X1 port map( D => n9734, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_941_port, QN => 
                           n_2621);
   DataPath_RF_BLOCKi_37_Q_reg_14_inst : DFF_X1 port map( D => n9733, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_942_port, QN => 
                           n_2622);
   DataPath_RF_BLOCKi_37_Q_reg_15_inst : DFF_X1 port map( D => n9732, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_943_port, QN => 
                           n_2623);
   DataPath_RF_BLOCKi_37_Q_reg_16_inst : DFF_X1 port map( D => n9731, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_944_port, QN => 
                           n_2624);
   DataPath_RF_BLOCKi_37_Q_reg_17_inst : DFF_X1 port map( D => n9730, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_945_port, QN => 
                           n_2625);
   DataPath_RF_BLOCKi_37_Q_reg_18_inst : DFF_X1 port map( D => n9729, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_946_port, QN => 
                           n_2626);
   DataPath_RF_BLOCKi_37_Q_reg_19_inst : DFF_X1 port map( D => n9728, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_947_port, QN => 
                           n_2627);
   DataPath_RF_BLOCKi_37_Q_reg_20_inst : DFF_X1 port map( D => n9727, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_948_port, QN => 
                           n_2628);
   DataPath_RF_BLOCKi_37_Q_reg_21_inst : DFF_X1 port map( D => n9726, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_949_port, QN => 
                           n_2629);
   DataPath_RF_BLOCKi_37_Q_reg_22_inst : DFF_X1 port map( D => n9725, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_950_port, QN => 
                           n_2630);
   DataPath_RF_BLOCKi_37_Q_reg_23_inst : DFF_X1 port map( D => n9724, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_951_port, QN => 
                           n_2631);
   DataPath_RF_BLOCKi_37_Q_reg_24_inst : DFF_X1 port map( D => n9723, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_952_port, QN => 
                           n_2632);
   DataPath_RF_BLOCKi_37_Q_reg_25_inst : DFF_X1 port map( D => n9722, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_953_port, QN => 
                           n_2633);
   DataPath_RF_BLOCKi_37_Q_reg_26_inst : DFF_X1 port map( D => n9721, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_954_port, QN => 
                           n_2634);
   DataPath_RF_BLOCKi_37_Q_reg_27_inst : DFF_X1 port map( D => n9720, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_955_port, QN => 
                           n_2635);
   DataPath_RF_BLOCKi_37_Q_reg_28_inst : DFF_X1 port map( D => n9719, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_956_port, QN => 
                           n_2636);
   DataPath_RF_BLOCKi_37_Q_reg_29_inst : DFF_X1 port map( D => n9718, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_957_port, QN => 
                           n_2637);
   DataPath_RF_BLOCKi_37_Q_reg_30_inst : DFF_X1 port map( D => n9717, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_958_port, QN => 
                           n_2638);
   DataPath_RF_BLOCKi_37_Q_reg_31_inst : DFF_X1 port map( D => n9716, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_959_port, QN => 
                           n_2639);
   DataPath_RF_BLOCKi_36_Q_reg_0_inst : DFF_X1 port map( D => n9715, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_896_port, QN => 
                           n_2640);
   DataPath_RF_BLOCKi_36_Q_reg_1_inst : DFF_X1 port map( D => n9714, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_897_port, QN => 
                           n_2641);
   DataPath_RF_BLOCKi_36_Q_reg_2_inst : DFF_X1 port map( D => n9713, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_898_port, QN => 
                           n_2642);
   DataPath_RF_BLOCKi_36_Q_reg_3_inst : DFF_X1 port map( D => n9712, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_899_port, QN => 
                           n_2643);
   DataPath_RF_BLOCKi_36_Q_reg_4_inst : DFF_X1 port map( D => n9711, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_900_port, QN => 
                           n_2644);
   DataPath_RF_BLOCKi_36_Q_reg_5_inst : DFF_X1 port map( D => n9710, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_901_port, QN => 
                           n_2645);
   DataPath_RF_BLOCKi_36_Q_reg_6_inst : DFF_X1 port map( D => n9709, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_902_port, QN => 
                           n_2646);
   DataPath_RF_BLOCKi_36_Q_reg_7_inst : DFF_X1 port map( D => n9708, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_903_port, QN => 
                           n_2647);
   DataPath_RF_BLOCKi_36_Q_reg_8_inst : DFF_X1 port map( D => n9707, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_904_port, QN => 
                           n_2648);
   DataPath_RF_BLOCKi_36_Q_reg_9_inst : DFF_X1 port map( D => n9706, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_905_port, QN => 
                           n_2649);
   DataPath_RF_BLOCKi_36_Q_reg_10_inst : DFF_X1 port map( D => n9705, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_906_port, QN => 
                           n_2650);
   DataPath_RF_BLOCKi_36_Q_reg_11_inst : DFF_X1 port map( D => n9704, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_907_port, QN => 
                           n_2651);
   DataPath_RF_BLOCKi_36_Q_reg_12_inst : DFF_X1 port map( D => n9703, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_908_port, QN => 
                           n_2652);
   DataPath_RF_BLOCKi_36_Q_reg_13_inst : DFF_X1 port map( D => n9702, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_909_port, QN => 
                           n_2653);
   DataPath_RF_BLOCKi_36_Q_reg_14_inst : DFF_X1 port map( D => n9701, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_910_port, QN => 
                           n_2654);
   DataPath_RF_BLOCKi_36_Q_reg_15_inst : DFF_X1 port map( D => n9700, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_911_port, QN => 
                           n_2655);
   DataPath_RF_BLOCKi_36_Q_reg_16_inst : DFF_X1 port map( D => n9699, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_912_port, QN => 
                           n_2656);
   DataPath_RF_BLOCKi_36_Q_reg_17_inst : DFF_X1 port map( D => n9698, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_913_port, QN => 
                           n_2657);
   DataPath_RF_BLOCKi_36_Q_reg_18_inst : DFF_X1 port map( D => n9697, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_914_port, QN => 
                           n_2658);
   DataPath_RF_BLOCKi_36_Q_reg_19_inst : DFF_X1 port map( D => n9696, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_915_port, QN => 
                           n_2659);
   DataPath_RF_BLOCKi_36_Q_reg_20_inst : DFF_X1 port map( D => n9695, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_916_port, QN => 
                           n_2660);
   DataPath_RF_BLOCKi_36_Q_reg_21_inst : DFF_X1 port map( D => n9694, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_917_port, QN => 
                           n_2661);
   DataPath_RF_BLOCKi_36_Q_reg_22_inst : DFF_X1 port map( D => n9693, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_918_port, QN => 
                           n_2662);
   DataPath_RF_BLOCKi_36_Q_reg_23_inst : DFF_X1 port map( D => n9692, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_919_port, QN => 
                           n_2663);
   DataPath_RF_BLOCKi_36_Q_reg_24_inst : DFF_X1 port map( D => n9691, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_920_port, QN => 
                           n_2664);
   DataPath_RF_BLOCKi_36_Q_reg_25_inst : DFF_X1 port map( D => n9690, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_921_port, QN => 
                           n_2665);
   DataPath_RF_BLOCKi_36_Q_reg_26_inst : DFF_X1 port map( D => n9689, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_922_port, QN => 
                           n_2666);
   DataPath_RF_BLOCKi_36_Q_reg_27_inst : DFF_X1 port map( D => n9688, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_923_port, QN => 
                           n_2667);
   DataPath_RF_BLOCKi_36_Q_reg_28_inst : DFF_X1 port map( D => n9687, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_924_port, QN => 
                           n_2668);
   DataPath_RF_BLOCKi_36_Q_reg_29_inst : DFF_X1 port map( D => n9686, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_925_port, QN => 
                           n_2669);
   DataPath_RF_BLOCKi_36_Q_reg_30_inst : DFF_X1 port map( D => n9685, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_926_port, QN => 
                           n_2670);
   DataPath_RF_BLOCKi_36_Q_reg_31_inst : DFF_X1 port map( D => n9684, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_927_port, QN => 
                           n_2671);
   DataPath_RF_BLOCKi_35_Q_reg_0_inst : DFF_X1 port map( D => n9683, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_864_port, QN => 
                           n_2672);
   DataPath_RF_BLOCKi_35_Q_reg_1_inst : DFF_X1 port map( D => n9682, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_865_port, QN => 
                           n_2673);
   DataPath_RF_BLOCKi_35_Q_reg_2_inst : DFF_X1 port map( D => n9681, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_866_port, QN => 
                           n_2674);
   DataPath_RF_BLOCKi_35_Q_reg_3_inst : DFF_X1 port map( D => n9680, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_867_port, QN => 
                           n_2675);
   DataPath_RF_BLOCKi_35_Q_reg_4_inst : DFF_X1 port map( D => n9679, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_868_port, QN => 
                           n_2676);
   DataPath_RF_BLOCKi_35_Q_reg_5_inst : DFF_X1 port map( D => n9678, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_869_port, QN => 
                           n_2677);
   DataPath_RF_BLOCKi_35_Q_reg_6_inst : DFF_X1 port map( D => n9677, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_870_port, QN => 
                           n_2678);
   DataPath_RF_BLOCKi_35_Q_reg_7_inst : DFF_X1 port map( D => n9676, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_871_port, QN => 
                           n_2679);
   DataPath_RF_BLOCKi_35_Q_reg_8_inst : DFF_X1 port map( D => n9675, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_872_port, QN => 
                           n_2680);
   DataPath_RF_BLOCKi_35_Q_reg_9_inst : DFF_X1 port map( D => n9674, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_873_port, QN => 
                           n_2681);
   DataPath_RF_BLOCKi_35_Q_reg_10_inst : DFF_X1 port map( D => n9673, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_874_port, QN => 
                           n_2682);
   DataPath_RF_BLOCKi_35_Q_reg_11_inst : DFF_X1 port map( D => n9672, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_875_port, QN => 
                           n_2683);
   DataPath_RF_BLOCKi_35_Q_reg_12_inst : DFF_X1 port map( D => n9671, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_876_port, QN => 
                           n_2684);
   DataPath_RF_BLOCKi_35_Q_reg_13_inst : DFF_X1 port map( D => n9670, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_877_port, QN => 
                           n_2685);
   DataPath_RF_BLOCKi_35_Q_reg_14_inst : DFF_X1 port map( D => n9669, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_878_port, QN => 
                           n_2686);
   DataPath_RF_BLOCKi_35_Q_reg_15_inst : DFF_X1 port map( D => n9668, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_879_port, QN => 
                           n_2687);
   DataPath_RF_BLOCKi_35_Q_reg_16_inst : DFF_X1 port map( D => n9667, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_880_port, QN => 
                           n_2688);
   DataPath_RF_BLOCKi_35_Q_reg_17_inst : DFF_X1 port map( D => n9666, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_881_port, QN => 
                           n_2689);
   DataPath_RF_BLOCKi_35_Q_reg_18_inst : DFF_X1 port map( D => n9665, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_882_port, QN => 
                           n_2690);
   DataPath_RF_BLOCKi_35_Q_reg_19_inst : DFF_X1 port map( D => n9664, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_883_port, QN => 
                           n_2691);
   DataPath_RF_BLOCKi_35_Q_reg_20_inst : DFF_X1 port map( D => n9663, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_884_port, QN => 
                           n_2692);
   DataPath_RF_BLOCKi_35_Q_reg_21_inst : DFF_X1 port map( D => n9662, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_885_port, QN => 
                           n_2693);
   DataPath_RF_BLOCKi_35_Q_reg_22_inst : DFF_X1 port map( D => n9661, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_886_port, QN => 
                           n_2694);
   DataPath_RF_BLOCKi_35_Q_reg_23_inst : DFF_X1 port map( D => n9660, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_887_port, QN => 
                           n_2695);
   DataPath_RF_BLOCKi_35_Q_reg_24_inst : DFF_X1 port map( D => n9659, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_888_port, QN => 
                           n_2696);
   DataPath_RF_BLOCKi_35_Q_reg_25_inst : DFF_X1 port map( D => n9658, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_889_port, QN => 
                           n_2697);
   DataPath_RF_BLOCKi_35_Q_reg_26_inst : DFF_X1 port map( D => n9657, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_890_port, QN => 
                           n_2698);
   DataPath_RF_BLOCKi_35_Q_reg_27_inst : DFF_X1 port map( D => n9656, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_891_port, QN => 
                           n_2699);
   DataPath_RF_BLOCKi_35_Q_reg_28_inst : DFF_X1 port map( D => n9655, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_892_port, QN => 
                           n_2700);
   DataPath_RF_BLOCKi_35_Q_reg_29_inst : DFF_X1 port map( D => n9654, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_893_port, QN => 
                           n_2701);
   DataPath_RF_BLOCKi_35_Q_reg_30_inst : DFF_X1 port map( D => n9653, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_894_port, QN => 
                           n_2702);
   DataPath_RF_BLOCKi_35_Q_reg_31_inst : DFF_X1 port map( D => n9652, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_895_port, QN => 
                           n_2703);
   DataPath_RF_BLOCKi_34_Q_reg_0_inst : DFF_X1 port map( D => n9651, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_832_port, QN => 
                           n_2704);
   DataPath_RF_BLOCKi_34_Q_reg_1_inst : DFF_X1 port map( D => n9650, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_833_port, QN => 
                           n_2705);
   DataPath_RF_BLOCKi_34_Q_reg_2_inst : DFF_X1 port map( D => n9649, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_834_port, QN => 
                           n_2706);
   DataPath_RF_BLOCKi_34_Q_reg_3_inst : DFF_X1 port map( D => n9648, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_835_port, QN => 
                           n_2707);
   DataPath_RF_BLOCKi_34_Q_reg_4_inst : DFF_X1 port map( D => n9647, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_836_port, QN => 
                           n_2708);
   DataPath_RF_BLOCKi_34_Q_reg_5_inst : DFF_X1 port map( D => n9646, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_837_port, QN => 
                           n_2709);
   DataPath_RF_BLOCKi_34_Q_reg_6_inst : DFF_X1 port map( D => n9645, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_838_port, QN => 
                           n_2710);
   DataPath_RF_BLOCKi_34_Q_reg_7_inst : DFF_X1 port map( D => n9644, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_839_port, QN => 
                           n_2711);
   DataPath_RF_BLOCKi_34_Q_reg_8_inst : DFF_X1 port map( D => n9643, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_840_port, QN => 
                           n_2712);
   DataPath_RF_BLOCKi_34_Q_reg_9_inst : DFF_X1 port map( D => n9642, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_841_port, QN => 
                           n_2713);
   DataPath_RF_BLOCKi_34_Q_reg_10_inst : DFF_X1 port map( D => n9641, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_842_port, QN => 
                           n_2714);
   DataPath_RF_BLOCKi_34_Q_reg_11_inst : DFF_X1 port map( D => n9640, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_843_port, QN => 
                           n_2715);
   DataPath_RF_BLOCKi_34_Q_reg_12_inst : DFF_X1 port map( D => n9639, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_844_port, QN => 
                           n_2716);
   DataPath_RF_BLOCKi_34_Q_reg_13_inst : DFF_X1 port map( D => n9638, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_845_port, QN => 
                           n_2717);
   DataPath_RF_BLOCKi_34_Q_reg_14_inst : DFF_X1 port map( D => n9637, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_846_port, QN => 
                           n_2718);
   DataPath_RF_BLOCKi_34_Q_reg_15_inst : DFF_X1 port map( D => n9636, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_847_port, QN => 
                           n_2719);
   DataPath_RF_BLOCKi_34_Q_reg_16_inst : DFF_X1 port map( D => n9635, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_848_port, QN => 
                           n_2720);
   DataPath_RF_BLOCKi_34_Q_reg_17_inst : DFF_X1 port map( D => n9634, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_849_port, QN => 
                           n_2721);
   DataPath_RF_BLOCKi_34_Q_reg_18_inst : DFF_X1 port map( D => n9633, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_850_port, QN => 
                           n_2722);
   DataPath_RF_BLOCKi_34_Q_reg_19_inst : DFF_X1 port map( D => n9632, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_851_port, QN => 
                           n_2723);
   DataPath_RF_BLOCKi_34_Q_reg_20_inst : DFF_X1 port map( D => n9631, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_852_port, QN => 
                           n_2724);
   DataPath_RF_BLOCKi_34_Q_reg_21_inst : DFF_X1 port map( D => n9630, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_853_port, QN => 
                           n_2725);
   DataPath_RF_BLOCKi_34_Q_reg_22_inst : DFF_X1 port map( D => n9629, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_854_port, QN => 
                           n_2726);
   DataPath_RF_BLOCKi_34_Q_reg_23_inst : DFF_X1 port map( D => n9628, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_855_port, QN => 
                           n_2727);
   DataPath_RF_BLOCKi_34_Q_reg_24_inst : DFF_X1 port map( D => n9627, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_856_port, QN => 
                           n_2728);
   DataPath_RF_BLOCKi_34_Q_reg_25_inst : DFF_X1 port map( D => n9626, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_857_port, QN => 
                           n_2729);
   DataPath_RF_BLOCKi_34_Q_reg_26_inst : DFF_X1 port map( D => n9625, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_858_port, QN => 
                           n_2730);
   DataPath_RF_BLOCKi_34_Q_reg_27_inst : DFF_X1 port map( D => n9624, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_859_port, QN => 
                           n_2731);
   DataPath_RF_BLOCKi_34_Q_reg_28_inst : DFF_X1 port map( D => n9623, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_860_port, QN => 
                           n_2732);
   DataPath_RF_BLOCKi_34_Q_reg_29_inst : DFF_X1 port map( D => n9622, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_861_port, QN => 
                           n_2733);
   DataPath_RF_BLOCKi_34_Q_reg_30_inst : DFF_X1 port map( D => n9621, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_862_port, QN => 
                           n_2734);
   DataPath_RF_BLOCKi_34_Q_reg_31_inst : DFF_X1 port map( D => n9620, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_863_port, QN => 
                           n_2735);
   DataPath_RF_BLOCKi_33_Q_reg_0_inst : DFF_X1 port map( D => n9619, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_800_port, QN => 
                           n_2736);
   DataPath_RF_BLOCKi_33_Q_reg_1_inst : DFF_X1 port map( D => n9618, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_801_port, QN => 
                           n_2737);
   DataPath_RF_BLOCKi_33_Q_reg_2_inst : DFF_X1 port map( D => n9617, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_802_port, QN => 
                           n_2738);
   DataPath_RF_BLOCKi_33_Q_reg_3_inst : DFF_X1 port map( D => n9616, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_803_port, QN => 
                           n_2739);
   DataPath_RF_BLOCKi_33_Q_reg_4_inst : DFF_X1 port map( D => n9615, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_804_port, QN => 
                           n_2740);
   DataPath_RF_BLOCKi_33_Q_reg_5_inst : DFF_X1 port map( D => n9614, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_805_port, QN => 
                           n_2741);
   DataPath_RF_BLOCKi_33_Q_reg_6_inst : DFF_X1 port map( D => n9613, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_806_port, QN => 
                           n_2742);
   DataPath_RF_BLOCKi_33_Q_reg_7_inst : DFF_X1 port map( D => n9612, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_807_port, QN => 
                           n_2743);
   DataPath_RF_BLOCKi_33_Q_reg_8_inst : DFF_X1 port map( D => n9611, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_808_port, QN => 
                           n_2744);
   DataPath_RF_BLOCKi_33_Q_reg_9_inst : DFF_X1 port map( D => n9610, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_809_port, QN => 
                           n_2745);
   DataPath_RF_BLOCKi_33_Q_reg_10_inst : DFF_X1 port map( D => n9609, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_810_port, QN => 
                           n_2746);
   DataPath_RF_BLOCKi_33_Q_reg_11_inst : DFF_X1 port map( D => n9608, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_811_port, QN => 
                           n_2747);
   DataPath_RF_BLOCKi_33_Q_reg_12_inst : DFF_X1 port map( D => n9607, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_812_port, QN => 
                           n_2748);
   DataPath_RF_BLOCKi_33_Q_reg_13_inst : DFF_X1 port map( D => n9606, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_813_port, QN => 
                           n_2749);
   DataPath_RF_BLOCKi_33_Q_reg_14_inst : DFF_X1 port map( D => n9605, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_814_port, QN => 
                           n_2750);
   DataPath_RF_BLOCKi_33_Q_reg_15_inst : DFF_X1 port map( D => n9604, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_815_port, QN => 
                           n_2751);
   DataPath_RF_BLOCKi_33_Q_reg_16_inst : DFF_X1 port map( D => n9603, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_816_port, QN => 
                           n_2752);
   DataPath_RF_BLOCKi_33_Q_reg_17_inst : DFF_X1 port map( D => n9602, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_817_port, QN => 
                           n_2753);
   DataPath_RF_BLOCKi_33_Q_reg_18_inst : DFF_X1 port map( D => n9601, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_818_port, QN => 
                           n_2754);
   DataPath_RF_BLOCKi_33_Q_reg_19_inst : DFF_X1 port map( D => n9600, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_819_port, QN => 
                           n_2755);
   DataPath_RF_BLOCKi_33_Q_reg_20_inst : DFF_X1 port map( D => n9599, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_820_port, QN => 
                           n_2756);
   DataPath_RF_BLOCKi_33_Q_reg_21_inst : DFF_X1 port map( D => n9598, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_821_port, QN => 
                           n_2757);
   DataPath_RF_BLOCKi_33_Q_reg_22_inst : DFF_X1 port map( D => n9597, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_822_port, QN => 
                           n_2758);
   DataPath_RF_BLOCKi_33_Q_reg_23_inst : DFF_X1 port map( D => n9596, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_823_port, QN => 
                           n_2759);
   DataPath_RF_BLOCKi_33_Q_reg_24_inst : DFF_X1 port map( D => n9595, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_824_port, QN => 
                           n_2760);
   DataPath_RF_BLOCKi_33_Q_reg_25_inst : DFF_X1 port map( D => n9594, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_825_port, QN => 
                           n_2761);
   DataPath_RF_BLOCKi_33_Q_reg_26_inst : DFF_X1 port map( D => n9593, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_826_port, QN => 
                           n_2762);
   DataPath_RF_BLOCKi_33_Q_reg_27_inst : DFF_X1 port map( D => n9592, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_827_port, QN => 
                           n_2763);
   DataPath_RF_BLOCKi_33_Q_reg_28_inst : DFF_X1 port map( D => n9591, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_828_port, QN => 
                           n_2764);
   DataPath_RF_BLOCKi_33_Q_reg_29_inst : DFF_X1 port map( D => n9590, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_829_port, QN => 
                           n_2765);
   DataPath_RF_BLOCKi_33_Q_reg_30_inst : DFF_X1 port map( D => n9589, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_830_port, QN => 
                           n_2766);
   DataPath_RF_BLOCKi_33_Q_reg_31_inst : DFF_X1 port map( D => n9588, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_831_port, QN => 
                           n_2767);
   DataPath_RF_BLOCKi_32_Q_reg_0_inst : DFF_X1 port map( D => n9587, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_768_port, QN => 
                           n_2768);
   DataPath_RF_BLOCKi_32_Q_reg_1_inst : DFF_X1 port map( D => n9586, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_769_port, QN => 
                           n_2769);
   DataPath_RF_BLOCKi_32_Q_reg_2_inst : DFF_X1 port map( D => n9585, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_770_port, QN => 
                           n_2770);
   DataPath_RF_BLOCKi_32_Q_reg_3_inst : DFF_X1 port map( D => n9584, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_771_port, QN => 
                           n_2771);
   DataPath_RF_BLOCKi_32_Q_reg_4_inst : DFF_X1 port map( D => n9583, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_772_port, QN => 
                           n_2772);
   DataPath_RF_BLOCKi_32_Q_reg_5_inst : DFF_X1 port map( D => n9582, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_773_port, QN => 
                           n_2773);
   DataPath_RF_BLOCKi_32_Q_reg_6_inst : DFF_X1 port map( D => n9581, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_774_port, QN => 
                           n_2774);
   DataPath_RF_BLOCKi_32_Q_reg_7_inst : DFF_X1 port map( D => n9580, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_775_port, QN => 
                           n_2775);
   DataPath_RF_BLOCKi_32_Q_reg_8_inst : DFF_X1 port map( D => n9579, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_776_port, QN => 
                           n_2776);
   DataPath_RF_BLOCKi_32_Q_reg_9_inst : DFF_X1 port map( D => n9578, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_777_port, QN => 
                           n_2777);
   DataPath_RF_BLOCKi_32_Q_reg_10_inst : DFF_X1 port map( D => n9577, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_778_port, QN => 
                           n_2778);
   DataPath_RF_BLOCKi_32_Q_reg_11_inst : DFF_X1 port map( D => n9576, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_779_port, QN => 
                           n_2779);
   DataPath_RF_BLOCKi_32_Q_reg_12_inst : DFF_X1 port map( D => n9575, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_780_port, QN => 
                           n_2780);
   DataPath_RF_BLOCKi_32_Q_reg_13_inst : DFF_X1 port map( D => n9574, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_781_port, QN => 
                           n_2781);
   DataPath_RF_BLOCKi_32_Q_reg_14_inst : DFF_X1 port map( D => n9573, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_782_port, QN => 
                           n_2782);
   DataPath_RF_BLOCKi_32_Q_reg_15_inst : DFF_X1 port map( D => n9572, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_783_port, QN => 
                           n_2783);
   DataPath_RF_BLOCKi_32_Q_reg_16_inst : DFF_X1 port map( D => n9571, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_784_port, QN => 
                           n_2784);
   DataPath_RF_BLOCKi_32_Q_reg_17_inst : DFF_X1 port map( D => n9570, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_785_port, QN => 
                           n_2785);
   DataPath_RF_BLOCKi_32_Q_reg_18_inst : DFF_X1 port map( D => n9569, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_786_port, QN => 
                           n_2786);
   DataPath_RF_BLOCKi_32_Q_reg_19_inst : DFF_X1 port map( D => n9568, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_787_port, QN => 
                           n_2787);
   DataPath_RF_BLOCKi_32_Q_reg_20_inst : DFF_X1 port map( D => n9567, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_788_port, QN => 
                           n_2788);
   DataPath_RF_BLOCKi_32_Q_reg_21_inst : DFF_X1 port map( D => n9566, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_789_port, QN => 
                           n_2789);
   DataPath_RF_BLOCKi_32_Q_reg_22_inst : DFF_X1 port map( D => n9565, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_790_port, QN => 
                           n_2790);
   DataPath_RF_BLOCKi_32_Q_reg_23_inst : DFF_X1 port map( D => n9564, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_791_port, QN => 
                           n_2791);
   DataPath_RF_BLOCKi_32_Q_reg_24_inst : DFF_X1 port map( D => n9563, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_792_port, QN => 
                           n_2792);
   DataPath_RF_BLOCKi_32_Q_reg_25_inst : DFF_X1 port map( D => n9562, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_793_port, QN => 
                           n_2793);
   DataPath_RF_BLOCKi_32_Q_reg_26_inst : DFF_X1 port map( D => n9561, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_794_port, QN => 
                           n_2794);
   DataPath_RF_BLOCKi_32_Q_reg_27_inst : DFF_X1 port map( D => n9560, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_795_port, QN => 
                           n_2795);
   DataPath_RF_BLOCKi_32_Q_reg_28_inst : DFF_X1 port map( D => n9559, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_796_port, QN => 
                           n_2796);
   DataPath_RF_BLOCKi_32_Q_reg_29_inst : DFF_X1 port map( D => n9558, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_797_port, QN => 
                           n_2797);
   DataPath_RF_BLOCKi_32_Q_reg_30_inst : DFF_X1 port map( D => n9557, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_798_port, QN => 
                           n_2798);
   DataPath_RF_BLOCKi_32_Q_reg_31_inst : DFF_X1 port map( D => n9556, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_799_port, QN => 
                           n_2799);
   DataPath_RF_BLOCKi_31_Q_reg_0_inst : DFF_X1 port map( D => n9555, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_736_port, QN => 
                           n_2800);
   DataPath_RF_BLOCKi_31_Q_reg_1_inst : DFF_X1 port map( D => n9554, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_737_port, QN => 
                           n_2801);
   DataPath_RF_BLOCKi_31_Q_reg_2_inst : DFF_X1 port map( D => n9553, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_738_port, QN => 
                           n_2802);
   DataPath_RF_BLOCKi_31_Q_reg_3_inst : DFF_X1 port map( D => n9552, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_739_port, QN => 
                           n_2803);
   DataPath_RF_BLOCKi_31_Q_reg_4_inst : DFF_X1 port map( D => n9551, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_740_port, QN => 
                           n_2804);
   DataPath_RF_BLOCKi_31_Q_reg_5_inst : DFF_X1 port map( D => n9550, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_741_port, QN => 
                           n_2805);
   DataPath_RF_BLOCKi_31_Q_reg_6_inst : DFF_X1 port map( D => n9549, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_742_port, QN => 
                           n_2806);
   DataPath_RF_BLOCKi_31_Q_reg_7_inst : DFF_X1 port map( D => n9548, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_743_port, QN => 
                           n_2807);
   DataPath_RF_BLOCKi_31_Q_reg_8_inst : DFF_X1 port map( D => n9547, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_744_port, QN => 
                           n_2808);
   DataPath_RF_BLOCKi_31_Q_reg_9_inst : DFF_X1 port map( D => n9546, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_745_port, QN => 
                           n_2809);
   DataPath_RF_BLOCKi_31_Q_reg_10_inst : DFF_X1 port map( D => n9545, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_746_port, QN => 
                           n_2810);
   DataPath_RF_BLOCKi_31_Q_reg_11_inst : DFF_X1 port map( D => n9544, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_747_port, QN => 
                           n_2811);
   DataPath_RF_BLOCKi_31_Q_reg_12_inst : DFF_X1 port map( D => n9543, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_748_port, QN => 
                           n_2812);
   DataPath_RF_BLOCKi_31_Q_reg_13_inst : DFF_X1 port map( D => n9542, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_749_port, QN => 
                           n_2813);
   DataPath_RF_BLOCKi_31_Q_reg_14_inst : DFF_X1 port map( D => n9541, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_750_port, QN => 
                           n_2814);
   DataPath_RF_BLOCKi_31_Q_reg_15_inst : DFF_X1 port map( D => n9540, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_751_port, QN => 
                           n_2815);
   DataPath_RF_BLOCKi_31_Q_reg_16_inst : DFF_X1 port map( D => n9539, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_752_port, QN => 
                           n_2816);
   DataPath_RF_BLOCKi_31_Q_reg_17_inst : DFF_X1 port map( D => n9538, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_753_port, QN => 
                           n_2817);
   DataPath_RF_BLOCKi_31_Q_reg_18_inst : DFF_X1 port map( D => n9537, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_754_port, QN => 
                           n_2818);
   DataPath_RF_BLOCKi_31_Q_reg_19_inst : DFF_X1 port map( D => n9536, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_755_port, QN => 
                           n_2819);
   DataPath_RF_BLOCKi_31_Q_reg_20_inst : DFF_X1 port map( D => n9535, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_756_port, QN => 
                           n_2820);
   DataPath_RF_BLOCKi_31_Q_reg_21_inst : DFF_X1 port map( D => n9534, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_757_port, QN => 
                           n_2821);
   DataPath_RF_BLOCKi_31_Q_reg_22_inst : DFF_X1 port map( D => n9533, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_758_port, QN => 
                           n_2822);
   DataPath_RF_BLOCKi_31_Q_reg_23_inst : DFF_X1 port map( D => n9532, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_759_port, QN => 
                           n_2823);
   DataPath_RF_BLOCKi_31_Q_reg_24_inst : DFF_X1 port map( D => n9531, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_760_port, QN => 
                           n_2824);
   DataPath_RF_BLOCKi_31_Q_reg_25_inst : DFF_X1 port map( D => n9530, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_761_port, QN => 
                           n_2825);
   DataPath_RF_BLOCKi_31_Q_reg_26_inst : DFF_X1 port map( D => n9529, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_762_port, QN => 
                           n_2826);
   DataPath_RF_BLOCKi_31_Q_reg_27_inst : DFF_X1 port map( D => n9528, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_763_port, QN => 
                           n_2827);
   DataPath_RF_BLOCKi_31_Q_reg_28_inst : DFF_X1 port map( D => n9527, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_764_port, QN => 
                           n_2828);
   DataPath_RF_BLOCKi_31_Q_reg_29_inst : DFF_X1 port map( D => n9526, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_765_port, QN => 
                           n_2829);
   DataPath_RF_BLOCKi_31_Q_reg_30_inst : DFF_X1 port map( D => n9525, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_766_port, QN => 
                           n_2830);
   DataPath_RF_BLOCKi_31_Q_reg_31_inst : DFF_X1 port map( D => n9524, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_767_port, QN => 
                           n_2831);
   DataPath_RF_BLOCKi_30_Q_reg_0_inst : DFF_X1 port map( D => n9523, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_704_port, QN => 
                           n_2832);
   DataPath_RF_BLOCKi_30_Q_reg_1_inst : DFF_X1 port map( D => n9522, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_705_port, QN => 
                           n_2833);
   DataPath_RF_BLOCKi_30_Q_reg_2_inst : DFF_X1 port map( D => n9521, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_706_port, QN => 
                           n_2834);
   DataPath_RF_BLOCKi_30_Q_reg_3_inst : DFF_X1 port map( D => n9520, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_707_port, QN => 
                           n_2835);
   DataPath_RF_BLOCKi_30_Q_reg_4_inst : DFF_X1 port map( D => n9519, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_708_port, QN => 
                           n_2836);
   DataPath_RF_BLOCKi_30_Q_reg_5_inst : DFF_X1 port map( D => n9518, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_709_port, QN => 
                           n_2837);
   DataPath_RF_BLOCKi_30_Q_reg_6_inst : DFF_X1 port map( D => n9517, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_710_port, QN => 
                           n_2838);
   DataPath_RF_BLOCKi_30_Q_reg_7_inst : DFF_X1 port map( D => n9516, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_711_port, QN => 
                           n_2839);
   DataPath_RF_BLOCKi_30_Q_reg_8_inst : DFF_X1 port map( D => n9515, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_712_port, QN => 
                           n_2840);
   DataPath_RF_BLOCKi_30_Q_reg_9_inst : DFF_X1 port map( D => n9514, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_713_port, QN => 
                           n_2841);
   DataPath_RF_BLOCKi_30_Q_reg_10_inst : DFF_X1 port map( D => n9513, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_714_port, QN => 
                           n_2842);
   DataPath_RF_BLOCKi_30_Q_reg_11_inst : DFF_X1 port map( D => n9512, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_715_port, QN => 
                           n_2843);
   DataPath_RF_BLOCKi_30_Q_reg_12_inst : DFF_X1 port map( D => n9511, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_716_port, QN => 
                           n_2844);
   DataPath_RF_BLOCKi_30_Q_reg_13_inst : DFF_X1 port map( D => n9510, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_717_port, QN => 
                           n_2845);
   DataPath_RF_BLOCKi_30_Q_reg_14_inst : DFF_X1 port map( D => n9509, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_718_port, QN => 
                           n_2846);
   DataPath_RF_BLOCKi_30_Q_reg_15_inst : DFF_X1 port map( D => n9508, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_719_port, QN => 
                           n_2847);
   DataPath_RF_BLOCKi_30_Q_reg_16_inst : DFF_X1 port map( D => n9507, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_720_port, QN => 
                           n_2848);
   DataPath_RF_BLOCKi_30_Q_reg_17_inst : DFF_X1 port map( D => n9506, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_721_port, QN => 
                           n_2849);
   DataPath_RF_BLOCKi_30_Q_reg_18_inst : DFF_X1 port map( D => n9505, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_722_port, QN => 
                           n_2850);
   DataPath_RF_BLOCKi_30_Q_reg_19_inst : DFF_X1 port map( D => n9504, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_723_port, QN => 
                           n_2851);
   DataPath_RF_BLOCKi_30_Q_reg_20_inst : DFF_X1 port map( D => n9503, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_724_port, QN => 
                           n_2852);
   DataPath_RF_BLOCKi_30_Q_reg_21_inst : DFF_X1 port map( D => n9502, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_725_port, QN => 
                           n_2853);
   DataPath_RF_BLOCKi_30_Q_reg_22_inst : DFF_X1 port map( D => n9501, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_726_port, QN => 
                           n_2854);
   DataPath_RF_BLOCKi_30_Q_reg_23_inst : DFF_X1 port map( D => n9500, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_727_port, QN => 
                           n_2855);
   DataPath_RF_BLOCKi_30_Q_reg_24_inst : DFF_X1 port map( D => n9499, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_728_port, QN => 
                           n_2856);
   DataPath_RF_BLOCKi_30_Q_reg_25_inst : DFF_X1 port map( D => n9498, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_729_port, QN => 
                           n_2857);
   DataPath_RF_BLOCKi_30_Q_reg_26_inst : DFF_X1 port map( D => n9497, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_730_port, QN => 
                           n_2858);
   DataPath_RF_BLOCKi_30_Q_reg_27_inst : DFF_X1 port map( D => n9496, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_731_port, QN => 
                           n_2859);
   DataPath_RF_BLOCKi_30_Q_reg_28_inst : DFF_X1 port map( D => n9495, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_732_port, QN => 
                           n_2860);
   DataPath_RF_BLOCKi_30_Q_reg_29_inst : DFF_X1 port map( D => n9494, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_733_port, QN => 
                           n_2861);
   DataPath_RF_BLOCKi_30_Q_reg_30_inst : DFF_X1 port map( D => n9493, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_734_port, QN => 
                           n_2862);
   DataPath_RF_BLOCKi_30_Q_reg_31_inst : DFF_X1 port map( D => n9492, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_735_port, QN => 
                           n_2863);
   DataPath_RF_BLOCKi_29_Q_reg_0_inst : DFF_X1 port map( D => n9491, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_672_port, QN => 
                           n_2864);
   DataPath_RF_BLOCKi_29_Q_reg_1_inst : DFF_X1 port map( D => n9490, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_673_port, QN => 
                           n_2865);
   DataPath_RF_BLOCKi_29_Q_reg_2_inst : DFF_X1 port map( D => n9489, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_674_port, QN => 
                           n_2866);
   DataPath_RF_BLOCKi_29_Q_reg_3_inst : DFF_X1 port map( D => n9488, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_675_port, QN => 
                           n_2867);
   DataPath_RF_BLOCKi_29_Q_reg_4_inst : DFF_X1 port map( D => n9487, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_676_port, QN => 
                           n_2868);
   DataPath_RF_BLOCKi_29_Q_reg_5_inst : DFF_X1 port map( D => n9486, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_677_port, QN => 
                           n_2869);
   DataPath_RF_BLOCKi_29_Q_reg_6_inst : DFF_X1 port map( D => n9485, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_678_port, QN => 
                           n_2870);
   DataPath_RF_BLOCKi_29_Q_reg_7_inst : DFF_X1 port map( D => n9484, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_679_port, QN => 
                           n_2871);
   DataPath_RF_BLOCKi_29_Q_reg_8_inst : DFF_X1 port map( D => n9483, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_680_port, QN => 
                           n_2872);
   DataPath_RF_BLOCKi_29_Q_reg_9_inst : DFF_X1 port map( D => n9482, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_681_port, QN => 
                           n_2873);
   DataPath_RF_BLOCKi_29_Q_reg_10_inst : DFF_X1 port map( D => n9481, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_682_port, QN => 
                           n_2874);
   DataPath_RF_BLOCKi_29_Q_reg_11_inst : DFF_X1 port map( D => n9480, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_683_port, QN => 
                           n_2875);
   DataPath_RF_BLOCKi_29_Q_reg_12_inst : DFF_X1 port map( D => n9479, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_684_port, QN => 
                           n_2876);
   DataPath_RF_BLOCKi_29_Q_reg_13_inst : DFF_X1 port map( D => n9478, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_685_port, QN => 
                           n_2877);
   DataPath_RF_BLOCKi_29_Q_reg_14_inst : DFF_X1 port map( D => n9477, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_686_port, QN => 
                           n_2878);
   DataPath_RF_BLOCKi_29_Q_reg_15_inst : DFF_X1 port map( D => n9476, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_687_port, QN => 
                           n_2879);
   DataPath_RF_BLOCKi_29_Q_reg_16_inst : DFF_X1 port map( D => n9475, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_688_port, QN => 
                           n_2880);
   DataPath_RF_BLOCKi_29_Q_reg_17_inst : DFF_X1 port map( D => n9474, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_689_port, QN => 
                           n_2881);
   DataPath_RF_BLOCKi_29_Q_reg_18_inst : DFF_X1 port map( D => n9473, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_690_port, QN => 
                           n_2882);
   DataPath_RF_BLOCKi_29_Q_reg_19_inst : DFF_X1 port map( D => n9472, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_691_port, QN => 
                           n_2883);
   DataPath_RF_BLOCKi_29_Q_reg_20_inst : DFF_X1 port map( D => n9471, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_692_port, QN => 
                           n_2884);
   DataPath_RF_BLOCKi_29_Q_reg_21_inst : DFF_X1 port map( D => n9470, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_693_port, QN => 
                           n_2885);
   DataPath_RF_BLOCKi_29_Q_reg_22_inst : DFF_X1 port map( D => n9469, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_694_port, QN => 
                           n_2886);
   DataPath_RF_BLOCKi_29_Q_reg_23_inst : DFF_X1 port map( D => n9468, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_695_port, QN => 
                           n_2887);
   DataPath_RF_BLOCKi_29_Q_reg_24_inst : DFF_X1 port map( D => n9467, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_696_port, QN => 
                           n_2888);
   DataPath_RF_BLOCKi_29_Q_reg_25_inst : DFF_X1 port map( D => n9466, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_697_port, QN => 
                           n_2889);
   DataPath_RF_BLOCKi_29_Q_reg_26_inst : DFF_X1 port map( D => n9465, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_698_port, QN => 
                           n_2890);
   DataPath_RF_BLOCKi_29_Q_reg_27_inst : DFF_X1 port map( D => n9464, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_699_port, QN => 
                           n_2891);
   DataPath_RF_BLOCKi_29_Q_reg_28_inst : DFF_X1 port map( D => n9463, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_700_port, QN => 
                           n_2892);
   DataPath_RF_BLOCKi_29_Q_reg_29_inst : DFF_X1 port map( D => n9462, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_701_port, QN => 
                           n_2893);
   DataPath_RF_BLOCKi_29_Q_reg_30_inst : DFF_X1 port map( D => n9461, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_702_port, QN => 
                           n_2894);
   DataPath_RF_BLOCKi_29_Q_reg_31_inst : DFF_X1 port map( D => n9460, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_703_port, QN => 
                           n_2895);
   DataPath_RF_BLOCKi_28_Q_reg_0_inst : DFF_X1 port map( D => n9459, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_640_port, QN => 
                           n_2896);
   DataPath_RF_BLOCKi_28_Q_reg_1_inst : DFF_X1 port map( D => n9458, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_641_port, QN => 
                           n_2897);
   DataPath_RF_BLOCKi_28_Q_reg_2_inst : DFF_X1 port map( D => n9457, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_642_port, QN => 
                           n_2898);
   DataPath_RF_BLOCKi_28_Q_reg_3_inst : DFF_X1 port map( D => n9456, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_643_port, QN => 
                           n_2899);
   DataPath_RF_BLOCKi_28_Q_reg_4_inst : DFF_X1 port map( D => n9455, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_644_port, QN => 
                           n_2900);
   DataPath_RF_BLOCKi_28_Q_reg_5_inst : DFF_X1 port map( D => n9454, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_645_port, QN => 
                           n_2901);
   DataPath_RF_BLOCKi_28_Q_reg_6_inst : DFF_X1 port map( D => n9453, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_646_port, QN => 
                           n_2902);
   DataPath_RF_BLOCKi_28_Q_reg_7_inst : DFF_X1 port map( D => n9452, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_647_port, QN => 
                           n_2903);
   DataPath_RF_BLOCKi_28_Q_reg_8_inst : DFF_X1 port map( D => n9451, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_648_port, QN => 
                           n_2904);
   DataPath_RF_BLOCKi_28_Q_reg_9_inst : DFF_X1 port map( D => n9450, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_649_port, QN => 
                           n_2905);
   DataPath_RF_BLOCKi_28_Q_reg_10_inst : DFF_X1 port map( D => n9449, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_650_port, QN => 
                           n_2906);
   DataPath_RF_BLOCKi_28_Q_reg_11_inst : DFF_X1 port map( D => n9448, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_651_port, QN => 
                           n_2907);
   DataPath_RF_BLOCKi_28_Q_reg_12_inst : DFF_X1 port map( D => n9447, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_652_port, QN => 
                           n_2908);
   DataPath_RF_BLOCKi_28_Q_reg_13_inst : DFF_X1 port map( D => n9446, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_653_port, QN => 
                           n_2909);
   DataPath_RF_BLOCKi_28_Q_reg_14_inst : DFF_X1 port map( D => n9445, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_654_port, QN => 
                           n_2910);
   DataPath_RF_BLOCKi_28_Q_reg_15_inst : DFF_X1 port map( D => n9444, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_655_port, QN => 
                           n_2911);
   DataPath_RF_BLOCKi_28_Q_reg_16_inst : DFF_X1 port map( D => n9443, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_656_port, QN => 
                           n_2912);
   DataPath_RF_BLOCKi_28_Q_reg_17_inst : DFF_X1 port map( D => n9442, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_657_port, QN => 
                           n_2913);
   DataPath_RF_BLOCKi_28_Q_reg_18_inst : DFF_X1 port map( D => n9441, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_658_port, QN => 
                           n_2914);
   DataPath_RF_BLOCKi_28_Q_reg_19_inst : DFF_X1 port map( D => n9440, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_659_port, QN => 
                           n_2915);
   DataPath_RF_BLOCKi_28_Q_reg_20_inst : DFF_X1 port map( D => n9439, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_660_port, QN => 
                           n_2916);
   DataPath_RF_BLOCKi_28_Q_reg_21_inst : DFF_X1 port map( D => n9438, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_661_port, QN => 
                           n_2917);
   DataPath_RF_BLOCKi_28_Q_reg_22_inst : DFF_X1 port map( D => n9437, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_662_port, QN => 
                           n_2918);
   DataPath_RF_BLOCKi_28_Q_reg_23_inst : DFF_X1 port map( D => n9436, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_663_port, QN => 
                           n_2919);
   DataPath_RF_BLOCKi_28_Q_reg_24_inst : DFF_X1 port map( D => n9435, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_664_port, QN => 
                           n_2920);
   DataPath_RF_BLOCKi_28_Q_reg_25_inst : DFF_X1 port map( D => n9434, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_665_port, QN => 
                           n_2921);
   DataPath_RF_BLOCKi_28_Q_reg_26_inst : DFF_X1 port map( D => n9433, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_666_port, QN => 
                           n_2922);
   DataPath_RF_BLOCKi_28_Q_reg_27_inst : DFF_X1 port map( D => n9432, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_667_port, QN => 
                           n_2923);
   DataPath_RF_BLOCKi_28_Q_reg_28_inst : DFF_X1 port map( D => n9431, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_668_port, QN => 
                           n_2924);
   DataPath_RF_BLOCKi_28_Q_reg_29_inst : DFF_X1 port map( D => n9430, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_669_port, QN => 
                           n_2925);
   DataPath_RF_BLOCKi_28_Q_reg_30_inst : DFF_X1 port map( D => n9429, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_670_port, QN => 
                           n_2926);
   DataPath_RF_BLOCKi_28_Q_reg_31_inst : DFF_X1 port map( D => n9428, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_671_port, QN => 
                           n_2927);
   DataPath_RF_BLOCKi_27_Q_reg_0_inst : DFF_X1 port map( D => n9427, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_608_port, QN => 
                           n_2928);
   DataPath_RF_BLOCKi_27_Q_reg_1_inst : DFF_X1 port map( D => n9426, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_609_port, QN => 
                           n_2929);
   DataPath_RF_BLOCKi_27_Q_reg_2_inst : DFF_X1 port map( D => n9425, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_610_port, QN => 
                           n_2930);
   DataPath_RF_BLOCKi_27_Q_reg_3_inst : DFF_X1 port map( D => n9424, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_611_port, QN => 
                           n_2931);
   DataPath_RF_BLOCKi_27_Q_reg_4_inst : DFF_X1 port map( D => n9423, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_612_port, QN => 
                           n_2932);
   DataPath_RF_BLOCKi_27_Q_reg_5_inst : DFF_X1 port map( D => n9422, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_613_port, QN => 
                           n_2933);
   DataPath_RF_BLOCKi_27_Q_reg_6_inst : DFF_X1 port map( D => n9421, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_614_port, QN => 
                           n_2934);
   DataPath_RF_BLOCKi_27_Q_reg_7_inst : DFF_X1 port map( D => n9420, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_615_port, QN => 
                           n_2935);
   DataPath_RF_BLOCKi_27_Q_reg_8_inst : DFF_X1 port map( D => n9419, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_616_port, QN => 
                           n_2936);
   DataPath_RF_BLOCKi_27_Q_reg_9_inst : DFF_X1 port map( D => n9418, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_617_port, QN => 
                           n_2937);
   DataPath_RF_BLOCKi_27_Q_reg_10_inst : DFF_X1 port map( D => n9417, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_618_port, QN => 
                           n_2938);
   DataPath_RF_BLOCKi_27_Q_reg_11_inst : DFF_X1 port map( D => n9416, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_619_port, QN => 
                           n_2939);
   DataPath_RF_BLOCKi_27_Q_reg_12_inst : DFF_X1 port map( D => n9415, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_620_port, QN => 
                           n_2940);
   DataPath_RF_BLOCKi_27_Q_reg_13_inst : DFF_X1 port map( D => n9414, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_621_port, QN => 
                           n_2941);
   DataPath_RF_BLOCKi_27_Q_reg_14_inst : DFF_X1 port map( D => n9413, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_622_port, QN => 
                           n_2942);
   DataPath_RF_BLOCKi_27_Q_reg_15_inst : DFF_X1 port map( D => n9412, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_623_port, QN => 
                           n_2943);
   DataPath_RF_BLOCKi_27_Q_reg_16_inst : DFF_X1 port map( D => n9411, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_624_port, QN => 
                           n_2944);
   DataPath_RF_BLOCKi_27_Q_reg_17_inst : DFF_X1 port map( D => n9410, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_625_port, QN => 
                           n_2945);
   DataPath_RF_BLOCKi_27_Q_reg_18_inst : DFF_X1 port map( D => n9409, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_626_port, QN => 
                           n_2946);
   DataPath_RF_BLOCKi_27_Q_reg_19_inst : DFF_X1 port map( D => n9408, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_627_port, QN => 
                           n_2947);
   DataPath_RF_BLOCKi_27_Q_reg_20_inst : DFF_X1 port map( D => n9407, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_628_port, QN => 
                           n_2948);
   DataPath_RF_BLOCKi_27_Q_reg_21_inst : DFF_X1 port map( D => n9406, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_629_port, QN => 
                           n_2949);
   DataPath_RF_BLOCKi_27_Q_reg_22_inst : DFF_X1 port map( D => n9405, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_630_port, QN => 
                           n_2950);
   DataPath_RF_BLOCKi_27_Q_reg_23_inst : DFF_X1 port map( D => n9404, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_631_port, QN => 
                           n_2951);
   DataPath_RF_BLOCKi_27_Q_reg_24_inst : DFF_X1 port map( D => n9403, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_632_port, QN => 
                           n_2952);
   DataPath_RF_BLOCKi_27_Q_reg_25_inst : DFF_X1 port map( D => n9402, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_633_port, QN => 
                           n_2953);
   DataPath_RF_BLOCKi_27_Q_reg_26_inst : DFF_X1 port map( D => n9401, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_634_port, QN => 
                           n_2954);
   DataPath_RF_BLOCKi_27_Q_reg_27_inst : DFF_X1 port map( D => n9400, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_635_port, QN => 
                           n_2955);
   DataPath_RF_BLOCKi_27_Q_reg_28_inst : DFF_X1 port map( D => n9399, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_636_port, QN => 
                           n_2956);
   DataPath_RF_BLOCKi_27_Q_reg_29_inst : DFF_X1 port map( D => n9398, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_637_port, QN => 
                           n_2957);
   DataPath_RF_BLOCKi_27_Q_reg_30_inst : DFF_X1 port map( D => n9397, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_638_port, QN => 
                           n_2958);
   DataPath_RF_BLOCKi_27_Q_reg_31_inst : DFF_X1 port map( D => n9396, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_639_port, QN => 
                           n_2959);
   DataPath_RF_BLOCKi_26_Q_reg_0_inst : DFF_X1 port map( D => n9395, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_576_port, QN => 
                           n_2960);
   DataPath_RF_BLOCKi_26_Q_reg_1_inst : DFF_X1 port map( D => n9394, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_577_port, QN => 
                           n_2961);
   DataPath_RF_BLOCKi_26_Q_reg_2_inst : DFF_X1 port map( D => n9393, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_578_port, QN => 
                           n_2962);
   DataPath_RF_BLOCKi_26_Q_reg_3_inst : DFF_X1 port map( D => n9392, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_579_port, QN => 
                           n_2963);
   DataPath_RF_BLOCKi_26_Q_reg_4_inst : DFF_X1 port map( D => n9391, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_580_port, QN => 
                           n_2964);
   DataPath_RF_BLOCKi_26_Q_reg_5_inst : DFF_X1 port map( D => n9390, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_581_port, QN => 
                           n_2965);
   DataPath_RF_BLOCKi_26_Q_reg_6_inst : DFF_X1 port map( D => n9389, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_582_port, QN => 
                           n_2966);
   DataPath_RF_BLOCKi_26_Q_reg_7_inst : DFF_X1 port map( D => n9388, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_583_port, QN => 
                           n_2967);
   DataPath_RF_BLOCKi_26_Q_reg_8_inst : DFF_X1 port map( D => n9387, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_584_port, QN => 
                           n_2968);
   DataPath_RF_BLOCKi_26_Q_reg_9_inst : DFF_X1 port map( D => n9386, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_585_port, QN => 
                           n_2969);
   DataPath_RF_BLOCKi_26_Q_reg_10_inst : DFF_X1 port map( D => n9385, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_586_port, QN => 
                           n_2970);
   DataPath_RF_BLOCKi_26_Q_reg_11_inst : DFF_X1 port map( D => n9384, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_587_port, QN => 
                           n_2971);
   DataPath_RF_BLOCKi_26_Q_reg_12_inst : DFF_X1 port map( D => n9383, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_588_port, QN => 
                           n_2972);
   DataPath_RF_BLOCKi_26_Q_reg_13_inst : DFF_X1 port map( D => n9382, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_589_port, QN => 
                           n_2973);
   DataPath_RF_BLOCKi_26_Q_reg_14_inst : DFF_X1 port map( D => n9381, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_590_port, QN => 
                           n_2974);
   DataPath_RF_BLOCKi_26_Q_reg_15_inst : DFF_X1 port map( D => n9380, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_591_port, QN => 
                           n_2975);
   DataPath_RF_BLOCKi_26_Q_reg_16_inst : DFF_X1 port map( D => n9379, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_592_port, QN => 
                           n_2976);
   DataPath_RF_BLOCKi_26_Q_reg_17_inst : DFF_X1 port map( D => n9378, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_593_port, QN => 
                           n_2977);
   DataPath_RF_BLOCKi_26_Q_reg_18_inst : DFF_X1 port map( D => n9377, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_594_port, QN => 
                           n_2978);
   DataPath_RF_BLOCKi_26_Q_reg_19_inst : DFF_X1 port map( D => n9376, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_595_port, QN => 
                           n_2979);
   DataPath_RF_BLOCKi_26_Q_reg_20_inst : DFF_X1 port map( D => n9375, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_596_port, QN => 
                           n_2980);
   DataPath_RF_BLOCKi_26_Q_reg_21_inst : DFF_X1 port map( D => n9374, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_597_port, QN => 
                           n_2981);
   DataPath_RF_BLOCKi_26_Q_reg_22_inst : DFF_X1 port map( D => n9373, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_598_port, QN => 
                           n_2982);
   DataPath_RF_BLOCKi_26_Q_reg_23_inst : DFF_X1 port map( D => n9372, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_599_port, QN => 
                           n_2983);
   DataPath_RF_BLOCKi_26_Q_reg_24_inst : DFF_X1 port map( D => n9371, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_600_port, QN => 
                           n_2984);
   DataPath_RF_BLOCKi_26_Q_reg_25_inst : DFF_X1 port map( D => n9370, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_601_port, QN => 
                           n_2985);
   DataPath_RF_BLOCKi_26_Q_reg_26_inst : DFF_X1 port map( D => n9369, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_602_port, QN => 
                           n_2986);
   DataPath_RF_BLOCKi_26_Q_reg_27_inst : DFF_X1 port map( D => n9368, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_603_port, QN => 
                           n_2987);
   DataPath_RF_BLOCKi_26_Q_reg_28_inst : DFF_X1 port map( D => n9367, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_604_port, QN => 
                           n_2988);
   DataPath_RF_BLOCKi_26_Q_reg_29_inst : DFF_X1 port map( D => n9366, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_605_port, QN => 
                           n_2989);
   DataPath_RF_BLOCKi_26_Q_reg_30_inst : DFF_X1 port map( D => n9365, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_606_port, QN => 
                           n_2990);
   DataPath_RF_BLOCKi_26_Q_reg_31_inst : DFF_X1 port map( D => n9364, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_607_port, QN => 
                           n_2991);
   DataPath_RF_BLOCKi_25_Q_reg_0_inst : DFF_X1 port map( D => n9363, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_544_port, QN => 
                           n_2992);
   DataPath_RF_BLOCKi_25_Q_reg_1_inst : DFF_X1 port map( D => n9362, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_545_port, QN => 
                           n_2993);
   DataPath_RF_BLOCKi_25_Q_reg_2_inst : DFF_X1 port map( D => n9361, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_546_port, QN => 
                           n_2994);
   DataPath_RF_BLOCKi_25_Q_reg_3_inst : DFF_X1 port map( D => n9360, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_547_port, QN => 
                           n_2995);
   DataPath_RF_BLOCKi_25_Q_reg_4_inst : DFF_X1 port map( D => n9359, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_548_port, QN => 
                           n_2996);
   DataPath_RF_BLOCKi_25_Q_reg_5_inst : DFF_X1 port map( D => n9358, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_549_port, QN => 
                           n_2997);
   DataPath_RF_BLOCKi_25_Q_reg_6_inst : DFF_X1 port map( D => n9357, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_550_port, QN => 
                           n_2998);
   DataPath_RF_BLOCKi_25_Q_reg_7_inst : DFF_X1 port map( D => n9356, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_551_port, QN => 
                           n_2999);
   DataPath_RF_BLOCKi_25_Q_reg_8_inst : DFF_X1 port map( D => n9355, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_552_port, QN => 
                           n_3000);
   DataPath_RF_BLOCKi_25_Q_reg_9_inst : DFF_X1 port map( D => n9354, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_553_port, QN => 
                           n_3001);
   DataPath_RF_BLOCKi_25_Q_reg_10_inst : DFF_X1 port map( D => n9353, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_554_port, QN => 
                           n_3002);
   DataPath_RF_BLOCKi_25_Q_reg_11_inst : DFF_X1 port map( D => n9352, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_555_port, QN => 
                           n_3003);
   DataPath_RF_BLOCKi_25_Q_reg_12_inst : DFF_X1 port map( D => n9351, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_556_port, QN => 
                           n_3004);
   DataPath_RF_BLOCKi_25_Q_reg_13_inst : DFF_X1 port map( D => n9350, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_557_port, QN => 
                           n_3005);
   DataPath_RF_BLOCKi_25_Q_reg_14_inst : DFF_X1 port map( D => n9349, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_558_port, QN => 
                           n_3006);
   DataPath_RF_BLOCKi_25_Q_reg_15_inst : DFF_X1 port map( D => n9348, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_559_port, QN => 
                           n_3007);
   DataPath_RF_BLOCKi_25_Q_reg_16_inst : DFF_X1 port map( D => n9347, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_560_port, QN => 
                           n_3008);
   DataPath_RF_BLOCKi_25_Q_reg_17_inst : DFF_X1 port map( D => n9346, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_561_port, QN => 
                           n_3009);
   DataPath_RF_BLOCKi_25_Q_reg_18_inst : DFF_X1 port map( D => n9345, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_562_port, QN => 
                           n_3010);
   DataPath_RF_BLOCKi_25_Q_reg_19_inst : DFF_X1 port map( D => n9344, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_563_port, QN => 
                           n_3011);
   DataPath_RF_BLOCKi_25_Q_reg_20_inst : DFF_X1 port map( D => n9343, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_564_port, QN => 
                           n_3012);
   DataPath_RF_BLOCKi_25_Q_reg_21_inst : DFF_X1 port map( D => n9342, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_565_port, QN => 
                           n_3013);
   DataPath_RF_BLOCKi_25_Q_reg_22_inst : DFF_X1 port map( D => n9341, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_566_port, QN => 
                           n_3014);
   DataPath_RF_BLOCKi_25_Q_reg_23_inst : DFF_X1 port map( D => n9340, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_567_port, QN => 
                           n_3015);
   DataPath_RF_BLOCKi_25_Q_reg_24_inst : DFF_X1 port map( D => n9339, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_568_port, QN => 
                           n_3016);
   DataPath_RF_BLOCKi_25_Q_reg_25_inst : DFF_X1 port map( D => n9338, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_569_port, QN => 
                           n_3017);
   DataPath_RF_BLOCKi_25_Q_reg_26_inst : DFF_X1 port map( D => n9337, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_570_port, QN => 
                           n_3018);
   DataPath_RF_BLOCKi_25_Q_reg_27_inst : DFF_X1 port map( D => n9336, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_571_port, QN => 
                           n_3019);
   DataPath_RF_BLOCKi_25_Q_reg_28_inst : DFF_X1 port map( D => n9335, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_572_port, QN => 
                           n_3020);
   DataPath_RF_BLOCKi_25_Q_reg_29_inst : DFF_X1 port map( D => n9334, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_573_port, QN => 
                           n_3021);
   DataPath_RF_BLOCKi_25_Q_reg_30_inst : DFF_X1 port map( D => n9333, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_574_port, QN => 
                           n_3022);
   DataPath_RF_BLOCKi_25_Q_reg_31_inst : DFF_X1 port map( D => n9332, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_575_port, QN => 
                           n_3023);
   DataPath_RF_BLOCKi_24_Q_reg_0_inst : DFF_X1 port map( D => n9331, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_512_port, QN => 
                           n_3024);
   DataPath_RF_BLOCKi_24_Q_reg_1_inst : DFF_X1 port map( D => n9330, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_513_port, QN => 
                           n_3025);
   DataPath_RF_BLOCKi_24_Q_reg_2_inst : DFF_X1 port map( D => n9329, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_514_port, QN => 
                           n_3026);
   DataPath_RF_BLOCKi_24_Q_reg_3_inst : DFF_X1 port map( D => n9328, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_515_port, QN => 
                           n_3027);
   DataPath_RF_BLOCKi_24_Q_reg_4_inst : DFF_X1 port map( D => n9327, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_516_port, QN => 
                           n_3028);
   DataPath_RF_BLOCKi_24_Q_reg_5_inst : DFF_X1 port map( D => n9326, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_517_port, QN => 
                           n_3029);
   DataPath_RF_BLOCKi_24_Q_reg_6_inst : DFF_X1 port map( D => n9325, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_518_port, QN => 
                           n_3030);
   DataPath_RF_BLOCKi_24_Q_reg_7_inst : DFF_X1 port map( D => n9324, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_519_port, QN => 
                           n_3031);
   DataPath_RF_BLOCKi_24_Q_reg_8_inst : DFF_X1 port map( D => n9323, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_520_port, QN => 
                           n_3032);
   DataPath_RF_BLOCKi_24_Q_reg_9_inst : DFF_X1 port map( D => n9322, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_521_port, QN => 
                           n_3033);
   DataPath_RF_BLOCKi_24_Q_reg_10_inst : DFF_X1 port map( D => n9321, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_522_port, QN => 
                           n_3034);
   DataPath_RF_BLOCKi_24_Q_reg_11_inst : DFF_X1 port map( D => n9320, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_523_port, QN => 
                           n_3035);
   DataPath_RF_BLOCKi_24_Q_reg_12_inst : DFF_X1 port map( D => n9319, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_524_port, QN => 
                           n_3036);
   DataPath_RF_BLOCKi_24_Q_reg_13_inst : DFF_X1 port map( D => n9318, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_525_port, QN => 
                           n_3037);
   DataPath_RF_BLOCKi_24_Q_reg_14_inst : DFF_X1 port map( D => n9317, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_526_port, QN => 
                           n_3038);
   DataPath_RF_BLOCKi_24_Q_reg_15_inst : DFF_X1 port map( D => n9316, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_527_port, QN => 
                           n_3039);
   DataPath_RF_BLOCKi_24_Q_reg_16_inst : DFF_X1 port map( D => n9315, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_528_port, QN => 
                           n_3040);
   DataPath_RF_BLOCKi_24_Q_reg_17_inst : DFF_X1 port map( D => n9314, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_529_port, QN => 
                           n_3041);
   DataPath_RF_BLOCKi_24_Q_reg_18_inst : DFF_X1 port map( D => n9313, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_530_port, QN => 
                           n_3042);
   DataPath_RF_BLOCKi_24_Q_reg_19_inst : DFF_X1 port map( D => n9312, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_531_port, QN => 
                           n_3043);
   DataPath_RF_BLOCKi_24_Q_reg_20_inst : DFF_X1 port map( D => n9311, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_532_port, QN => 
                           n_3044);
   DataPath_RF_BLOCKi_24_Q_reg_21_inst : DFF_X1 port map( D => n9310, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_533_port, QN => 
                           n_3045);
   DataPath_RF_BLOCKi_24_Q_reg_22_inst : DFF_X1 port map( D => n9309, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_534_port, QN => 
                           n_3046);
   DataPath_RF_BLOCKi_24_Q_reg_23_inst : DFF_X1 port map( D => n9308, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_535_port, QN => 
                           n_3047);
   DataPath_RF_BLOCKi_24_Q_reg_24_inst : DFF_X1 port map( D => n9307, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_536_port, QN => 
                           n_3048);
   DataPath_RF_BLOCKi_24_Q_reg_25_inst : DFF_X1 port map( D => n9306, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_537_port, QN => 
                           n_3049);
   DataPath_RF_BLOCKi_24_Q_reg_26_inst : DFF_X1 port map( D => n9305, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_538_port, QN => 
                           n_3050);
   DataPath_RF_BLOCKi_24_Q_reg_27_inst : DFF_X1 port map( D => n9304, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_539_port, QN => 
                           n_3051);
   DataPath_RF_BLOCKi_24_Q_reg_28_inst : DFF_X1 port map( D => n9303, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_540_port, QN => 
                           n_3052);
   DataPath_RF_BLOCKi_24_Q_reg_29_inst : DFF_X1 port map( D => n9302, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_541_port, QN => 
                           n_3053);
   DataPath_RF_BLOCKi_24_Q_reg_30_inst : DFF_X1 port map( D => n9301, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_542_port, QN => 
                           n_3054);
   DataPath_RF_BLOCKi_24_Q_reg_31_inst : DFF_X1 port map( D => n9300, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_543_port, QN => 
                           n_3055);
   DataPath_RF_BLOCKi_23_Q_reg_0_inst : DFF_X1 port map( D => n9299, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_480_port, QN => 
                           n_3056);
   DataPath_RF_BLOCKi_23_Q_reg_1_inst : DFF_X1 port map( D => n9298, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_481_port, QN => 
                           n_3057);
   DataPath_RF_BLOCKi_23_Q_reg_2_inst : DFF_X1 port map( D => n9297, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_482_port, QN => 
                           n_3058);
   DataPath_RF_BLOCKi_23_Q_reg_3_inst : DFF_X1 port map( D => n9296, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_483_port, QN => 
                           n_3059);
   DataPath_RF_BLOCKi_23_Q_reg_4_inst : DFF_X1 port map( D => n9295, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_484_port, QN => 
                           n_3060);
   DataPath_RF_BLOCKi_23_Q_reg_5_inst : DFF_X1 port map( D => n9294, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_485_port, QN => 
                           n_3061);
   DataPath_RF_BLOCKi_23_Q_reg_6_inst : DFF_X1 port map( D => n9293, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_486_port, QN => 
                           n_3062);
   DataPath_RF_BLOCKi_23_Q_reg_7_inst : DFF_X1 port map( D => n9292, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_487_port, QN => 
                           n_3063);
   DataPath_RF_BLOCKi_23_Q_reg_8_inst : DFF_X1 port map( D => n9291, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_488_port, QN => 
                           n_3064);
   DataPath_RF_BLOCKi_23_Q_reg_9_inst : DFF_X1 port map( D => n9290, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_489_port, QN => 
                           n_3065);
   DataPath_RF_BLOCKi_23_Q_reg_10_inst : DFF_X1 port map( D => n9289, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_490_port, QN => 
                           n_3066);
   DataPath_RF_BLOCKi_23_Q_reg_11_inst : DFF_X1 port map( D => n9288, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_491_port, QN => 
                           n_3067);
   DataPath_RF_BLOCKi_23_Q_reg_12_inst : DFF_X1 port map( D => n9287, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_492_port, QN => 
                           n_3068);
   DataPath_RF_BLOCKi_23_Q_reg_13_inst : DFF_X1 port map( D => n9286, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_493_port, QN => 
                           n_3069);
   DataPath_RF_BLOCKi_23_Q_reg_14_inst : DFF_X1 port map( D => n9285, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_494_port, QN => 
                           n_3070);
   DataPath_RF_BLOCKi_23_Q_reg_15_inst : DFF_X1 port map( D => n9284, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_495_port, QN => 
                           n_3071);
   DataPath_RF_BLOCKi_23_Q_reg_16_inst : DFF_X1 port map( D => n9283, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_496_port, QN => 
                           n_3072);
   DataPath_RF_BLOCKi_23_Q_reg_17_inst : DFF_X1 port map( D => n9282, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_497_port, QN => 
                           n_3073);
   DataPath_RF_BLOCKi_23_Q_reg_18_inst : DFF_X1 port map( D => n9281, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_498_port, QN => 
                           n_3074);
   DataPath_RF_BLOCKi_23_Q_reg_19_inst : DFF_X1 port map( D => n9280, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_499_port, QN => 
                           n_3075);
   DataPath_RF_BLOCKi_23_Q_reg_20_inst : DFF_X1 port map( D => n9279, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_500_port, QN => 
                           n_3076);
   DataPath_RF_BLOCKi_23_Q_reg_21_inst : DFF_X1 port map( D => n9278, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_501_port, QN => 
                           n_3077);
   DataPath_RF_BLOCKi_23_Q_reg_22_inst : DFF_X1 port map( D => n9277, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_502_port, QN => 
                           n_3078);
   DataPath_RF_BLOCKi_23_Q_reg_23_inst : DFF_X1 port map( D => n9276, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_503_port, QN => 
                           n_3079);
   DataPath_RF_BLOCKi_23_Q_reg_24_inst : DFF_X1 port map( D => n9275, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_504_port, QN => 
                           n_3080);
   DataPath_RF_BLOCKi_23_Q_reg_25_inst : DFF_X1 port map( D => n9274, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_505_port, QN => 
                           n_3081);
   DataPath_RF_BLOCKi_23_Q_reg_26_inst : DFF_X1 port map( D => n9273, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_506_port, QN => 
                           n_3082);
   DataPath_RF_BLOCKi_23_Q_reg_27_inst : DFF_X1 port map( D => n9272, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_507_port, QN => 
                           n_3083);
   DataPath_RF_BLOCKi_23_Q_reg_28_inst : DFF_X1 port map( D => n9271, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_508_port, QN => 
                           n_3084);
   DataPath_RF_BLOCKi_23_Q_reg_29_inst : DFF_X1 port map( D => n9270, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_509_port, QN => 
                           n_3085);
   DataPath_RF_BLOCKi_23_Q_reg_30_inst : DFF_X1 port map( D => n9269, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_510_port, QN => 
                           n_3086);
   DataPath_RF_BLOCKi_23_Q_reg_31_inst : DFF_X1 port map( D => n9268, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_511_port, QN => 
                           n_3087);
   DataPath_RF_BLOCKi_22_Q_reg_0_inst : DFF_X1 port map( D => n9267, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_448_port, QN => 
                           n_3088);
   DataPath_RF_BLOCKi_22_Q_reg_1_inst : DFF_X1 port map( D => n9266, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_449_port, QN => 
                           n_3089);
   DataPath_RF_BLOCKi_22_Q_reg_2_inst : DFF_X1 port map( D => n9265, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_450_port, QN => 
                           n_3090);
   DataPath_RF_BLOCKi_22_Q_reg_3_inst : DFF_X1 port map( D => n9264, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_451_port, QN => 
                           n_3091);
   DataPath_RF_BLOCKi_22_Q_reg_4_inst : DFF_X1 port map( D => n9263, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_452_port, QN => 
                           n_3092);
   DataPath_RF_BLOCKi_22_Q_reg_5_inst : DFF_X1 port map( D => n9262, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_453_port, QN => 
                           n_3093);
   DataPath_RF_BLOCKi_22_Q_reg_6_inst : DFF_X1 port map( D => n9261, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_454_port, QN => 
                           n_3094);
   DataPath_RF_BLOCKi_22_Q_reg_7_inst : DFF_X1 port map( D => n9260, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_455_port, QN => 
                           n_3095);
   DataPath_RF_BLOCKi_22_Q_reg_8_inst : DFF_X1 port map( D => n9259, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_456_port, QN => 
                           n_3096);
   DataPath_RF_BLOCKi_22_Q_reg_9_inst : DFF_X1 port map( D => n9258, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_457_port, QN => 
                           n_3097);
   DataPath_RF_BLOCKi_22_Q_reg_10_inst : DFF_X1 port map( D => n9257, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_458_port, QN => 
                           n_3098);
   DataPath_RF_BLOCKi_22_Q_reg_11_inst : DFF_X1 port map( D => n9256, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_459_port, QN => 
                           n_3099);
   DataPath_RF_BLOCKi_22_Q_reg_12_inst : DFF_X1 port map( D => n9255, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_460_port, QN => 
                           n_3100);
   DataPath_RF_BLOCKi_22_Q_reg_13_inst : DFF_X1 port map( D => n9254, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_461_port, QN => 
                           n_3101);
   DataPath_RF_BLOCKi_22_Q_reg_14_inst : DFF_X1 port map( D => n9253, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_462_port, QN => 
                           n_3102);
   DataPath_RF_BLOCKi_22_Q_reg_15_inst : DFF_X1 port map( D => n9252, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_463_port, QN => 
                           n_3103);
   DataPath_RF_BLOCKi_22_Q_reg_16_inst : DFF_X1 port map( D => n9251, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_464_port, QN => 
                           n_3104);
   DataPath_RF_BLOCKi_22_Q_reg_17_inst : DFF_X1 port map( D => n9250, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_465_port, QN => 
                           n_3105);
   DataPath_RF_BLOCKi_22_Q_reg_18_inst : DFF_X1 port map( D => n9249, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_466_port, QN => 
                           n_3106);
   DataPath_RF_BLOCKi_22_Q_reg_19_inst : DFF_X1 port map( D => n9248, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_467_port, QN => 
                           n_3107);
   DataPath_RF_BLOCKi_22_Q_reg_20_inst : DFF_X1 port map( D => n9247, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_468_port, QN => 
                           n_3108);
   DataPath_RF_BLOCKi_22_Q_reg_21_inst : DFF_X1 port map( D => n9246, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_469_port, QN => 
                           n_3109);
   DataPath_RF_BLOCKi_22_Q_reg_22_inst : DFF_X1 port map( D => n9245, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_470_port, QN => 
                           n_3110);
   DataPath_RF_BLOCKi_22_Q_reg_23_inst : DFF_X1 port map( D => n9244, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_471_port, QN => 
                           n_3111);
   DataPath_RF_BLOCKi_22_Q_reg_24_inst : DFF_X1 port map( D => n9243, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_472_port, QN => 
                           n_3112);
   DataPath_RF_BLOCKi_22_Q_reg_25_inst : DFF_X1 port map( D => n9242, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_473_port, QN => 
                           n_3113);
   DataPath_RF_BLOCKi_22_Q_reg_26_inst : DFF_X1 port map( D => n9241, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_474_port, QN => 
                           n_3114);
   DataPath_RF_BLOCKi_22_Q_reg_27_inst : DFF_X1 port map( D => n9240, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_475_port, QN => 
                           n_3115);
   DataPath_RF_BLOCKi_22_Q_reg_28_inst : DFF_X1 port map( D => n9239, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_476_port, QN => 
                           n_3116);
   DataPath_RF_BLOCKi_22_Q_reg_29_inst : DFF_X1 port map( D => n9238, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_477_port, QN => 
                           n_3117);
   DataPath_RF_BLOCKi_22_Q_reg_30_inst : DFF_X1 port map( D => n9237, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_478_port, QN => 
                           n_3118);
   DataPath_RF_BLOCKi_22_Q_reg_31_inst : DFF_X1 port map( D => n9236, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_479_port, QN => 
                           n_3119);
   DataPath_RF_BLOCKi_21_Q_reg_0_inst : DFF_X1 port map( D => n9235, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_416_port, QN => 
                           n_3120);
   DataPath_RF_BLOCKi_21_Q_reg_1_inst : DFF_X1 port map( D => n9234, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_417_port, QN => 
                           n_3121);
   DataPath_RF_BLOCKi_21_Q_reg_2_inst : DFF_X1 port map( D => n9233, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_418_port, QN => 
                           n_3122);
   DataPath_RF_BLOCKi_21_Q_reg_3_inst : DFF_X1 port map( D => n9232, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_419_port, QN => 
                           n_3123);
   DataPath_RF_BLOCKi_21_Q_reg_4_inst : DFF_X1 port map( D => n9231, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_420_port, QN => 
                           n_3124);
   DataPath_RF_BLOCKi_21_Q_reg_5_inst : DFF_X1 port map( D => n9230, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_421_port, QN => 
                           n_3125);
   DataPath_RF_BLOCKi_21_Q_reg_6_inst : DFF_X1 port map( D => n9229, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_422_port, QN => 
                           n_3126);
   DataPath_RF_BLOCKi_21_Q_reg_7_inst : DFF_X1 port map( D => n9228, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_423_port, QN => 
                           n_3127);
   DataPath_RF_BLOCKi_21_Q_reg_8_inst : DFF_X1 port map( D => n9227, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_424_port, QN => 
                           n_3128);
   DataPath_RF_BLOCKi_21_Q_reg_9_inst : DFF_X1 port map( D => n9226, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_425_port, QN => 
                           n_3129);
   DataPath_RF_BLOCKi_21_Q_reg_10_inst : DFF_X1 port map( D => n9225, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_426_port, QN => 
                           n_3130);
   DataPath_RF_BLOCKi_21_Q_reg_11_inst : DFF_X1 port map( D => n9224, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_427_port, QN => 
                           n_3131);
   DataPath_RF_BLOCKi_21_Q_reg_12_inst : DFF_X1 port map( D => n9223, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_428_port, QN => 
                           n_3132);
   DataPath_RF_BLOCKi_21_Q_reg_13_inst : DFF_X1 port map( D => n9222, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_429_port, QN => 
                           n_3133);
   DataPath_RF_BLOCKi_21_Q_reg_14_inst : DFF_X1 port map( D => n9221, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_430_port, QN => 
                           n_3134);
   DataPath_RF_BLOCKi_21_Q_reg_15_inst : DFF_X1 port map( D => n9220, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_431_port, QN => 
                           n_3135);
   DataPath_RF_BLOCKi_21_Q_reg_16_inst : DFF_X1 port map( D => n9219, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_432_port, QN => 
                           n_3136);
   DataPath_RF_BLOCKi_21_Q_reg_17_inst : DFF_X1 port map( D => n9218, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_433_port, QN => 
                           n_3137);
   DataPath_RF_BLOCKi_21_Q_reg_18_inst : DFF_X1 port map( D => n9217, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_434_port, QN => 
                           n_3138);
   DataPath_RF_BLOCKi_21_Q_reg_19_inst : DFF_X1 port map( D => n9216, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_435_port, QN => 
                           n_3139);
   DataPath_RF_BLOCKi_21_Q_reg_20_inst : DFF_X1 port map( D => n9215, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_436_port, QN => 
                           n_3140);
   DataPath_RF_BLOCKi_21_Q_reg_21_inst : DFF_X1 port map( D => n9214, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_437_port, QN => 
                           n_3141);
   DataPath_RF_BLOCKi_21_Q_reg_22_inst : DFF_X1 port map( D => n9213, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_438_port, QN => 
                           n_3142);
   DataPath_RF_BLOCKi_21_Q_reg_23_inst : DFF_X1 port map( D => n9212, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_439_port, QN => 
                           n_3143);
   DataPath_RF_BLOCKi_21_Q_reg_24_inst : DFF_X1 port map( D => n9211, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_440_port, QN => 
                           n_3144);
   DataPath_RF_BLOCKi_21_Q_reg_25_inst : DFF_X1 port map( D => n9210, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_441_port, QN => 
                           n_3145);
   DataPath_RF_BLOCKi_21_Q_reg_26_inst : DFF_X1 port map( D => n9209, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_442_port, QN => 
                           n_3146);
   DataPath_RF_BLOCKi_21_Q_reg_27_inst : DFF_X1 port map( D => n9208, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_443_port, QN => 
                           n_3147);
   DataPath_RF_BLOCKi_21_Q_reg_28_inst : DFF_X1 port map( D => n9207, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_444_port, QN => 
                           n_3148);
   DataPath_RF_BLOCKi_21_Q_reg_29_inst : DFF_X1 port map( D => n9206, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_445_port, QN => 
                           n_3149);
   DataPath_RF_BLOCKi_21_Q_reg_30_inst : DFF_X1 port map( D => n9205, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_446_port, QN => 
                           n_3150);
   DataPath_RF_BLOCKi_21_Q_reg_31_inst : DFF_X1 port map( D => n9204, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_447_port, QN => 
                           n_3151);
   DataPath_RF_BLOCKi_20_Q_reg_0_inst : DFF_X1 port map( D => n9203, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_384_port, QN => 
                           n_3152);
   DataPath_RF_BLOCKi_20_Q_reg_1_inst : DFF_X1 port map( D => n9202, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_385_port, QN => 
                           n_3153);
   DataPath_RF_BLOCKi_20_Q_reg_2_inst : DFF_X1 port map( D => n9201, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_386_port, QN => 
                           n_3154);
   DataPath_RF_BLOCKi_20_Q_reg_3_inst : DFF_X1 port map( D => n9200, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_387_port, QN => 
                           n_3155);
   DataPath_RF_BLOCKi_20_Q_reg_4_inst : DFF_X1 port map( D => n9199, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_388_port, QN => 
                           n_3156);
   DataPath_RF_BLOCKi_20_Q_reg_5_inst : DFF_X1 port map( D => n9198, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_389_port, QN => 
                           n_3157);
   DataPath_RF_BLOCKi_20_Q_reg_6_inst : DFF_X1 port map( D => n9197, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_390_port, QN => 
                           n_3158);
   DataPath_RF_BLOCKi_20_Q_reg_7_inst : DFF_X1 port map( D => n9196, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_391_port, QN => 
                           n_3159);
   DataPath_RF_BLOCKi_20_Q_reg_8_inst : DFF_X1 port map( D => n9195, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_392_port, QN => 
                           n_3160);
   DataPath_RF_BLOCKi_20_Q_reg_9_inst : DFF_X1 port map( D => n9194, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_393_port, QN => 
                           n_3161);
   DataPath_RF_BLOCKi_20_Q_reg_10_inst : DFF_X1 port map( D => n9193, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_394_port, QN => 
                           n_3162);
   DataPath_RF_BLOCKi_20_Q_reg_11_inst : DFF_X1 port map( D => n9192, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_395_port, QN => 
                           n_3163);
   DataPath_RF_BLOCKi_20_Q_reg_12_inst : DFF_X1 port map( D => n9191, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_396_port, QN => 
                           n_3164);
   DataPath_RF_BLOCKi_20_Q_reg_13_inst : DFF_X1 port map( D => n9190, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_397_port, QN => 
                           n_3165);
   DataPath_RF_BLOCKi_20_Q_reg_14_inst : DFF_X1 port map( D => n9189, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_398_port, QN => 
                           n_3166);
   DataPath_RF_BLOCKi_20_Q_reg_15_inst : DFF_X1 port map( D => n9188, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_399_port, QN => 
                           n_3167);
   DataPath_RF_BLOCKi_20_Q_reg_16_inst : DFF_X1 port map( D => n9187, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_400_port, QN => 
                           n_3168);
   DataPath_RF_BLOCKi_20_Q_reg_17_inst : DFF_X1 port map( D => n9186, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_401_port, QN => 
                           n_3169);
   DataPath_RF_BLOCKi_20_Q_reg_18_inst : DFF_X1 port map( D => n9185, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_402_port, QN => 
                           n_3170);
   DataPath_RF_BLOCKi_20_Q_reg_19_inst : DFF_X1 port map( D => n9184, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_403_port, QN => 
                           n_3171);
   DataPath_RF_BLOCKi_20_Q_reg_20_inst : DFF_X1 port map( D => n9183, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_404_port, QN => 
                           n_3172);
   DataPath_RF_BLOCKi_20_Q_reg_21_inst : DFF_X1 port map( D => n9182, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_405_port, QN => 
                           n_3173);
   DataPath_RF_BLOCKi_20_Q_reg_22_inst : DFF_X1 port map( D => n9181, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_406_port, QN => 
                           n_3174);
   DataPath_RF_BLOCKi_20_Q_reg_23_inst : DFF_X1 port map( D => n9180, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_407_port, QN => 
                           n_3175);
   DataPath_RF_BLOCKi_20_Q_reg_24_inst : DFF_X1 port map( D => n9179, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_408_port, QN => 
                           n_3176);
   DataPath_RF_BLOCKi_20_Q_reg_25_inst : DFF_X1 port map( D => n9178, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_409_port, QN => 
                           n_3177);
   DataPath_RF_BLOCKi_20_Q_reg_26_inst : DFF_X1 port map( D => n9177, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_410_port, QN => 
                           n_3178);
   DataPath_RF_BLOCKi_20_Q_reg_27_inst : DFF_X1 port map( D => n9176, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_411_port, QN => 
                           n_3179);
   DataPath_RF_BLOCKi_20_Q_reg_28_inst : DFF_X1 port map( D => n9175, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_412_port, QN => 
                           n_3180);
   DataPath_RF_BLOCKi_20_Q_reg_29_inst : DFF_X1 port map( D => n9174, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_413_port, QN => 
                           n_3181);
   DataPath_RF_BLOCKi_20_Q_reg_30_inst : DFF_X1 port map( D => n9173, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_414_port, QN => 
                           n_3182);
   DataPath_RF_BLOCKi_20_Q_reg_31_inst : DFF_X1 port map( D => n9172, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_415_port, QN => 
                           n_3183);
   DataPath_RF_BLOCKi_19_Q_reg_0_inst : DFF_X1 port map( D => n9171, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_352_port, QN => 
                           n_3184);
   DataPath_RF_BLOCKi_19_Q_reg_1_inst : DFF_X1 port map( D => n9170, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_353_port, QN => 
                           n_3185);
   DataPath_RF_BLOCKi_19_Q_reg_2_inst : DFF_X1 port map( D => n9169, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_354_port, QN => 
                           n_3186);
   DataPath_RF_BLOCKi_19_Q_reg_3_inst : DFF_X1 port map( D => n9168, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_355_port, QN => 
                           n_3187);
   DataPath_RF_BLOCKi_19_Q_reg_4_inst : DFF_X1 port map( D => n9167, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_356_port, QN => 
                           n_3188);
   DataPath_RF_BLOCKi_19_Q_reg_5_inst : DFF_X1 port map( D => n9166, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_357_port, QN => 
                           n_3189);
   DataPath_RF_BLOCKi_19_Q_reg_6_inst : DFF_X1 port map( D => n9165, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_358_port, QN => 
                           n_3190);
   DataPath_RF_BLOCKi_19_Q_reg_7_inst : DFF_X1 port map( D => n9164, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_359_port, QN => 
                           n_3191);
   DataPath_RF_BLOCKi_19_Q_reg_8_inst : DFF_X1 port map( D => n9163, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_360_port, QN => 
                           n_3192);
   DataPath_RF_BLOCKi_19_Q_reg_9_inst : DFF_X1 port map( D => n9162, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_361_port, QN => 
                           n_3193);
   DataPath_RF_BLOCKi_19_Q_reg_10_inst : DFF_X1 port map( D => n9161, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_362_port, QN => 
                           n_3194);
   DataPath_RF_BLOCKi_19_Q_reg_11_inst : DFF_X1 port map( D => n9160, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_363_port, QN => 
                           n_3195);
   DataPath_RF_BLOCKi_19_Q_reg_12_inst : DFF_X1 port map( D => n9159, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_364_port, QN => 
                           n_3196);
   DataPath_RF_BLOCKi_19_Q_reg_13_inst : DFF_X1 port map( D => n9158, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_365_port, QN => 
                           n_3197);
   DataPath_RF_BLOCKi_19_Q_reg_14_inst : DFF_X1 port map( D => n9157, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_366_port, QN => 
                           n_3198);
   DataPath_RF_BLOCKi_19_Q_reg_15_inst : DFF_X1 port map( D => n9156, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_367_port, QN => 
                           n_3199);
   DataPath_RF_BLOCKi_19_Q_reg_16_inst : DFF_X1 port map( D => n9155, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_368_port, QN => 
                           n_3200);
   DataPath_RF_BLOCKi_19_Q_reg_17_inst : DFF_X1 port map( D => n9154, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_369_port, QN => 
                           n_3201);
   DataPath_RF_BLOCKi_19_Q_reg_18_inst : DFF_X1 port map( D => n9153, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_370_port, QN => 
                           n_3202);
   DataPath_RF_BLOCKi_19_Q_reg_19_inst : DFF_X1 port map( D => n9152, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_371_port, QN => 
                           n_3203);
   DataPath_RF_BLOCKi_19_Q_reg_20_inst : DFF_X1 port map( D => n9151, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_372_port, QN => 
                           n_3204);
   DataPath_RF_BLOCKi_19_Q_reg_21_inst : DFF_X1 port map( D => n9150, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_373_port, QN => 
                           n_3205);
   DataPath_RF_BLOCKi_19_Q_reg_22_inst : DFF_X1 port map( D => n9149, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_374_port, QN => 
                           n_3206);
   DataPath_RF_BLOCKi_19_Q_reg_23_inst : DFF_X1 port map( D => n9148, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_375_port, QN => 
                           n_3207);
   DataPath_RF_BLOCKi_19_Q_reg_24_inst : DFF_X1 port map( D => n9147, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_376_port, QN => 
                           n_3208);
   DataPath_RF_BLOCKi_19_Q_reg_25_inst : DFF_X1 port map( D => n9146, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_377_port, QN => 
                           n_3209);
   DataPath_RF_BLOCKi_19_Q_reg_26_inst : DFF_X1 port map( D => n9145, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_378_port, QN => 
                           n_3210);
   DataPath_RF_BLOCKi_19_Q_reg_27_inst : DFF_X1 port map( D => n9144, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_379_port, QN => 
                           n_3211);
   DataPath_RF_BLOCKi_19_Q_reg_28_inst : DFF_X1 port map( D => n9143, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_380_port, QN => 
                           n_3212);
   DataPath_RF_BLOCKi_19_Q_reg_29_inst : DFF_X1 port map( D => n9142, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_381_port, QN => 
                           n_3213);
   DataPath_RF_BLOCKi_19_Q_reg_30_inst : DFF_X1 port map( D => n9141, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_382_port, QN => 
                           n_3214);
   DataPath_RF_BLOCKi_19_Q_reg_31_inst : DFF_X1 port map( D => n9140, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_383_port, QN => 
                           n_3215);
   DataPath_RF_BLOCKi_18_Q_reg_0_inst : DFF_X1 port map( D => n9139, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_320_port, QN => 
                           n_3216);
   DataPath_RF_BLOCKi_18_Q_reg_1_inst : DFF_X1 port map( D => n9138, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_321_port, QN => 
                           n_3217);
   DataPath_RF_BLOCKi_18_Q_reg_2_inst : DFF_X1 port map( D => n9137, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_322_port, QN => 
                           n_3218);
   DataPath_RF_BLOCKi_18_Q_reg_3_inst : DFF_X1 port map( D => n9136, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_323_port, QN => 
                           n_3219);
   DataPath_RF_BLOCKi_18_Q_reg_4_inst : DFF_X1 port map( D => n9135, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_324_port, QN => 
                           n_3220);
   DataPath_RF_BLOCKi_18_Q_reg_5_inst : DFF_X1 port map( D => n9134, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_325_port, QN => 
                           n_3221);
   DataPath_RF_BLOCKi_18_Q_reg_6_inst : DFF_X1 port map( D => n9133, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_326_port, QN => 
                           n_3222);
   DataPath_RF_BLOCKi_18_Q_reg_7_inst : DFF_X1 port map( D => n9132, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_327_port, QN => 
                           n_3223);
   DataPath_RF_BLOCKi_18_Q_reg_8_inst : DFF_X1 port map( D => n9131, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_328_port, QN => 
                           n_3224);
   DataPath_RF_BLOCKi_18_Q_reg_9_inst : DFF_X1 port map( D => n9130, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_329_port, QN => 
                           n_3225);
   DataPath_RF_BLOCKi_18_Q_reg_10_inst : DFF_X1 port map( D => n9129, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_330_port, QN => 
                           n_3226);
   DataPath_RF_BLOCKi_18_Q_reg_11_inst : DFF_X1 port map( D => n9128, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_331_port, QN => 
                           n_3227);
   DataPath_RF_BLOCKi_18_Q_reg_12_inst : DFF_X1 port map( D => n9127, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_332_port, QN => 
                           n_3228);
   DataPath_RF_BLOCKi_18_Q_reg_13_inst : DFF_X1 port map( D => n9126, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_333_port, QN => 
                           n_3229);
   DataPath_RF_BLOCKi_18_Q_reg_14_inst : DFF_X1 port map( D => n9125, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_334_port, QN => 
                           n_3230);
   DataPath_RF_BLOCKi_18_Q_reg_15_inst : DFF_X1 port map( D => n9124, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_335_port, QN => 
                           n_3231);
   DataPath_RF_BLOCKi_18_Q_reg_16_inst : DFF_X1 port map( D => n9123, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_336_port, QN => 
                           n_3232);
   DataPath_RF_BLOCKi_18_Q_reg_17_inst : DFF_X1 port map( D => n9122, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_337_port, QN => 
                           n_3233);
   DataPath_RF_BLOCKi_18_Q_reg_18_inst : DFF_X1 port map( D => n9121, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_338_port, QN => 
                           n_3234);
   DataPath_RF_BLOCKi_18_Q_reg_19_inst : DFF_X1 port map( D => n9120, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_339_port, QN => 
                           n_3235);
   DataPath_RF_BLOCKi_18_Q_reg_20_inst : DFF_X1 port map( D => n9119, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_340_port, QN => 
                           n_3236);
   DataPath_RF_BLOCKi_18_Q_reg_21_inst : DFF_X1 port map( D => n9118, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_341_port, QN => 
                           n_3237);
   DataPath_RF_BLOCKi_18_Q_reg_22_inst : DFF_X1 port map( D => n9117, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_342_port, QN => 
                           n_3238);
   DataPath_RF_BLOCKi_18_Q_reg_23_inst : DFF_X1 port map( D => n9116, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_343_port, QN => 
                           n_3239);
   DataPath_RF_BLOCKi_18_Q_reg_24_inst : DFF_X1 port map( D => n9115, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_344_port, QN => 
                           n_3240);
   DataPath_RF_BLOCKi_18_Q_reg_25_inst : DFF_X1 port map( D => n9114, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_345_port, QN => 
                           n_3241);
   DataPath_RF_BLOCKi_18_Q_reg_26_inst : DFF_X1 port map( D => n9113, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_346_port, QN => 
                           n_3242);
   DataPath_RF_BLOCKi_18_Q_reg_27_inst : DFF_X1 port map( D => n9112, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_347_port, QN => 
                           n_3243);
   DataPath_RF_BLOCKi_18_Q_reg_28_inst : DFF_X1 port map( D => n9111, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_348_port, QN => 
                           n_3244);
   DataPath_RF_BLOCKi_18_Q_reg_29_inst : DFF_X1 port map( D => n9110, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_349_port, QN => 
                           n_3245);
   DataPath_RF_BLOCKi_18_Q_reg_30_inst : DFF_X1 port map( D => n9109, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_350_port, QN => 
                           n_3246);
   DataPath_RF_BLOCKi_18_Q_reg_31_inst : DFF_X1 port map( D => n9108, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_351_port, QN => 
                           n_3247);
   DataPath_RF_BLOCKi_17_Q_reg_0_inst : DFF_X1 port map( D => n9107, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_288_port, QN => 
                           n_3248);
   DataPath_RF_BLOCKi_17_Q_reg_1_inst : DFF_X1 port map( D => n9106, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_289_port, QN => 
                           n_3249);
   DataPath_RF_BLOCKi_17_Q_reg_2_inst : DFF_X1 port map( D => n9105, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_290_port, QN => 
                           n_3250);
   DataPath_RF_BLOCKi_17_Q_reg_3_inst : DFF_X1 port map( D => n9104, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_291_port, QN => 
                           n_3251);
   DataPath_RF_BLOCKi_17_Q_reg_4_inst : DFF_X1 port map( D => n9103, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_292_port, QN => 
                           n_3252);
   DataPath_RF_BLOCKi_17_Q_reg_5_inst : DFF_X1 port map( D => n9102, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_293_port, QN => 
                           n_3253);
   DataPath_RF_BLOCKi_17_Q_reg_6_inst : DFF_X1 port map( D => n9101, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_294_port, QN => 
                           n_3254);
   DataPath_RF_BLOCKi_17_Q_reg_7_inst : DFF_X1 port map( D => n9100, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_295_port, QN => 
                           n_3255);
   DataPath_RF_BLOCKi_17_Q_reg_8_inst : DFF_X1 port map( D => n9099, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_296_port, QN => 
                           n_3256);
   DataPath_RF_BLOCKi_17_Q_reg_9_inst : DFF_X1 port map( D => n9098, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_297_port, QN => 
                           n_3257);
   DataPath_RF_BLOCKi_17_Q_reg_10_inst : DFF_X1 port map( D => n9097, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_298_port, QN => 
                           n_3258);
   DataPath_RF_BLOCKi_17_Q_reg_11_inst : DFF_X1 port map( D => n9096, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_299_port, QN => 
                           n_3259);
   DataPath_RF_BLOCKi_17_Q_reg_12_inst : DFF_X1 port map( D => n9095, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_300_port, QN => 
                           n_3260);
   DataPath_RF_BLOCKi_17_Q_reg_13_inst : DFF_X1 port map( D => n9094, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_301_port, QN => 
                           n_3261);
   DataPath_RF_BLOCKi_17_Q_reg_14_inst : DFF_X1 port map( D => n9093, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_302_port, QN => 
                           n_3262);
   DataPath_RF_BLOCKi_17_Q_reg_15_inst : DFF_X1 port map( D => n9092, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_303_port, QN => 
                           n_3263);
   DataPath_RF_BLOCKi_17_Q_reg_16_inst : DFF_X1 port map( D => n9091, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_304_port, QN => 
                           n_3264);
   DataPath_RF_BLOCKi_17_Q_reg_17_inst : DFF_X1 port map( D => n9090, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_305_port, QN => 
                           n_3265);
   DataPath_RF_BLOCKi_17_Q_reg_18_inst : DFF_X1 port map( D => n9089, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_306_port, QN => 
                           n_3266);
   DataPath_RF_BLOCKi_17_Q_reg_19_inst : DFF_X1 port map( D => n9088, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_307_port, QN => 
                           n_3267);
   DataPath_RF_BLOCKi_17_Q_reg_20_inst : DFF_X1 port map( D => n9087, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_308_port, QN => 
                           n_3268);
   DataPath_RF_BLOCKi_17_Q_reg_21_inst : DFF_X1 port map( D => n9086, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_309_port, QN => 
                           n_3269);
   DataPath_RF_BLOCKi_17_Q_reg_22_inst : DFF_X1 port map( D => n9085, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_310_port, QN => 
                           n_3270);
   DataPath_RF_BLOCKi_17_Q_reg_23_inst : DFF_X1 port map( D => n9084, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_311_port, QN => 
                           n_3271);
   DataPath_RF_BLOCKi_17_Q_reg_24_inst : DFF_X1 port map( D => n9083, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_312_port, QN => 
                           n_3272);
   DataPath_RF_BLOCKi_17_Q_reg_25_inst : DFF_X1 port map( D => n9082, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_313_port, QN => 
                           n_3273);
   DataPath_RF_BLOCKi_17_Q_reg_26_inst : DFF_X1 port map( D => n9081, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_314_port, QN => 
                           n_3274);
   DataPath_RF_BLOCKi_17_Q_reg_27_inst : DFF_X1 port map( D => n9080, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_315_port, QN => 
                           n_3275);
   DataPath_RF_BLOCKi_17_Q_reg_28_inst : DFF_X1 port map( D => n9079, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_316_port, QN => 
                           n_3276);
   DataPath_RF_BLOCKi_17_Q_reg_29_inst : DFF_X1 port map( D => n9078, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_317_port, QN => 
                           n_3277);
   DataPath_RF_BLOCKi_17_Q_reg_30_inst : DFF_X1 port map( D => n9077, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_318_port, QN => 
                           n_3278);
   DataPath_RF_BLOCKi_17_Q_reg_31_inst : DFF_X1 port map( D => n9076, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_319_port, QN => 
                           n_3279);
   DataPath_RF_BLOCKi_16_Q_reg_0_inst : DFF_X1 port map( D => n9075, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_256_port, QN => 
                           n_3280);
   DataPath_RF_BLOCKi_16_Q_reg_1_inst : DFF_X1 port map( D => n9074, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_257_port, QN => 
                           n_3281);
   DataPath_RF_BLOCKi_16_Q_reg_2_inst : DFF_X1 port map( D => n9073, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_258_port, QN => 
                           n_3282);
   DataPath_RF_BLOCKi_16_Q_reg_3_inst : DFF_X1 port map( D => n9072, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_259_port, QN => 
                           n_3283);
   DataPath_RF_BLOCKi_16_Q_reg_4_inst : DFF_X1 port map( D => n9071, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_260_port, QN => 
                           n_3284);
   DataPath_RF_BLOCKi_16_Q_reg_5_inst : DFF_X1 port map( D => n9070, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_261_port, QN => 
                           n_3285);
   DataPath_RF_BLOCKi_16_Q_reg_6_inst : DFF_X1 port map( D => n9069, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_262_port, QN => 
                           n_3286);
   DataPath_RF_BLOCKi_16_Q_reg_7_inst : DFF_X1 port map( D => n9068, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_263_port, QN => 
                           n_3287);
   DataPath_RF_BLOCKi_16_Q_reg_8_inst : DFF_X1 port map( D => n9067, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_264_port, QN => 
                           n_3288);
   DataPath_RF_BLOCKi_16_Q_reg_9_inst : DFF_X1 port map( D => n9066, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_265_port, QN => 
                           n_3289);
   DataPath_RF_BLOCKi_16_Q_reg_10_inst : DFF_X1 port map( D => n9065, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_266_port, QN => 
                           n_3290);
   DataPath_RF_BLOCKi_16_Q_reg_11_inst : DFF_X1 port map( D => n9064, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_267_port, QN => 
                           n_3291);
   DataPath_RF_BLOCKi_16_Q_reg_12_inst : DFF_X1 port map( D => n9063, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_268_port, QN => 
                           n_3292);
   DataPath_RF_BLOCKi_16_Q_reg_13_inst : DFF_X1 port map( D => n9062, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_269_port, QN => 
                           n_3293);
   DataPath_RF_BLOCKi_16_Q_reg_14_inst : DFF_X1 port map( D => n9061, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_270_port, QN => 
                           n_3294);
   DataPath_RF_BLOCKi_16_Q_reg_15_inst : DFF_X1 port map( D => n9060, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_271_port, QN => 
                           n_3295);
   DataPath_RF_BLOCKi_16_Q_reg_16_inst : DFF_X1 port map( D => n9059, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_272_port, QN => 
                           n_3296);
   DataPath_RF_BLOCKi_16_Q_reg_17_inst : DFF_X1 port map( D => n9058, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_273_port, QN => 
                           n_3297);
   DataPath_RF_BLOCKi_16_Q_reg_18_inst : DFF_X1 port map( D => n9057, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_274_port, QN => 
                           n_3298);
   DataPath_RF_BLOCKi_16_Q_reg_19_inst : DFF_X1 port map( D => n9056, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_275_port, QN => 
                           n_3299);
   DataPath_RF_BLOCKi_16_Q_reg_20_inst : DFF_X1 port map( D => n9055, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_276_port, QN => 
                           n_3300);
   DataPath_RF_BLOCKi_16_Q_reg_21_inst : DFF_X1 port map( D => n9054, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_277_port, QN => 
                           n_3301);
   DataPath_RF_BLOCKi_16_Q_reg_22_inst : DFF_X1 port map( D => n9053, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_278_port, QN => 
                           n_3302);
   DataPath_RF_BLOCKi_16_Q_reg_23_inst : DFF_X1 port map( D => n9052, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_279_port, QN => 
                           n_3303);
   DataPath_RF_BLOCKi_16_Q_reg_24_inst : DFF_X1 port map( D => n9051, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_280_port, QN => 
                           n_3304);
   DataPath_RF_BLOCKi_16_Q_reg_25_inst : DFF_X1 port map( D => n9050, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_281_port, QN => 
                           n_3305);
   DataPath_RF_BLOCKi_16_Q_reg_26_inst : DFF_X1 port map( D => n9049, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_282_port, QN => 
                           n_3306);
   DataPath_RF_BLOCKi_16_Q_reg_27_inst : DFF_X1 port map( D => n9048, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_283_port, QN => 
                           n_3307);
   DataPath_RF_BLOCKi_16_Q_reg_28_inst : DFF_X1 port map( D => n9047, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_284_port, QN => 
                           n_3308);
   DataPath_RF_BLOCKi_16_Q_reg_29_inst : DFF_X1 port map( D => n9046, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_285_port, QN => 
                           n_3309);
   DataPath_RF_BLOCKi_16_Q_reg_30_inst : DFF_X1 port map( D => n9045, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_286_port, QN => 
                           n_3310);
   DataPath_RF_BLOCKi_16_Q_reg_31_inst : DFF_X1 port map( D => n9044, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_287_port, QN => 
                           n_3311);
   DataPath_RF_BLOCKi_15_Q_reg_0_inst : DFF_X1 port map( D => n9043, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_224_port, QN => 
                           n_3312);
   DataPath_RF_BLOCKi_15_Q_reg_1_inst : DFF_X1 port map( D => n9042, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_225_port, QN => 
                           n_3313);
   DataPath_RF_BLOCKi_15_Q_reg_2_inst : DFF_X1 port map( D => n9041, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_226_port, QN => 
                           n_3314);
   DataPath_RF_BLOCKi_15_Q_reg_3_inst : DFF_X1 port map( D => n9040, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_227_port, QN => 
                           n_3315);
   DataPath_RF_BLOCKi_15_Q_reg_4_inst : DFF_X1 port map( D => n9039, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_228_port, QN => 
                           n_3316);
   DataPath_RF_BLOCKi_15_Q_reg_5_inst : DFF_X1 port map( D => n9038, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_229_port, QN => 
                           n_3317);
   DataPath_RF_BLOCKi_15_Q_reg_6_inst : DFF_X1 port map( D => n9037, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_230_port, QN => 
                           n_3318);
   DataPath_RF_BLOCKi_15_Q_reg_7_inst : DFF_X1 port map( D => n9036, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_231_port, QN => 
                           n_3319);
   DataPath_RF_BLOCKi_15_Q_reg_8_inst : DFF_X1 port map( D => n9035, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_232_port, QN => 
                           n_3320);
   DataPath_RF_BLOCKi_15_Q_reg_9_inst : DFF_X1 port map( D => n9034, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_233_port, QN => 
                           n_3321);
   DataPath_RF_BLOCKi_15_Q_reg_10_inst : DFF_X1 port map( D => n9033, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_234_port, QN => 
                           n_3322);
   DataPath_RF_BLOCKi_15_Q_reg_11_inst : DFF_X1 port map( D => n9032, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_235_port, QN => 
                           n_3323);
   DataPath_RF_BLOCKi_15_Q_reg_12_inst : DFF_X1 port map( D => n9031, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_236_port, QN => 
                           n_3324);
   DataPath_RF_BLOCKi_15_Q_reg_13_inst : DFF_X1 port map( D => n9030, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_237_port, QN => 
                           n_3325);
   DataPath_RF_BLOCKi_15_Q_reg_14_inst : DFF_X1 port map( D => n9029, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_238_port, QN => 
                           n_3326);
   DataPath_RF_BLOCKi_15_Q_reg_15_inst : DFF_X1 port map( D => n9028, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_239_port, QN => 
                           n_3327);
   DataPath_RF_BLOCKi_15_Q_reg_16_inst : DFF_X1 port map( D => n9027, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_240_port, QN => 
                           n_3328);
   DataPath_RF_BLOCKi_15_Q_reg_17_inst : DFF_X1 port map( D => n9026, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_241_port, QN => 
                           n_3329);
   DataPath_RF_BLOCKi_15_Q_reg_18_inst : DFF_X1 port map( D => n9025, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_242_port, QN => 
                           n_3330);
   DataPath_RF_BLOCKi_15_Q_reg_19_inst : DFF_X1 port map( D => n9024, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_243_port, QN => 
                           n_3331);
   DataPath_RF_BLOCKi_15_Q_reg_20_inst : DFF_X1 port map( D => n9023, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_244_port, QN => 
                           n_3332);
   DataPath_RF_BLOCKi_15_Q_reg_21_inst : DFF_X1 port map( D => n9022, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_245_port, QN => 
                           n_3333);
   DataPath_RF_BLOCKi_15_Q_reg_22_inst : DFF_X1 port map( D => n9021, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_246_port, QN => 
                           n_3334);
   DataPath_RF_BLOCKi_15_Q_reg_23_inst : DFF_X1 port map( D => n9020, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_247_port, QN => 
                           n_3335);
   DataPath_RF_BLOCKi_15_Q_reg_24_inst : DFF_X1 port map( D => n9019, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_248_port, QN => 
                           n_3336);
   DataPath_RF_BLOCKi_15_Q_reg_25_inst : DFF_X1 port map( D => n9018, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_249_port, QN => 
                           n_3337);
   DataPath_RF_BLOCKi_15_Q_reg_26_inst : DFF_X1 port map( D => n9017, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_250_port, QN => 
                           n_3338);
   DataPath_RF_BLOCKi_15_Q_reg_27_inst : DFF_X1 port map( D => n9016, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_251_port, QN => 
                           n_3339);
   DataPath_RF_BLOCKi_15_Q_reg_28_inst : DFF_X1 port map( D => n9015, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_252_port, QN => 
                           n_3340);
   DataPath_RF_BLOCKi_15_Q_reg_29_inst : DFF_X1 port map( D => n9014, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_253_port, QN => 
                           n_3341);
   DataPath_RF_BLOCKi_15_Q_reg_30_inst : DFF_X1 port map( D => n9013, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_254_port, QN => 
                           n_3342);
   DataPath_RF_BLOCKi_15_Q_reg_31_inst : DFF_X1 port map( D => n9012, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_255_port, QN => 
                           n_3343);
   DataPath_RF_BLOCKi_14_Q_reg_0_inst : DFF_X1 port map( D => n9011, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_192_port, QN => 
                           n_3344);
   DataPath_RF_BLOCKi_14_Q_reg_1_inst : DFF_X1 port map( D => n9010, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_193_port, QN => 
                           n_3345);
   DataPath_RF_BLOCKi_14_Q_reg_2_inst : DFF_X1 port map( D => n9009, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_194_port, QN => 
                           n_3346);
   DataPath_RF_BLOCKi_14_Q_reg_3_inst : DFF_X1 port map( D => n9008, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_195_port, QN => 
                           n_3347);
   DataPath_RF_BLOCKi_14_Q_reg_4_inst : DFF_X1 port map( D => n9007, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_196_port, QN => 
                           n_3348);
   DataPath_RF_BLOCKi_14_Q_reg_5_inst : DFF_X1 port map( D => n9006, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_197_port, QN => 
                           n_3349);
   DataPath_RF_BLOCKi_14_Q_reg_6_inst : DFF_X1 port map( D => n9005, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_198_port, QN => 
                           n_3350);
   DataPath_RF_BLOCKi_14_Q_reg_7_inst : DFF_X1 port map( D => n9004, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_199_port, QN => 
                           n_3351);
   DataPath_RF_BLOCKi_14_Q_reg_8_inst : DFF_X1 port map( D => n9003, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_200_port, QN => 
                           n_3352);
   DataPath_RF_BLOCKi_14_Q_reg_9_inst : DFF_X1 port map( D => n9002, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_201_port, QN => 
                           n_3353);
   DataPath_RF_BLOCKi_14_Q_reg_10_inst : DFF_X1 port map( D => n9001, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_202_port, QN => 
                           n_3354);
   DataPath_RF_BLOCKi_14_Q_reg_11_inst : DFF_X1 port map( D => n9000, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_203_port, QN => 
                           n_3355);
   DataPath_RF_BLOCKi_14_Q_reg_12_inst : DFF_X1 port map( D => n8999, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_204_port, QN => 
                           n_3356);
   DataPath_RF_BLOCKi_14_Q_reg_13_inst : DFF_X1 port map( D => n8998, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_205_port, QN => 
                           n_3357);
   DataPath_RF_BLOCKi_14_Q_reg_14_inst : DFF_X1 port map( D => n8997, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_206_port, QN => 
                           n_3358);
   DataPath_RF_BLOCKi_14_Q_reg_15_inst : DFF_X1 port map( D => n8996, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_207_port, QN => 
                           n_3359);
   DataPath_RF_BLOCKi_14_Q_reg_16_inst : DFF_X1 port map( D => n8995, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_208_port, QN => 
                           n_3360);
   DataPath_RF_BLOCKi_14_Q_reg_17_inst : DFF_X1 port map( D => n8994, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_209_port, QN => 
                           n_3361);
   DataPath_RF_BLOCKi_14_Q_reg_18_inst : DFF_X1 port map( D => n8993, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_210_port, QN => 
                           n_3362);
   DataPath_RF_BLOCKi_14_Q_reg_19_inst : DFF_X1 port map( D => n8992, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_211_port, QN => 
                           n_3363);
   DataPath_RF_BLOCKi_14_Q_reg_20_inst : DFF_X1 port map( D => n8991, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_212_port, QN => 
                           n_3364);
   DataPath_RF_BLOCKi_14_Q_reg_21_inst : DFF_X1 port map( D => n8990, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_213_port, QN => 
                           n_3365);
   DataPath_RF_BLOCKi_14_Q_reg_22_inst : DFF_X1 port map( D => n8989, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_214_port, QN => 
                           n_3366);
   DataPath_RF_BLOCKi_14_Q_reg_23_inst : DFF_X1 port map( D => n8988, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_215_port, QN => 
                           n_3367);
   DataPath_RF_BLOCKi_14_Q_reg_24_inst : DFF_X1 port map( D => n8987, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_216_port, QN => 
                           n_3368);
   DataPath_RF_BLOCKi_14_Q_reg_25_inst : DFF_X1 port map( D => n8986, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_217_port, QN => 
                           n_3369);
   DataPath_RF_BLOCKi_14_Q_reg_26_inst : DFF_X1 port map( D => n8985, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_218_port, QN => 
                           n_3370);
   DataPath_RF_BLOCKi_14_Q_reg_27_inst : DFF_X1 port map( D => n8984, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_219_port, QN => 
                           n_3371);
   DataPath_RF_BLOCKi_14_Q_reg_28_inst : DFF_X1 port map( D => n8983, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_220_port, QN => 
                           n_3372);
   DataPath_RF_BLOCKi_14_Q_reg_29_inst : DFF_X1 port map( D => n8982, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_221_port, QN => 
                           n_3373);
   DataPath_RF_BLOCKi_14_Q_reg_30_inst : DFF_X1 port map( D => n8981, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_222_port, QN => 
                           n_3374);
   DataPath_RF_BLOCKi_14_Q_reg_31_inst : DFF_X1 port map( D => n8980, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_223_port, QN => 
                           n_3375);
   DataPath_RF_BLOCKi_13_Q_reg_0_inst : DFF_X1 port map( D => n8979, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_160_port, QN => 
                           n_3376);
   DataPath_RF_BLOCKi_13_Q_reg_1_inst : DFF_X1 port map( D => n8978, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_161_port, QN => 
                           n_3377);
   DataPath_RF_BLOCKi_13_Q_reg_2_inst : DFF_X1 port map( D => n8977, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_162_port, QN => 
                           n_3378);
   DataPath_RF_BLOCKi_13_Q_reg_3_inst : DFF_X1 port map( D => n8976, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_163_port, QN => 
                           n_3379);
   DataPath_RF_BLOCKi_13_Q_reg_4_inst : DFF_X1 port map( D => n8975, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_164_port, QN => 
                           n_3380);
   DataPath_RF_BLOCKi_13_Q_reg_5_inst : DFF_X1 port map( D => n8974, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_165_port, QN => 
                           n_3381);
   DataPath_RF_BLOCKi_13_Q_reg_6_inst : DFF_X1 port map( D => n8973, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_166_port, QN => 
                           n_3382);
   DataPath_RF_BLOCKi_13_Q_reg_7_inst : DFF_X1 port map( D => n8972, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_167_port, QN => 
                           n_3383);
   DataPath_RF_BLOCKi_13_Q_reg_8_inst : DFF_X1 port map( D => n8971, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_168_port, QN => 
                           n_3384);
   DataPath_RF_BLOCKi_13_Q_reg_9_inst : DFF_X1 port map( D => n8970, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_169_port, QN => 
                           n_3385);
   DataPath_RF_BLOCKi_13_Q_reg_10_inst : DFF_X1 port map( D => n8969, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_170_port, QN => 
                           n_3386);
   DataPath_RF_BLOCKi_13_Q_reg_11_inst : DFF_X1 port map( D => n8968, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_171_port, QN => 
                           n_3387);
   DataPath_RF_BLOCKi_13_Q_reg_12_inst : DFF_X1 port map( D => n8967, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_172_port, QN => 
                           n_3388);
   DataPath_RF_BLOCKi_13_Q_reg_13_inst : DFF_X1 port map( D => n8966, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_173_port, QN => 
                           n_3389);
   DataPath_RF_BLOCKi_13_Q_reg_14_inst : DFF_X1 port map( D => n8965, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_174_port, QN => 
                           n_3390);
   DataPath_RF_BLOCKi_13_Q_reg_15_inst : DFF_X1 port map( D => n8964, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_175_port, QN => 
                           n_3391);
   DataPath_RF_BLOCKi_13_Q_reg_16_inst : DFF_X1 port map( D => n8963, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_176_port, QN => 
                           n_3392);
   DataPath_RF_BLOCKi_13_Q_reg_17_inst : DFF_X1 port map( D => n8962, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_177_port, QN => 
                           n_3393);
   DataPath_RF_BLOCKi_13_Q_reg_18_inst : DFF_X1 port map( D => n8961, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_178_port, QN => 
                           n_3394);
   DataPath_RF_BLOCKi_13_Q_reg_19_inst : DFF_X1 port map( D => n8960, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_179_port, QN => 
                           n_3395);
   DataPath_RF_BLOCKi_13_Q_reg_20_inst : DFF_X1 port map( D => n8959, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_180_port, QN => 
                           n_3396);
   DataPath_RF_BLOCKi_13_Q_reg_21_inst : DFF_X1 port map( D => n8958, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_181_port, QN => 
                           n_3397);
   DataPath_RF_BLOCKi_13_Q_reg_22_inst : DFF_X1 port map( D => n8957, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_182_port, QN => 
                           n_3398);
   DataPath_RF_BLOCKi_13_Q_reg_23_inst : DFF_X1 port map( D => n8956, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_183_port, QN => 
                           n_3399);
   DataPath_RF_BLOCKi_13_Q_reg_24_inst : DFF_X1 port map( D => n8955, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_184_port, QN => 
                           n_3400);
   DataPath_RF_BLOCKi_13_Q_reg_25_inst : DFF_X1 port map( D => n8954, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_185_port, QN => 
                           n_3401);
   DataPath_RF_BLOCKi_13_Q_reg_26_inst : DFF_X1 port map( D => n8953, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_186_port, QN => 
                           n_3402);
   DataPath_RF_BLOCKi_13_Q_reg_27_inst : DFF_X1 port map( D => n8952, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_187_port, QN => 
                           n_3403);
   DataPath_RF_BLOCKi_13_Q_reg_28_inst : DFF_X1 port map( D => n8951, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_188_port, QN => 
                           n_3404);
   DataPath_RF_BLOCKi_13_Q_reg_29_inst : DFF_X1 port map( D => n8950, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_189_port, QN => 
                           n_3405);
   DataPath_RF_BLOCKi_13_Q_reg_30_inst : DFF_X1 port map( D => n8949, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_190_port, QN => 
                           n_3406);
   DataPath_RF_BLOCKi_13_Q_reg_31_inst : DFF_X1 port map( D => n8948, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_191_port, QN => 
                           n_3407);
   DataPath_RF_BLOCKi_12_Q_reg_0_inst : DFF_X1 port map( D => n8947, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_128_port, QN => 
                           n_3408);
   DataPath_RF_BLOCKi_12_Q_reg_1_inst : DFF_X1 port map( D => n8946, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_129_port, QN => 
                           n_3409);
   DataPath_RF_BLOCKi_12_Q_reg_2_inst : DFF_X1 port map( D => n8945, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_130_port, QN => 
                           n_3410);
   DataPath_RF_BLOCKi_12_Q_reg_3_inst : DFF_X1 port map( D => n8944, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_131_port, QN => 
                           n_3411);
   DataPath_RF_BLOCKi_12_Q_reg_4_inst : DFF_X1 port map( D => n8943, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_132_port, QN => 
                           n_3412);
   DataPath_RF_BLOCKi_12_Q_reg_5_inst : DFF_X1 port map( D => n8942, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_133_port, QN => 
                           n_3413);
   DataPath_RF_BLOCKi_12_Q_reg_6_inst : DFF_X1 port map( D => n8941, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_134_port, QN => 
                           n_3414);
   DataPath_RF_BLOCKi_12_Q_reg_7_inst : DFF_X1 port map( D => n8940, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_135_port, QN => 
                           n_3415);
   DataPath_RF_BLOCKi_12_Q_reg_8_inst : DFF_X1 port map( D => n8939, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_136_port, QN => 
                           n_3416);
   DataPath_RF_BLOCKi_12_Q_reg_9_inst : DFF_X1 port map( D => n8938, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_137_port, QN => 
                           n_3417);
   DataPath_RF_BLOCKi_12_Q_reg_10_inst : DFF_X1 port map( D => n8937, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_138_port, QN => 
                           n_3418);
   DataPath_RF_BLOCKi_12_Q_reg_11_inst : DFF_X1 port map( D => n8936, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_139_port, QN => 
                           n_3419);
   DataPath_RF_BLOCKi_12_Q_reg_12_inst : DFF_X1 port map( D => n8935, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_140_port, QN => 
                           n_3420);
   DataPath_RF_BLOCKi_12_Q_reg_13_inst : DFF_X1 port map( D => n8934, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_141_port, QN => 
                           n_3421);
   DataPath_RF_BLOCKi_12_Q_reg_14_inst : DFF_X1 port map( D => n8933, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_142_port, QN => 
                           n_3422);
   DataPath_RF_BLOCKi_12_Q_reg_15_inst : DFF_X1 port map( D => n8932, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_143_port, QN => 
                           n_3423);
   DataPath_RF_BLOCKi_12_Q_reg_16_inst : DFF_X1 port map( D => n8931, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_144_port, QN => 
                           n_3424);
   DataPath_RF_BLOCKi_12_Q_reg_17_inst : DFF_X1 port map( D => n8930, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_145_port, QN => 
                           n_3425);
   DataPath_RF_BLOCKi_12_Q_reg_18_inst : DFF_X1 port map( D => n8929, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_146_port, QN => 
                           n_3426);
   DataPath_RF_BLOCKi_12_Q_reg_19_inst : DFF_X1 port map( D => n8928, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_147_port, QN => 
                           n_3427);
   DataPath_RF_BLOCKi_12_Q_reg_20_inst : DFF_X1 port map( D => n8927, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_148_port, QN => 
                           n_3428);
   DataPath_RF_BLOCKi_12_Q_reg_21_inst : DFF_X1 port map( D => n8926, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_149_port, QN => 
                           n_3429);
   DataPath_RF_BLOCKi_12_Q_reg_22_inst : DFF_X1 port map( D => n8925, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_150_port, QN => 
                           n_3430);
   DataPath_RF_BLOCKi_12_Q_reg_23_inst : DFF_X1 port map( D => n8924, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_151_port, QN => 
                           n_3431);
   DataPath_RF_BLOCKi_12_Q_reg_24_inst : DFF_X1 port map( D => n8923, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_152_port, QN => 
                           n_3432);
   DataPath_RF_BLOCKi_12_Q_reg_25_inst : DFF_X1 port map( D => n8922, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_153_port, QN => 
                           n_3433);
   DataPath_RF_BLOCKi_12_Q_reg_26_inst : DFF_X1 port map( D => n8921, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_154_port, QN => 
                           n_3434);
   DataPath_RF_BLOCKi_12_Q_reg_27_inst : DFF_X1 port map( D => n8920, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_155_port, QN => 
                           n_3435);
   DataPath_RF_BLOCKi_12_Q_reg_28_inst : DFF_X1 port map( D => n8919, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_156_port, QN => 
                           n_3436);
   DataPath_RF_BLOCKi_12_Q_reg_29_inst : DFF_X1 port map( D => n8918, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_157_port, QN => 
                           n_3437);
   DataPath_RF_BLOCKi_12_Q_reg_30_inst : DFF_X1 port map( D => n8917, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_158_port, QN => 
                           n_3438);
   DataPath_RF_BLOCKi_12_Q_reg_31_inst : DFF_X1 port map( D => n8916, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_159_port, QN => 
                           n_3439);
   DataPath_RF_BLOCKi_11_Q_reg_0_inst : DFF_X1 port map( D => n8915, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_96_port, QN => 
                           n_3440);
   DataPath_RF_BLOCKi_11_Q_reg_1_inst : DFF_X1 port map( D => n8914, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_97_port, QN => 
                           n_3441);
   DataPath_RF_BLOCKi_11_Q_reg_2_inst : DFF_X1 port map( D => n8913, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_98_port, QN => 
                           n_3442);
   DataPath_RF_BLOCKi_11_Q_reg_3_inst : DFF_X1 port map( D => n8912, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_99_port, QN => 
                           n_3443);
   DataPath_RF_BLOCKi_11_Q_reg_4_inst : DFF_X1 port map( D => n8911, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_100_port, QN => 
                           n_3444);
   DataPath_RF_BLOCKi_11_Q_reg_5_inst : DFF_X1 port map( D => n8910, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_101_port, QN => 
                           n_3445);
   DataPath_RF_BLOCKi_11_Q_reg_6_inst : DFF_X1 port map( D => n8909, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_102_port, QN => 
                           n_3446);
   DataPath_RF_BLOCKi_11_Q_reg_7_inst : DFF_X1 port map( D => n8908, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_103_port, QN => 
                           n_3447);
   DataPath_RF_BLOCKi_11_Q_reg_8_inst : DFF_X1 port map( D => n8907, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_104_port, QN => 
                           n_3448);
   DataPath_RF_BLOCKi_11_Q_reg_9_inst : DFF_X1 port map( D => n8906, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_105_port, QN => 
                           n_3449);
   DataPath_RF_BLOCKi_11_Q_reg_10_inst : DFF_X1 port map( D => n8905, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_106_port, QN => 
                           n_3450);
   DataPath_RF_BLOCKi_11_Q_reg_11_inst : DFF_X1 port map( D => n8904, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_107_port, QN => 
                           n_3451);
   DataPath_RF_BLOCKi_11_Q_reg_12_inst : DFF_X1 port map( D => n8903, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_108_port, QN => 
                           n_3452);
   DataPath_RF_BLOCKi_11_Q_reg_13_inst : DFF_X1 port map( D => n8902, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_109_port, QN => 
                           n_3453);
   DataPath_RF_BLOCKi_11_Q_reg_14_inst : DFF_X1 port map( D => n8901, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_110_port, QN => 
                           n_3454);
   DataPath_RF_BLOCKi_11_Q_reg_15_inst : DFF_X1 port map( D => n8900, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_111_port, QN => 
                           n_3455);
   DataPath_RF_BLOCKi_11_Q_reg_16_inst : DFF_X1 port map( D => n8899, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_112_port, QN => 
                           n_3456);
   DataPath_RF_BLOCKi_11_Q_reg_17_inst : DFF_X1 port map( D => n8898, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_113_port, QN => 
                           n_3457);
   DataPath_RF_BLOCKi_11_Q_reg_18_inst : DFF_X1 port map( D => n8897, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_114_port, QN => 
                           n_3458);
   DataPath_RF_BLOCKi_11_Q_reg_19_inst : DFF_X1 port map( D => n8896, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_115_port, QN => 
                           n_3459);
   DataPath_RF_BLOCKi_11_Q_reg_20_inst : DFF_X1 port map( D => n8895, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_116_port, QN => 
                           n_3460);
   DataPath_RF_BLOCKi_11_Q_reg_21_inst : DFF_X1 port map( D => n8894, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_117_port, QN => 
                           n_3461);
   DataPath_RF_BLOCKi_11_Q_reg_22_inst : DFF_X1 port map( D => n8893, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_118_port, QN => 
                           n_3462);
   DataPath_RF_BLOCKi_11_Q_reg_23_inst : DFF_X1 port map( D => n8892, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_119_port, QN => 
                           n_3463);
   DataPath_RF_BLOCKi_11_Q_reg_24_inst : DFF_X1 port map( D => n8891, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_120_port, QN => 
                           n_3464);
   DataPath_RF_BLOCKi_11_Q_reg_25_inst : DFF_X1 port map( D => n8890, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_121_port, QN => 
                           n_3465);
   DataPath_RF_BLOCKi_11_Q_reg_26_inst : DFF_X1 port map( D => n8889, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_122_port, QN => 
                           n_3466);
   DataPath_RF_BLOCKi_11_Q_reg_27_inst : DFF_X1 port map( D => n8888, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_123_port, QN => 
                           n_3467);
   DataPath_RF_BLOCKi_11_Q_reg_28_inst : DFF_X1 port map( D => n8887, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_124_port, QN => 
                           n_3468);
   DataPath_RF_BLOCKi_11_Q_reg_29_inst : DFF_X1 port map( D => n8886, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_125_port, QN => 
                           n_3469);
   DataPath_RF_BLOCKi_11_Q_reg_30_inst : DFF_X1 port map( D => n8885, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_126_port, QN => 
                           n_3470);
   DataPath_RF_BLOCKi_11_Q_reg_31_inst : DFF_X1 port map( D => n8884, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_127_port, QN => 
                           n_3471);
   DataPath_RF_BLOCKi_10_Q_reg_0_inst : DFF_X1 port map( D => n8883, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_64_port, QN => 
                           n_3472);
   DataPath_RF_BLOCKi_10_Q_reg_1_inst : DFF_X1 port map( D => n8882, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_65_port, QN => 
                           n_3473);
   DataPath_RF_BLOCKi_10_Q_reg_2_inst : DFF_X1 port map( D => n8881, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_66_port, QN => 
                           n_3474);
   DataPath_RF_BLOCKi_10_Q_reg_3_inst : DFF_X1 port map( D => n8880, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_67_port, QN => 
                           n_3475);
   DataPath_RF_BLOCKi_10_Q_reg_4_inst : DFF_X1 port map( D => n8879, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_68_port, QN => 
                           n_3476);
   DataPath_RF_BLOCKi_10_Q_reg_5_inst : DFF_X1 port map( D => n8878, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_69_port, QN => 
                           n_3477);
   DataPath_RF_BLOCKi_10_Q_reg_6_inst : DFF_X1 port map( D => n8877, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_70_port, QN => 
                           n_3478);
   DataPath_RF_BLOCKi_10_Q_reg_7_inst : DFF_X1 port map( D => n8876, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_71_port, QN => 
                           n_3479);
   DataPath_RF_BLOCKi_10_Q_reg_8_inst : DFF_X1 port map( D => n8875, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_72_port, QN => 
                           n_3480);
   DataPath_RF_BLOCKi_10_Q_reg_9_inst : DFF_X1 port map( D => n8874, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_73_port, QN => 
                           n_3481);
   DataPath_RF_BLOCKi_10_Q_reg_10_inst : DFF_X1 port map( D => n8873, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_74_port, QN => 
                           n_3482);
   DataPath_RF_BLOCKi_10_Q_reg_11_inst : DFF_X1 port map( D => n8872, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_75_port, QN => 
                           n_3483);
   DataPath_RF_BLOCKi_10_Q_reg_12_inst : DFF_X1 port map( D => n8871, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_76_port, QN => 
                           n_3484);
   DataPath_RF_BLOCKi_10_Q_reg_13_inst : DFF_X1 port map( D => n8870, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_77_port, QN => 
                           n_3485);
   DataPath_RF_BLOCKi_10_Q_reg_14_inst : DFF_X1 port map( D => n8869, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_78_port, QN => 
                           n_3486);
   DataPath_RF_BLOCKi_10_Q_reg_15_inst : DFF_X1 port map( D => n8868, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_79_port, QN => 
                           n_3487);
   DataPath_RF_BLOCKi_10_Q_reg_16_inst : DFF_X1 port map( D => n8867, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_80_port, QN => 
                           n_3488);
   DataPath_RF_BLOCKi_10_Q_reg_17_inst : DFF_X1 port map( D => n8866, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_81_port, QN => 
                           n_3489);
   DataPath_RF_BLOCKi_10_Q_reg_18_inst : DFF_X1 port map( D => n8865, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_82_port, QN => 
                           n_3490);
   DataPath_RF_BLOCKi_10_Q_reg_19_inst : DFF_X1 port map( D => n8864, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_83_port, QN => 
                           n_3491);
   DataPath_RF_BLOCKi_10_Q_reg_20_inst : DFF_X1 port map( D => n8863, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_84_port, QN => 
                           n_3492);
   DataPath_RF_BLOCKi_10_Q_reg_21_inst : DFF_X1 port map( D => n8862, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_85_port, QN => 
                           n_3493);
   DataPath_RF_BLOCKi_10_Q_reg_22_inst : DFF_X1 port map( D => n8861, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_86_port, QN => 
                           n_3494);
   DataPath_RF_BLOCKi_10_Q_reg_23_inst : DFF_X1 port map( D => n8860, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_87_port, QN => 
                           n_3495);
   DataPath_RF_BLOCKi_10_Q_reg_24_inst : DFF_X1 port map( D => n8859, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_88_port, QN => 
                           n_3496);
   DataPath_RF_BLOCKi_10_Q_reg_25_inst : DFF_X1 port map( D => n8858, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_89_port, QN => 
                           n_3497);
   DataPath_RF_BLOCKi_10_Q_reg_26_inst : DFF_X1 port map( D => n8857, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_90_port, QN => 
                           n_3498);
   DataPath_RF_BLOCKi_10_Q_reg_27_inst : DFF_X1 port map( D => n8856, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_91_port, QN => 
                           n_3499);
   DataPath_RF_BLOCKi_10_Q_reg_28_inst : DFF_X1 port map( D => n8855, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_92_port, QN => 
                           n_3500);
   DataPath_RF_BLOCKi_10_Q_reg_29_inst : DFF_X1 port map( D => n8854, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_93_port, QN => 
                           n_3501);
   DataPath_RF_BLOCKi_10_Q_reg_30_inst : DFF_X1 port map( D => n8853, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_94_port, QN => 
                           n_3502);
   DataPath_RF_BLOCKi_10_Q_reg_31_inst : DFF_X1 port map( D => n8852, CK => CLK
                           , Q => DataPath_RF_bus_reg_dataout_95_port, QN => 
                           n_3503);
   DataPath_RF_BLOCKi_9_Q_reg_0_inst : DFF_X1 port map( D => n8851, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_32_port, QN => 
                           n_3504);
   DataPath_RF_BLOCKi_9_Q_reg_1_inst : DFF_X1 port map( D => n8850, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_33_port, QN => 
                           n_3505);
   DataPath_RF_BLOCKi_9_Q_reg_2_inst : DFF_X1 port map( D => n8849, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_34_port, QN => 
                           n_3506);
   DataPath_RF_BLOCKi_9_Q_reg_3_inst : DFF_X1 port map( D => n8848, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_35_port, QN => 
                           n_3507);
   DataPath_RF_BLOCKi_9_Q_reg_4_inst : DFF_X1 port map( D => n8847, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_36_port, QN => 
                           n_3508);
   DataPath_RF_BLOCKi_9_Q_reg_5_inst : DFF_X1 port map( D => n8846, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_37_port, QN => 
                           n_3509);
   DataPath_RF_BLOCKi_9_Q_reg_6_inst : DFF_X1 port map( D => n8845, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_38_port, QN => 
                           n_3510);
   DataPath_RF_BLOCKi_9_Q_reg_7_inst : DFF_X1 port map( D => n8844, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_39_port, QN => 
                           n_3511);
   DataPath_RF_BLOCKi_9_Q_reg_8_inst : DFF_X1 port map( D => n8843, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_40_port, QN => 
                           n_3512);
   DataPath_RF_BLOCKi_9_Q_reg_9_inst : DFF_X1 port map( D => n8842, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_41_port, QN => 
                           n_3513);
   DataPath_RF_BLOCKi_9_Q_reg_10_inst : DFF_X1 port map( D => n8841, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_42_port, QN => 
                           n_3514);
   DataPath_RF_BLOCKi_9_Q_reg_11_inst : DFF_X1 port map( D => n8840, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_43_port, QN => 
                           n_3515);
   DataPath_RF_BLOCKi_9_Q_reg_12_inst : DFF_X1 port map( D => n8839, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_44_port, QN => 
                           n_3516);
   DataPath_RF_BLOCKi_9_Q_reg_13_inst : DFF_X1 port map( D => n8838, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_45_port, QN => 
                           n_3517);
   DataPath_RF_BLOCKi_9_Q_reg_14_inst : DFF_X1 port map( D => n8837, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_46_port, QN => 
                           n_3518);
   DataPath_RF_BLOCKi_9_Q_reg_15_inst : DFF_X1 port map( D => n8836, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_47_port, QN => 
                           n_3519);
   DataPath_RF_BLOCKi_9_Q_reg_16_inst : DFF_X1 port map( D => n8835, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_48_port, QN => 
                           n_3520);
   DataPath_RF_BLOCKi_9_Q_reg_17_inst : DFF_X1 port map( D => n8834, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_49_port, QN => 
                           n_3521);
   DataPath_RF_BLOCKi_9_Q_reg_18_inst : DFF_X1 port map( D => n8833, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_50_port, QN => 
                           n_3522);
   DataPath_RF_BLOCKi_9_Q_reg_19_inst : DFF_X1 port map( D => n8832, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_51_port, QN => 
                           n_3523);
   DataPath_RF_BLOCKi_9_Q_reg_20_inst : DFF_X1 port map( D => n8831, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_52_port, QN => 
                           n_3524);
   DataPath_RF_BLOCKi_9_Q_reg_21_inst : DFF_X1 port map( D => n8830, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_53_port, QN => 
                           n_3525);
   DataPath_RF_BLOCKi_9_Q_reg_22_inst : DFF_X1 port map( D => n8829, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_54_port, QN => 
                           n_3526);
   DataPath_RF_BLOCKi_9_Q_reg_23_inst : DFF_X1 port map( D => n8828, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_55_port, QN => 
                           n_3527);
   DataPath_RF_BLOCKi_9_Q_reg_24_inst : DFF_X1 port map( D => n8827, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_56_port, QN => 
                           n_3528);
   DataPath_RF_BLOCKi_9_Q_reg_25_inst : DFF_X1 port map( D => n8826, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_57_port, QN => 
                           n_3529);
   DataPath_RF_BLOCKi_9_Q_reg_26_inst : DFF_X1 port map( D => n8825, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_58_port, QN => 
                           n_3530);
   DataPath_RF_BLOCKi_9_Q_reg_27_inst : DFF_X1 port map( D => n8824, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_59_port, QN => 
                           n_3531);
   DataPath_RF_BLOCKi_9_Q_reg_28_inst : DFF_X1 port map( D => n8823, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_60_port, QN => 
                           n_3532);
   DataPath_RF_BLOCKi_9_Q_reg_29_inst : DFF_X1 port map( D => n8822, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_61_port, QN => 
                           n_3533);
   DataPath_RF_BLOCKi_9_Q_reg_30_inst : DFF_X1 port map( D => n8821, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_62_port, QN => 
                           n_3534);
   DataPath_RF_BLOCKi_9_Q_reg_31_inst : DFF_X1 port map( D => n8820, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_63_port, QN => 
                           n_3535);
   DataPath_RF_BLOCKi_8_Q_reg_0_inst : DFF_X1 port map( D => n8819, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_0_port, QN => 
                           n_3536);
   DataPath_RF_BLOCKi_8_Q_reg_1_inst : DFF_X1 port map( D => n8818, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_1_port, QN => 
                           n_3537);
   DataPath_RF_BLOCKi_8_Q_reg_2_inst : DFF_X1 port map( D => n8817, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_2_port, QN => 
                           n_3538);
   DataPath_RF_BLOCKi_8_Q_reg_3_inst : DFF_X1 port map( D => n8816, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_3_port, QN => 
                           n_3539);
   DataPath_RF_BLOCKi_8_Q_reg_4_inst : DFF_X1 port map( D => n8815, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_4_port, QN => 
                           n_3540);
   DataPath_RF_BLOCKi_8_Q_reg_5_inst : DFF_X1 port map( D => n8814, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_5_port, QN => 
                           n_3541);
   DataPath_RF_BLOCKi_8_Q_reg_6_inst : DFF_X1 port map( D => n8813, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_6_port, QN => 
                           n_3542);
   DataPath_RF_BLOCKi_8_Q_reg_7_inst : DFF_X1 port map( D => n8812, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_7_port, QN => 
                           n_3543);
   DataPath_RF_BLOCKi_8_Q_reg_8_inst : DFF_X1 port map( D => n8811, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_8_port, QN => 
                           n_3544);
   DataPath_RF_BLOCKi_8_Q_reg_9_inst : DFF_X1 port map( D => n8810, CK => CLK, 
                           Q => DataPath_RF_bus_reg_dataout_9_port, QN => 
                           n_3545);
   DataPath_RF_BLOCKi_8_Q_reg_10_inst : DFF_X1 port map( D => n8809, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_10_port, QN => 
                           n_3546);
   DataPath_RF_BLOCKi_8_Q_reg_11_inst : DFF_X1 port map( D => n8808, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_11_port, QN => 
                           n_3547);
   DataPath_RF_BLOCKi_8_Q_reg_12_inst : DFF_X1 port map( D => n8807, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_12_port, QN => 
                           n_3548);
   DataPath_RF_BLOCKi_8_Q_reg_13_inst : DFF_X1 port map( D => n8806, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_13_port, QN => 
                           n_3549);
   DataPath_RF_BLOCKi_8_Q_reg_14_inst : DFF_X1 port map( D => n8805, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_14_port, QN => 
                           n_3550);
   DataPath_RF_BLOCKi_8_Q_reg_15_inst : DFF_X1 port map( D => n8804, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_15_port, QN => 
                           n_3551);
   DataPath_RF_BLOCKi_8_Q_reg_16_inst : DFF_X1 port map( D => n8803, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_16_port, QN => 
                           n_3552);
   DataPath_RF_BLOCKi_8_Q_reg_17_inst : DFF_X1 port map( D => n8802, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_17_port, QN => 
                           n_3553);
   DataPath_RF_BLOCKi_8_Q_reg_18_inst : DFF_X1 port map( D => n8801, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_18_port, QN => 
                           n_3554);
   DataPath_RF_BLOCKi_8_Q_reg_19_inst : DFF_X1 port map( D => n8800, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_19_port, QN => 
                           n_3555);
   DataPath_RF_BLOCKi_8_Q_reg_20_inst : DFF_X1 port map( D => n8799, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_20_port, QN => 
                           n_3556);
   DataPath_RF_BLOCKi_8_Q_reg_21_inst : DFF_X1 port map( D => n8798, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_21_port, QN => 
                           n_3557);
   DataPath_RF_BLOCKi_8_Q_reg_22_inst : DFF_X1 port map( D => n8797, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_22_port, QN => 
                           n_3558);
   DataPath_RF_BLOCKi_8_Q_reg_23_inst : DFF_X1 port map( D => n8796, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_23_port, QN => 
                           n_3559);
   DataPath_RF_BLOCKi_8_Q_reg_24_inst : DFF_X1 port map( D => n8795, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_24_port, QN => 
                           n_3560);
   DataPath_RF_BLOCKi_8_Q_reg_25_inst : DFF_X1 port map( D => n8794, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_25_port, QN => 
                           n_3561);
   DataPath_RF_BLOCKi_8_Q_reg_26_inst : DFF_X1 port map( D => n8793, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_26_port, QN => 
                           n_3562);
   DataPath_RF_BLOCKi_8_Q_reg_27_inst : DFF_X1 port map( D => n8792, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_27_port, QN => 
                           n_3563);
   DataPath_RF_BLOCKi_8_Q_reg_28_inst : DFF_X1 port map( D => n8791, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_28_port, QN => 
                           n_3564);
   DataPath_RF_BLOCKi_8_Q_reg_29_inst : DFF_X1 port map( D => n8790, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_29_port, QN => 
                           n_3565);
   DataPath_RF_BLOCKi_8_Q_reg_30_inst : DFF_X1 port map( D => n8789, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_30_port, QN => 
                           n_3566);
   DataPath_RF_BLOCKi_8_Q_reg_31_inst : DFF_X1 port map( D => n8788, CK => CLK,
                           Q => DataPath_RF_bus_reg_dataout_31_port, QN => 
                           n_3567);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_0_inst : DFF_X1 port map( D => n8755, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_0_port, QN => 
                           n_3568);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_1_inst : DFF_X1 port map( D => n8754, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_1_port, QN => 
                           n_3569);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_2_inst : DFF_X1 port map( D => n8753, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_2_port, QN => 
                           n_3570);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_3_inst : DFF_X1 port map( D => n8752, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_3_port, QN => 
                           n_3571);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_4_inst : DFF_X1 port map( D => n8751, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_4_port, QN => 
                           n_3572);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_5_inst : DFF_X1 port map( D => n8750, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_5_port, QN => 
                           n_3573);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_6_inst : DFF_X1 port map( D => n8749, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_6_port, QN => 
                           n_3574);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_7_inst : DFF_X1 port map( D => n8748, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_7_port, QN => 
                           n_3575);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_8_inst : DFF_X1 port map( D => n8747, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_8_port, QN => 
                           n_3576);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_9_inst : DFF_X1 port map( D => n8746, CK =>
                           CLK, Q => DataPath_i_REG_LDSTR_OUT_9_port, QN => 
                           n_3577);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_10_inst : DFF_X1 port map( D => n8745, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_10_port, QN =>
                           n_3578);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_11_inst : DFF_X1 port map( D => n8744, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_11_port, QN =>
                           n_3579);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_12_inst : DFF_X1 port map( D => n8743, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_12_port, QN =>
                           n_3580);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_13_inst : DFF_X1 port map( D => n8742, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_13_port, QN =>
                           n_3581);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_14_inst : DFF_X1 port map( D => n8741, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_14_port, QN =>
                           n_3582);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_15_inst : DFF_X1 port map( D => n8740, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_15_port, QN =>
                           n_3583);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_16_inst : DFF_X1 port map( D => n8739, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_16_port, QN =>
                           n_3584);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_17_inst : DFF_X1 port map( D => n8738, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_17_port, QN =>
                           n_3585);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_18_inst : DFF_X1 port map( D => n8737, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_18_port, QN =>
                           n_3586);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_19_inst : DFF_X1 port map( D => n8736, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_19_port, QN =>
                           n_3587);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_20_inst : DFF_X1 port map( D => n8735, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_20_port, QN =>
                           n_3588);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_21_inst : DFF_X1 port map( D => n8734, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_21_port, QN =>
                           n_3589);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_22_inst : DFF_X1 port map( D => n8733, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_22_port, QN =>
                           n_3590);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_23_inst : DFF_X1 port map( D => n8732, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_23_port, QN =>
                           n_3591);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_24_inst : DFF_X1 port map( D => n8731, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_24_port, QN =>
                           n_3592);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_25_inst : DFF_X1 port map( D => n8730, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_25_port, QN =>
                           n_3593);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_26_inst : DFF_X1 port map( D => n8729, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_26_port, QN =>
                           n_3594);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_27_inst : DFF_X1 port map( D => n8728, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_27_port, QN =>
                           n_3595);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_28_inst : DFF_X1 port map( D => n8727, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_28_port, QN =>
                           n_3596);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_29_inst : DFF_X1 port map( D => n8726, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_29_port, QN =>
                           n_3597);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_30_inst : DFF_X1 port map( D => n8725, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_30_port, QN =>
                           n_3598);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_31_inst : DFF_X1 port map( D => n8724, CK 
                           => CLK, Q => DataPath_i_REG_LDSTR_OUT_31_port, QN =>
                           n_3599);
   DataPath_REG_ALU_OUT_Q_reg_0_inst : DFF_X1 port map( D => n8691, CK => CLK, 
                           Q => DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_0_port, 
                           QN => n_3600);
   DataPath_REG_ALU_OUT_Q_reg_1_inst : DFF_X1 port map( D => n8690, CK => CLK, 
                           Q => DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_1_port, 
                           QN => n408);
   DataPath_REG_ALU_OUT_Q_reg_2_inst : DFF_X1 port map( D => n8689, CK => CLK, 
                           Q => DRAM_ADDRESS_2_port, QN => n_3601);
   DataPath_REG_ALU_OUT_Q_reg_3_inst : DFF_X1 port map( D => n8688, CK => CLK, 
                           Q => DRAM_ADDRESS_3_port, QN => n_3602);
   DataPath_REG_ALU_OUT_Q_reg_4_inst : DFF_X1 port map( D => n8687, CK => CLK, 
                           Q => DRAM_ADDRESS_4_port, QN => n_3603);
   DataPath_REG_ALU_OUT_Q_reg_5_inst : DFF_X1 port map( D => n8686, CK => CLK, 
                           Q => DRAM_ADDRESS_5_port, QN => n_3604);
   DataPath_REG_ALU_OUT_Q_reg_6_inst : DFF_X1 port map( D => n8685, CK => CLK, 
                           Q => DRAM_ADDRESS_6_port, QN => n_3605);
   DataPath_REG_ALU_OUT_Q_reg_7_inst : DFF_X1 port map( D => n8684, CK => CLK, 
                           Q => DRAM_ADDRESS_7_port, QN => n_3606);
   DataPath_REG_ALU_OUT_Q_reg_8_inst : DFF_X1 port map( D => n8683, CK => CLK, 
                           Q => DRAM_ADDRESS_8_port, QN => n_3607);
   DataPath_REG_ALU_OUT_Q_reg_9_inst : DFF_X1 port map( D => n8682, CK => CLK, 
                           Q => DRAM_ADDRESS_9_port, QN => n_3608);
   DataPath_REG_ALU_OUT_Q_reg_10_inst : DFF_X1 port map( D => n8681, CK => CLK,
                           Q => DRAM_ADDRESS_10_port, QN => n_3609);
   DataPath_REG_ALU_OUT_Q_reg_11_inst : DFF_X1 port map( D => n8680, CK => CLK,
                           Q => DRAM_ADDRESS_11_port, QN => n_3610);
   DataPath_REG_ALU_OUT_Q_reg_12_inst : DFF_X1 port map( D => n8679, CK => CLK,
                           Q => DRAM_ADDRESS_12_port, QN => n_3611);
   DataPath_REG_ALU_OUT_Q_reg_13_inst : DFF_X1 port map( D => n8678, CK => CLK,
                           Q => DRAM_ADDRESS_13_port, QN => n_3612);
   DataPath_REG_ALU_OUT_Q_reg_14_inst : DFF_X1 port map( D => n8677, CK => CLK,
                           Q => DRAM_ADDRESS_14_port, QN => n_3613);
   DataPath_REG_ALU_OUT_Q_reg_15_inst : DFF_X1 port map( D => n8676, CK => CLK,
                           Q => DRAM_ADDRESS_15_port, QN => n_3614);
   DataPath_REG_ALU_OUT_Q_reg_16_inst : DFF_X1 port map( D => n8675, CK => CLK,
                           Q => DRAM_ADDRESS_16_port, QN => n_3615);
   DataPath_REG_ALU_OUT_Q_reg_17_inst : DFF_X1 port map( D => n8674, CK => CLK,
                           Q => DRAM_ADDRESS_17_port, QN => n424);
   DataPath_REG_ALU_OUT_Q_reg_31_inst : DFF_X1 port map( D => n8660, CK => CLK,
                           Q => DRAM_ADDRESS_31_port, QN => n7497);
   DataPath_REG_IN2_Q_reg_0_inst : DFF_X1 port map( D => n2028, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_0_port, QN => n1745);
   DataPath_REG_IN2_Q_reg_1_inst : DFF_X1 port map( D => n2027, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_1_port, QN => n2139);
   DataPath_REG_IN2_Q_reg_3_inst : DFF_X1 port map( D => n2116, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_3_port, QN => n_3616);
   DataPath_REG_IN2_Q_reg_4_inst : DFF_X1 port map( D => n2115, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_4_port, QN => n324);
   DataPath_REG_IN2_Q_reg_5_inst : DFF_X1 port map( D => n2114, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_5_port, QN => n_3617);
   DataPath_REG_IN2_Q_reg_6_inst : DFF_X1 port map( D => n2113, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_6_port, QN => n323);
   DataPath_REG_IN2_Q_reg_7_inst : DFF_X1 port map( D => n2014, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_7_port, QN => n254);
   DataPath_REG_IN2_Q_reg_8_inst : DFF_X1 port map( D => n2013, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_8_port, QN => n327);
   DataPath_REG_IN2_Q_reg_9_inst : DFF_X1 port map( D => n2012, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_9_port, QN => n261);
   DataPath_REG_IN2_Q_reg_10_inst : DFF_X1 port map( D => n2011, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_10_port, QN => n325);
   DataPath_REG_IN2_Q_reg_11_inst : DFF_X1 port map( D => n2010, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_11_port, QN => n281);
   DataPath_REG_IN2_Q_reg_12_inst : DFF_X1 port map( D => n2009, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_12_port, QN => n352);
   DataPath_REG_IN2_Q_reg_13_inst : DFF_X1 port map( D => n2008, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_13_port, QN => n255);
   DataPath_REG_IN2_Q_reg_14_inst : DFF_X1 port map( D => n2007, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_14_port, QN => n351);
   DataPath_REG_IN2_Q_reg_15_inst : DFF_X1 port map( D => n2006, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_15_port, QN => n353);
   DataPath_REG_IN2_Q_reg_16_inst : DFF_X1 port map( D => n2005, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_16_port, QN => n358);
   DataPath_REG_IN2_Q_reg_17_inst : DFF_X1 port map( D => n2004, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_17_port, QN => n350);
   DataPath_REG_IN2_Q_reg_19_inst : DFF_X1 port map( D => n2002, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_19_port, QN => n357);
   DataPath_REG_IN1_Q_reg_1_inst : DFF_X1 port map( D => n2091, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_1_port, QN => n542);
   DataPath_REG_IN1_Q_reg_3_inst : DFF_X1 port map( D => n2089, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_3_port, QN => n318);
   DataPath_REG_IN1_Q_reg_4_inst : DFF_X1 port map( D => n2055, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_4_port, QN => n1543);
   DataPath_REG_IN1_Q_reg_6_inst : DFF_X1 port map( D => n2053, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_6_port, QN => n810);
   DataPath_REG_IN1_Q_reg_7_inst : DFF_X1 port map( D => n2052, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_7_port, QN => n265);
   DataPath_REG_IN1_Q_reg_9_inst : DFF_X1 port map( D => n2050, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_9_port, QN => n_3618);
   DataPath_REG_IN1_Q_reg_10_inst : DFF_X1 port map( D => n2049, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_10_port, QN => n326);
   DataPath_REG_IN1_Q_reg_11_inst : DFF_X1 port map( D => n2048, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_11_port, QN => n_3619);
   DataPath_REG_IN1_Q_reg_12_inst : DFF_X1 port map( D => n2047, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_12_port, QN => n_3620);
   DataPath_REG_IN1_Q_reg_13_inst : DFF_X1 port map( D => n2046, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_13_port, QN => n_3621);
   DataPath_REG_IN1_Q_reg_14_inst : DFF_X1 port map( D => n2045, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_14_port, QN => n329);
   DataPath_REG_IN1_Q_reg_15_inst : DFF_X1 port map( D => n2026, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_15_port, QN => n330);
   DataPath_REG_IN1_Q_reg_16_inst : DFF_X1 port map( D => n2025, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_16_port, QN => n333);
   DataPath_REG_IN1_Q_reg_17_inst : DFF_X1 port map( D => n2024, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_17_port, QN => n334);
   DataPath_REG_IN1_Q_reg_18_inst : DFF_X1 port map( D => n2023, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_18_port, QN => n332);
   DataPath_REG_IN1_Q_reg_19_inst : DFF_X1 port map( D => n2022, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_19_port, QN => n331);
   DataPath_REG_IN1_Q_reg_20_inst : DFF_X1 port map( D => n2021, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_20_port, QN => n336);
   DataPath_REG_IN1_Q_reg_21_inst : DFF_X1 port map( D => n2020, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_21_port, QN => n337);
   DataPath_REG_IN1_Q_reg_22_inst : DFF_X1 port map( D => n2019, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_22_port, QN => n335);
   DataPath_REG_IN1_Q_reg_23_inst : DFF_X1 port map( D => n2018, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_23_port, QN => n359);
   DataPath_REG_IN1_Q_reg_24_inst : DFF_X1 port map( D => n2017, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_24_port, QN => n355);
   DataPath_REG_IN1_Q_reg_25_inst : DFF_X1 port map( D => n2016, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_25_port, QN => n354);
   DataPath_REG_IN1_Q_reg_26_inst : DFF_X1 port map( D => n2015, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_26_port, QN => n356);
   DataPath_REG_IN1_Q_reg_28_inst : DFF_X1 port map( D => n2111, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_28_port, QN => n360);
   DataPath_REG_IN1_Q_reg_29_inst : DFF_X1 port map( D => n2110, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_29_port, QN => n361);
   DataPath_REG_IN1_Q_reg_30_inst : DFF_X1 port map( D => n2109, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_30_port, QN => n362);
   DataPath_REG_IN1_Q_reg_31_inst : DFF_X1 port map( D => n2108, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_31_port, QN => n363);
   DataPath_REG_B_Q_reg_0_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_0_port, QN => n1716);
   DataPath_REG_B_Q_reg_1_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_1_port, QN => n2140);
   DataPath_REG_B_Q_reg_4_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_4_port, QN => n4293);
   DataPath_REG_B_Q_reg_5_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_5_port, QN => n_3622);
   DataPath_REG_B_Q_reg_6_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_6_port, QN => n263);
   DataPath_REG_B_Q_reg_8_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_8_port, QN => n264);
   DataPath_REG_B_Q_reg_9_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_9_port, QN => n257);
   DataPath_REG_B_Q_reg_10_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_10_port, QN => n272);
   DataPath_REG_B_Q_reg_11_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_11_port, QN => n258);
   DataPath_REG_B_Q_reg_12_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_12_port, QN => n274);
   DataPath_REG_B_Q_reg_13_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_13_port, QN => n253);
   DataPath_REG_B_Q_reg_14_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_14_port, QN => n273);
   DataPath_REG_B_Q_reg_15_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_15_port, QN => n275);
   DataPath_REG_B_Q_reg_16_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_16_port, QN => n277);
   DataPath_REG_B_Q_reg_17_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_17_port, QN => n271);
   DataPath_REG_B_Q_reg_19_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_19_port, QN => n276);
   DataPath_RF_POP_ADDRGEN_curr_state_reg_1_inst : DFF_X1 port map( D => n12978
                           , CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_state_1_port, QN => 
                           n12949);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N61, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, QN => 
                           n12933);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_14_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N60, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_14_port, QN => 
                           n12934);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_13_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N59, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_13_port, QN => 
                           n12935);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_12_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N58, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_12_port, QN => 
                           n12936);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_11_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N57, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_11_port, QN => 
                           n12937);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_10_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N56, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_10_port, QN => 
                           n12938);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_9_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N55, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_9_port, QN => 
                           n12939);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_8_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N54, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_8_port, QN => 
                           n12940);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_7_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N53, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_7_port, QN => 
                           n12941);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_6_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N52, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_6_port, QN => 
                           n12942);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_5_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N51, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_5_port, QN => 
                           n12943);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_4_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N50, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_4_port, QN => 
                           n12944);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_3_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N49, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_3_port, QN => 
                           n12945);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_2_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N48, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_2_port, QN => 
                           n12946);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N47, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_1_port, QN => 
                           n12947);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N46, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_0_port, QN => 
                           n12948);
   DataPath_RF_POP_ADDRGEN_curr_state_reg_0_inst : DFF_X1 port map( D => n12979
                           , CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_state_0_port, QN => 
                           n12950);
   DataPath_WRF_CUhw_curr_data_reg_7_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n163, CK => CLK, Q => n_3623, QN 
                           => DataPath_WRF_CUhw_n31);
   DataPath_WRF_CUhw_curr_data_reg_6_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n162, CK => CLK, Q => n_3624, QN 
                           => DataPath_WRF_CUhw_n32);
   DataPath_WRF_CUhw_curr_data_reg_5_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n161, CK => CLK, Q => n_3625, QN 
                           => DataPath_WRF_CUhw_n33);
   DataPath_WRF_CUhw_curr_data_reg_4_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n160, CK => CLK, Q => n_3626, QN 
                           => DataPath_WRF_CUhw_n34);
   DataPath_WRF_CUhw_curr_data_reg_3_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n159, CK => CLK, Q => n_3627, QN 
                           => DataPath_WRF_CUhw_n35);
   DataPath_WRF_CUhw_curr_data_reg_2_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n158, CK => CLK, Q => n_3628, QN 
                           => DataPath_WRF_CUhw_n36);
   DataPath_WRF_CUhw_curr_data_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n157, CK => CLK, Q => n_3629, QN 
                           => DataPath_WRF_CUhw_n37);
   DataPath_WRF_CUhw_curr_data_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n156, CK => CLK, Q => n_3630, QN 
                           => DataPath_WRF_CUhw_n38);
   DataPath_WRF_CUhw_curr_data_reg_31_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n187, CK => CLK, Q => n_3631, QN 
                           => DataPath_WRF_CUhw_n7);
   DataPath_WRF_CUhw_curr_data_reg_30_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n186, CK => CLK, Q => n_3632, QN 
                           => DataPath_WRF_CUhw_n8);
   DataPath_WRF_CUhw_curr_data_reg_29_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n185, CK => CLK, Q => n_3633, QN 
                           => DataPath_WRF_CUhw_n9);
   DataPath_WRF_CUhw_curr_data_reg_28_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n184, CK => CLK, Q => n_3634, QN 
                           => DataPath_WRF_CUhw_n10);
   DataPath_WRF_CUhw_curr_data_reg_27_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n183, CK => CLK, Q => n_3635, QN 
                           => DataPath_WRF_CUhw_n11);
   DataPath_WRF_CUhw_curr_data_reg_26_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n182, CK => CLK, Q => n_3636, QN 
                           => DataPath_WRF_CUhw_n12);
   DataPath_WRF_CUhw_curr_data_reg_25_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n181, CK => CLK, Q => n_3637, QN 
                           => DataPath_WRF_CUhw_n13);
   DataPath_WRF_CUhw_curr_data_reg_24_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n180, CK => CLK, Q => n_3638, QN 
                           => DataPath_WRF_CUhw_n14);
   DataPath_WRF_CUhw_curr_data_reg_23_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n179, CK => CLK, Q => n_3639, QN 
                           => DataPath_WRF_CUhw_n15);
   DataPath_WRF_CUhw_curr_data_reg_22_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n178, CK => CLK, Q => n_3640, QN 
                           => DataPath_WRF_CUhw_n16);
   DataPath_WRF_CUhw_curr_data_reg_21_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n177, CK => CLK, Q => n_3641, QN 
                           => DataPath_WRF_CUhw_n17);
   DataPath_WRF_CUhw_curr_data_reg_20_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n176, CK => CLK, Q => n_3642, QN 
                           => DataPath_WRF_CUhw_n18);
   DataPath_WRF_CUhw_curr_data_reg_19_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n175, CK => CLK, Q => n_3643, QN 
                           => DataPath_WRF_CUhw_n19);
   DataPath_WRF_CUhw_curr_data_reg_18_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n174, CK => CLK, Q => n_3644, QN 
                           => DataPath_WRF_CUhw_n20);
   DataPath_WRF_CUhw_curr_data_reg_17_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n173, CK => CLK, Q => n_3645, QN 
                           => DataPath_WRF_CUhw_n21);
   DataPath_WRF_CUhw_curr_data_reg_16_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n172, CK => CLK, Q => n_3646, QN 
                           => DataPath_WRF_CUhw_n22);
   DataPath_WRF_CUhw_curr_data_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n171, CK => CLK, Q => n_3647, QN 
                           => DataPath_WRF_CUhw_n23);
   DataPath_WRF_CUhw_curr_data_reg_14_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n170, CK => CLK, Q => n_3648, QN 
                           => DataPath_WRF_CUhw_n24);
   DataPath_WRF_CUhw_curr_data_reg_13_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n169, CK => CLK, Q => n_3649, QN 
                           => DataPath_WRF_CUhw_n25);
   DataPath_WRF_CUhw_curr_data_reg_12_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n168, CK => CLK, Q => n_3650, QN 
                           => DataPath_WRF_CUhw_n26);
   DataPath_WRF_CUhw_curr_data_reg_11_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n167, CK => CLK, Q => n_3651, QN 
                           => DataPath_WRF_CUhw_n27);
   DataPath_WRF_CUhw_curr_data_reg_10_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n166, CK => CLK, Q => n_3652, QN 
                           => DataPath_WRF_CUhw_n28);
   DataPath_WRF_CUhw_curr_data_reg_9_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n165, CK => CLK, Q => n_3653, QN 
                           => DataPath_WRF_CUhw_n29);
   DataPath_WRF_CUhw_curr_data_reg_8_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_n164, CK => CLK, Q => n_3654, QN 
                           => DataPath_WRF_CUhw_n30);
   CU_I_CW_EX_reg_6_inst : DFF_X1 port map( D => CU_I_n129, CK => CLK, Q => 
                           n_3655, QN => CU_I_n105);
   CU_I_CW_EX_reg_5_inst : DFF_X1 port map( D => CU_I_n130, CK => CLK, Q => 
                           n_3656, QN => CU_I_n103);
   CU_I_CW_EX_reg_4_inst : DFF_X1 port map( D => CU_I_n131, CK => CLK, Q => 
                           n_3657, QN => CU_I_n101);
   CU_I_CW_EX_reg_3_inst : DFF_X1 port map( D => CU_I_n132, CK => CLK, Q => 
                           n_3658, QN => CU_I_n99);
   CU_I_CW_EX_reg_2_inst : DFF_X1 port map( D => CU_I_n133, CK => CLK, Q => 
                           n_3659, QN => CU_I_n140);
   CU_I_CW_EX_reg_1_inst : DFF_X1 port map( D => CU_I_n134, CK => CLK, Q => 
                           n_3660, QN => CU_I_n110);
   CU_I_CW_EX_reg_0_inst : DFF_X1 port map( D => CU_I_n135, CK => CLK, Q => 
                           n_3661, QN => CU_I_n112);
   CU_I_CW_MEM_reg_2_inst : DFF_X1 port map( D => CU_I_n157, CK => CLK, Q => 
                           n_3662, QN => CU_I_n98);
   CU_I_CW_MEM_reg_1_inst : DFF_X1 port map( D => CU_I_n141, CK => CLK, Q => 
                           n_3663, QN => CU_I_n111);
   CU_I_CW_MEM_reg_0_inst : DFF_X1 port map( D => CU_I_n142, CK => CLK, Q => 
                           n_3664, QN => CU_I_n113);
   CU_I_setcmp_1_reg_2_inst : DFF_X1 port map( D => CU_I_n145, CK => CLK, Q => 
                           n_3665, QN => n11484);
   CU_I_CW_MEM_reg_6_inst : DFF_X1 port map( D => CU_I_n136, CK => CLK, Q => 
                           n_3666, QN => DRAM_READNOTWRITE_port);
   DataPath_RF_PUSH_ADDRGEN_curr_state_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_n54, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n22);
   DataPath_WRF_CUhw_curr_state_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N144_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_state_0_port, QN => 
                           DataPath_WRF_CUhw_n73);
   DataPath_REG_IN2_Q_reg_30_inst : DFF_X1 port map( D => n2056, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_30_port, QN => n7075);
   DataPath_REG_IN2_Q_reg_29_inst : DFF_X1 port map( D => n1992, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_29_port, QN => n4431);
   DataPath_REG_IN2_Q_reg_28_inst : DFF_X1 port map( D => n1993, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_28_port, QN => n4433);
   DataPath_REG_IN2_Q_reg_27_inst : DFF_X1 port map( D => n1994, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_27_port, QN => n4364);
   DataPath_REG_IN2_Q_reg_26_inst : DFF_X1 port map( D => n1995, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_26_port, QN => n4368);
   DataPath_REG_IN2_Q_reg_25_inst : DFF_X1 port map( D => n1996, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_25_port, QN => n4354);
   DataPath_REG_IN2_Q_reg_24_inst : DFF_X1 port map( D => n1997, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_24_port, QN => n4357);
   DataPath_REG_IN2_Q_reg_23_inst : DFF_X1 port map( D => n1998, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_23_port, QN => n4406);
   DataPath_REG_IN2_Q_reg_22_inst : DFF_X1 port map( D => n1999, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_22_port, QN => n4409);
   DataPath_REG_IN2_Q_reg_21_inst : DFF_X1 port map( D => n2000, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_21_port, QN => n4415);
   DataPath_REG_IN2_Q_reg_20_inst : DFF_X1 port map( D => n2001, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_20_port, QN => n4412);
   DataPath_REG_IN2_Q_reg_31_inst : DFF_X1 port map( D => n2107, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_31_port, QN => n7078);
   DataPath_REG_B_Q_reg_31_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_31_port, QN => n7079);
   DataPath_REG_B_Q_reg_30_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_30_port, QN => n7076);
   DataPath_REG_B_Q_reg_29_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_29_port, QN => n4432);
   DataPath_REG_B_Q_reg_28_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_28_port, QN => n4434);
   DataPath_REG_B_Q_reg_27_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_27_port, QN => n4365);
   DataPath_REG_B_Q_reg_26_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_26_port, QN => n4369);
   DataPath_REG_B_Q_reg_25_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_25_port, QN => n4355);
   DataPath_REG_B_Q_reg_24_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_24_port, QN => n4358);
   DataPath_REG_B_Q_reg_23_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_23_port, QN => n4407);
   DataPath_REG_B_Q_reg_22_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_22_port, QN => n4410);
   DataPath_REG_B_Q_reg_21_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_21_port, QN => n4416);
   DataPath_REG_B_Q_reg_20_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_20_port, QN => n4413);
   DataPath_WRB3_Q_reg_4_inst : DFF_X1 port map( D => n8655, CK => CLK, Q => 
                           i_ADD_WB_4_port, QN => n11602);
   DataPath_WRB3_Q_reg_3_inst : DFF_X1 port map( D => n8656, CK => CLK, Q => 
                           i_ADD_WB_3_port, QN => n11601);
   DataPath_WRB3_Q_reg_2_inst : DFF_X1 port map( D => n8657, CK => CLK, Q => 
                           i_ADD_WB_2_port, QN => n11600);
   DataPath_WRB3_Q_reg_1_inst : DFF_X1 port map( D => n8658, CK => CLK, Q => 
                           i_ADD_WB_1_port, QN => n11599);
   DataPath_WRB3_Q_reg_0_inst : DFF_X1 port map( D => n8659, CK => CLK, Q => 
                           i_ADD_WB_0_port, QN => n11598);
   DataPath_WRB2_Q_reg_4_inst : DFF_X1 port map( D => n8650, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB2_4_port, QN => n_3667);
   DataPath_WRB2_Q_reg_3_inst : DFF_X1 port map( D => n8651, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB2_3_port, QN => n_3668);
   DataPath_WRB2_Q_reg_2_inst : DFF_X1 port map( D => n8652, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB2_2_port, QN => n_3669);
   DataPath_WRB2_Q_reg_1_inst : DFF_X1 port map( D => n8653, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB2_1_port, QN => n_3670);
   DataPath_WRB2_Q_reg_0_inst : DFF_X1 port map( D => n8654, CK => CLK, Q => 
                           DataPath_i_PIPLIN_WRB2_0_port, QN => n_3671);
   DataPath_RF_SWP_Q_reg_0_inst : DFF_X1 port map( D => n430, CK => CLK, Q => 
                           DataPath_RF_c_swin_0_port, QN => n_3672);
   DataPath_REG_MEM_ALUOUT_Q_reg_7_inst : DFF_X1 port map( D => n8780, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_7_port, QN => 
                           n_3673);
   DataPath_REG_MEM_ALUOUT_Q_reg_6_inst : DFF_X1 port map( D => n8781, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_6_port, QN => 
                           n_3674);
   DataPath_REG_MEM_ALUOUT_Q_reg_5_inst : DFF_X1 port map( D => n8782, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_5_port, QN => 
                           n_3675);
   DataPath_REG_MEM_ALUOUT_Q_reg_4_inst : DFF_X1 port map( D => n8783, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_4_port, QN => 
                           n_3676);
   DataPath_REG_MEM_ALUOUT_Q_reg_3_inst : DFF_X1 port map( D => n8784, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_3_port, QN => 
                           n_3677);
   DataPath_REG_MEM_ALUOUT_Q_reg_2_inst : DFF_X1 port map( D => n8785, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_2_port, QN => 
                           n_3678);
   DataPath_REG_MEM_ALUOUT_Q_reg_1_inst : DFF_X1 port map( D => n8786, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_1_port, QN => 
                           n_3679);
   DataPath_REG_MEM_ALUOUT_Q_reg_0_inst : DFF_X1 port map( D => n8787, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_0_port, QN => 
                           n_3680);
   DataPath_RF_SWP_Q_reg_2_inst : DFF_X1 port map( D => n428, CK => CLK, Q => 
                           DataPath_RF_c_swin_2_port, QN => n11604);
   DataPath_RF_SWP_Q_reg_1_inst : DFF_X1 port map( D => n427, CK => CLK, Q => 
                           DataPath_RF_c_swin_1_port, QN => n11603);
   DataPath_RF_SWP_Q_reg_3_inst : DFF_X1 port map( D => n426, CK => CLK, Q => 
                           DataPath_RF_c_swin_3_port, QN => n11605);
   DataPath_RF_SWP_Q_reg_4_inst : DFF_X1 port map( D => n425, CK => CLK, Q => 
                           DataPath_RF_c_swin_4_port, QN => n_3681);
   DataPath_REG_MEM_ALUOUT_Q_reg_31_inst : DFF_X1 port map( D => n8756, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_31_port, QN => 
                           n_3682);
   DataPath_REG_MEM_ALUOUT_Q_reg_30_inst : DFF_X1 port map( D => n8757, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_30_port, QN => 
                           n_3683);
   DataPath_REG_MEM_ALUOUT_Q_reg_29_inst : DFF_X1 port map( D => n8758, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_29_port, QN => 
                           n_3684);
   DataPath_REG_MEM_ALUOUT_Q_reg_28_inst : DFF_X1 port map( D => n8759, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_28_port, QN => 
                           n_3685);
   DataPath_REG_MEM_ALUOUT_Q_reg_27_inst : DFF_X1 port map( D => n8760, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_27_port, QN => 
                           n_3686);
   DataPath_REG_MEM_ALUOUT_Q_reg_26_inst : DFF_X1 port map( D => n8761, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_26_port, QN => 
                           n_3687);
   DataPath_REG_MEM_ALUOUT_Q_reg_25_inst : DFF_X1 port map( D => n8762, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_25_port, QN => 
                           n_3688);
   DataPath_REG_MEM_ALUOUT_Q_reg_24_inst : DFF_X1 port map( D => n8763, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_24_port, QN => 
                           n_3689);
   DataPath_REG_MEM_ALUOUT_Q_reg_23_inst : DFF_X1 port map( D => n8764, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_23_port, QN => 
                           n_3690);
   DataPath_REG_MEM_ALUOUT_Q_reg_22_inst : DFF_X1 port map( D => n8765, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_22_port, QN => 
                           n_3691);
   DataPath_REG_MEM_ALUOUT_Q_reg_21_inst : DFF_X1 port map( D => n8766, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_21_port, QN => 
                           n_3692);
   DataPath_REG_MEM_ALUOUT_Q_reg_20_inst : DFF_X1 port map( D => n8767, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_20_port, QN => 
                           n_3693);
   DataPath_REG_MEM_ALUOUT_Q_reg_19_inst : DFF_X1 port map( D => n8768, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_19_port, QN => 
                           n_3694);
   DataPath_REG_MEM_ALUOUT_Q_reg_18_inst : DFF_X1 port map( D => n8769, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_18_port, QN => 
                           n_3695);
   DataPath_REG_MEM_ALUOUT_Q_reg_17_inst : DFF_X1 port map( D => n8770, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_17_port, QN => 
                           n_3696);
   DataPath_REG_MEM_ALUOUT_Q_reg_16_inst : DFF_X1 port map( D => n8771, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_16_port, QN => 
                           n_3697);
   DataPath_REG_MEM_ALUOUT_Q_reg_15_inst : DFF_X1 port map( D => n8772, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_15_port, QN => 
                           n_3698);
   DataPath_REG_MEM_ALUOUT_Q_reg_14_inst : DFF_X1 port map( D => n8773, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_14_port, QN => 
                           n_3699);
   DataPath_REG_MEM_ALUOUT_Q_reg_13_inst : DFF_X1 port map( D => n8774, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_13_port, QN => 
                           n_3700);
   DataPath_REG_MEM_ALUOUT_Q_reg_12_inst : DFF_X1 port map( D => n8775, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_12_port, QN => 
                           n_3701);
   DataPath_REG_MEM_ALUOUT_Q_reg_11_inst : DFF_X1 port map( D => n8776, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_11_port, QN => 
                           n_3702);
   DataPath_REG_MEM_ALUOUT_Q_reg_10_inst : DFF_X1 port map( D => n8777, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_10_port, QN => 
                           n_3703);
   DataPath_REG_MEM_ALUOUT_Q_reg_9_inst : DFF_X1 port map( D => n8778, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_9_port, QN => 
                           n_3704);
   DataPath_REG_MEM_ALUOUT_Q_reg_8_inst : DFF_X1 port map( D => n8779, CK => 
                           CLK, Q => DataPath_i_REG_MEM_ALUOUT_8_port, QN => 
                           n_3705);
   DataPath_REG_ME_Q_reg_7_inst : DFF_X1 port map( D => n8716, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_7_port, QN => n_3706)
                           ;
   DataPath_REG_ME_Q_reg_6_inst : DFF_X1 port map( D => n8717, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_6_port, QN => n_3707)
                           ;
   DataPath_REG_ME_Q_reg_5_inst : DFF_X1 port map( D => n8718, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_5_port, QN => n_3708)
                           ;
   DataPath_REG_ME_Q_reg_4_inst : DFF_X1 port map( D => n8719, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_4_port, QN => n_3709)
                           ;
   DataPath_REG_ME_Q_reg_3_inst : DFF_X1 port map( D => n8720, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_3_port, QN => n_3710)
                           ;
   DataPath_REG_ME_Q_reg_2_inst : DFF_X1 port map( D => n8721, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_2_port, QN => n_3711)
                           ;
   DataPath_REG_ME_Q_reg_1_inst : DFF_X1 port map( D => n8722, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_1_port, QN => n_3712)
                           ;
   DataPath_REG_ME_Q_reg_0_inst : DFF_X1 port map( D => n8723, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_0_port, QN => n_3713)
                           ;
   DataPath_REG_ME_Q_reg_31_inst : DFF_X1 port map( D => n8692, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_31_port, QN => n_3714
                           );
   DataPath_REG_ME_Q_reg_30_inst : DFF_X1 port map( D => n8693, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_30_port, QN => n_3715
                           );
   DataPath_REG_ME_Q_reg_29_inst : DFF_X1 port map( D => n8694, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_29_port, QN => n_3716
                           );
   DataPath_REG_ME_Q_reg_28_inst : DFF_X1 port map( D => n8695, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_28_port, QN => n_3717
                           );
   DataPath_REG_ME_Q_reg_27_inst : DFF_X1 port map( D => n8696, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_27_port, QN => n_3718
                           );
   DataPath_REG_ME_Q_reg_26_inst : DFF_X1 port map( D => n8697, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_26_port, QN => n_3719
                           );
   DataPath_REG_ME_Q_reg_25_inst : DFF_X1 port map( D => n8698, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_25_port, QN => n_3720
                           );
   DataPath_REG_ME_Q_reg_24_inst : DFF_X1 port map( D => n8699, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_24_port, QN => n_3721
                           );
   DataPath_REG_ME_Q_reg_23_inst : DFF_X1 port map( D => n8700, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_23_port, QN => n_3722
                           );
   DataPath_REG_ME_Q_reg_22_inst : DFF_X1 port map( D => n8701, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_22_port, QN => n_3723
                           );
   DataPath_REG_ME_Q_reg_21_inst : DFF_X1 port map( D => n8702, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_21_port, QN => n_3724
                           );
   DataPath_REG_ME_Q_reg_20_inst : DFF_X1 port map( D => n8703, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_20_port, QN => n_3725
                           );
   DataPath_REG_ME_Q_reg_19_inst : DFF_X1 port map( D => n8704, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_19_port, QN => n_3726
                           );
   DataPath_REG_ME_Q_reg_18_inst : DFF_X1 port map( D => n8705, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_18_port, QN => n_3727
                           );
   DataPath_REG_ME_Q_reg_17_inst : DFF_X1 port map( D => n8706, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_17_port, QN => n_3728
                           );
   DataPath_REG_ME_Q_reg_16_inst : DFF_X1 port map( D => n8707, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_16_port, QN => n_3729
                           );
   DataPath_REG_ME_Q_reg_15_inst : DFF_X1 port map( D => n8708, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_15_port, QN => n_3730
                           );
   DataPath_REG_ME_Q_reg_14_inst : DFF_X1 port map( D => n8709, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_14_port, QN => n_3731
                           );
   DataPath_REG_ME_Q_reg_13_inst : DFF_X1 port map( D => n8710, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_13_port, QN => n_3732
                           );
   DataPath_REG_ME_Q_reg_12_inst : DFF_X1 port map( D => n8711, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_12_port, QN => n_3733
                           );
   DataPath_REG_ME_Q_reg_11_inst : DFF_X1 port map( D => n8712, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_11_port, QN => n_3734
                           );
   DataPath_REG_ME_Q_reg_10_inst : DFF_X1 port map( D => n8713, CK => CLK, Q =>
                           DataPath_i_REG_ME_DATA_DATAMEM_10_port, QN => n_3735
                           );
   DataPath_REG_ME_Q_reg_9_inst : DFF_X1 port map( D => n8714, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_9_port, QN => n_3736)
                           ;
   DataPath_REG_ME_Q_reg_8_inst : DFF_X1 port map( D => n8715, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_8_port, QN => n_3737)
                           ;
   DataPath_REG_CMP_Q_reg_1_inst : DFF_X1 port map( D => n2098, CK => CLK, Q =>
                           DataPath_i_LGET_1_port, QN => n_3738);
   CU_I_CW_WB_reg_0_inst : DFF_X1 port map( D => CU_I_N49, CK => CLK, Q => 
                           n_3739, QN => n11541);
   DataPath_WRF_CUhw_curr_addr_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N147_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_1_port, QN => n_3740);
   DataPath_WRF_CUhw_curr_addr_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N146_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_N109, QN => n_3741);
   CU_I_unsigned_1_reg : DFF_X1 port map( D => CU_I_n151, CK => CLK, Q => 
                           n_3742, QN => n11481);
   DataPath_WRF_CUhw_curr_state_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N145_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_state_1_port, QN => n_3743);
   DataPath_RF_CWP_Q_reg_4_inst : DFF_X1 port map( D => n8649, CK => CLK, Q => 
                           DataPath_RF_c_win_4_port, QN => n_3744);
   DataPath_WRF_CUhw_curr_addr_reg_2_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N148_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_2_port, QN => n_3745);
   DataPath_WRF_CUhw_curr_addr_reg_3_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N149_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_3_port, QN => n_3746);
   DataPath_WRF_CUhw_curr_addr_reg_4_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N150_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_4_port, QN => n_3747);
   DataPath_WRF_CUhw_curr_addr_reg_5_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N151, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_5_port, QN => n_3748);
   DataPath_WRF_CUhw_curr_addr_reg_6_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N152_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_6_port, QN => n_3749);
   DataPath_WRF_CUhw_curr_addr_reg_7_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N153_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_7_port, QN => n_3750);
   DataPath_WRF_CUhw_curr_addr_reg_8_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N154_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_8_port, QN => n_3751);
   DataPath_WRF_CUhw_curr_addr_reg_9_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N155_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_9_port, QN => n_3752);
   DataPath_WRF_CUhw_curr_addr_reg_10_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N156_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_10_port, QN => n_3753);
   DataPath_WRF_CUhw_curr_addr_reg_11_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N157_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_11_port, QN => n_3754);
   DataPath_WRF_CUhw_curr_addr_reg_12_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N158_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_12_port, QN => n_3755);
   DataPath_WRF_CUhw_curr_addr_reg_13_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N159_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_13_port, QN => n_3756);
   DataPath_WRF_CUhw_curr_addr_reg_14_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N160_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_14_port, QN => n_3757);
   DataPath_WRF_CUhw_curr_addr_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N161_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_15_port, QN => n_3758);
   DataPath_WRF_CUhw_curr_addr_reg_16_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N162_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_16_port, QN => n_3759);
   DataPath_WRF_CUhw_curr_addr_reg_17_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N163_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_17_port, QN => n_3760);
   DataPath_WRF_CUhw_curr_addr_reg_18_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N164_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_18_port, QN => n_3761);
   DataPath_WRF_CUhw_curr_addr_reg_19_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N165_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_19_port, QN => n_3762);
   DataPath_WRF_CUhw_curr_addr_reg_20_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N166_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_20_port, QN => n_3763);
   DataPath_WRF_CUhw_curr_addr_reg_21_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N167_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_21_port, QN => n_3764);
   DataPath_WRF_CUhw_curr_addr_reg_22_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N168_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_22_port, QN => n_3765);
   DataPath_WRF_CUhw_curr_addr_reg_23_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N169_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_23_port, QN => n_3766);
   DataPath_WRF_CUhw_curr_addr_reg_24_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N170_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_24_port, QN => n_3767);
   DataPath_WRF_CUhw_curr_addr_reg_25_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N171_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_25_port, QN => n_3768);
   DataPath_WRF_CUhw_curr_addr_reg_26_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N172_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_26_port, QN => n_3769);
   DataPath_WRF_CUhw_curr_addr_reg_27_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N173_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_27_port, QN => n_3770);
   DataPath_WRF_CUhw_curr_addr_reg_28_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N174_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_28_port, QN => n_3771);
   DataPath_WRF_CUhw_curr_addr_reg_29_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N175_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_29_port, QN => n_3772);
   DataPath_WRF_CUhw_curr_addr_reg_30_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N176_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_30_port, QN => n_3773);
   DataPath_WRF_CUhw_curr_addr_reg_31_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N177_port, CK => CLK, Q => 
                           DataPath_WRF_CUhw_curr_addr_31_port, QN => n_3774);
   DataPath_REG_IN2_Q_reg_18_inst : DFF_X1 port map( D => n2003, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_18_port, QN => n4393);
   DataPath_REG_B_Q_reg_18_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_18_port, QN => n4394);
   DataPath_REG_ALU_OUT_Q_reg_18_inst : DFF_X1 port map( D => n8673, CK => CLK,
                           Q => DRAM_ADDRESS_18_port, QN => n7942);
   DataPath_REG_ALU_OUT_Q_reg_19_inst : DFF_X1 port map( D => n8672, CK => CLK,
                           Q => DRAM_ADDRESS_19_port, QN => n7907);
   DataPath_REG_ALU_OUT_Q_reg_20_inst : DFF_X1 port map( D => n8671, CK => CLK,
                           Q => DRAM_ADDRESS_20_port, QN => n7872);
   DataPath_REG_ALU_OUT_Q_reg_21_inst : DFF_X1 port map( D => n8670, CK => CLK,
                           Q => DRAM_ADDRESS_21_port, QN => n7841);
   DataPath_REG_IN1_Q_reg_27_inst : DFF_X1 port map( D => n2112, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN1_27_port, QN => n4366);
   DataPath_REG_B_Q_reg_7_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_7_port, QN => n4302);
   DataPath_REG_IN2_Q_reg_2_inst : DFF_X1 port map( D => n2117, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_2_port, QN => n4441);
   DataPath_REG_A_Q_reg_12_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_12_port, QN => n_3775);
   DataPath_REG_A_Q_reg_13_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_13_port, QN => n_3776);
   DataPath_REG_A_Q_reg_9_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_9_port, QN => n_3777);
   DataPath_REG_B_Q_reg_2_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_2_port, QN => n4442);
   DataPath_REG_IN1_Q_reg_2_inst : DFF_X1 port map( D => n2090, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_2_port, QN => n4272);
   DataPath_REG_IN1_Q_reg_0_inst : DFF_X1 port map( D => n2092, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_0_port, QN => n4268);
   U137 : NOR2_X2 port map( A1 => n8325, A2 => n4106, ZN => CU_I_n152);
   U138 : NOR2_X2 port map( A1 => n11483, A2 => n4106, ZN => CU_I_n147);
   U139 : NOR2_X2 port map( A1 => CU_I_n118, A2 => n4106, ZN => CU_I_n146);
   U140 : NOR2_X2 port map( A1 => n4140, A2 => n4106, ZN => CU_I_n144);
   U141 : INV_X2 port map( A => CU_I_n58, ZN => CU_I_n154);
   U142 : NOR2_X2 port map( A1 => n7081, A2 => n4107, ZN => CU_I_n153);
   U143 : NOR2_X2 port map( A1 => CU_I_n114, A2 => n4107, ZN => CU_I_n155);
   U144 : NOR2_X2 port map( A1 => n11484, A2 => n4106, ZN => CU_I_n145);
   U145 : NOR2_X2 port map( A1 => n11540, A2 => n4107, ZN => CU_I_n156);
   U178 : NAND2_X2 port map( A1 => n1932, A2 => i_ALU_OP_1_port, ZN => CU_I_n58
                           );
   U179 : INV_X2 port map( A => DataPath_i_DONE_SPILL_EX, ZN => DataPath_RF_n9)
                           ;
   U180 : INV_X2 port map( A => n11597, ZN => DataPath_RF_n10);
   WS1_4_port <= '0';
   U182 : MUX2_X2 port map( A => n6593, B => n6592, S => n7835, Z => n616);
   U183 : MUX2_X1 port map( A => n6628, B => n6627, S => n246, Z => n6654);
   U185 : MUX2_X1 port map( A => n5347, B => n5346, S => n2246, Z => n5579);
   U186 : XNOR2_X1 port map( A => n200, B => n912, ZN => n1392);
   U187 : XOR2_X1 port map( A => n6585, B => n6629, Z => n200);
   U188 : NAND2_X1 port map( A1 => n6816, A2 => n1065, ZN => n201);
   U190 : XNOR2_X1 port map( A => n6604, B => n6603, ZN => n236);
   U191 : XNOR2_X1 port map( A => n568, B => n7003, ZN => n202);
   U192 : OAI21_X1 port map( B1 => n7895, B2 => n1517, A => n1783, ZN => n203);
   U193 : MUX2_X1 port map( A => n1690, B => n1691, S => n1702, Z => n1069);
   U194 : BUF_X1 port map( A => n6956, Z => n574);
   U195 : MUX2_X1 port map( A => n6517, B => n6518, S => n6369, Z => n6604);
   U196 : OAI21_X1 port map( B1 => n1097, B2 => n1847, A => n6510, ZN => n204);
   U197 : OAI21_X1 port map( B1 => n1445, B2 => n5990, A => n17153, ZN => n205)
                           ;
   U199 : CLKBUF_X1 port map( A => n6826, Z => n207);
   U200 : AND2_X2 port map( A1 => n7936, A2 => n6470, ZN => n1783);
   U201 : NAND3_X1 port map( A1 => n6273, A2 => n6301, A3 => n6274, ZN => n208)
                           ;
   U203 : MUX2_X1 port map( A => n6431, B => n6432, S => n529, Z => n708);
   U204 : MUX2_X1 port map( A => n6239, B => n6240, S => n6839, Z => n897);
   U205 : NAND2_X1 port map( A1 => n5886, A2 => n210, ZN => n211);
   U206 : NAND2_X1 port map( A1 => n5885, A2 => n1571, ZN => n212);
   U207 : NAND2_X1 port map( A1 => n211, A2 => n212, ZN => n892);
   U208 : INV_X1 port map( A => n1571, ZN => n210);
   U209 : MUX2_X1 port map( A => n5454, B => n5455, S => n213, Z => n704);
   U210 : INV_X32 port map( A => n2245, ZN => n213);
   U212 : AND2_X1 port map( A1 => n6458, A2 => n1195, ZN => n214);
   U213 : AND2_X1 port map( A1 => n6458, A2 => n1195, ZN => n1104);
   U214 : OAI21_X1 port map( B1 => n6252, B2 => n747, A => n6193, ZN => n215);
   U215 : XOR2_X1 port map( A => n4552, B => n1906, Z => n216);
   U216 : MUX2_X1 port map( A => n6321, B => n6322, S => n6839, Z => n780);
   U218 : OR2_X1 port map( A1 => n5197, A2 => n5453, ZN => n5440);
   U219 : NAND2_X1 port map( A1 => n5176, A2 => n2247, ZN => n217);
   U220 : OR2_X1 port map( A1 => n5499, A2 => n5284, ZN => n218);
   U221 : NAND2_X1 port map( A1 => n218, A2 => n5201, ZN => n5399);
   U222 : NAND2_X1 port map( A1 => n5536, A2 => n1224, ZN => n219);
   U224 : INV_X1 port map( A => n6378, ZN => n220);
   U225 : NAND2_X1 port map( A1 => n6335, A2 => n1555, ZN => n221);
   U226 : NAND2_X1 port map( A1 => n6335, A2 => n1555, ZN => n222);
   U227 : CLKBUF_X1 port map( A => n6551, Z => n1540);
   U228 : NAND2_X1 port map( A1 => n1752, A2 => n223, ZN => n224);
   U229 : NAND2_X1 port map( A1 => n1751, A2 => n6369, ZN => n225);
   U230 : NAND2_X1 port map( A1 => n225, A2 => n224, ZN => n585);
   U231 : INV_X1 port map( A => n6369, ZN => n223);
   U232 : MUX2_X2 port map( A => n276, B => n357, S => n526, Z => n6369);
   U233 : MUX2_X1 port map( A => n1869, B => n1868, S => n6495, Z => n1263);
   U234 : OR2_X1 port map( A1 => n5222, A2 => n5225, ZN => n226);
   U235 : NAND2_X1 port map( A1 => n226, A2 => n5218, ZN => n5219);
   U236 : OR2_X1 port map( A1 => n4721, A2 => n4722, ZN => n227);
   U237 : NAND2_X1 port map( A1 => n227, A2 => n4723, ZN => n4616);
   U238 : OR2_X1 port map( A1 => n251, A2 => n4715, ZN => n228);
   U239 : NAND2_X1 port map( A1 => n228, A2 => n4716, ZN => n4617);
   U240 : OR2_X1 port map( A1 => n6868, A2 => n6871, ZN => n229);
   U241 : NAND2_X1 port map( A1 => n229, A2 => n6866, ZN => n7322);
   U243 : NAND2_X1 port map( A1 => n5275, A2 => n5274, ZN => n230);
   U245 : MUX2_X1 port map( A => n1348, B => n1349, S => n4436, Z => n1347);
   U246 : AND2_X1 port map( A1 => n963, A2 => n964, ZN => n231);
   U247 : NOR2_X1 port map( A1 => n7679, A2 => n1699, ZN => n1305);
   U248 : XNOR2_X1 port map( A => n6397, B => n232, ZN => n235);
   U249 : INV_X32 port map( A => n1511, ZN => n232);
   U252 : BUF_X1 port map( A => n6177, Z => n911);
   U253 : BUF_X4 port map( A => n8158, Z => n2246);
   U254 : BUF_X4 port map( A => n8158, Z => n2245);
   U255 : BUF_X4 port map( A => n8245, Z => n2266);
   U256 : AND2_X2 port map( A1 => n8089, A2 => n8023, ZN => n1242);
   U257 : BUF_X4 port map( A => n1242, Z => n2224);
   U258 : INV_X2 port map( A => n1859, ZN => n2242);
   U259 : INV_X2 port map( A => n260, ZN => n2984);
   U260 : AND2_X2 port map( A1 => n6899, A2 => n6898, ZN => n1126);
   U262 : MUX2_X2 port map( A => n6953, B => n6952, S => n2267, Z => n725);
   U263 : MUX2_X2 port map( A => n6315, B => n6314, S => n8229, Z => n6354);
   U264 : MUX2_X2 port map( A => n7422, B => n7421, S => n7973, Z => n7423);
   U265 : CLKBUF_X1 port map( A => n5568, Z => n233);
   U266 : XNOR2_X1 port map( A => n1112, B => n5997, ZN => n6097);
   U267 : XNOR2_X1 port map( A => n234, B => n235, ZN => n6401);
   U268 : NAND2_X1 port map( A1 => n6399, A2 => n6400, ZN => n234);
   U270 : MUX2_X1 port map( A => n2259, B => n4498, S => n4462, Z => n4500);
   U271 : MUX2_X1 port map( A => n5727, B => n5726, S => n2243, Z => n698);
   U272 : XNOR2_X1 port map( A => n236, B => n6608, ZN => n6615);
   U273 : NAND2_X1 port map( A1 => n1167, A2 => n1341, ZN => n237);
   U274 : OR2_X1 port map( A1 => n6500, A2 => n6501, ZN => n238);
   U275 : NAND2_X1 port map( A1 => n238, A2 => n6499, ZN => n6489);
   U277 : NAND2_X1 port map( A1 => n1052, A2 => n239, ZN => n240);
   U278 : NAND2_X1 port map( A1 => n1051, A2 => n1407, ZN => n241);
   U279 : NAND2_X1 port map( A1 => n240, A2 => n241, ZN => n953);
   U280 : INV_X1 port map( A => n1407, ZN => n239);
   U281 : MUX2_X1 port map( A => n6377, B => n6376, S => n986, Z => n1094);
   U282 : AND2_X2 port map( A1 => n5717, A2 => n1893, ZN => n1826);
   U283 : MUX2_X1 port map( A => n6593, B => n6592, S => n7835, Z => n6823);
   U284 : MUX2_X1 port map( A => n6493, B => n6494, S => n6369, Z => n6810);
   U285 : NAND2_X1 port map( A1 => n1362, A2 => n6317, ZN => n242);
   U286 : OR2_X1 port map( A1 => n743, A2 => n6323, ZN => n243);
   U287 : NAND2_X1 port map( A1 => n243, A2 => n564, ZN => n603);
   U288 : MUX2_X1 port map( A => n6504, B => n6503, S => n1702, Z => n1182);
   U289 : NOR2_X1 port map( A1 => n6204, A2 => n6205, ZN => n244);
   U290 : NAND2_X1 port map( A1 => n1733, A2 => n6495, ZN => n245);
   U291 : NAND2_X1 port map( A1 => n245, A2 => n247, ZN => n1301);
   U292 : INV_X2 port map( A => n6369, ZN => n1702);
   U293 : MUX2_X1 port map( A => n5663, B => n5662, S => n2244, Z => n660);
   U294 : MUX2_X1 port map( A => n6601, B => n6602, S => n6495, Z => n6661);
   U295 : NAND2_X1 port map( A1 => n1734, A2 => n246, ZN => n247);
   U296 : NAND2_X1 port map( A1 => n1733, A2 => n6495, ZN => n248);
   U297 : NAND2_X1 port map( A1 => n247, A2 => n248, ZN => n568);
   U298 : INV_X1 port map( A => n6495, ZN => n246);
   U299 : CLKBUF_X1 port map( A => n5164, Z => n249);
   U303 : CLKBUF_X1 port map( A => n897, Z => n250);
   U304 : BUF_X1 port map( A => n5501, Z => n1318);
   U307 : MUX2_X2 port map( A => n5340, B => n5339, S => n2246, Z => n5570);
   U308 : OR2_X1 port map( A1 => n1312, A2 => n1311, ZN => n5576);
   U309 : MUX2_X1 port map( A => DataPath_i_PIPLIN_IN1_11_port, B => 
                           DataPath_i_PIPLIN_A_11_port, S => n4142, Z => n252);
   U310 : INV_X4 port map( A => n252, ZN => n7257);
   U311 : INV_X2 port map( A => n7257, ZN => n2207);
   U312 : OR2_X2 port map( A1 => n5523, A2 => n5579, ZN => n5568);
   U313 : CLKBUF_X1 port map( A => n5380, Z => n801);
   U314 : MUX2_X1 port map( A => n5340, B => n5339, S => n2246, Z => n471);
   U316 : OR2_X1 port map( A1 => n4702, A2 => n4687, ZN => n1205);
   U317 : INV_X1 port map( A => n6730, ZN => n1376);
   U318 : OAI22_X1 port map( A1 => n2179, A2 => n2142, B1 => n2188, B2 => n7283
                           , ZN => n4729);
   U319 : INV_X1 port map( A => n1377, ZN => n6752);
   U320 : AND2_X1 port map( A1 => n6921, A2 => n6905, ZN => n1850);
   U321 : OAI22_X1 port map( A1 => n2215, A2 => n2181, B1 => n2218, B2 => n2213
                           , ZN => n5549);
   U322 : OAI22_X1 port map( A1 => n2178, A2 => n2183, B1 => n2182, B2 => n2179
                           , ZN => n5845);
   U323 : INV_X1 port map( A => n1500, ZN => n6043);
   U324 : INV_X1 port map( A => n979, ZN => n6074);
   U325 : OR2_X1 port map( A1 => n504, A2 => n5529, ZN => n5612);
   U326 : OR2_X1 port map( A1 => n4966, A2 => n5059, ZN => n1496);
   U327 : OAI22_X1 port map( A1 => n2209, A2 => n7285, B1 => n2205, B2 => n7284
                           , ZN => n6221);
   U328 : INV_X1 port map( A => n5807, ZN => n5896);
   U329 : INV_X1 port map( A => n6793, ZN => n6797);
   U330 : INV_X1 port map( A => n6343, ZN => n6396);
   U331 : INV_X1 port map( A => n941, ZN => n4805);
   U332 : INV_X1 port map( A => n6396, ZN => n1511);
   U334 : INV_X1 port map( A => n2268, ZN => n1584);
   U335 : INV_X1 port map( A => n5281, ZN => n5426);
   U337 : INV_X1 port map( A => n2245, ZN => n1092);
   U338 : INV_X1 port map( A => n827, ZN => n4589);
   U339 : OAI22_X1 port map( A1 => n2227, A2 => n7244, B1 => n2240, B2 => n7243
                           , ZN => n7005);
   U340 : INV_X1 port map( A => n744, ZN => n5949);
   U341 : AND2_X1 port map( A1 => n955, A2 => n954, ZN => n743);
   U342 : AND2_X1 port map( A1 => n4940, A2 => n1568, ZN => n1350);
   U343 : AND2_X1 port map( A1 => n4870, A2 => n4871, ZN => n1795);
   U345 : NAND2_X1 port map( A1 => n6595, A2 => n7247, ZN => n7248);
   U346 : INV_X1 port map( A => n2245, ZN => n700);
   U347 : AND2_X1 port map( A1 => n8165, A2 => n501, ZN => n1790);
   U348 : NOR4_X1 port map( A1 => DataPath_RF_SPILLADDR_ENC_n12, A2 => 
                           DataPath_RF_SPILLADDR_ENC_n13, A3 => 
                           DataPath_RF_spill_address_ext_4_port, A4 => 
                           DataPath_RF_SPILLADDR_ENC_n14, ZN => 
                           DataPath_RF_spill_address_3_port);
   U349 : OR2_X1 port map( A1 => n789, A2 => n7242, ZN => n562);
   U350 : AND2_X1 port map( A1 => n916, A2 => n7007, ZN => n1781);
   U351 : XOR2_X1 port map( A => n7800, B => n7835, Z => n7247);
   U352 : INV_X1 port map( A => n1894, ZN => n907);
   U353 : INV_X1 port map( A => n1872, ZN => n1091);
   U354 : OAI211_X1 port map( C1 => n8052, C2 => n8082, A => n8051, B => n8050,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n179);
   U355 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n7, A2 => DataPath_RF_DEC_n15
                           , ZN => DataPath_RF_dec_output_8_port);
   U356 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n7, A2 => DataPath_RF_DEC_n17
                           , ZN => DataPath_RF_dec_output_24_port);
   U357 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n8, A2 => DataPath_RF_DEC_n15
                           , ZN => DataPath_RF_dec_output_9_port);
   U358 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n8, A2 => DataPath_RF_DEC_n17
                           , ZN => DataPath_RF_dec_output_25_port);
   U359 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n9, A2 => DataPath_RF_DEC_n17
                           , ZN => DataPath_RF_dec_output_26_port);
   U360 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n9, A2 => DataPath_RF_DEC_n15
                           , ZN => DataPath_RF_dec_output_10_port);
   U361 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n10, A2 => 
                           DataPath_RF_DEC_n17, ZN => 
                           DataPath_RF_dec_output_27_port);
   U362 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n10, A2 => 
                           DataPath_RF_DEC_n15, ZN => 
                           DataPath_RF_dec_output_11_port);
   U363 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n11, A2 => 
                           DataPath_RF_DEC_n17, ZN => 
                           DataPath_RF_dec_output_28_port);
   U364 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n11, A2 => 
                           DataPath_RF_DEC_n15, ZN => 
                           DataPath_RF_dec_output_12_port);
   U365 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n12, A2 => 
                           DataPath_RF_DEC_n17, ZN => 
                           DataPath_RF_dec_output_29_port);
   U366 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n12, A2 => 
                           DataPath_RF_DEC_n15, ZN => 
                           DataPath_RF_dec_output_13_port);
   U367 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n13, A2 => 
                           DataPath_RF_DEC_n17, ZN => 
                           DataPath_RF_dec_output_30_port);
   U368 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n13, A2 => 
                           DataPath_RF_DEC_n15, ZN => 
                           DataPath_RF_dec_output_14_port);
   U369 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n14, A2 => 
                           DataPath_RF_DEC_n17, ZN => 
                           DataPath_RF_dec_output_31_port);
   U370 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n14, A2 => 
                           DataPath_RF_DEC_n15, ZN => 
                           DataPath_RF_dec_output_15_port);
   U371 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n7, A2 => DataPath_RF_DEC_n16
                           , ZN => DataPath_RF_dec_output_16_port);
   U372 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n8, A2 => DataPath_RF_DEC_n16
                           , ZN => DataPath_RF_dec_output_17_port);
   U373 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n9, A2 => DataPath_RF_DEC_n16
                           , ZN => DataPath_RF_dec_output_18_port);
   U374 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n10, A2 => 
                           DataPath_RF_DEC_n16, ZN => 
                           DataPath_RF_dec_output_19_port);
   U375 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n11, A2 => 
                           DataPath_RF_DEC_n16, ZN => 
                           DataPath_RF_dec_output_20_port);
   U376 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n12, A2 => 
                           DataPath_RF_DEC_n16, ZN => 
                           DataPath_RF_dec_output_21_port);
   U377 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n13, A2 => 
                           DataPath_RF_DEC_n16, ZN => 
                           DataPath_RF_dec_output_22_port);
   U378 : NOR2_X1 port map( A1 => DataPath_RF_DEC_n14, A2 => 
                           DataPath_RF_DEC_n16, ZN => 
                           DataPath_RF_dec_output_23_port);
   U379 : NOR3_X1 port map( A1 => n12957, A2 => n12960, A3 => n4155, ZN => 
                           DataPath_i_DONE_FILL_EX);
   U380 : NOR2_X1 port map( A1 => DataPath_LDSTR_n80, A2 => n4118, ZN => 
                           DataPath_LDSTR_n47);
   U381 : CLKBUF_X3 port map( A => n8245, Z => n2265);
   U382 : BUF_X2 port map( A => n8263, Z => n2267);
   U383 : INV_X2 port map( A => n6839, ZN => n8229);
   U384 : BUF_X2 port map( A => n8263, Z => n2268);
   U385 : INV_X2 port map( A => n528, ZN => n529);
   U386 : CLKBUF_X3 port map( A => n799, Z => n2247);
   U387 : INV_X2 port map( A => n529, ZN => n7973);
   U388 : INV_X1 port map( A => n8229, ZN => n1407);
   U389 : AND2_X1 port map( A1 => n1907, A2 => n1861, ZN => n260);
   U390 : INV_X1 port map( A => n2267, ZN => n1731);
   U391 : INV_X1 port map( A => n6594, ZN => n7771);
   U392 : MUX2_X1 port map( A => n4416, B => n4415, S => n527, Z => n6495);
   U393 : INV_X1 port map( A => n1006, ZN => n960);
   U394 : INV_X1 port map( A => n6316, ZN => n6319);
   U395 : INV_X1 port map( A => n799, ZN => n6890);
   U396 : AND2_X1 port map( A1 => n6096, A2 => n6073, ZN => n262);
   U397 : OR2_X1 port map( A1 => n2273, A2 => n4129, ZN => n266);
   U398 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_30_port, B => 
                           n1987, Z => n267);
   U399 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_29_port, B => 
                           n1984, Z => n268);
   U400 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_28_port, B => 
                           n1981, Z => n269);
   U401 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_31_port, B => 
                           n2127, ZN => n270);
   U402 : AND2_X1 port map( A1 => n8042, A2 => n11498, ZN => n282);
   U403 : INV_X1 port map( A => n6495, ZN => n7835);
   U404 : MUX2_X1 port map( A => n4365, B => n4364, S => n526, Z => n7471);
   U405 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_25_port, B => 
                           n1974, Z => n283);
   U406 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_26_port, B => 
                           n1977, Z => n284);
   U407 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_27_port, B => 
                           n1979, Z => n285);
   U408 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_17_port, B => 
                           n1957, Z => n286);
   U409 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_18_port, B => 
                           n1958, Z => n287);
   U410 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_19_port, B => 
                           n1936, Z => n288);
   U411 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_20_port, B => 
                           n1937, Z => n289);
   U412 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_21_port, B => 
                           n1938, Z => n290);
   U413 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_22_port, B => 
                           n1939, Z => n291);
   U414 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_23_port, B => 
                           n1940, Z => n292);
   U415 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_24_port, B => 
                           n1971, Z => n293);
   U416 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_16_port, B => 
                           n1956, Z => n294);
   U417 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_8_port, B => n1947
                           , Z => n295);
   U418 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_9_port, B => n1948
                           , Z => n296);
   U419 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_10_port, B => 
                           n1949, Z => n297);
   U420 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_11_port, B => 
                           n1950, Z => n298);
   U421 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_12_port, B => 
                           n1951, Z => n299);
   U422 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_13_port, B => 
                           n1952, Z => n300);
   U423 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_14_port, B => 
                           n1953, Z => n301);
   U424 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_15_port, B => 
                           n1954, Z => n302);
   U425 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_n73, A2 => 
                           DataPath_WRF_CUhw_curr_state_1_port, ZN => n303);
   U426 : XOR2_X1 port map( A => DataPath_WRF_CUhw_N26_port, B => 
                           DataPath_WRF_CUhw_curr_addr_2_port, Z => n304);
   U427 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_4_port, B => n1955
                           , Z => n305);
   U428 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_5_port, B => n1944
                           , Z => n306);
   U429 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_6_port, B => n1945
                           , Z => n307);
   U430 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_7_port, B => n1946
                           , Z => n308);
   U431 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_3_port, B => n1991
                           , Z => n309);
   U432 : AND2_X1 port map( A1 => n1053, A2 => n6855, ZN => n310);
   U433 : XNOR2_X1 port map( A => n4729, B => n4728, ZN => n311);
   U434 : INV_X1 port map( A => n5811, ZN => n5955);
   U435 : INV_X1 port map( A => n5523, ZN => n5588);
   U436 : INV_X1 port map( A => n5829, ZN => n5868);
   U437 : INV_X1 port map( A => n5537, ZN => n5679);
   U438 : INV_X1 port map( A => n5299, ZN => n5348);
   U439 : AND2_X1 port map( A1 => n4802, A2 => n4822, ZN => n312);
   U440 : AND2_X1 port map( A1 => n5460, A2 => n8165, ZN => n313);
   U441 : OR2_X1 port map( A1 => n6775, A2 => n6776, ZN => n314);
   U442 : AND2_X1 port map( A1 => n6957, A2 => n2266, ZN => n315);
   U444 : AND3_X1 port map( A1 => n4823, A2 => n4822, A3 => n2251, ZN => n316);
   U445 : INV_X1 port map( A => n7624, ZN => n2228);
   U446 : AND2_X1 port map( A1 => n4835, A2 => n818, ZN => n317);
   U447 : AND2_X1 port map( A1 => n4669, A2 => n4765, ZN => n319);
   U448 : AND2_X1 port map( A1 => n4735, A2 => n4736, ZN => n320);
   U449 : OR2_X1 port map( A1 => n637, A2 => n774, ZN => n321);
   U450 : MUX2_X1 port map( A => n6423, B => n6424, S => n529, Z => n1070);
   U451 : AND2_X1 port map( A1 => n6764, A2 => n6762, ZN => n322);
   U452 : INV_X1 port map( A => n5526, ZN => n5562);
   U453 : INV_X1 port map( A => n5562, ZN => n1603);
   U454 : INV_X1 port map( A => n6488, ZN => n6515);
   U455 : AND2_X1 port map( A1 => n6085, A2 => n2266, ZN => n338);
   U456 : OAI22_X1 port map( A1 => n2240, A2 => n7291, B1 => n2239, B2 => n2185
                           , ZN => n6142);
   U457 : INV_X1 port map( A => n6589, ZN => n6603);
   U458 : AND2_X1 port map( A1 => n6057, A2 => n2266, ZN => n339);
   U459 : INV_X1 port map( A => n6355, ZN => n6436);
   U460 : INV_X1 port map( A => n6468, ZN => n6522);
   U461 : INV_X1 port map( A => n6222, ZN => n6241);
   U462 : INV_X1 port map( A => n6200, ZN => n6292);
   U463 : INV_X1 port map( A => n5805, ZN => n5860);
   U464 : INV_X1 port map( A => n6765, ZN => n6774);
   U465 : INV_X1 port map( A => n6574, ZN => n6619);
   U466 : INV_X1 port map( A => n6484, ZN => n6523);
   U467 : OAI22_X1 port map( A1 => n2199, A2 => n7285, B1 => n2197, B2 => n7284
                           , ZN => n6217);
   U468 : AND2_X1 port map( A1 => n6079, A2 => n6967, ZN => n340);
   U469 : AND2_X1 port map( A1 => n6160, A2 => n6967, ZN => n341);
   U470 : OR2_X1 port map( A1 => n6089, A2 => n2266, ZN => n342);
   U471 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_16_port, A2 => n8325, ZN 
                           => n343);
   U472 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_15_port, A2 => n8325, ZN 
                           => n344);
   U473 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_12_port, A2 => n8325, ZN 
                           => n345);
   U474 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_11_port, A2 => n8325, ZN 
                           => n346);
   U475 : OR2_X1 port map( A1 => n5845, A2 => n6776, ZN => n347);
   U476 : OR2_X1 port map( A1 => n6060, A2 => n2266, ZN => n348);
   U477 : INV_X1 port map( A => n6802, ZN => n6806);
   U478 : OR2_X1 port map( A1 => n6057, A2 => n6967, ZN => n349);
   U479 : OAI22_X1 port map( A1 => n2199, A2 => n7248, B1 => n2197, B2 => n7247
                           , ZN => n7449);
   U480 : INV_X1 port map( A => n2268, ZN => n1211);
   U481 : INV_X1 port map( A => n6984, ZN => n6982);
   U482 : XNOR2_X1 port map( A => n4373, B => n7644, ZN => n364);
   U483 : AND2_X1 port map( A1 => n2272, A2 => n7617, ZN => n365);
   U484 : AND2_X1 port map( A1 => n2272, A2 => n7748, ZN => n366);
   U485 : AND2_X1 port map( A1 => n2272, A2 => n8326, ZN => n367);
   U486 : AND2_X1 port map( A1 => n7210, A2 => n11539, ZN => n368);
   U487 : AND2_X1 port map( A1 => n7603, A2 => n7567, ZN => n369);
   U488 : AND2_X1 port map( A1 => n1860, A2 => n4284, ZN => n370);
   U489 : XNOR2_X1 port map( A => n7516, B => n7581, ZN => n371);
   U490 : AND2_X1 port map( A1 => n4387, A2 => n4386, ZN => n372);
   U491 : AND2_X1 port map( A1 => n4381, A2 => n4380, ZN => n373);
   U492 : AND2_X1 port map( A1 => n4375, A2 => n4374, ZN => n374);
   U493 : AND2_X1 port map( A1 => n7761, A2 => n7787, ZN => n375);
   U494 : AND2_X1 port map( A1 => n7892, A2 => n7918, ZN => n376);
   U497 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_10_port, A2 => n8325, ZN 
                           => n377);
   U498 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_9_port, A2 => n8325, ZN =>
                           n378);
   U499 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_8_port, A2 => n8325, ZN =>
                           n379);
   U500 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_7_port, A2 => n8325, ZN =>
                           n380);
   U501 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_6_port, A2 => n8325, ZN =>
                           n381);
   U502 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_5_port, A2 => n8325, ZN =>
                           n382);
   U503 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_4_port, A2 => n8325, ZN =>
                           n383);
   U504 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_3_port, A2 => n8325, ZN =>
                           n384);
   U505 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_2_port, A2 => n8325, ZN =>
                           n385);
   U506 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_1_port, A2 => n8325, ZN =>
                           n386);
   U507 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_30_port, B => 
                           n1989, Z => n387);
   U508 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_25_port, B => 
                           n1982, Z => n388);
   U509 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_26_port, B => 
                           n1983, Z => n389);
   U510 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_29_port, B => 
                           n1988, Z => n390);
   U511 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_28_port, B => 
                           n1986, Z => n391);
   U512 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_27_port, B => 
                           n1985, Z => n392);
   U513 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_17_port, B => 
                           n1972, Z => n393);
   U514 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_18_port, B => 
                           n1973, Z => n394);
   U515 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_19_port, B => 
                           n1975, Z => n395);
   U516 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_20_port, B => 
                           n1976, Z => n396);
   U517 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_21_port, B => 
                           n1941, Z => n397);
   U518 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_22_port, B => 
                           n1942, Z => n398);
   U519 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_23_port, B => 
                           n1943, Z => n399);
   U520 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_24_port, B => 
                           n1980, Z => n400);
   U521 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_16_port, B => 
                           n1970, Z => n401);
   U522 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_11_port, B => 
                           n1965, Z => n402);
   U523 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_12_port, B => 
                           n1966, Z => n403);
   U524 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_13_port, B => 
                           n1967, Z => n404);
   U525 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_14_port, B => 
                           n1968, Z => n405);
   U526 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_15_port, B => 
                           n1969, Z => n406);
   U527 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_31_port, B => 
                           n2128, ZN => n407);
   U528 : INV_X1 port map( A => n7471, ZN => n7647);
   U529 : AND3_X1 port map( A1 => n2253, A2 => n8140, A3 => n7083, ZN => n410);
   U530 : AND2_X1 port map( A1 => n7550, A2 => n2258, ZN => n411);
   U531 : XOR2_X1 port map( A => DataPath_WRF_CUhw_N217, B => 
                           DataPath_WRF_CUhw_curr_addr_2_port, Z => n412);
   U532 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_4_port, B => n1978
                           , Z => n413);
   U533 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_5_port, B => n1959
                           , Z => n414);
   U534 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_6_port, B => n1960
                           , Z => n415);
   U535 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_7_port, B => n1961
                           , Z => n416);
   U536 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_8_port, B => n1962
                           , Z => n417);
   U537 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_9_port, B => n1963
                           , Z => n418);
   U538 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_10_port, B => 
                           n1964, Z => n419);
   U539 : XOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_3_port, B => n1990
                           , Z => n420);
   U540 : AND2_X1 port map( A1 => DataPath_RF_next_cwp_1_port, A2 => n4262, ZN 
                           => n421);
   U541 : AND2_X1 port map( A1 => DataPath_RF_next_cwp_2_port, A2 => n4261, ZN 
                           => n422);
   U542 : AND2_X1 port map( A1 => DataPath_RF_next_cwp_3_port, A2 => n4257, ZN 
                           => n423);
   U543 : AND2_X1 port map( A1 => DataPath_RF_next_swp_4_port, A2 => n4260, ZN 
                           => n425);
   U544 : AND2_X1 port map( A1 => DataPath_RF_next_swp_3_port, A2 => n4260, ZN 
                           => n426);
   U545 : AND2_X1 port map( A1 => DataPath_RF_next_swp_1_port, A2 => n4260, ZN 
                           => n427);
   U546 : AND2_X1 port map( A1 => DataPath_RF_next_swp_2_port, A2 => n4260, ZN 
                           => n428);
   U547 : OR2_X1 port map( A1 => DataPath_RF_next_cwp_0_port, A2 => n4184, ZN 
                           => n429);
   U548 : OR2_X1 port map( A1 => DataPath_RF_next_swp_0_port, A2 => n4183, ZN 
                           => n430);
   U549 : XNOR2_X1 port map( A => n17209, B => n7641, ZN => n431);
   U550 : NAND2_X1 port map( A1 => n7060, A2 => n432, ZN => n593);
   U551 : NOR2_X1 port map( A1 => n7471, A2 => n7588, ZN => n432);
   U552 : NAND2_X1 port map( A1 => n593, A2 => n592, ZN => n433);
   U553 : CLKBUF_X1 port map( A => n1796, Z => n434);
   U554 : NOR2_X1 port map( A1 => n4624, A2 => n4733, ZN => n435);
   U555 : OR2_X2 port map( A1 => n6345, A2 => n1031, ZN => n6416);
   U556 : MUX2_X2 port map( A => n6875, B => n6874, S => n804, Z => n7342);
   U557 : MUX2_X2 port map( A => n4714, B => n4713, S => n2250, Z => n5012);
   U558 : MUX2_X2 port map( A => n7334, B => n7333, S => n2250, Z => n7335);
   U559 : XNOR2_X1 port map( A => n6824, B => n599, ZN => n436);
   U561 : AND2_X1 port map( A1 => n5072, A2 => n4963, ZN => n438);
   U562 : CLKBUF_X1 port map( A => n6066, Z => n439);
   U563 : MUX2_X1 port map( A => n6111, B => n6110, S => n2266, Z => n6272);
   U564 : INV_X1 port map( A => n6366, ZN => n440);
   U565 : XNOR2_X1 port map( A => n1822, B => n5431, ZN => n441);
   U567 : BUF_X1 port map( A => n608, Z => n1141);
   U568 : AND2_X1 port map( A1 => n5472, A2 => n5473, ZN => n1785);
   U569 : NAND2_X1 port map( A1 => n5162, A2 => n17197, ZN => n443);
   U570 : OR2_X1 port map( A1 => n251, A2 => n4679, ZN => n444);
   U571 : NAND2_X1 port map( A1 => n444, A2 => n4717, ZN => n4680);
   U572 : OR2_X1 port map( A1 => n4695, A2 => n4690, ZN => n445);
   U573 : NAND2_X1 port map( A1 => n445, A2 => n4689, ZN => n5220);
   U574 : AND2_X1 port map( A1 => n6917, A2 => n6916, ZN => n446);
   U575 : AND2_X1 port map( A1 => n6915, A2 => n6914, ZN => n447);
   U576 : NOR3_X1 port map( A1 => n17218, A2 => n447, A3 => n446, ZN => n7379);
   U577 : MUX2_X1 port map( A => n6409, B => n6408, S => n7973, Z => n6526);
   U578 : XNOR2_X1 port map( A => n1357, B => n5127, ZN => n448);
   U579 : MUX2_X2 port map( A => n5371, B => n5372, S => n1092, Z => n975);
   U580 : BUF_X1 port map( A => n4813, Z => n449);
   U581 : INV_X1 port map( A => n4630, ZN => n450);
   U582 : XNOR2_X1 port map( A => n4798, B => n4797, ZN => n4813);
   U583 : XNOR2_X1 port map( A => n5593, B => n5521, ZN => n451);
   U584 : XNOR2_X1 port map( A => n1603, B => n5561, ZN => n1604);
   U585 : NAND2_X1 port map( A1 => n555, A2 => n772, ZN => n452);
   U586 : MUX2_X1 port map( A => n6137, B => n6138, S => n750, Z => n6203);
   U587 : MUX2_X1 port map( A => n5869, B => n5870, S => n1211, Z => n6095);
   U588 : NOR2_X1 port map( A1 => n5609, A2 => n5549, ZN => n1791);
   U589 : XNOR2_X1 port map( A => n1416, B => n6461, ZN => n1073);
   U590 : CLKBUF_X1 port map( A => n1354, Z => n453);
   U591 : AND2_X1 port map( A1 => n787, A2 => n6857, ZN => n454);
   U592 : OR2_X1 port map( A1 => n6733, A2 => n6736, ZN => n455);
   U593 : NAND2_X1 port map( A1 => n455, A2 => n6712, ZN => n6856);
   U594 : CLKBUF_X1 port map( A => n6263, Z => n1194);
   U595 : NAND2_X1 port map( A1 => n480, A2 => n481, ZN => n456);
   U596 : INV_X1 port map( A => n1193, ZN => n457);
   U597 : MUX2_X2 port map( A => n6659, B => n6658, S => n7771, Z => n1193);
   U598 : MUX2_X1 port map( A => n5384, B => n5383, S => n2246, Z => n664);
   U599 : MUX2_X1 port map( A => n5454, B => n5455, S => n936, Z => n5697);
   U601 : MUX2_X1 port map( A => n5923, B => n5922, S => n464, Z => n6008);
   U602 : MUX2_X2 port map( A => n6130, B => n6131, S => n750, Z => n6296);
   U603 : AND2_X1 port map( A1 => n1403, A2 => n458, ZN => n1829);
   U604 : AND2_X1 port map( A1 => n1402, A2 => n6577, ZN => n458);
   U605 : OR2_X1 port map( A1 => n6405, A2 => n6360, ZN => n459);
   U606 : NAND2_X1 port map( A1 => n459, A2 => n640, ZN => n6338);
   U607 : NOR2_X1 port map( A1 => n929, A2 => n960, ZN => n460);
   U608 : NAND2_X1 port map( A1 => n586, A2 => n710, ZN => n461);
   U609 : INV_X1 port map( A => n5771, ZN => n462);
   U610 : AND2_X1 port map( A1 => n4757, A2 => n4756, ZN => n463);
   U611 : INV_X1 port map( A => n749, ZN => n6933);
   U612 : NAND2_X1 port map( A1 => n5890, A2 => n464, ZN => n465);
   U613 : NAND2_X1 port map( A1 => n5891, A2 => n1743, ZN => n466);
   U614 : NAND2_X1 port map( A1 => n465, A2 => n466, ZN => n1533);
   U615 : INV_X1 port map( A => n1743, ZN => n464);
   U616 : INV_X1 port map( A => n2268, ZN => n1743);
   U617 : CLKBUF_X1 port map( A => n1403, Z => n467);
   U618 : XNOR2_X1 port map( A => n468, B => n7399, ZN => n7409);
   U619 : XOR2_X1 port map( A => n7397, B => n7398, Z => n468);
   U620 : MUX2_X2 port map( A => n5238, B => n5239, S => n6890, Z => n5326);
   U621 : NAND2_X1 port map( A1 => n6588, A2 => n628, ZN => n469);
   U623 : NAND2_X1 port map( A1 => n1089, A2 => n5673, ZN => n1378);
   U624 : MUX2_X1 port map( A => n6614, B => n6615, S => n6495, Z => n1175);
   U625 : AND2_X1 port map( A1 => n6892, A2 => n6891, ZN => n749);
   U626 : INV_X1 port map( A => n4659, ZN => n472);
   U627 : OR2_X1 port map( A1 => n6203, A2 => n6312, ZN => n6299);
   U628 : NAND2_X1 port map( A1 => n6587, A2 => n6589, ZN => n473);
   U629 : NAND2_X1 port map( A1 => n473, A2 => n6571, ZN => n6597);
   U630 : MUX2_X2 port map( A => n5378, B => n5377, S => n2246, Z => n504);
   U631 : MUX2_X2 port map( A => n4727, B => n4726, S => n2250, Z => n5037);
   U632 : MUX2_X1 port map( A => n5870, B => n5869, S => n1571, Z => n1112);
   U633 : OR2_X1 port map( A1 => n5697, A2 => n5683, ZN => n5681);
   U634 : MUX2_X1 port map( A => n6395, B => n6394, S => n7973, Z => n6505);
   U635 : OR2_X2 port map( A1 => n4499, A2 => n4463, ZN => n4496);
   U637 : AND3_X1 port map( A1 => n4834, A2 => n4844, A3 => n4831, ZN => n474);
   U638 : OAI21_X1 port map( B1 => n4594, B2 => n4860, A => n4865, ZN => n475);
   U639 : INV_X1 port map( A => n5723, ZN => n476);
   U640 : OAI211_X1 port map( C1 => n648, C2 => n1834, A => n5974, B => n690, 
                           ZN => n477);
   U641 : MUX2_X2 port map( A => n5516, B => n5515, S => n2245, Z => n5723);
   U642 : XNOR2_X1 port map( A => n5041, B => n4933, ZN => n5042);
   U643 : MUX2_X2 port map( A => n5258, B => n5257, S => n2129, Z => n5773);
   U644 : MUX2_X2 port map( A => n6269, B => n6270, S => n859, Z => n6403);
   U645 : NAND2_X1 port map( A1 => n1325, A2 => n6369, ZN => n478);
   U646 : NAND2_X1 port map( A1 => n1326, A2 => n1702, ZN => n479);
   U647 : NAND2_X1 port map( A1 => n479, A2 => n478, ZN => n1324);
   U648 : NAND2_X1 port map( A1 => n1754, A2 => n1121, ZN => n480);
   U649 : NAND2_X1 port map( A1 => n1755, A2 => n2244, ZN => n481);
   U650 : NAND2_X1 port map( A1 => n480, A2 => n481, ZN => n551);
   U651 : AND2_X1 port map( A1 => n4514, A2 => n4756, ZN => n1060);
   U652 : INV_X1 port map( A => n1060, ZN => n4609);
   U653 : NAND2_X1 port map( A1 => n6653, A2 => n1637, ZN => n482);
   U654 : OAI211_X1 port map( C1 => n4644, C2 => n792, A => n4642, B => n4643, 
                           ZN => n483);
   U655 : MUX2_X2 port map( A => n5463, B => n5462, S => n2246, Z => n8142);
   U657 : OR2_X1 port map( A1 => n4593, A2 => n804, ZN => n4905);
   U658 : OR2_X1 port map( A1 => n2163, A2 => n5812, ZN => n484);
   U659 : MUX2_X2 port map( A => n4782, B => n4781, S => n804, Z => n4937);
   U660 : NAND2_X1 port map( A1 => n17180, A2 => n1465, ZN => n485);
   U661 : OR2_X1 port map( A1 => n5019, A2 => n5020, ZN => n486);
   U662 : NAND2_X1 port map( A1 => n5021, A2 => n486, ZN => n4927);
   U663 : MUX2_X1 port map( A => n5133, B => n5132, S => n799, Z => n5458);
   U664 : XNOR2_X1 port map( A => n487, B => n488, ZN => n1051);
   U665 : XNOR2_X1 port map( A => n6326, B => n6323, ZN => n487);
   U666 : AND2_X1 port map( A1 => n886, A2 => n6185, ZN => n488);
   U667 : OR2_X2 port map( A1 => n4496, A2 => n4464, ZN => n4493);
   U669 : AND2_X1 port map( A1 => n1704, A2 => n4667, ZN => n489);
   U670 : NAND2_X1 port map( A1 => n5177, A2 => n6890, ZN => n490);
   U671 : NAND2_X1 port map( A1 => n490, A2 => n217, ZN => n5276);
   U672 : INV_X1 port map( A => n8208, ZN => n2262);
   U673 : XNOR2_X1 port map( A => n874, B => n491, ZN => n7408);
   U674 : AND2_X1 port map( A1 => n1021, A2 => n7405, ZN => n491);
   U675 : XNOR2_X1 port map( A => n492, B => n7449, ZN => n1881);
   U676 : NAND2_X1 port map( A1 => n1018, A2 => n1017, ZN => n492);
   U677 : AND2_X1 port map( A1 => n4875, A2 => n2250, ZN => n1386);
   U678 : CLKBUF_X1 port map( A => n550, Z => n1552);
   U679 : OAI22_X1 port map( A1 => n2191, A2 => n17195, B1 => n2230, B2 => n494
                           , ZN => n493);
   U680 : BUF_X1 port map( A => n4558, Z => n494);
   U681 : XNOR2_X1 port map( A => n6773, B => n6765, ZN => n5840);
   U682 : OR2_X2 port map( A1 => n4489, A2 => n4466, ZN => n4485);
   U684 : NOR2_X1 port map( A1 => n979, A2 => n342, ZN => n6090);
   U685 : AND2_X1 port map( A1 => n5706, A2 => n5707, ZN => n495);
   U686 : MUX2_X2 port map( A => n1661, B => n1662, S => n7771, Z => n1660);
   U687 : NAND2_X1 port map( A1 => n5177, A2 => n6890, ZN => n496);
   U688 : NAND2_X1 port map( A1 => n5176, A2 => n2247, ZN => n497);
   U689 : NAND2_X1 port map( A1 => n496, A2 => n497, ZN => n678);
   U690 : OR2_X1 port map( A1 => n5045, A2 => n4967, ZN => n498);
   U691 : NAND2_X1 port map( A1 => n498, A2 => n5048, ZN => n4968);
   U692 : MUX2_X1 port map( A => n5396, B => n5395, S => n2245, Z => n5638);
   U693 : XNOR2_X1 port map( A => n499, B => n5769, ZN => n5267);
   U694 : XOR2_X1 port map( A => n5774, B => n5773, Z => n499);
   U695 : XNOR2_X1 port map( A => n500, B => n7439, ZN => n7448);
   U696 : XOR2_X1 port map( A => n7437, B => n7438, Z => n500);
   U697 : MUX2_X1 port map( A => n5403, B => n5404, S => n1092, Z => n5735);
   U698 : MUX2_X1 port map( A => n5565, B => n5564, S => n2244, Z => n5833);
   U699 : MUX2_X2 port map( A => n5044, B => n5043, S => n2248, Z => n778);
   U700 : NAND2_X1 port map( A1 => n839, A2 => n7705, ZN => n1614);
   U701 : INV_X1 port map( A => n699, ZN => n501);
   U702 : OR2_X1 port map( A1 => n8129, A2 => n5456, ZN => n5709);
   U703 : XOR2_X1 port map( A => n1379, B => n5101, Z => n5103);
   U704 : OR2_X2 port map( A1 => n4485, A2 => n4467, ZN => n4481);
   U705 : CLKBUF_X1 port map( A => n6350, Z => n950);
   U706 : XNOR2_X1 port map( A => n6745, B => n6710, ZN => n5792);
   U707 : MUX2_X1 port map( A => n5663, B => n5662, S => n2244, Z => n5924);
   U708 : CLKBUF_X1 port map( A => n8163, Z => n1149);
   U709 : MUX2_X2 port map( A => n5403, B => n5404, S => n1092, Z => n929);
   U710 : MUX2_X2 port map( A => n4720, B => n4719, S => n2250, Z => n4976);
   U711 : AND3_X1 port map( A1 => n502, A2 => n2249, A3 => n5029, ZN => n5035);
   U712 : NAND2_X1 port map( A1 => n1024, A2 => n4968, ZN => n502);
   U713 : NAND2_X1 port map( A1 => n5273, A2 => n5162, ZN => n503);
   U714 : NAND3_X1 port map( A1 => n658, A2 => n659, A3 => n5203, ZN => n505);
   U715 : MUX2_X1 port map( A => n5377, B => n5378, S => n936, Z => n5617);
   U716 : AND3_X1 port map( A1 => n1079, A2 => n1080, A3 => n6071, ZN => n506);
   U717 : MUX2_X2 port map( A => n5677, B => n5678, S => n1351, Z => n1275);
   U718 : MUX2_X2 port map( A => n2165, B => n2164, S => n1369, Z => n2163);
   U719 : MUX2_X2 port map( A => n5493, B => n5494, S => n1092, Z => n942);
   U720 : XNOR2_X1 port map( A => n507, B => n5690, ZN => n2165);
   U721 : XOR2_X1 port map( A => n1157, B => n5537, Z => n507);
   U722 : MUX2_X2 port map( A => n4755, B => n4754, S => n2250, Z => n5052);
   U723 : CLKBUF_X1 port map( A => n6157, Z => n508);
   U724 : INV_X1 port map( A => n731, ZN => n509);
   U726 : MUX2_X1 port map( A => n5474, B => n5475, S => n700, Z => n510);
   U727 : MUX2_X2 port map( A => n1754, B => n1755, S => n2244, Z => n1753);
   U728 : CLKBUF_X1 port map( A => n1271, Z => n511);
   U729 : NAND2_X1 port map( A1 => n1573, A2 => n1572, ZN => n512);
   U731 : NAND3_X1 port map( A1 => n4840, A2 => n4838, A3 => n4839, ZN => n513)
                           ;
   U732 : MUX2_X2 port map( A => n5428, B => n5427, S => n2245, Z => n790);
   U734 : XNOR2_X1 port map( A => n5058, B => n5062, ZN => n5063);
   U735 : XNOR2_X1 port map( A => n5643, B => n514, ZN => n5651);
   U736 : XNOR2_X1 port map( A => n5638, B => n5637, ZN => n514);
   U737 : AND2_X1 port map( A1 => n4741, A2 => n4743, ZN => n515);
   U738 : AND3_X1 port map( A1 => n4670, A2 => n4742, A3 => n515, ZN => n837);
   U739 : OR2_X1 port map( A1 => n4708, A2 => n4682, ZN => n516);
   U740 : NAND2_X1 port map( A1 => n516, A2 => n4711, ZN => n4683);
   U741 : NAND2_X1 port map( A1 => n937, A2 => n938, ZN => n517);
   U742 : NAND2_X1 port map( A1 => n937, A2 => n938, ZN => n518);
   U743 : CLKBUF_X1 port map( A => n8276, Z => n519);
   U744 : NAND2_X1 port map( A1 => n937, A2 => n938, ZN => n6904);
   U745 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n147, ZN => n520);
   U746 : INV_X1 port map( A => n520, ZN => n521);
   U747 : OAI22_X1 port map( A1 => n2138, A2 => n2184, B1 => n2238, B2 => n2182
                           , ZN => n5919);
   U748 : INV_X1 port map( A => n6646, ZN => n6681);
   U749 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n170, ZN => n522);
   U750 : INV_X1 port map( A => n522, ZN => n523);
   U751 : INV_X1 port map( A => n7453, ZN => n1717);
   U752 : INV_X1 port map( A => n7465, ZN => n1726);
   U753 : INV_X1 port map( A => n509, ZN => n524);
   U754 : INV_X1 port map( A => n509, ZN => n525);
   U755 : INV_X1 port map( A => n509, ZN => n526);
   U756 : INV_X1 port map( A => n509, ZN => n527);
   U757 : INV_X1 port map( A => n6231, ZN => n528);
   U758 : MUX2_X1 port map( A => n271, B => n350, S => n526, Z => n6231);
   U759 : INV_X1 port map( A => n7446, ZN => n763);
   U760 : INV_X1 port map( A => n7022, ZN => n1630);
   U761 : NAND2_X1 port map( A1 => n530, A2 => n5734, ZN => n5646);
   U762 : INV_X1 port map( A => n5735, ZN => n530);
   U763 : OAI211_X1 port map( C1 => n5535, C2 => n5537, A => n5681, B => n5495,
                           ZN => n5496);
   U764 : AND2_X1 port map( A1 => n5539, A2 => n1041, ZN => n5725);
   U765 : OAI21_X1 port map( B1 => n1789, B2 => n17208, A => n6150, ZN => n6165
                           );
   U766 : AOI22_X1 port map( A1 => n531, A2 => n6325, B1 => n6185, B2 => n886, 
                           ZN => n532);
   U767 : INV_X1 port map( A => n743, ZN => n531);
   U768 : INV_X1 port map( A => n532, ZN => n6186);
   U769 : MUX2_X1 port map( A => n5133, B => n5132, S => n799, Z => n1170);
   U771 : XNOR2_X1 port map( A => n5672, B => n5673, ZN => n1473);
   U772 : XNOR2_X1 port map( A => n791, B => n5664, ZN => n5668);
   U773 : OAI21_X1 port map( B1 => n5150, B2 => n5151, A => n5149, ZN => n5152)
                           ;
   U774 : AOI22_X1 port map( A1 => n17197, A2 => n5162, B1 => n8150, B2 => 
                           n8163, ZN => n5178);
   U775 : AOI22_X1 port map( A1 => n5388, A2 => n5398, B1 => n5400, B2 => n5270
                           , ZN => n5389);
   U776 : OAI211_X1 port map( C1 => n1822, C2 => n5431, A => n5429, B => n5430,
                           ZN => n5406);
   U777 : NAND2_X1 port map( A1 => n4556, A2 => n4452, ZN => n4641);
   U778 : AOI21_X1 port map( B1 => n5883, B2 => n5882, A => n1885, ZN => n5884)
                           ;
   U779 : OAI22_X1 port map( A1 => n630, A2 => n6210, B1 => n995, B2 => n6328, 
                           ZN => n6324);
   U780 : XNOR2_X1 port map( A => n4937, B => n5084, ZN => n5087);
   U781 : AOI22_X1 port map( A1 => n5954, A2 => n5959, B1 => n5812, B2 => n1290
                           , ZN => n5956);
   U782 : OR2_X1 port map( A1 => n2163, A2 => n5812, ZN => n1492);
   U783 : XNOR2_X1 port map( A => n5595, B => n1088, ZN => n5597);
   U784 : XNOR2_X1 port map( A => n5235, B => n5236, ZN => n4982);
   U785 : AND2_X1 port map( A1 => n4556, A2 => n1215, ZN => n1891);
   U786 : XNOR2_X1 port map( A => n4570, B => n1760, ZN => n4440);
   U787 : OAI22_X1 port map( A1 => n6194, A2 => n6195, B1 => n6241, B2 => n6223
                           , ZN => n6235);
   U788 : XNOR2_X1 port map( A => n664, B => n5548, ZN => n1430);
   U789 : XNOR2_X1 port map( A => n6139, B => n6012, ZN => n1596);
   U790 : OAI22_X1 port map( A1 => n4633, A2 => n4829, B1 => n4825, B2 => n4653
                           , ZN => n4806);
   U791 : AND2_X1 port map( A1 => n5872, A2 => n5871, ZN => n5874);
   U792 : OAI21_X1 port map( B1 => n262, B2 => n979, A => n6075, ZN => n6077);
   U793 : NAND3_X1 port map( A1 => n4839, A2 => n4838, A3 => n4840, ZN => n4946
                           );
   U794 : OAI21_X1 port map( B1 => n6168, B2 => n6151, A => n6006, ZN => n6007)
                           ;
   U795 : AOI21_X1 port map( B1 => n5689, B2 => n5688, A => n5687, ZN => n5690)
                           ;
   U796 : XNOR2_X1 port map( A => n5945, B => n5944, ZN => n5946);
   U797 : OR2_X1 port map( A1 => n1275, A2 => n5955, ZN => n824);
   U799 : XNOR2_X1 port map( A => n5895, B => n876, ZN => n5902);
   U800 : XNOR2_X1 port map( A => n5905, B => n1538, ZN => n5912);
   U801 : MUX2_X1 port map( A => n5626, B => n5627, S => n6912, Z => n933);
   U802 : AND2_X1 port map( A1 => n5412, A2 => n5413, ZN => n5416);
   U803 : NOR2_X1 port map( A1 => n6114, A2 => n6115, ZN => n6020);
   U804 : OAI22_X1 port map( A1 => n533, A2 => n534, B1 => n5298, B2 => n5348, 
                           ZN => n5210);
   U805 : INV_X1 port map( A => n1365, ZN => n533);
   U806 : INV_X1 port map( A => n5209, ZN => n534);
   U807 : OAI211_X1 port map( C1 => n1514, C2 => n5807, A => n5892, B => n5893,
                           ZN => n5871);
   U808 : OAI211_X1 port map( C1 => n5576, C2 => n1809, A => n5575, B => n5574,
                           ZN => n5577);
   U809 : NAND3_X1 port map( A1 => n8165, A2 => n5272, A3 => n5460, ZN => n5467
                           );
   U810 : MUX2_X1 port map( A => n5454, B => n5455, S => n6920, Z => n535);
   U811 : INV_X1 port map( A => n535, ZN => n5694);
   U812 : NAND2_X1 port map( A1 => n824, A2 => n823, ZN => n1623);
   U813 : MUX2_X1 port map( A => n5704, B => n5705, S => n6912, Z => n536);
   U814 : INV_X1 port map( A => n536, ZN => n8257);
   U815 : OAI22_X1 port map( A1 => n537, A2 => n538, B1 => n6529, B2 => n6530, 
                           ZN => n6481);
   U816 : INV_X1 port map( A => n721, ZN => n537);
   U817 : INV_X1 port map( A => n6479, ZN => n538);
   U818 : XNOR2_X1 port map( A => n6497, B => n6490, ZN => n1468);
   U819 : OAI21_X1 port map( B1 => n6471, B2 => n6473, A => n6447, ZN => n6535)
                           ;
   U820 : AND2_X1 port map( A1 => n5675, A2 => n1089, ZN => n539);
   U821 : INV_X1 port map( A => n539, ZN => n1382);
   U822 : AOI22_X1 port map( A1 => n5291, A2 => n1033, B1 => n540, B2 => n5373,
                           ZN => n694);
   U823 : INV_X1 port map( A => n1370, ZN => n540);
   U824 : NAND2_X1 port map( A1 => n5052, A2 => n5053, ZN => n4964);
   U825 : OR2_X1 port map( A1 => n793, A2 => n4943, ZN => n5155);
   U826 : OAI211_X1 port map( C1 => n1064, C2 => n5072, A => n5073, B => n923, 
                           ZN => n4917);
   U827 : OAI22_X1 port map( A1 => n830, A2 => n2198, B1 => n2195, B2 => n7249,
                           ZN => n4453);
   U828 : NOR2_X1 port map( A1 => n541, A2 => n8180, ZN => n1002);
   U829 : INV_X1 port map( A => n1875, ZN => n541);
   U830 : MUX2_X1 port map( A => n4267, B => n542, S => i_S1, Z => n7688);
   U831 : OAI21_X1 port map( B1 => n1212, B2 => n5868, A => n5866, ZN => n5828)
                           ;
   U832 : OAI211_X1 port map( C1 => n5535, C2 => n5679, A => n5534, B => n5688,
                           ZN => n5536);
   U833 : XOR2_X1 port map( A => n5353, B => n5352, Z => n5354);
   U834 : OAI21_X1 port map( B1 => n7012, B2 => n7032, A => n7011, ZN => n7029)
                           ;
   U835 : XNOR2_X1 port map( A => n892, B => n6022, ZN => n6105);
   U836 : OAI21_X1 port map( B1 => n1445, B2 => n5990, A => n713, ZN => n5830);
   U837 : OAI211_X1 port map( C1 => n1567, C2 => n5145, A => n543, B => n4941, 
                           ZN => n5164);
   U838 : INV_X1 port map( A => n4911, ZN => n543);
   U839 : CLKBUF_X1 port map( A => CU_I_n108, Z => n544);
   U840 : INV_X1 port map( A => n2131, ZN => n545);
   U842 : XNOR2_X1 port map( A => n17168, B => n6016, ZN => n1296);
   U843 : OAI21_X1 port map( B1 => n4594, B2 => n4860, A => n4865, ZN => n1569)
                           ;
   U844 : OR2_X1 port map( A1 => n1132, A2 => n6619, ZN => n6612);
   U845 : BUF_X2 port map( A => n8276, Z => n2270);
   U847 : OAI211_X1 port map( C1 => n17195, C2 => n216, A => n4554, B => n4553,
                           ZN => n546);
   U849 : AND2_X1 port map( A1 => n4439, A2 => n4440, ZN => n548);
   U850 : AND2_X1 port map( A1 => n4439, A2 => n4440, ZN => n2167);
   U851 : OR2_X1 port map( A1 => n5821, A2 => n5920, ZN => n5913);
   U852 : XNOR2_X1 port map( A => n7411, B => n7410, ZN => n549);
   U853 : MUX2_X2 port map( A => n7408, B => n7409, S => n859, Z => n7410);
   U854 : OAI211_X1 port map( C1 => n807, C2 => n4447, A => n4446, B => n4445, 
                           ZN => n550);
   U856 : MUX2_X1 port map( A => n5120, B => n5119, S => n2248, Z => n5476);
   U858 : NOR3_X1 port map( A1 => n8204, A2 => n8280, A3 => n2262, ZN => n554);
   U862 : XNOR2_X1 port map( A => n1747, B => n7465, ZN => n569);
   U863 : AND2_X1 port map( A1 => n6080, A2 => n1340, ZN => n557);
   U864 : XOR2_X1 port map( A => n5638, B => n5637, Z => n558);
   U865 : MUX2_X1 port map( A => n6239, B => n6240, S => n859, Z => n6371);
   U866 : MUX2_X2 port map( A => n1757, B => n1756, S => n6369, Z => n1133);
   U867 : MUX2_X1 port map( A => n1757, B => n1756, S => n6369, Z => n1132);
   U868 : INV_X1 port map( A => n7440, ZN => n559);
   U869 : INV_X1 port map( A => n1035, ZN => n7440);
   U870 : AND2_X1 port map( A1 => n6812, A2 => n6811, ZN => n1035);
   U871 : OAI21_X1 port map( B1 => n6733, B2 => n6736, A => n6712, ZN => n560);
   U872 : XNOR2_X1 port map( A => n6296, B => n6202, ZN => n561);
   U873 : XNOR2_X1 port map( A => n1882, B => n562, ZN => n7468);
   U874 : AND2_X1 port map( A1 => n751, A2 => n752, ZN => n563);
   U875 : NAND2_X1 port map( A1 => n886, A2 => n6185, ZN => n564);
   U877 : NAND2_X1 port map( A1 => n650, A2 => n651, ZN => n566);
   U878 : NAND2_X1 port map( A1 => n860, A2 => n861, ZN => n567);
   U880 : XNOR2_X1 port map( A => n569, B => n7016, ZN => n7017);
   U881 : MUX2_X1 port map( A => n5930, B => n5931, S => n1584, Z => n2159);
   U882 : NAND2_X1 port map( A1 => n6021, A2 => n1304, ZN => n571);
   U884 : MUX2_X1 port map( A => n6368, B => n6367, S => n986, Z => n6491);
   U885 : OAI21_X1 port map( B1 => n6599, B2 => n6598, A => n469, ZN => n572);
   U886 : INV_X2 port map( A => n2232, ZN => n2229);
   U887 : OAI21_X1 port map( B1 => n1155, B2 => n703, A => n550, ZN => n573);
   U888 : NAND2_X1 port map( A1 => n4444, A2 => n4443, ZN => n8208);
   U889 : XNOR2_X1 port map( A => n575, B => n7434, ZN => n7435);
   U890 : XOR2_X1 port map( A => n7423, B => n7424, Z => n575);
   U891 : CLKBUF_X1 port map( A => n1466, Z => n576);
   U892 : XNOR2_X1 port map( A => n7379, B => n7378, ZN => n6951);
   U893 : MUX2_X1 port map( A => n6799, B => n6798, S => n986, Z => n1415);
   U894 : INV_X1 port map( A => n529, ZN => n986);
   U895 : CLKBUF_X1 port map( A => n4645, Z => n577);
   U896 : CLKBUF_X1 port map( A => n1082, Z => n1681);
   U897 : MUX2_X2 port map( A => n1724, B => n1725, S => n4436, Z => n578);
   U898 : MUX2_X1 port map( A => n1724, B => n1725, S => n4436, Z => n1723);
   U899 : XNOR2_X1 port map( A => n996, B => n6589, ZN => n580);
   U900 : MUX2_X1 port map( A => n5435, B => n5434, S => n2246, Z => n1089);
   U901 : OAI22_X1 port map( A1 => n731, A2 => n4442, B1 => n4441, B2 => n838, 
                           ZN => n581);
   U902 : CLKBUF_X1 port map( A => n6685, Z => n582);
   U903 : CLKBUF_X1 port map( A => n6326, Z => n583);
   U904 : CLKBUF_X1 port map( A => n5310, Z => n584);
   U905 : MUX2_X1 port map( A => n1751, B => n1752, S => n1702, Z => n1750);
   U906 : NAND2_X1 port map( A1 => n5912, A2 => n1584, ZN => n586);
   U907 : NAND2_X1 port map( A1 => n901, A2 => n1138, ZN => n587);
   U908 : OAI211_X1 port map( C1 => n1514, C2 => n5807, A => n5893, B => n5892,
                           ZN => n588);
   U909 : OAI222_X1 port map( A1 => n6848, A2 => n1449, B1 => n1862, B2 => 
                           n6847, C1 => n1862, C2 => n6846, ZN => n589);
   U910 : XNOR2_X1 port map( A => n1763, B => n7453, ZN => n607);
   U911 : AND2_X1 port map( A1 => n1548, A2 => n1235, ZN => n590);
   U912 : XNOR2_X1 port map( A => n1416, B => n6344, ZN => n1036);
   U913 : XNOR2_X1 port map( A => n1682, B => n5805, ZN => n591);
   U914 : NAND2_X1 port map( A1 => n7061, A2 => n594, ZN => n592);
   U915 : NAND2_X1 port map( A1 => n593, A2 => n592, ZN => n1808);
   U916 : AND2_X1 port map( A1 => n7471, A2 => n7069, ZN => n594);
   U917 : NAND2_X1 port map( A1 => n7013, A2 => n1488, ZN => n595);
   U918 : OAI22_X1 port map( A1 => n1146, A2 => n6858, B1 => n2270, B2 => n809,
                           ZN => n596);
   U920 : BUF_X1 port map( A => n4547, Z => n761);
   U921 : INV_X1 port map( A => n548, ZN => n2142);
   U922 : INV_X1 port map( A => n1710, ZN => n598);
   U923 : NAND2_X1 port map( A1 => n6821, A2 => n904, ZN => n599);
   U924 : OAI22_X1 port map( A1 => n2244, A2 => n5616, B1 => n5615, B2 => n6912
                           , ZN => n600);
   U925 : MUX2_X1 port map( A => n5516, B => n5515, S => n2245, Z => n601);
   U926 : NOR2_X1 port map( A1 => n6252, A2 => n1395, ZN => n602);
   U927 : XNOR2_X1 port map( A => n1156, B => n1777, ZN => n604);
   U928 : OAI211_X1 port map( C1 => n5979, C2 => n5978, A => n477, B => n5977, 
                           ZN => n605);
   U929 : NAND2_X1 port map( A1 => n6460, A2 => n6344, ZN => n606);
   U930 : OAI222_X1 port map( A1 => n2132, A2 => n8102, B1 => n8090, B2 => 
                           n8089, C1 => DataPath_ALUhw_SHIFTER_HW_n600, C2 => 
                           n8088, ZN => n8096);
   U931 : XNOR2_X1 port map( A => n607, B => n7245, ZN => n1749);
   U932 : BUF_X1 port map( A => n4884, Z => n608);
   U933 : INV_X2 port map( A => n7110, ZN => n804);
   U934 : BUF_X4 port map( A => n2155, Z => n2250);
   U935 : BUF_X1 port map( A => n804, Z => n2251);
   U936 : CLKBUF_X1 port map( A => n2250, Z => n2129);
   U937 : INV_X1 port map( A => n804, ZN => n818);
   U938 : CLKBUF_X1 port map( A => n1810, Z => n1219);
   U939 : INV_X1 port map( A => n6388, ZN => n610);
   U940 : NAND2_X1 port map( A1 => n6190, A2 => n633, ZN => n611);
   U941 : OR2_X1 port map( A1 => n6950, A2 => n6949, ZN => n612);
   U942 : NAND2_X1 port map( A1 => n612, A2 => n6948, ZN => n7377);
   U943 : MUX2_X1 port map( A => n5363, B => n5362, S => n2246, Z => n613);
   U944 : MUX2_X1 port map( A => n5363, B => n5362, S => n2246, Z => n5600);
   U945 : XNOR2_X1 port map( A => n451, B => n614, ZN => n5596);
   U946 : AND2_X1 port map( A1 => n5552, A2 => n1310, ZN => n614);
   U948 : CLKBUF_X1 port map( A => n6686, Z => n615);
   U949 : AND3_X1 port map( A1 => n1593, A2 => n6066, A3 => n1432, ZN => n617);
   U950 : NAND2_X1 port map( A1 => n6489, A2 => n927, ZN => n618);
   U951 : NAND2_X1 port map( A1 => n672, A2 => n673, ZN => n619);
   U952 : NAND2_X1 port map( A1 => n4661, A2 => n1529, ZN => n621);
   U953 : AND2_X1 port map( A1 => n910, A2 => n4923, ZN => n622);
   U954 : OR2_X1 port map( A1 => n5341, A2 => n5303, ZN => n623);
   U955 : NAND2_X1 port map( A1 => n623, A2 => n5344, ZN => n5337);
   U956 : NOR2_X1 port map( A1 => n1566, A2 => n321, ZN => n4602);
   U957 : CLKBUF_X1 port map( A => n6327, Z => n624);
   U958 : INV_X1 port map( A => n1422, ZN => n7253);
   U959 : MUX2_X1 port map( A => n1052, B => n1051, S => n1407, Z => n1050);
   U960 : AND2_X1 port map( A1 => n1132, A2 => n6574, ZN => n625);
   U961 : AND2_X1 port map( A1 => n6656, A2 => n1185, ZN => n626);
   U962 : OR2_X1 port map( A1 => n5815, A2 => n8258, ZN => n627);
   U963 : NAND2_X1 port map( A1 => n5814, A2 => n627, ZN => n5959);
   U964 : OR2_X1 port map( A1 => n996, A2 => n6589, ZN => n628);
   U966 : CLKBUF_X1 port map( A => n839, Z => n629);
   U967 : INV_X1 port map( A => n6329, ZN => n630);
   U968 : AND2_X1 port map( A1 => n724, A2 => n723, ZN => n632);
   U969 : OR2_X1 port map( A1 => n1003, A2 => n6267, ZN => n633);
   U970 : NAND2_X1 port map( A1 => n6190, A2 => n633, ZN => n1013);
   U971 : NAND2_X1 port map( A1 => n991, A2 => n735, ZN => n634);
   U972 : NAND3_X1 port map( A1 => n1366, A2 => n1367, A3 => n4971, ZN => n635)
                           ;
   U973 : OR2_X1 port map( A1 => n5019, A2 => n4974, ZN => n636);
   U974 : NAND2_X1 port map( A1 => n636, A2 => n5022, ZN => n4975);
   U975 : INV_X1 port map( A => n4543, ZN => n637);
   U976 : OR2_X1 port map( A1 => n1416, A2 => n6344, ZN => n6400);
   U977 : OR2_X1 port map( A1 => n5928, A2 => n5925, ZN => n638);
   U978 : NAND2_X1 port map( A1 => n638, A2 => n5926, ZN => n5721);
   U979 : XNOR2_X1 port map( A => n933, B => n5896, ZN => n1272);
   U980 : MUX2_X1 port map( A => n1662, B => n1661, S => n6594, Z => n1536);
   U981 : MUX2_X1 port map( A => n6614, B => n6615, S => n6495, Z => n6677);
   U982 : BUF_X1 port map( A => n855, Z => n1007);
   U983 : XNOR2_X1 port map( A => n5349, B => n5299, ZN => n5352);
   U984 : NAND2_X1 port map( A1 => n6337, A2 => n1489, ZN => n640);
   U986 : OAI22_X1 port map( A1 => n6209, A2 => n244, B1 => n995, B2 => n6328, 
                           ZN => n642);
   U987 : XNOR2_X1 port map( A => n6922, B => n6903, ZN => n6934);
   U988 : INV_X2 port map( A => n252, ZN => n2204);
   U989 : NAND2_X1 port map( A1 => n1004, A2 => n1005, ZN => n643);
   U990 : NAND2_X1 port map( A1 => n5567, A2 => n471, ZN => n644);
   U991 : NAND2_X1 port map( A1 => n5576, A2 => n233, ZN => n645);
   U993 : AND2_X1 port map( A1 => n4801, A2 => n312, ZN => n646);
   U994 : INV_X1 port map( A => n1934, ZN => n2216);
   U995 : MUX2_X1 port map( A => n6051, B => n6052, S => n750, Z => n1389);
   U997 : INV_X1 port map( A => n1317, ZN => n647);
   U998 : XOR2_X1 port map( A => n6403, B => n6406, Z => n1560);
   U999 : AND2_X1 port map( A1 => n5819, A2 => n1218, ZN => n648);
   U1000 : XNOR2_X1 port map( A => n4977, B => n5012, ZN => n5016);
   U1001 : CLKBUF_X1 port map( A => n5923, Z => n649);
   U1002 : NAND2_X1 port map( A1 => n1868, A2 => n6495, ZN => n650);
   U1003 : NAND2_X1 port map( A1 => n1869, A2 => n7835, ZN => n651);
   U1004 : NAND2_X1 port map( A1 => n650, A2 => n651, ZN => n1867);
   U1005 : NAND2_X1 port map( A1 => n6380, A2 => n6379, ZN => n652);
   U1006 : AND2_X1 port map( A1 => n6338, A2 => n1486, ZN => n653);
   U1007 : CLKBUF_X1 port map( A => n5922, Z => n654);
   U1008 : NAND2_X1 port map( A1 => n221, A2 => n1556, ZN => n655);
   U1009 : BUF_X1 port map( A => n5969, Z => n656);
   U1010 : CLKBUF_X1 port map( A => n552, Z => n657);
   U1011 : XNOR2_X1 port map( A => n5507, B => n5514, ZN => n5515);
   U1012 : OR2_X1 port map( A1 => n5204, A2 => n5391, ZN => n658);
   U1013 : OR2_X1 port map( A1 => n437, A2 => n5269, ZN => n659);
   U1014 : NAND3_X1 port map( A1 => n658, A2 => n659, A3 => n5203, ZN => n5381)
                           ;
   U1015 : NAND2_X1 port map( A1 => n5698, A2 => n5707, ZN => n1321);
   U1016 : OR3_X1 port map( A1 => n1526, A2 => n1525, A3 => n1524, ZN => n5692)
                           ;
   U1017 : XOR2_X1 port map( A => n552, B => n5490, Z => n5491);
   U1018 : INV_X1 port map( A => n770, ZN => n661);
   U1019 : BUF_X1 port map( A => n1891, Z => n1730);
   U1020 : OR2_X1 port map( A1 => n4534, A2 => n4456, ZN => n4526);
   U1021 : NAND2_X1 port map( A1 => n5718, A2 => n1363, ZN => n662);
   U1022 : MUX2_X2 port map( A => n5428, B => n5427, S => n2245, Z => n791);
   U1023 : MUX2_X1 port map( A => n5474, B => n5475, S => n700, Z => n663);
   U1024 : MUX2_X1 port map( A => n5474, B => n5475, S => n700, Z => n8129);
   U1025 : XNOR2_X1 port map( A => n842, B => n669, ZN => n995);
   U1026 : MUX2_X1 port map( A => n6432, B => n6431, S => n986, Z => n6551);
   U1027 : MUX2_X1 port map( A => n5384, B => n5383, S => n2246, Z => n5628);
   U1028 : AND2_X1 port map( A1 => n1704, A2 => n1284, ZN => n665);
   U1029 : OR2_X1 port map( A1 => n5263, A2 => n5266, ZN => n666);
   U1030 : NAND2_X1 port map( A1 => n5259, A2 => n666, ZN => n5260);
   U1031 : NAND2_X1 port map( A1 => n7046, A2 => n1230, ZN => n667);
   U1032 : NAND2_X1 port map( A1 => n482, A2 => n1638, ZN => n668);
   U1033 : MUX2_X1 port map( A => n654, B => n649, S => n1731, Z => n669);
   U1034 : MUX2_X1 port map( A => n5922, B => n5923, S => n1211, Z => n670);
   U1035 : MUX2_X1 port map( A => n5493, B => n5494, S => n936, Z => n5698);
   U1036 : MUX2_X1 port map( A => n6174, B => n6173, S => n2266, Z => n6208);
   U1037 : NOR2_X1 port map( A1 => n2156, A2 => n512, ZN => n671);
   U1038 : NAND2_X1 port map( A1 => n6248, A2 => n859, ZN => n672);
   U1039 : NAND2_X1 port map( A1 => n6247, A2 => n881, ZN => n673);
   U1040 : NAND2_X1 port map( A1 => n672, A2 => n673, ZN => n958);
   U1041 : INV_X1 port map( A => n1407, ZN => n881);
   U1042 : OR2_X1 port map( A1 => n5233, A2 => n5236, ZN => n674);
   U1043 : NAND2_X1 port map( A1 => n674, A2 => n5229, ZN => n5230);
   U1044 : OR2_X1 port map( A1 => n4979, A2 => n4981, ZN => n675);
   U1045 : NAND2_X1 port map( A1 => n675, A2 => n4929, ZN => n5229);
   U1046 : OR2_X1 port map( A1 => n6737, A2 => n6736, ZN => n676);
   U1047 : NAND2_X1 port map( A1 => n676, A2 => n6735, ZN => n6878);
   U1048 : XNOR2_X1 port map( A => n17164, B => n6319, ZN => n914);
   U1049 : XNOR2_X1 port map( A => n780, B => n6440, ZN => n6443);
   U1051 : INV_X1 port map( A => n2142, ZN => n677);
   U1052 : OR2_X1 port map( A1 => n2156, A2 => n6132, ZN => n6125);
   U1053 : OR2_X1 port map( A1 => n6529, A2 => n6482, ZN => n679);
   U1054 : NAND2_X1 port map( A1 => n679, A2 => n6527, ZN => n6458);
   U1055 : NOR3_X1 port map( A1 => n6913, A2 => n447, A3 => n446, ZN => n1466);
   U1056 : AND2_X1 port map( A1 => n905, A2 => n4630, ZN => n680);
   U1057 : OR2_X1 port map( A1 => n4721, A2 => n4676, ZN => n681);
   U1058 : NAND2_X1 port map( A1 => n4724, A2 => n681, ZN => n4677);
   U1059 : AND2_X1 port map( A1 => n4500, A2 => n4499, ZN => n682);
   U1060 : AND2_X1 port map( A1 => n1085, A2 => n1086, ZN => n683);
   U1061 : NAND2_X1 port map( A1 => n7387, A2 => n7386, ZN => n686);
   U1062 : NAND2_X1 port map( A1 => n684, A2 => n685, ZN => n687);
   U1063 : NAND2_X1 port map( A1 => n686, A2 => n687, ZN => n1900);
   U1064 : INV_X1 port map( A => n7387, ZN => n684);
   U1065 : INV_X1 port map( A => n7386, ZN => n685);
   U1066 : XNOR2_X1 port map( A => n5236, B => n5235, ZN => n688);
   U1067 : AND2_X1 port map( A1 => n905, A2 => n4630, ZN => n1617);
   U1068 : MUX2_X1 port map( A => n7385, B => n7384, S => n2267, Z => n7386);
   U1069 : MUX2_X2 port map( A => n5434, B => n5435, S => n1092, Z => n5672);
   U1070 : MUX2_X1 port map( A => n5143, B => n5142, S => n2248, Z => n8164);
   U1071 : INV_X1 port map( A => n5672, ZN => n689);
   U1072 : CLKBUF_X1 port map( A => n546, Z => n691);
   U1073 : NAND2_X1 port map( A1 => n6007, A2 => n1554, ZN => n692);
   U1074 : XNOR2_X1 port map( A => n5282, B => n5405, ZN => n798);
   U1075 : OR2_X2 port map( A1 => n4503, A2 => n4462, ZN => n4499);
   U1076 : OR2_X1 port map( A1 => n1594, A2 => n6488, ZN => n693);
   U1077 : NAND2_X1 port map( A1 => n6487, A2 => n693, ZN => n6499);
   U1078 : NOR2_X1 port map( A1 => n348, A2 => n1810, ZN => n6061);
   U1079 : OAI22_X1 port map( A1 => n809, A2 => n2195, B1 => n2270, B2 => n8045
                           , ZN => n4857);
   U1080 : NAND2_X1 port map( A1 => n668, A2 => n6668, ZN => n695);
   U1081 : NAND2_X1 port map( A1 => n1707, A2 => n1708, ZN => n696);
   U1083 : OR2_X1 port map( A1 => n4655, A2 => n4842, ZN => n4825);
   U1084 : OR2_X1 port map( A1 => n4930, A2 => n5006, ZN => n4998);
   U1086 : MUX2_X1 port map( A => n5143, B => n5142, S => n2248, Z => n699);
   U1087 : OR2_X1 port map( A1 => n6165, A2 => n6164, ZN => n701);
   U1088 : OR2_X1 port map( A1 => n6162, A2 => n6163, ZN => n702);
   U1089 : NAND3_X1 port map( A1 => n701, A2 => n702, A3 => n6161, ZN => n6166)
                           ;
   U1090 : AND2_X2 port map( A1 => n4429, A2 => n4430, ZN => n703);
   U1091 : AND2_X1 port map( A1 => n5819, A2 => n1218, ZN => n705);
   U1093 : MUX2_X1 port map( A => n5396, B => n5395, S => n2245, Z => n706);
   U1094 : NAND2_X1 port map( A1 => n5205, A2 => n887, ZN => n707);
   U1095 : OR2_X1 port map( A1 => n5608, A2 => n5609, ZN => n709);
   U1096 : NAND2_X1 port map( A1 => n5520, A2 => n709, ZN => n5598);
   U1097 : NAND2_X1 port map( A1 => n5911, A2 => n1571, ZN => n710);
   U1098 : MUX2_X2 port map( A => n4700, B => n4699, S => n2250, Z => n4981);
   U1100 : OR2_X1 port map( A1 => n6107, A2 => n6022, ZN => n1515);
   U1101 : AND2_X1 port map( A1 => n712, A2 => n7547, ZN => n1145);
   U1102 : NAND2_X1 port map( A1 => n7074, A2 => n7579, ZN => n712);
   U1103 : NAND2_X1 port map( A1 => n5828, A2 => n1483, ZN => n713);
   U1104 : CLKBUF_X1 port map( A => n1829, Z => n714);
   U1105 : XOR2_X1 port map( A => n715, B => n6372, Z => n6377);
   U1106 : XNOR2_X1 port map( A => n6371, B => n6374, ZN => n715);
   U1107 : NAND2_X1 port map( A1 => n991, A2 => n735, ZN => n716);
   U1108 : CLKBUF_X1 port map( A => n6094, Z => n1087);
   U1109 : XNOR2_X1 port map( A => n1178, B => n6200, ZN => n1248);
   U1110 : NAND2_X1 port map( A1 => n720, A2 => n719, ZN => n717);
   U1111 : NAND2_X1 port map( A1 => n6644, A2 => n940, ZN => n718);
   U1112 : AND2_X1 port map( A1 => n4828, A2 => n4829, ZN => n941);
   U1113 : NAND2_X1 port map( A1 => n6627, A2 => n7835, ZN => n719);
   U1114 : NAND2_X1 port map( A1 => n6628, A2 => n6495, ZN => n720);
   U1115 : NAND2_X1 port map( A1 => n720, A2 => n719, ZN => n1537);
   U1116 : NAND2_X1 port map( A1 => n245, A2 => n247, ZN => n1732);
   U1118 : MUX2_X2 port map( A => n6986, B => n6987, S => n6369, Z => n922);
   U1119 : OR2_X1 port map( A1 => n6534, A2 => n6480, ZN => n721);
   U1120 : NAND2_X1 port map( A1 => n6479, A2 => n721, ZN => n6528);
   U1121 : AND2_X1 port map( A1 => n6619, A2 => n1132, ZN => n722);
   U1122 : MUX2_X1 port map( A => n6423, B => n6424, S => n529, Z => n6534);
   U1123 : NAND2_X1 port map( A1 => n1640, A2 => n7771, ZN => n723);
   U1124 : NAND2_X1 port map( A1 => n1641, A2 => n6594, ZN => n724);
   U1125 : NAND2_X1 port map( A1 => n724, A2 => n723, ZN => n1639);
   U1127 : MUX2_X1 port map( A => n5421, B => n5420, S => n2245, Z => n726);
   U1128 : NOR2_X1 port map( A1 => n5105, A2 => n4949, ZN => n727);
   U1129 : INV_X1 port map( A => n727, ZN => n5191);
   U1130 : XNOR2_X1 port map( A => n17256, B => n5537, ZN => n728);
   U1131 : XOR2_X1 port map( A => n1293, B => n1777, Z => n729);
   U1132 : NAND2_X1 port map( A1 => n5092, A2 => n1587, ZN => n730);
   U1133 : INV_X1 port map( A => n838, ZN => n731);
   U1135 : BUF_X1 port map( A => CU_I_n107, Z => n838);
   U1137 : XNOR2_X1 port map( A => n5100, B => n4954, ZN => n5101);
   U1138 : NAND2_X1 port map( A1 => n732, A2 => n6267, ZN => n733);
   U1139 : NAND2_X1 port map( A1 => n6216, A2 => n733, ZN => n6259);
   U1140 : INV_X1 port map( A => n6262, ZN => n732);
   U1142 : OR2_X1 port map( A1 => n1867, A2 => n6682, ZN => n735);
   U1143 : OR2_X1 port map( A1 => n6355, A2 => n6354, ZN => n736);
   U1144 : NAND2_X1 port map( A1 => n6353, A2 => n736, ZN => n6450);
   U1145 : MUX2_X2 port map( A => n5981, B => n5982, S => n1211, Z => n1134);
   U1146 : XNOR2_X1 port map( A => n5782, B => n6747, ZN => n741);
   U1147 : XNOR2_X1 port map( A => n6253, B => n737, ZN => n6254);
   U1148 : XNOR2_X1 port map( A => n17172, B => n6252, ZN => n737);
   U1149 : MUX2_X1 port map( A => n5863, B => n5862, S => n1571, Z => n6024);
   U1150 : MUX2_X1 port map( A => n6322, B => n6321, S => n8229, Z => n6350);
   U1151 : NAND2_X1 port map( A1 => n5986, A2 => n1034, ZN => n738);
   U1152 : MUX2_X2 port map( A => n5025, B => n5024, S => n2248, Z => n5365);
   U1153 : MUX2_X1 port map( A => n6137, B => n6138, S => n750, Z => n739);
   U1154 : MUX2_X1 port map( A => n6137, B => n6138, S => n750, Z => n740);
   U1155 : XNOR2_X1 port map( A => n6706, B => n741, ZN => n5794);
   U1156 : CLKBUF_X1 port map( A => n8220, Z => n742);
   U1157 : AND2_X1 port map( A1 => n2163, A2 => n5957, ZN => n744);
   U1158 : XNOR2_X1 port map( A => n922, B => n7446, ZN => n6997);
   U1159 : NAND2_X1 port map( A1 => n6453, A2 => n986, ZN => n745);
   U1160 : NAND2_X1 port map( A1 => n6454, A2 => n754, ZN => n746);
   U1161 : NAND2_X1 port map( A1 => n745, A2 => n746, ZN => n6474);
   U1162 : INV_X1 port map( A => n7973, ZN => n754);
   U1163 : XNOR2_X1 port map( A => n7338, B => n7340, ZN => n6877);
   U1164 : AND2_X2 port map( A1 => n1531, A2 => n1649, ZN => n1647);
   U1165 : MUX2_X2 port map( A => n6331, B => n6330, S => n8229, Z => n8221);
   U1166 : OAI211_X2 port map( C1 => n6743, C2 => n6890, A => n6742, B => n6741
                           , ZN => n6922);
   U1167 : OR2_X1 port map( A1 => n933, A2 => n5807, ZN => n5881);
   U1168 : XOR2_X1 port map( A => n6253, B => n1398, Z => n747);
   U1170 : XNOR2_X1 port map( A => n471, B => n5569, ZN => n748);
   U1171 : NAND2_X1 port map( A1 => n6111, A2 => n750, ZN => n751);
   U1172 : NAND2_X1 port map( A1 => n6110, A2 => n2266, ZN => n752);
   U1173 : NAND2_X1 port map( A1 => n751, A2 => n752, ZN => n868);
   U1174 : INV_X1 port map( A => n2266, ZN => n750);
   U1176 : NAND2_X1 port map( A1 => n6034, A2 => n2266, ZN => n755);
   U1177 : MUX2_X2 port map( A => n5268, B => n5267, S => n2247, Z => n5790);
   U1178 : AOI22_X1 port map( A1 => n338, A2 => n6069, B1 => n6094, B2 => n6090
                           , ZN => n757);
   U1179 : NAND2_X1 port map( A1 => n1175, A2 => n6681, ZN => n759);
   U1180 : NAND2_X1 port map( A1 => n758, A2 => n6646, ZN => n760);
   U1181 : NAND2_X1 port map( A1 => n760, A2 => n759, ZN => n1171);
   U1182 : INV_X1 port map( A => n1175, ZN => n758);
   U1183 : XNOR2_X1 port map( A => n567, B => n6797, ZN => n781);
   U1184 : NAND2_X1 port map( A1 => n5275, A2 => n5274, ZN => n762);
   U1185 : INV_X1 port map( A => n6483, ZN => n764);
   U1186 : CLKBUF_X1 port map( A => n953, Z => n765);
   U1187 : NAND2_X1 port map( A1 => n6825, A2 => n7771, ZN => n766);
   U1188 : XNOR2_X1 port map( A => n767, B => n768, ZN => n6315);
   U1189 : XNOR2_X1 port map( A => n6309, B => n739, ZN => n767);
   U1190 : NAND2_X1 port map( A1 => n6298, A2 => n242, ZN => n768);
   U1191 : NAND2_X1 port map( A1 => n965, A2 => n966, ZN => n769);
   U1192 : CLKBUF_X1 port map( A => n8280, Z => n770);
   U1193 : MUX2_X2 port map( A => n7278, B => n7277, S => n2265, Z => n7407);
   U1194 : INV_X1 port map( A => n2154, ZN => n771);
   U1196 : INV_X1 port map( A => n4896, ZN => n772);
   U1198 : CLKBUF_X1 port map( A => n1830, Z => n773);
   U1199 : INV_X1 port map( A => n4538, ZN => n774);
   U1200 : AND2_X1 port map( A1 => n5531, A2 => n5532, ZN => n775);
   U1201 : XNOR2_X1 port map( A => n6938, B => n6937, ZN => n6940);
   U1202 : MUX2_X1 port map( A => n4789, B => n4788, S => n2250, Z => n4960);
   U1204 : CLKBUF_X1 port map( A => n8204, Z => n777);
   U1205 : BUF_X1 port map( A => CU_I_n107, Z => n1302);
   U1206 : XNOR2_X1 port map( A => n4722, B => n4678, ZN => n4725);
   U1207 : INV_X1 port map( A => n4933, ZN => n779);
   U1208 : MUX2_X1 port map( A => n2259, B => n4495, S => n4463, Z => n4497);
   U1210 : XNOR2_X1 port map( A => n6795, B => n781, ZN => n6367);
   U1211 : MUX2_X2 port map( A => n6493, B => n6494, S => n6369, Z => n1159);
   U1212 : XNOR2_X1 port map( A => n17164, B => n6316, ZN => n6320);
   U1213 : XNOR2_X1 port map( A => n704, B => n5683, ZN => n1736);
   U1214 : AND2_X1 port map( A1 => n6018, A2 => n6017, ZN => n782);
   U1215 : INV_X1 port map( A => n850, ZN => n783);
   U1216 : AND2_X1 port map( A1 => n1241, A2 => n1240, ZN => n784);
   U1217 : NAND2_X1 port map( A1 => n6029, A2 => n806, ZN => n785);
   U1218 : NAND2_X1 port map( A1 => n1202, A2 => n4674, ZN => n786);
   U1219 : OR2_X1 port map( A1 => n6879, A2 => n6882, ZN => n787);
   U1220 : NAND2_X1 port map( A1 => n787, A2 => n6857, ZN => n7338);
   U1221 : INV_X1 port map( A => n1146, ZN => n788);
   U1223 : AND2_X1 port map( A1 => n1420, A2 => n7465, ZN => n789);
   U1224 : MUX2_X1 port map( A => n6229, B => n6230, S => n859, Z => n6366);
   U1225 : NAND3_X1 port map( A1 => n4568, A2 => n4569, A3 => n1355, ZN => n792
                           );
   U1226 : MUX2_X1 port map( A => n4888, B => n4887, S => n2250, Z => n793);
   U1227 : MUX2_X1 port map( A => n4888, B => n4887, S => n804, Z => n794);
   U1228 : OR2_X1 port map( A1 => n4694, A2 => n4688, ZN => n795);
   U1229 : NAND2_X1 port map( A1 => n795, A2 => n4697, ZN => n4689);
   U1230 : INV_X1 port map( A => n6706, ZN => n796);
   U1231 : INV_X1 port map( A => n2196, ZN => n797);
   U1232 : INV_X2 port map( A => n1374, ZN => n2196);
   U1233 : XNOR2_X1 port map( A => n798, B => n5419, ZN => n5420);
   U1234 : MUX2_X1 port map( A => DataPath_i_PIPLIN_B_5_port, B => 
                           DataPath_i_PIPLIN_IN2_5_port, S => n2152, Z => n799)
                           ;
   U1235 : XNOR2_X1 port map( A => n441, B => n800, ZN => n5435);
   U1236 : NAND2_X1 port map( A1 => n5430, A2 => n5429, ZN => n800);
   U1237 : BUF_X1 port map( A => i_S1, Z => n2148);
   U1238 : CLKBUF_X1 port map( A => n7298, Z => n1329);
   U1239 : OAI221_X1 port map( B1 => n1319, B2 => n4943, C1 => n1358, C2 => 
                           n1319, A => n5155, ZN => n802);
   U1240 : XNOR2_X1 port map( A => n5411, B => n803, ZN => n5421);
   U1241 : XNOR2_X1 port map( A => n5405, B => n5418, ZN => n803);
   U1242 : MUX2_X1 port map( A => n1640, B => n1641, S => n6594, Z => n839);
   U1243 : CLKBUF_X1 port map( A => n6582, Z => n805);
   U1244 : OR2_X1 port map( A1 => n1082, A2 => n6057, ZN => n806);
   U1245 : NAND2_X1 port map( A1 => n806, A2 => n6029, ZN => n6050);
   U1246 : INV_X1 port map( A => n4448, ZN => n807);
   U1247 : OR2_X1 port map( A1 => n6406, A2 => n6405, ZN => n808);
   U1248 : NAND2_X1 port map( A1 => n6404, A2 => n808, ZN => n6359);
   U1249 : MUX2_X1 port map( A => n810, B => n811, S => n547, Z => n809);
   U1250 : INV_X1 port map( A => n809, ZN => n1933);
   U1251 : INV_X2 port map( A => n1933, ZN => n2238);
   U1252 : MUX2_X1 port map( A => DataPath_i_PIPLIN_IN1_3_port, B => 
                           DataPath_i_PIPLIN_A_3_port, S => CU_I_n108, Z => 
                           n812);
   U1253 : INV_X1 port map( A => n812, ZN => n7624);
   U1254 : XNOR2_X1 port map( A => n7437, B => n7438, ZN => n814);
   U1255 : MUX2_X1 port map( A => n7017, B => n7018, S => n4436, Z => n1693);
   U1256 : OAI22_X1 port map( A1 => n771, A2 => n7285, B1 => n2147, B2 => n7284
                           , ZN => n8227);
   U1257 : INV_X1 port map( A => n17186, ZN => n815);
   U1258 : AND2_X1 port map( A1 => n5286, A2 => n843, ZN => n816);
   U1259 : OR2_X1 port map( A1 => n4528, A2 => n4857, ZN => n817);
   U1260 : INV_X1 port map( A => n834, ZN => n1146);
   U1261 : INV_X1 port map( A => n2155, ZN => n7110);
   U1262 : INV_X1 port map( A => n4557, ZN => n819);
   U1264 : OR2_X1 port map( A1 => n4776, A2 => n4777, ZN => n820);
   U1265 : NAND2_X1 port map( A1 => n4778, A2 => n820, ZN => n4608);
   U1266 : MUX2_X1 port map( A => n4748, B => n4747, S => n2250, Z => n4969);
   U1267 : NAND3_X1 port map( A1 => n5166, A2 => n5163, A3 => n1621, ZN => n821
                           );
   U1268 : INV_X1 port map( A => n6209, ZN => n822);
   U1269 : NAND2_X1 port map( A1 => n1275, A2 => n5955, ZN => n823);
   U1270 : OAI21_X1 port map( B1 => n7025, B2 => n1291, A => n595, ZN => n825);
   U1271 : OR2_X2 port map( A1 => n4512, A2 => n4460, ZN => n4508);
   U1272 : AND2_X1 port map( A1 => n6021, A2 => n1304, ZN => n826);
   U1273 : AND2_X1 port map( A1 => n4883, A2 => n4592, ZN => n827);
   U1275 : CLKBUF_X1 port map( A => n8199, Z => n829);
   U1276 : INV_X1 port map( A => n7109, ZN => n8181);
   U1277 : INV_X1 port map( A => n2149, ZN => n830);
   U1278 : BUF_X2 port map( A => n7318, Z => n2149);
   U1279 : AND3_X2 port map( A1 => n4549, A2 => n4548, A3 => n4452, ZN => n831)
                           ;
   U1280 : INV_X1 port map( A => n793, ZN => n832);
   U1281 : OAI211_X1 port map( C1 => n4817, C2 => n4818, A => n4816, B => n4815
                           , ZN => n833);
   U1282 : XOR2_X1 port map( A => n5135, B => n4941, Z => n1456);
   U1284 : XNOR2_X1 port map( A => n5006, B => n4930, ZN => n5009);
   U1285 : MUX2_X1 port map( A => DataPath_i_PIPLIN_IN1_5_port, B => 
                           DataPath_i_PIPLIN_A_5_port, S => CU_I_n108, Z => 
                           n834);
   U1286 : NAND2_X1 port map( A1 => n5788, A2 => n5791, ZN => n6707);
   U1287 : OR2_X2 port map( A1 => n837, A2 => n836, ZN => n4730);
   U1288 : NOR2_X1 port map( A1 => n435, A2 => n4671, ZN => n836);
   U1289 : MUX2_X2 port map( A => n4732, B => n4731, S => n804, Z => n4933);
   U1290 : OR2_X1 port map( A1 => n4728, A2 => n4729, ZN => n1054);
   U1291 : CLKBUF_X1 port map( A => n6442, Z => n840);
   U1292 : XNOR2_X1 port map( A => n6526, B => n6482, ZN => n1626);
   U1293 : NAND2_X1 port map( A1 => n4429, A2 => n4430, ZN => n841);
   U1294 : NOR2_X1 port map( A1 => n6166, A2 => n6167, ZN => n842);
   U1295 : NAND2_X1 port map( A1 => n4429, A2 => n4430, ZN => n6858);
   U1296 : OR2_X1 port map( A1 => n5498, A2 => n5499, ZN => n843);
   U1297 : NAND2_X1 port map( A1 => n843, A2 => n5286, ZN => n5398);
   U1298 : AND2_X2 port map( A1 => n6755, A2 => n6702, ZN => n1852);
   U1299 : MUX2_X1 port map( A => n1325, B => n1326, S => n1702, Z => n913);
   U1300 : NAND2_X1 port map( A1 => n987, A2 => n844, ZN => n6507);
   U1301 : AND2_X1 port map( A1 => n988, A2 => n845, ZN => n844);
   U1302 : INV_X1 port map( A => n6522, ZN => n845);
   U1303 : MUX2_X1 port map( A => n1051, B => n1052, S => n881, Z => n846);
   U1304 : XNOR2_X1 port map( A => n5170, B => n5169, ZN => n5177);
   U1305 : NAND3_X1 port map( A1 => n1025, A2 => n1026, A3 => n4962, ZN => n847
                           );
   U1306 : CLKBUF_X1 port map( A => n1360, Z => n848);
   U1307 : XNOR2_X1 port map( A => n849, B => n7425, ZN => n7436);
   U1308 : XOR2_X1 port map( A => n7423, B => n7424, Z => n849);
   U1309 : AND3_X1 port map( A1 => n1079, A2 => n1080, A3 => n6071, ZN => n973)
                           ;
   U1311 : INV_X1 port map( A => n6025, ZN => n851);
   U1312 : INV_X1 port map( A => n838, ZN => n2152);
   U1313 : INV_X1 port map( A => n1578, ZN => n852);
   U1314 : CLKBUF_X1 port map( A => n8221, Z => n853);
   U1315 : MUX2_X1 port map( A => n5862, B => n5863, S => n1731, Z => n1297);
   U1316 : NAND2_X1 port map( A1 => n1410, A2 => n6804, ZN => n854);
   U1317 : MUX2_X2 port map( A => n5777, B => n5776, S => n2247, Z => n6706);
   U1318 : NAND2_X1 port map( A1 => n5496, A2 => n1099, ZN => n856);
   U1319 : XNOR2_X1 port map( A => n1721, B => n857, ZN => n6148);
   U1320 : AND2_X1 port map( A1 => n5967, A2 => n1523, ZN => n857);
   U1321 : XOR2_X1 port map( A => n6311, B => n2158, Z => n6314);
   U1322 : OAI22_X1 port map( A1 => n1646, A2 => n6020, B1 => n1008, B2 => 
                           n6019, ZN => n858);
   U1323 : XNOR2_X1 port map( A => n7058, B => n7045, ZN => n1191);
   U1324 : NAND2_X1 port map( A1 => n6230, A2 => n859, ZN => n860);
   U1325 : NAND2_X1 port map( A1 => n6229, A2 => n8229, ZN => n861);
   U1326 : NAND2_X1 port map( A1 => n861, A2 => n860, ZN => n880);
   U1327 : INV_X1 port map( A => n8229, ZN => n859);
   U1328 : OR2_X1 port map( A1 => n1415, A2 => n6984, ZN => n7426);
   U1329 : MUX2_X1 port map( A => n6799, B => n6798, S => n986, Z => n862);
   U1330 : MUX2_X1 port map( A => n6799, B => n6798, S => n986, Z => n6983);
   U1331 : XNOR2_X1 port map( A => n7034, B => n863, ZN => n1701);
   U1332 : AND2_X1 port map( A1 => n6691, A2 => n1614, ZN => n863);
   U1333 : XNOR2_X1 port map( A => n893, B => n864, ZN => n5474);
   U1334 : XOR2_X1 port map( A => n17191, B => n5484, Z => n864);
   U1335 : XNOR2_X1 port map( A => n5422, B => n5426, ZN => n1038);
   U1336 : AND2_X1 port map( A1 => n5887, A2 => n5806, ZN => n865);
   U1337 : OR2_X1 port map( A1 => n1082, A2 => n6060, ZN => n866);
   U1338 : NAND2_X1 port map( A1 => n5995, A2 => n866, ZN => n6037);
   U1339 : OAI22_X1 port map( A1 => n2244, A2 => n5616, B1 => n5615, B2 => 
                           n6912, ZN => n867);
   U1341 : INV_X1 port map( A => n5797, ZN => n869);
   U1342 : OR2_X1 port map( A1 => n4679, A2 => n4681, ZN => n870);
   U1343 : NAND2_X1 port map( A1 => n870, A2 => n4617, ZN => n4710);
   U1344 : OR2_X1 port map( A1 => n5251, A2 => n5254, ZN => n871);
   U1345 : NAND2_X1 port map( A1 => n871, A2 => n5249, ZN => n5756);
   U1346 : OR2_X1 port map( A1 => n4688, A2 => n4690, ZN => n872);
   U1347 : NAND2_X1 port map( A1 => n872, A2 => n4620, ZN => n5218);
   U1348 : OR2_X1 port map( A1 => n4673, A2 => n4675, ZN => n873);
   U1349 : NAND2_X1 port map( A1 => n873, A2 => n4615, ZN => n4723);
   U1350 : XNOR2_X1 port map( A => n7398, B => n7397, ZN => n874);
   U1351 : OAI21_X1 port map( B1 => n6920, B2 => n5316, A => n5315, ZN => n875)
                           ;
   U1352 : MUX2_X2 port map( A => n7396, B => n7395, S => n2266, Z => n7397);
   U1353 : NAND2_X1 port map( A1 => n5892, A2 => n5893, ZN => n876);
   U1354 : OAI22_X1 port map( A1 => n7066, A2 => n7577, B1 => n433, B2 => n7062
                           , ZN => n877);
   U1355 : OR2_X1 port map( A1 => n4922, A2 => n5054, ZN => n878);
   U1356 : OR2_X1 port map( A1 => n4921, A2 => n5052, ZN => n879);
   U1357 : NAND3_X1 port map( A1 => n4920, A2 => n879, A3 => n878, ZN => n5047)
                           ;
   U1358 : AND2_X1 port map( A1 => n1470, A2 => n17222, ZN => n882);
   U1359 : NAND2_X1 port map( A1 => n883, A2 => n884, ZN => n885);
   U1360 : NAND2_X1 port map( A1 => n885, A2 => n6184, ZN => n6327);
   U1361 : INV_X1 port map( A => n6206, ZN => n883);
   U1362 : INV_X1 port map( A => n915, ZN => n884);
   U1363 : OR2_X1 port map( A1 => n6204, A2 => n995, ZN => n886);
   U1364 : OR2_X1 port map( A1 => n971, A2 => n5289, ZN => n887);
   U1365 : NAND2_X1 port map( A1 => n5205, A2 => n887, ZN => n5375);
   U1366 : OR2_X1 port map( A1 => n5208, A2 => n5367, ZN => n888);
   U1367 : OR2_X1 port map( A1 => n5365, A2 => n5364, ZN => n889);
   U1368 : NAND3_X1 port map( A1 => n888, A2 => n889, A3 => n5207, ZN => n5360)
                           ;
   U1369 : NAND2_X1 port map( A1 => n5354, A2 => n2245, ZN => n890);
   U1372 : NOR2_X1 port map( A1 => n1785, A2 => n1011, ZN => n893);
   U1373 : AND2_X1 port map( A1 => n734, A2 => n5127, ZN => n894);
   U1374 : AND2_X1 port map( A1 => n1471, A2 => n1703, ZN => n895);
   U1375 : AND2_X1 port map( A1 => n1471, A2 => n1703, ZN => n1642);
   U1376 : MUX2_X2 port map( A => n5347, B => n5346, S => n2246, Z => n896);
   U1377 : MUX2_X1 port map( A => n1686, B => n1685, S => n1731, Z => n1106);
   U1378 : NAND2_X1 port map( A1 => n943, A2 => n1790, ZN => n898);
   U1379 : OR2_X1 port map( A1 => n6677, A2 => n6646, ZN => n6669);
   U1380 : OR2_X1 port map( A1 => n1133, A2 => n6574, ZN => n6607);
   U1381 : NAND2_X1 port map( A1 => n6186, A2 => n1361, ZN => n899);
   U1382 : OR2_X1 port map( A1 => n8226, A2 => n8227, ZN => n900);
   U1383 : NAND2_X1 port map( A1 => n900, A2 => n2166, ZN => n6184);
   U1384 : NAND2_X1 port map( A1 => n7050, A2 => n7471, ZN => n901);
   U1385 : NAND2_X1 port map( A1 => n7049, A2 => n7647, ZN => n902);
   U1386 : NAND2_X1 port map( A1 => n901, A2 => n902, ZN => n1507);
   U1387 : CLKBUF_X1 port map( A => n7479, Z => n903);
   U1388 : OR2_X1 port map( A1 => n616, A2 => n6822, ZN => n904);
   U1389 : AND3_X1 port map( A1 => n4454, A2 => n1730, A3 => n831, ZN => n905);
   U1390 : INV_X1 port map( A => n5326, ZN => n906);
   U1391 : AND3_X1 port map( A1 => n1730, A2 => n4454, A3 => n831, ZN => n1758)
                           ;
   U1392 : NOR2_X1 port map( A1 => n8221, A2 => n907, ZN => n1830);
   U1394 : NAND2_X1 port map( A1 => n1187, A2 => n5322, ZN => n908);
   U1395 : MUX2_X2 port map( A => n1890, B => n1889, S => n859, Z => n909);
   U1396 : OR2_X1 port map( A1 => n4967, A2 => n4969, ZN => n910);
   U1397 : NAND2_X1 port map( A1 => n910, A2 => n4923, ZN => n5026);
   U1398 : AND2_X1 port map( A1 => n805, A2 => n1397, ZN => n912);
   U1399 : XNOR2_X1 port map( A => n914, B => n899, ZN => n6322);
   U1400 : MUX2_X1 port map( A => n6173, B => n6174, S => n750, Z => n915);
   U1402 : XNOR2_X1 port map( A => n814, B => n917, ZN => n7447);
   U1403 : AND2_X1 port map( A1 => n7444, A2 => n928, ZN => n917);
   U1405 : XNOR2_X1 port map( A => n918, B => n640, ZN => n6409);
   U1406 : XOR2_X1 port map( A => n6403, B => n6406, Z => n918);
   U1407 : OR2_X1 port map( A1 => n855, A2 => n6343, ZN => n919);
   U1408 : XNOR2_X1 port map( A => n6123, B => n920, ZN => n6131);
   U1410 : AND2_X1 port map( A1 => n903, A2 => n7480, ZN => n921);
   U1411 : OAI211_X1 port map( C1 => n4936, C2 => n4937, A => n730, B => n5086,
                           ZN => n923);
   U1412 : MUX2_X1 port map( A => n6986, B => n6987, S => n6369, Z => n7445);
   U1413 : INV_X1 port map( A => n2190, ZN => n924);
   U1414 : OAI22_X1 port map( A1 => n5746, A2 => n1812, B1 => n5854, B2 => 
                           n5845, ZN => n925);
   U1415 : INV_X1 port map( A => n1873, ZN => n2189);
   U1416 : XNOR2_X1 port map( A => n581, B => n1906, ZN => n1873);
   U1417 : XNOR2_X1 port map( A => n604, B => n4949, ZN => n1300);
   U1418 : AND2_X1 port map( A1 => n4939, A2 => n5134, ZN => n926);
   U1419 : OR2_X1 port map( A1 => n6490, A2 => n1094, ZN => n927);
   U1420 : NAND2_X1 port map( A1 => n6489, A2 => n927, ZN => n6804);
   U1421 : OR2_X1 port map( A1 => n7446, A2 => n7445, ZN => n928);
   U1423 : OAI21_X1 port map( B1 => n1744, B2 => n5831, A => n205, ZN => n930);
   U1424 : NAND2_X1 port map( A1 => n699, A2 => n313, ZN => n5162);
   U1425 : XNOR2_X1 port map( A => n5087, B => n931, ZN => n5089);
   U1426 : NAND2_X1 port map( A1 => n5085, A2 => n5086, ZN => n931);
   U1427 : XNOR2_X1 port map( A => n932, B => n5470, ZN => n5475);
   U1428 : XOR2_X1 port map( A => n678, B => n5465, Z => n932);
   U1429 : MUX2_X1 port map( A => n5627, B => n5626, S => n2244, Z => n5897);
   U1430 : MUX2_X1 port map( A => n5651, B => n5650, S => n2244, Z => n934);
   U1431 : MUX2_X1 port map( A => n5651, B => n5650, S => n2244, Z => n935);
   U1432 : CLKBUF_X1 port map( A => n1170, Z => n1040);
   U1433 : NAND2_X1 port map( A1 => n6750, A2 => n936, ZN => n937);
   U1434 : NAND2_X1 port map( A1 => n6749, A2 => n2246, ZN => n938);
   U1435 : INV_X1 port map( A => n2246, ZN => n936);
   U1436 : NOR2_X1 port map( A1 => n1313, A2 => n6841, ZN => n1838);
   U1437 : NAND2_X1 port map( A1 => n1339, A2 => n1336, ZN => n939);
   U1438 : OR2_X1 port map( A1 => n6673, A2 => n711, ZN => n940);
   U1439 : NAND2_X1 port map( A1 => n6644, A2 => n940, ZN => n6815);
   U1440 : OAI222_X1 port map( A1 => n6848, A2 => n1449, B1 => n1862, B2 => 
                           n6847, C1 => n1862, C2 => n6846, ZN => n7287);
   U1441 : INV_X1 port map( A => n1532, ZN => n943);
   U1442 : INV_X1 port map( A => n2232, ZN => n2230);
   U1443 : XNOR2_X1 port map( A => n944, B => n1801, ZN => n4948);
   U1444 : AND2_X1 port map( A1 => n4852, A2 => n4853, ZN => n944);
   U1445 : CLKBUF_X1 port map( A => n7261, Z => n945);
   U1446 : XNOR2_X1 port map( A => n1314, B => n6765, ZN => n1078);
   U1447 : MUX2_X1 port map( A => n1749, B => n1748, S => n7771, Z => n1747);
   U1448 : NOR2_X1 port map( A1 => n1178, A2 => n6292, ZN => n946);
   U1449 : AND2_X1 port map( A1 => n854, A2 => n7427, ZN => n947);
   U1450 : XNOR2_X1 port map( A => n948, B => n782, ZN => n6116);
   U1451 : XOR2_X1 port map( A => n1533, B => n6115, Z => n948);
   U1453 : NAND2_X1 port map( A1 => n1122, A2 => n1123, ZN => n951);
   U1454 : NAND2_X1 port map( A1 => n1123, A2 => n1122, ZN => n952);
   U1455 : NAND2_X1 port map( A1 => n6148, A2 => n750, ZN => n954);
   U1456 : NAND2_X1 port map( A1 => n6147, A2 => n2265, ZN => n955);
   U1457 : NAND2_X1 port map( A1 => n954, A2 => n955, ZN => n6326);
   U1458 : CLKBUF_X1 port map( A => n17184, Z => n956);
   U1459 : OR2_X1 port map( A1 => n929, A2 => n5530, ZN => n957);
   U1460 : OR2_X1 port map( A1 => n5845, A2 => n5833, ZN => n959);
   U1461 : NAND2_X1 port map( A1 => n959, A2 => n5832, ZN => n5843);
   U1462 : XNOR2_X1 port map( A => n929, B => n960, ZN => n967);
   U1463 : XNOR2_X1 port map( A => n961, B => n5598, ZN => n5607);
   U1464 : XOR2_X1 port map( A => n769, B => n5599, Z => n961);
   U1465 : AND2_X1 port map( A1 => n6993, A2 => n6990, ZN => n962);
   U1466 : MUX2_X2 port map( A => n6260, B => n6261, S => n859, Z => n6459);
   U1467 : NAND2_X1 port map( A1 => n7060, A2 => n7647, ZN => n963);
   U1468 : NAND2_X1 port map( A1 => n7061, A2 => n7471, ZN => n964);
   U1470 : NAND2_X1 port map( A1 => n5363, A2 => n1092, ZN => n965);
   U1471 : NAND2_X1 port map( A1 => n5362, A2 => n2246, ZN => n966);
   U1472 : NAND2_X1 port map( A1 => n965, A2 => n966, ZN => n1198);
   U1473 : MUX2_X1 port map( A => n1691, B => n1690, S => n6369, Z => n1689);
   U1474 : XNOR2_X1 port map( A => n5733, B => n967, ZN => n5740);
   U1475 : XNOR2_X1 port map( A => n5555, B => n968, ZN => n5556);
   U1476 : XNOR2_X1 port map( A => n875, B => n1746, ZN => n968);
   U1477 : INV_X1 port map( A => n5734, ZN => n1006);
   U1478 : XNOR2_X1 port map( A => n748, B => n17146, ZN => n5578);
   U1479 : BUF_X1 port map( A => n5181, Z => n969);
   U1480 : OAI21_X1 port map( B1 => n1651, B2 => n6575, A => n6621, ZN => n970)
                           ;
   U1481 : INV_X1 port map( A => n5290, ZN => n971);
   U1482 : AND2_X1 port map( A1 => n1240, A2 => n1241, ZN => n972);
   U1483 : INV_X1 port map( A => n6198, ZN => n974);
   U1484 : MUX2_X1 port map( A => n5371, B => n5372, S => n936, Z => n5609);
   U1485 : OAI21_X1 port map( B1 => n1852, B2 => n1843, A => n6918, ZN => n976)
                           ;
   U1486 : OR2_X1 port map( A1 => n869, A2 => n5796, ZN => n977);
   U1487 : NAND2_X1 port map( A1 => n977, A2 => n5795, ZN => n6704);
   U1488 : OR2_X1 port map( A1 => n5632, A2 => n5633, ZN => n978);
   U1489 : NAND2_X1 port map( A1 => n978, A2 => n5631, ZN => n5547);
   U1490 : AND2_X2 port map( A1 => n6099, A2 => n5997, ZN => n979);
   U1491 : OAI21_X1 port map( B1 => n17186, B2 => n6363, A => n6362, ZN => n980
                           );
   U1492 : NAND2_X1 port map( A1 => n5835, A2 => n1509, ZN => n981);
   U1493 : AND2_X1 port map( A1 => n6223, A2 => n6241, ZN => n6195);
   U1494 : INV_X1 port map( A => n1580, ZN => n982);
   U1495 : AND2_X1 port map( A1 => n1101, A2 => n1102, ZN => n983);
   U1496 : AND2_X1 port map( A1 => n17188, A2 => n7007, ZN => n984);
   U1497 : OAI21_X1 port map( B1 => n1793, B2 => n1607, A => n6119, ZN => n985)
                           ;
   U1498 : NAND2_X1 port map( A1 => n6401, A2 => n986, ZN => n987);
   U1499 : NAND2_X1 port map( A1 => n6402, A2 => n529, ZN => n988);
   U1500 : NAND2_X1 port map( A1 => n987, A2 => n988, ZN => n6519);
   U1501 : INV_X1 port map( A => n6410, ZN => n6420);
   U1502 : NAND2_X1 port map( A1 => n6466, A2 => n1476, ZN => n989);
   U1503 : XNOR2_X1 port map( A => n7026, B => n990, ZN => n1724);
   U1504 : AND2_X1 port map( A1 => n7013, A2 => n1488, ZN => n990);
   U1505 : NAND2_X1 port map( A1 => n6642, A2 => n1384, ZN => n991);
   U1506 : AND2_X1 port map( A1 => n231, A2 => n7069, ZN => n992);
   U1507 : AND2_X1 port map( A1 => n6691, A2 => n1614, ZN => n993);
   U1508 : INV_X1 port map( A => n6354, ZN => n994);
   U1510 : AND2_X1 port map( A1 => n6359, A2 => n1409, ZN => n997);
   U1511 : NAND2_X1 port map( A1 => n639, A2 => n1033, ZN => n998);
   U1513 : XNOR2_X1 port map( A => n6977, B => n6978, ZN => n6794);
   U1514 : XNOR2_X1 port map( A => n6324, B => n6323, ZN => n1001);
   U1515 : XNOR2_X1 port map( A => n1408, B => n7054, ZN => n1188);
   U1516 : MUX2_X1 port map( A => n1752, B => n1751, S => n6369, Z => n1177);
   U1517 : XNOR2_X1 port map( A => n1001, B => n583, ZN => n1052);
   U1518 : AND2_X1 port map( A1 => n5190, A2 => n5189, ZN => n5193);
   U1520 : NAND2_X1 port map( A1 => n6376, A2 => n986, ZN => n1004);
   U1521 : NAND2_X1 port map( A1 => n6377, A2 => n529, ZN => n1005);
   U1522 : NAND2_X1 port map( A1 => n1004, A2 => n1005, ZN => n6497);
   U1523 : CLKBUF_X1 port map( A => n6112, Z => n1008);
   U1524 : MUX2_X1 port map( A => n5982, B => n5981, S => n2267, Z => n6139);
   U1525 : AND3_X1 port map( A1 => n6056, A2 => n851, A3 => n6055, ZN => n1009)
                           ;
   U1527 : AND2_X1 port map( A1 => n5531, A2 => n8128, ZN => n1010);
   U1528 : AND2_X1 port map( A1 => n1530, A2 => n5457, ZN => n1011);
   U1529 : XOR2_X1 port map( A => n5844, B => n1081, Z => n1685);
   U1530 : NAND2_X1 port map( A1 => n5547, A2 => n1444, ZN => n1012);
   U1531 : XNOR2_X1 port map( A => n5336, B => n1780, ZN => n5339);
   U1532 : OR2_X1 port map( A1 => n4654, A2 => n4850, ZN => n4837);
   U1533 : XNOR2_X1 port map( A => n1014, B => n1015, ZN => n1755);
   U1534 : AND2_X1 port map( A1 => n5669, A2 => n5670, ZN => n1014);
   U1535 : XNOR2_X1 port map( A => n791, B => n5671, ZN => n1015);
   U1536 : AND2_X1 port map( A1 => n6556, A2 => n6476, ZN => n1016);
   U1537 : XOR2_X1 port map( A => n5971, B => n5916, Z => n5918);
   U1538 : NAND2_X1 port map( A1 => n7447, A2 => n7835, ZN => n1017);
   U1539 : NAND2_X1 port map( A1 => n7448, A2 => n6495, ZN => n1018);
   U1540 : NOR2_X1 port map( A1 => n4529, A2 => n817, ZN => n4454);
   U1541 : OR2_X1 port map( A1 => n4682, A2 => n4684, ZN => n1019);
   U1542 : NAND2_X1 port map( A1 => n1019, A2 => n4618, ZN => n4703);
   U1543 : OR2_X1 port map( A1 => n4676, A2 => n4678, ZN => n1020);
   U1544 : NAND2_X1 port map( A1 => n1020, A2 => n4616, ZN => n4716);
   U1545 : OR2_X1 port map( A1 => n4598, A2 => n4453, ZN => n4529);
   U1546 : OR2_X1 port map( A1 => n7407, A2 => n7406, ZN => n1021);
   U1547 : OR2_X1 port map( A1 => n5624, A2 => n504, ZN => n1022);
   U1548 : NAND2_X1 port map( A1 => n5519, A2 => n1022, ZN => n5610);
   U1549 : OR2_X1 port map( A1 => n5551, A2 => n5553, ZN => n1023);
   U1550 : NAND2_X1 port map( A1 => n1023, A2 => n5598, ZN => n5580);
   U1551 : OR2_X1 port map( A1 => n5046, A2 => n4969, ZN => n1024);
   U1552 : NAND2_X1 port map( A1 => n1024, A2 => n4968, ZN => n5028);
   U1553 : OR2_X1 port map( A1 => n438, A2 => n5077, ZN => n1025);
   U1554 : OR2_X1 port map( A1 => n5072, A2 => n1611, ZN => n1026);
   U1555 : NAND3_X1 port map( A1 => n1025, A2 => n1026, A3 => n4962, ZN => 
                           n5068);
   U1556 : AND2_X1 port map( A1 => n467, A2 => n1402, ZN => n1027);
   U1557 : INV_X1 port map( A => n780, ZN => n1028);
   U1559 : AND2_X1 port map( A1 => n6178, A2 => n6149, ZN => n1789);
   U1560 : XNOR2_X1 port map( A => n219, B => n1029, ZN => n5677);
   U1561 : XNOR2_X1 port map( A => n5672, B => n5675, ZN => n1029);
   U1562 : NAND2_X1 port map( A1 => n7071, A2 => n7072, ZN => n1030);
   U1563 : MUX2_X2 port map( A => n6293, B => n6294, S => n859, Z => n1031);
   U1564 : MUX2_X1 port map( A => n6293, B => n6294, S => n859, Z => n1032);
   U1565 : OR2_X1 port map( A1 => n5379, A2 => n778, ZN => n1033);
   U1566 : OR2_X1 port map( A1 => n6108, A2 => n17150, ZN => n1034);
   U1567 : NAND2_X1 port map( A1 => n17215, A2 => n1034, ZN => n6096);
   U1568 : XNOR2_X1 port map( A => n1036, B => n997, ZN => n6462);
   U1569 : MUX2_X2 port map( A => n7435, B => n7436, S => n6369, Z => n7437);
   U1570 : OAI22_X1 port map( A1 => n1117, A2 => n602, B1 => n747, B2 => n6221,
                           ZN => n1037);
   U1571 : OR2_X1 port map( A1 => n6505, A2 => n6515, ZN => n1459);
   U1573 : BUF_X1 port map( A => n4910, Z => n1222);
   U1574 : XNOR2_X1 port map( A => n5424, B => n1038, ZN => n5427);
   U1575 : NAND2_X1 port map( A1 => n716, A2 => n6662, ZN => n1039);
   U1576 : OR2_X1 port map( A1 => n5658, A2 => n726, ZN => n1041);
   U1577 : NAND2_X1 port map( A1 => n5539, A2 => n1041, ZN => n5644);
   U1578 : XNOR2_X1 port map( A => n5328, B => n5211, ZN => n5329);
   U1579 : CLKBUF_X1 port map( A => n5174, Z => n1042);
   U1580 : NAND2_X1 port map( A1 => n4852, A2 => n4853, ZN => n1043);
   U1581 : OR2_X1 port map( A1 => n1576, A2 => n7014, ZN => n1488);
   U1582 : INV_X1 port map( A => n7498, ZN => n1044);
   U1583 : NOR2_X1 port map( A1 => n1046, A2 => n1045, ZN => n7493);
   U1584 : AND2_X1 port map( A1 => n7485, A2 => n7486, ZN => n1045);
   U1585 : NAND2_X1 port map( A1 => n7504, A2 => n1044, ZN => n1046);
   U1586 : AND2_X1 port map( A1 => n4843, A2 => n1569, ZN => n1047);
   U1587 : NAND4_X1 port map( A1 => n230, A2 => n5467, A3 => n5466, A4 => n898,
                           ZN => n1048);
   U1588 : XNOR2_X1 port map( A => n549, B => n1049, ZN => n7421);
   U1589 : AND2_X1 port map( A1 => n1331, A2 => n7419, ZN => n1049);
   U1590 : INV_X1 port map( A => n846, ZN => n6349);
   U1591 : OR2_X1 port map( A1 => n2246, A2 => n7308, ZN => n1053);
   U1592 : NAND2_X1 port map( A1 => n1742, A2 => n1054, ZN => n4615);
   U1593 : OR2_X1 port map( A1 => n5252, A2 => n5255, ZN => n1055);
   U1594 : NAND2_X1 port map( A1 => n1055, A2 => n5248, ZN => n5249);
   U1595 : MUX2_X2 port map( A => n1804, B => n1805, S => n2247, Z => n1803);
   U1596 : XNOR2_X1 port map( A => n5410, B => n1056, ZN => n5428);
   U1597 : XOR2_X1 port map( A => n5422, B => n5281, Z => n1056);
   U1598 : NAND2_X1 port map( A1 => n1283, A2 => n665, ZN => n1057);
   U1600 : AND2_X1 port map( A1 => n5156, A2 => n5129, ZN => n1059);
   U1601 : XNOR2_X1 port map( A => n1729, B => n7420, ZN => n1388);
   U1602 : NAND2_X1 port map( A1 => n5985, A2 => n1394, ZN => n1061);
   U1603 : AND2_X1 port map( A1 => n5547, A2 => n1444, ZN => n1062);
   U1604 : XNOR2_X1 port map( A => n5973, B => n1063, ZN => n5982);
   U1605 : XNOR2_X1 port map( A => n935, B => n5979, ZN => n1063);
   U1607 : OR2_X1 port map( A1 => n6820, A2 => n616, ZN => n1065);
   U1608 : NAND2_X1 port map( A1 => n6816, A2 => n1065, ZN => n6998);
   U1609 : OAI21_X1 port map( B1 => n6599, B2 => n1586, A => n6572, ZN => n1066
                           );
   U1611 : CLKBUF_X1 port map( A => n6568, Z => n1067);
   U1612 : XNOR2_X1 port map( A => n1068, B => n1516, ZN => n1393);
   U1613 : XNOR2_X1 port map( A => n6585, B => n6629, ZN => n1068);
   U1614 : INV_X1 port map( A => n794, ZN => n5140);
   U1615 : AND2_X1 port map( A1 => n6771, A2 => n6770, ZN => n1071);
   U1616 : AND2_X1 port map( A1 => n1841, A2 => n1210, ZN => n1072);
   U1617 : NOR3_X1 port map( A1 => n1071, A2 => n1072, A3 => n6769, ZN => n6780
                           );
   U1618 : XNOR2_X1 port map( A => n1073, B => n653, ZN => n6463);
   U1619 : XNOR2_X1 port map( A => n711, B => n6657, ZN => n1460);
   U1620 : XNOR2_X1 port map( A => n6422, B => n1074, ZN => n6423);
   U1621 : XOR2_X1 port map( A => n6410, B => n6421, Z => n1074);
   U1622 : OAI21_X1 port map( B1 => n6599, B2 => n1586, A => n6572, ZN => n6829
                           );
   U1623 : OR2_X1 port map( A1 => n725, A2 => n7393, ZN => n1075);
   U1624 : NAND2_X1 port map( A1 => n7392, A2 => n1075, ZN => n7394);
   U1625 : XNOR2_X1 port map( A => n6738, B => n6882, ZN => n6739);
   U1626 : OR2_X1 port map( A1 => n6484, A2 => n6524, ZN => n6510);
   U1627 : CLKBUF_X1 port map( A => n1782, Z => n1076);
   U1628 : XNOR2_X1 port map( A => n7343, B => n7342, ZN => n7305);
   U1629 : XNOR2_X1 port map( A => n7305, B => n7313, ZN => n7307);
   U1630 : NAND2_X1 port map( A1 => n6569, A2 => n1190, ZN => n1077);
   U1631 : NAND2_X1 port map( A1 => n7415, A2 => n7414, ZN => n1503);
   U1632 : XNOR2_X1 port map( A => n6945, B => n1078, ZN => n5839);
   U1633 : OR2_X1 port map( A1 => n6081, A2 => n6072, ZN => n1079);
   U1634 : OR2_X1 port map( A1 => n6078, A2 => n6076, ZN => n1080);
   U1635 : NAND2_X1 port map( A1 => n1330, A2 => n5747, ZN => n1081);
   U1636 : XOR2_X1 port map( A => n5855, B => n1671, Z => n1082);
   U1637 : NOR3_X1 port map( A1 => n1642, A2 => n1816, A3 => n347, ZN => n5846)
                           ;
   U1638 : INV_X1 port map( A => n6491, ZN => n1083);
   U1639 : INV_X1 port map( A => n6792, ZN => n1084);
   U1640 : NAND2_X1 port map( A1 => n5331, A2 => n2246, ZN => n1085);
   U1641 : NAND2_X1 port map( A1 => n5332, A2 => n936, ZN => n1086);
   U1642 : NAND2_X1 port map( A1 => n1085, A2 => n1086, ZN => n5561);
   U1643 : NAND2_X1 port map( A1 => n5580, A2 => n5581, ZN => n1088);
   U1644 : INV_X1 port map( A => n5464, ZN => n1090);
   U1645 : OR2_X2 port map( A1 => n8142, A2 => n1091, ZN => n8130);
   U1646 : AND2_X2 port map( A1 => n6704, A2 => n6703, ZN => n1843);
   U1647 : NOR3_X1 port map( A1 => n1841, A2 => n1877, A3 => n314, ZN => n6777)
                           ;
   U1648 : MUX2_X1 port map( A => n258, B => n281, S => n2152, Z => n6776);
   U1649 : XNOR2_X1 port map( A => n6443, B => n6351, ZN => n6444);
   U1650 : AND2_X1 port map( A1 => n4863, A2 => n1851, ZN => n1093);
   U1651 : NAND2_X1 port map( A1 => n972, A2 => n5812, ZN => n1095);
   U1652 : XNOR2_X1 port map( A => n1096, B => n6415, ZN => n6424);
   U1653 : XNOR2_X1 port map( A => n6410, B => n6421, ZN => n1096);
   U1654 : AND2_X1 port map( A1 => n6481, A2 => n1306, ZN => n1097);
   U1655 : XNOR2_X1 port map( A => n17210, B => n17155, ZN => n1326);
   U1656 : NAND2_X1 port map( A1 => n6558, A2 => n6557, ZN => n1098);
   U1657 : OR2_X1 port map( A1 => n5679, A2 => n17256, ZN => n1099);
   U1658 : NAND2_X1 port map( A1 => n5496, A2 => n1099, ZN => n5674);
   U1659 : NAND2_X1 port map( A1 => n1100, A2 => n4551, ZN => n1101);
   U1660 : NAND2_X1 port map( A1 => n17165, A2 => n1833, ZN => n1102);
   U1661 : NAND2_X1 port map( A1 => n1101, A2 => n1102, ZN => n4647);
   U1662 : INV_X1 port map( A => n1833, ZN => n1100);
   U1663 : INV_X1 port map( A => n6623, ZN => n1103);
   U1664 : OAI21_X1 port map( B1 => n5867, B2 => n5829, A => n5864, ZN => n1105
                           );
   U1665 : OR2_X1 port map( A1 => n5805, A2 => n5859, ZN => n1107);
   U1666 : NAND2_X1 port map( A1 => n1107, A2 => n5857, ZN => n5852);
   U1667 : MUX2_X1 port map( A => n1685, B => n1686, S => n2268, Z => n1684);
   U1668 : INV_X1 port map( A => n1333, ZN => n1108);
   U1669 : INV_X1 port map( A => n5788, ZN => n1109);
   U1670 : OR2_X1 port map( A1 => n5012, A2 => n5013, ZN => n1110);
   U1671 : NAND2_X1 port map( A1 => n1110, A2 => n5014, ZN => n4989);
   U1672 : OR2_X1 port map( A1 => n5262, A2 => n5265, ZN => n1111);
   U1673 : NAND2_X1 port map( A1 => n1111, A2 => n5260, ZN => n5767);
   U1674 : MUX2_X2 port map( A => n5228, B => n5227, S => n804, Z => n5265);
   U1675 : XNOR2_X1 port map( A => n1165, B => n1113, ZN => n1719);
   U1676 : XNOR2_X1 port map( A => n1134, B => n6141, ZN => n1113);
   U1677 : XNOR2_X1 port map( A => n1114, B => n6554, ZN => n1325);
   U1678 : AND2_X1 port map( A1 => n6553, A2 => n6552, ZN => n1114);
   U1679 : XOR2_X1 port map( A => n6205, B => n6328, Z => n2161);
   U1680 : OR2_X1 port map( A1 => n7003, A2 => n7002, ZN => n1115);
   U1681 : NAND2_X1 port map( A1 => n1115, A2 => n7001, ZN => n7451);
   U1682 : NAND2_X1 port map( A1 => n5958, A2 => n1095, ZN => n1116);
   U1683 : AND2_X1 port map( A1 => n1225, A2 => n6219, ZN => n1117);
   U1684 : CLKBUF_X1 port map( A => n8187, Z => n1118);
   U1685 : AND2_X1 port map( A1 => n7441, A2 => n7440, ZN => n1119);
   U1686 : NOR2_X1 port map( A1 => n1179, A2 => n1119, ZN => n7442);
   U1688 : NAND2_X1 port map( A1 => n5597, A2 => n1121, ZN => n1122);
   U1689 : NAND2_X1 port map( A1 => n5596, A2 => n2244, ZN => n1123);
   U1690 : INV_X1 port map( A => n2244, ZN => n1121);
   U1691 : BUF_X4 port map( A => n8135, Z => n2244);
   U1692 : MUX2_X2 port map( A => n6401, B => n6402, S => n529, Z => n1124);
   U1693 : INV_X1 port map( A => n1760, ZN => n7196);
   U1694 : NAND2_X1 port map( A1 => n7549, A2 => n411, ZN => n7551);
   U1695 : OAI22_X1 port map( A1 => n863, A2 => n6692, B1 => n7010, B2 => n7012
                           , ZN => n1125);
   U1696 : NAND2_X1 port map( A1 => n1201, A2 => n6753, ZN => n1127);
   U1697 : BUF_X2 port map( A => n1760, Z => n2130);
   U1698 : XNOR2_X1 port map( A => n5703, B => n1128, ZN => n5704);
   U1699 : XNOR2_X1 port map( A => n704, B => n5696, ZN => n1128);
   U1700 : INV_X1 port map( A => n1391, ZN => n6651);
   U1701 : XNOR2_X1 port map( A => n1124, B => n845, ZN => n1589);
   U1702 : OR2_X1 port map( A1 => n4685, A2 => n4687, ZN => n1129);
   U1703 : NAND2_X1 port map( A1 => n1129, A2 => n4619, ZN => n4696);
   U1704 : NAND2_X1 port map( A1 => n7491, A2 => n7581, ZN => n1130);
   U1705 : INV_X1 port map( A => n6024, ZN => n1131);
   U1706 : XNOR2_X1 port map( A => n5020, B => n4976, ZN => n5023);
   U1707 : XOR2_X1 port map( A => n4863, B => n4886, Z => n4887);
   U1708 : BUF_X1 port map( A => n7316, Z => n2225);
   U1709 : BUF_X2 port map( A => n7316, Z => n2226);
   U1710 : CLKBUF_X1 port map( A => n545, Z => n1135);
   U1711 : MUX2_X1 port map( A => n1666, B => n1665, S => n4436, Z => n1408);
   U1712 : XNOR2_X1 port map( A => n1881, B => n1136, ZN => n7454);
   U1713 : AND2_X1 port map( A1 => n1316, A2 => n7452, ZN => n1136);
   U1715 : NAND2_X1 port map( A1 => n7049, A2 => n7647, ZN => n1138);
   U1716 : OAI21_X1 port map( B1 => n8154, B2 => n5460, A => n443, ZN => n1139)
                           ;
   U1717 : OR2_X1 port map( A1 => n7054, A2 => n7047, ZN => n1140);
   U1718 : NAND2_X1 port map( A1 => n7038, A2 => n1140, ZN => n7472);
   U1720 : MUX2_X2 port map( A => n7373, B => n7372, S => n2244, Z => n7374);
   U1721 : MUX2_X1 port map( A => n1665, B => n1666, S => n7712, Z => n1142);
   U1722 : OR2_X1 port map( A1 => n6236, A2 => n6233, ZN => n1143);
   U1723 : NAND2_X1 port map( A1 => n6235, A2 => n1143, ZN => n6196);
   U1724 : XNOR2_X1 port map( A => n1664, B => n7051, ZN => n1299);
   U1725 : MUX2_X1 port map( A => n4984, B => n4983, S => n2247, Z => n5334);
   U1726 : XNOR2_X1 port map( A => n5445, B => n5446, ZN => n5447);
   U1727 : OR2_X1 port map( A1 => n929, A2 => n5734, ZN => n5640);
   U1728 : AND2_X1 port map( A1 => n4836, A2 => n1774, ZN => n1144);
   U1730 : NAND2_X1 port map( A1 => n1145, A2 => n7508, ZN => n7492);
   U1731 : INV_X2 port map( A => n834, ZN => n2239);
   U1732 : NAND2_X1 port map( A1 => n2174, A2 => n986, ZN => n1147);
   U1733 : NAND2_X1 port map( A1 => n2173, A2 => n529, ZN => n1148);
   U1734 : NAND2_X1 port map( A1 => n1148, A2 => n1147, ZN => n1517);
   U1735 : INV_X1 port map( A => n6288, ZN => n1150);
   U1736 : NOR3_X1 port map( A1 => n1233, A2 => n6086, A3 => n1234, ZN => n1151
                           );
   U1737 : CLKBUF_X1 port map( A => n1806, Z => n1152);
   U1738 : NOR3_X1 port map( A1 => n1234, A2 => n1233, A3 => n617, ZN => n6092)
                           ;
   U1739 : OR2_X1 port map( A1 => n6548, A2 => n1070, ZN => n1153);
   U1740 : NAND2_X1 port map( A1 => n6457, A2 => n1153, ZN => n6527);
   U1741 : AND2_X1 port map( A1 => n6196, A2 => n1687, ZN => n1154);
   U1742 : AND2_X1 port map( A1 => n6196, A2 => n1687, ZN => n1644);
   U1743 : INV_X1 port map( A => n807, ZN => n1155);
   U1744 : XNOR2_X1 port map( A => n1156, B => n1777, ZN => n5116);
   U1746 : OR2_X1 port map( A1 => n5878, A2 => n1058, ZN => n1158);
   U1747 : NAND2_X1 port map( A1 => n1158, A2 => n5744, ZN => n5864);
   U1748 : XNOR2_X1 port map( A => n5959, B => n1160, ZN => n5960);
   U1749 : AND2_X1 port map( A1 => n1492, A2 => n1493, ZN => n1160);
   U1750 : AND2_X1 port map( A1 => n6157, A2 => n6177, ZN => n1161);
   U1751 : INV_X1 port map( A => n1059, ZN => n1162);
   U1752 : NAND2_X1 port map( A1 => n6335, A2 => n1555, ZN => n1163);
   U1753 : XNOR2_X1 port map( A => n1164, B => n5724, ZN => n5727);
   U1754 : OR2_X1 port map( A1 => n17220, A2 => n1807, ZN => n1164);
   U1755 : NAND2_X1 port map( A1 => n5968, A2 => n1648, ZN => n1165);
   U1756 : MUX2_X2 port map( A => n6639, B => n6638, S => n7835, Z => n6647);
   U1757 : XNOR2_X1 port map( A => n17258, B => n5168, ZN => n5169);
   U1758 : XNOR2_X1 port map( A => n513, B => n1817, ZN => n1166);
   U1759 : XNOR2_X1 port map( A => n5998, B => n6169, ZN => n2160);
   U1760 : NAND2_X1 port map( A1 => n436, A2 => n7771, ZN => n1167);
   U1761 : CLKBUF_X1 port map( A => n6791, Z => n1332);
   U1762 : NAND2_X1 port map( A1 => n6504, A2 => n6369, ZN => n1168);
   U1763 : NAND2_X1 port map( A1 => n6503, A2 => n1702, ZN => n1169);
   U1764 : NAND2_X1 port map( A1 => n1168, A2 => n1169, ZN => n1181);
   U1765 : XNOR2_X1 port map( A => n6678, B => n1171, ZN => n1661);
   U1766 : NOR2_X1 port map( A1 => n6522, A2 => n1124, ZN => n1172);
   U1767 : OAI211_X1 port map( C1 => n1087, C2 => n6093, A => n757, B => n6092,
                           ZN => n1173);
   U1768 : AND2_X1 port map( A1 => n17190, A2 => n511, ZN => n1174);
   U1769 : XNOR2_X1 port map( A => n5436, B => n5437, ZN => n1176);
   U1770 : NAND3_X1 port map( A1 => n6077, A2 => n6078, A3 => n340, ZN => n6080
                           );
   U1771 : MUX2_X1 port map( A => n253, B => n255, S => n527, Z => n6967);
   U1772 : AND2_X1 port map( A1 => n6994, A2 => n6993, ZN => n1179);
   U1773 : XNOR2_X1 port map( A => n1180, B => n1820, ZN => n5434);
   U1774 : AND2_X1 port map( A1 => n5432, A2 => n5433, ZN => n1180);
   U1775 : AND2_X1 port map( A1 => n1816, A2 => n1858, ZN => n1183);
   U1776 : AND2_X1 port map( A1 => n1812, A2 => n5847, ZN => n1184);
   U1777 : NOR3_X1 port map( A1 => n5846, A2 => n1184, A3 => n1183, ZN => n5851
                           );
   U1778 : MUX2_X1 port map( A => n6504, B => n6503, S => n1702, Z => n6596);
   U1779 : XNOR2_X1 port map( A => n5401, B => n17214, ZN => n5402);
   U1780 : OR2_X1 port map( A1 => n711, A2 => n6657, ZN => n1185);
   U1781 : NAND2_X1 port map( A1 => n6656, A2 => n1185, ZN => n6818);
   U1782 : OR2_X1 port map( A1 => n6128, A2 => n17168, ZN => n1186);
   U1783 : NAND2_X1 port map( A1 => n5984, A2 => n1186, ZN => n6113);
   U1784 : NAND2_X1 port map( A1 => n5343, A2 => n5319, ZN => n1187);
   U1785 : XNOR2_X1 port map( A => n1188, B => n7052, ZN => n7053);
   U1786 : OR2_X1 port map( A1 => n5134, A2 => n4911, ZN => n1189);
   U1787 : OR2_X1 port map( A1 => n6632, A2 => n1580, ZN => n1190);
   U1788 : NAND2_X1 port map( A1 => n6569, A2 => n1190, ZN => n6621);
   U1789 : OR2_X1 port map( A1 => n855, A2 => n6396, ZN => n6382);
   U1790 : OR2_X1 port map( A1 => n6976, A2 => n6977, ZN => n7269);
   U1791 : XNOR2_X1 port map( A => n922, B => n763, ZN => n6988);
   U1792 : XNOR2_X1 port map( A => n1191, B => n578, ZN => n7060);
   U1793 : CLKBUF_X1 port map( A => n1142, Z => n1192);
   U1794 : MUX2_X1 port map( A => n6659, B => n6658, S => n7771, Z => n7023);
   U1795 : OR2_X1 port map( A1 => n6530, A2 => n1120, ZN => n1195);
   U1796 : AND2_X1 port map( A1 => n1707, A2 => n1708, ZN => n1196);
   U1797 : XOR2_X1 port map( A => n1360, B => n5145, Z => n1197);
   U1798 : XNOR2_X1 port map( A => n587, B => n7487, ZN => n1229);
   U1799 : AND2_X1 port map( A1 => n835, A2 => n4550, ZN => n1199);
   U1800 : XNOR2_X1 port map( A => n1200, B => n5359, ZN => n5363);
   U1801 : OR2_X1 port map( A1 => n5358, A2 => n1835, ZN => n1200);
   U1802 : OR2_X1 port map( A1 => n6755, A2 => n6754, ZN => n1201);
   U1803 : NAND2_X1 port map( A1 => n6753, A2 => n1201, ZN => n6899);
   U1804 : OR2_X1 port map( A1 => n4729, A2 => n4675, ZN => n1202);
   U1805 : NAND2_X1 port map( A1 => n1202, A2 => n4674, ZN => n4724);
   U1806 : OR2_X1 port map( A1 => n5255, A2 => n5254, ZN => n1203);
   U1807 : NAND2_X1 port map( A1 => n1203, A2 => n5253, ZN => n5758);
   U1808 : OR2_X1 port map( A1 => n5225, A2 => n5224, ZN => n1204);
   U1809 : NAND2_X1 port map( A1 => n1204, A2 => n5223, ZN => n5250);
   U1810 : NAND2_X1 port map( A1 => n1205, A2 => n4686, ZN => n4697);
   U1811 : OR2_X1 port map( A1 => n4722, A2 => n4678, ZN => n1206);
   U1812 : NAND2_X1 port map( A1 => n1206, A2 => n4677, ZN => n4717);
   U1813 : XNOR2_X1 port map( A => n518, B => n1798, ZN => n1207);
   U1814 : INV_X1 port map( A => n2135, ZN => n1208);
   U1815 : CLKBUF_X1 port map( A => n7389, Z => n1209);
   U1816 : AND2_X1 port map( A1 => n6775, A2 => n2268, ZN => n1210);
   U1817 : XNOR2_X1 port map( A => n611, B => n6220, ZN => n1380);
   U1818 : INV_X1 port map( A => n952, ZN => n1212);
   U1819 : INV_X1 port map( A => n6442, ZN => n1213);
   U1820 : INV_X1 port map( A => n704, ZN => n1214);
   U1821 : AND2_X1 port map( A1 => n4575, A2 => n4574, ZN => n1215);
   U1822 : NOR3_X1 port map( A1 => n1526, A2 => n1525, A3 => n1524, ZN => n1216
                           );
   U1823 : CLKBUF_X1 port map( A => n8130, Z => n1217);
   U1824 : NAND2_X1 port map( A1 => n5927, A2 => n5928, ZN => n1218);
   U1825 : NAND2_X1 port map( A1 => n5819, A2 => n1218, ZN => n5820);
   U1826 : INV_X1 port map( A => n6023, ZN => n1220);
   U1827 : AND2_X1 port map( A1 => n1530, A2 => n5274, ZN => n1221);
   U1829 : AND2_X1 port map( A1 => n6079, A2 => n1297, ZN => n1223);
   U1830 : OR2_X1 port map( A1 => n17256, A2 => n5537, ZN => n1224);
   U1831 : NAND2_X1 port map( A1 => n5536, A2 => n1224, ZN => n5676);
   U1832 : OR2_X1 port map( A1 => n1806, A2 => n6220, ZN => n1225);
   U1833 : NAND2_X1 port map( A1 => n1225, A2 => n6219, ZN => n6255);
   U1834 : MUX2_X1 port map( A => n6052, B => n6051, S => n2266, Z => n6234);
   U1835 : AND2_X1 port map( A1 => n6251, A2 => n6070, ZN => n1226);
   U1837 : NAND2_X1 port map( A1 => n821, A2 => n5108, ZN => n1227);
   U1838 : NAND2_X1 port map( A1 => n4915, A2 => n4914, ZN => n1228);
   U1839 : XNOR2_X1 port map( A => n6937, B => n1126, ZN => n6939);
   U1840 : XNOR2_X1 port map( A => n1229, B => n7488, ZN => n7064);
   U1841 : XNOR2_X1 port map( A => n568, B => n7003, ZN => n6824);
   U1842 : OR2_X1 port map( A1 => n7047, A2 => n7051, ZN => n1230);
   U1843 : NAND2_X1 port map( A1 => n1230, A2 => n7046, ZN => n7473);
   U1844 : OR2_X1 port map( A1 => n7478, A2 => n1693, ZN => n1231);
   U1845 : OR2_X1 port map( A1 => n7476, A2 => n7647, ZN => n1232);
   U1846 : NAND3_X1 port map( A1 => n7475, A2 => n1232, A3 => n1231, ZN => 
                           n7479);
   U1847 : AND2_X1 port map( A1 => n6088, A2 => n338, ZN => n1233);
   U1848 : AND2_X1 port map( A1 => n979, A2 => n6087, ZN => n1234);
   U1849 : NAND2_X1 port map( A1 => n7074, A2 => n7579, ZN => n1235);
   U1850 : NAND2_X1 port map( A1 => n5301, A2 => n5300, ZN => n1236);
   U1851 : XNOR2_X1 port map( A => n1238, B => n4904, ZN => n1567);
   U1852 : AND2_X1 port map( A1 => n4908, A2 => n4903, ZN => n1238);
   U1853 : NAND2_X1 port map( A1 => n2165, A2 => n1239, ZN => n1240);
   U1854 : NAND2_X1 port map( A1 => n2164, A2 => n1369, ZN => n1241);
   U1855 : NAND2_X1 port map( A1 => n1241, A2 => n1240, ZN => n1290);
   U1856 : INV_X1 port map( A => n1369, ZN => n1239);
   U1857 : INV_X1 port map( A => n2243, ZN => n1369);
   U1858 : OR2_X1 port map( A1 => n5760, A2 => n5759, ZN => n1243);
   U1859 : NAND2_X1 port map( A1 => n1243, A2 => n5758, ZN => n5761);
   U1860 : OR2_X1 port map( A1 => n4701, A2 => n4685, ZN => n1244);
   U1861 : NAND2_X1 port map( A1 => n4704, A2 => n1244, ZN => n4686);
   U1862 : OR2_X1 port map( A1 => n5252, A2 => n5251, ZN => n1245);
   U1863 : NAND2_X1 port map( A1 => n1245, A2 => n5250, ZN => n5253);
   U1864 : CLKBUF_X1 port map( A => n17230, Z => n1246);
   U1865 : XNOR2_X1 port map( A => n1247, B => n1248, ZN => n6293);
   U1866 : AND2_X1 port map( A1 => n6290, A2 => n6291, ZN => n1247);
   U1867 : XNOR2_X1 port map( A => n6524, B => n6484, ZN => n6525);
   U1868 : NAND2_X1 port map( A1 => n5677, A2 => n1249, ZN => n1250);
   U1869 : NAND2_X1 port map( A1 => n5678, A2 => n1351, ZN => n1251);
   U1870 : NAND2_X1 port map( A1 => n1250, A2 => n1251, ZN => n5948);
   U1871 : INV_X1 port map( A => n1351, ZN => n1249);
   U1872 : AND2_X1 port map( A1 => n6214, A2 => n1740, ZN => n1252);
   U1873 : INV_X1 port map( A => n2243, ZN => n1351);
   U1874 : MUX2_X1 port map( A => n4898, B => n4897, S => n804, Z => n1354);
   U1876 : AND2_X1 port map( A1 => n4940, A2 => n1568, ZN => n1253);
   U1877 : NAND2_X1 port map( A1 => n6616, A2 => n6619, ZN => n1254);
   U1878 : NAND2_X1 port map( A1 => n4544, A2 => n637, ZN => n1255);
   U1879 : NAND2_X1 port map( A1 => n2264, A2 => n4543, ZN => n1256);
   U1880 : NAND2_X1 port map( A1 => n1255, A2 => n1256, ZN => n4545);
   U1881 : AND2_X1 port map( A1 => n4635, A2 => n4651, ZN => n1257);
   U1882 : AND2_X1 port map( A1 => n1436, A2 => n1258, ZN => n1827);
   U1883 : AND2_X1 port map( A1 => n1437, A2 => n1892, ZN => n1258);
   U1884 : AND2_X1 port map( A1 => n1696, A2 => n1260, ZN => n1259);
   U1885 : NAND2_X1 port map( A1 => n1413, A2 => n6693, ZN => n1260);
   U1886 : NAND2_X1 port map( A1 => n1413, A2 => n6693, ZN => n1261);
   U1887 : XNOR2_X1 port map( A => n6136, B => n461, ZN => n1598);
   U1888 : NAND2_X1 port map( A1 => n484, A2 => n1493, ZN => n1262);
   U1889 : OR2_X1 port map( A1 => n7030, A2 => n7031, ZN => n1338);
   U1890 : NAND2_X1 port map( A1 => n4775, A2 => n818, ZN => n1264);
   U1891 : NAND2_X1 port map( A1 => n4774, A2 => n2250, ZN => n1265);
   U1892 : NAND2_X1 port map( A1 => n1265, A2 => n1264, ZN => n4963);
   U1893 : CLKBUF_X1 port map( A => DataPath_i_PIPLIN_B_0_port, Z => n1266);
   U1894 : OR2_X1 port map( A1 => n4666, A2 => n4668, ZN => n1267);
   U1895 : NAND2_X1 port map( A1 => n1267, A2 => n4608, ZN => n4772);
   U1896 : XNOR2_X1 port map( A => n1268, B => n5093, ZN => n1823);
   U1897 : AND2_X1 port map( A1 => n4916, A2 => n1461, ZN => n1268);
   U1898 : INV_X1 port map( A => n4851, ZN => n1269);
   U1899 : XNOR2_X1 port map( A => n1275, B => n2162, ZN => n5952);
   U1900 : NOR2_X1 port map( A1 => n4546, A2 => n4545, ZN => n1270);
   U1901 : NAND2_X1 port map( A1 => n6826, A2 => n6594, ZN => n1271);
   U1902 : NAND2_X1 port map( A1 => n1271, A2 => n766, ZN => n7019);
   U1903 : MUX2_X1 port map( A => n4407, B => n4406, S => n526, Z => n6594);
   U1904 : XNOR2_X1 port map( A => n5900, B => n1272, ZN => n5901);
   U1905 : XNOR2_X1 port map( A => n5109, B => n1273, ZN => n5120);
   U1906 : XNOR2_X1 port map( A => n604, B => n5117, ZN => n1273);
   U1907 : AND2_X1 port map( A1 => n4837, A2 => n4848, ZN => n1274);
   U1908 : INV_X1 port map( A => n17259, ZN => n1276);
   U1909 : AND2_X1 port map( A1 => n5826, A2 => n1457, ZN => n1277);
   U1910 : AND2_X1 port map( A1 => n1577, A2 => n8239, ZN => n1278);
   U1911 : OR2_X1 port map( A1 => n4694, A2 => n4695, ZN => n1279);
   U1912 : NAND2_X1 port map( A1 => n1279, A2 => n4696, ZN => n4620);
   U1913 : OR2_X1 port map( A1 => n4701, A2 => n4702, ZN => n1280);
   U1914 : NAND2_X1 port map( A1 => n1280, A2 => n4703, ZN => n4619);
   U1915 : OR2_X1 port map( A1 => n5221, A2 => n5224, ZN => n1281);
   U1916 : NAND2_X1 port map( A1 => n1281, A2 => n5219, ZN => n5248);
   U1917 : XNOR2_X1 port map( A => n5774, B => n5773, ZN => n1282);
   U1918 : INV_X1 port map( A => n5800, ZN => n1746);
   U1919 : MUX2_X1 port map( A => n6431, B => n6432, S => n529, Z => n1578);
   U1920 : NAND2_X1 port map( A1 => n4786, A2 => n1286, ZN => n1283);
   U1921 : AND2_X1 port map( A1 => n1283, A2 => n1284, ZN => n4667);
   U1922 : OR2_X1 port map( A1 => n1285, A2 => n1528, ZN => n1284);
   U1923 : INV_X1 port map( A => n1738, ZN => n1285);
   U1924 : AND2_X1 port map( A1 => n1737, A2 => n1738, ZN => n1286);
   U1925 : AND2_X1 port map( A1 => n755, A2 => n1670, ZN => n1287);
   U1926 : NAND2_X1 port map( A1 => n1047, A2 => n317, ZN => n4839);
   U1927 : AND3_X1 port map( A1 => n249, A2 => n5163, A3 => n1288, ZN => n5167)
                           ;
   U1929 : XNOR2_X1 port map( A => n6242, B => n1289, ZN => n6244);
   U1930 : XNOR2_X1 port map( A => n1681, B => n6241, ZN => n1289);
   U1931 : BUF_X1 port map( A => n5833, Z => n1671);
   U1932 : INV_X1 port map( A => n1193, ZN => n1291);
   U1933 : NAND2_X1 port map( A1 => n1130, A2 => n7503, ZN => n1292);
   U1934 : XNOR2_X1 port map( A => n1293, B => n1777, ZN => n5105);
   U1935 : AND2_X1 port map( A1 => n4826, A2 => n4827, ZN => n1293);
   U1936 : OR2_X2 port map( A1 => n4508, A2 => n4461, ZN => n4503);
   U1937 : XNOR2_X1 port map( A => n2153, B => n5135, ZN => n4911);
   U1938 : XNOR2_X1 port map( A => n5661, B => n1294, ZN => n5662);
   U1939 : XNOR2_X1 port map( A => n5657, B => n5658, ZN => n1294);
   U1940 : XNOR2_X1 port map( A => n6041, B => n5836, ZN => n5844);
   U1941 : XNOR2_X1 port map( A => n1295, B => n5451, ZN => n5455);
   U1942 : XOR2_X1 port map( A => n5197, B => n5453, Z => n1295);
   U1943 : XNOR2_X1 port map( A => n6129, B => n1296, ZN => n6130);
   U1944 : XOR2_X1 port map( A => n561, B => n6308, Z => n1890);
   U1945 : OR2_X1 port map( A1 => n5090, A2 => n4958, ZN => n1298);
   U1946 : NAND2_X1 port map( A1 => n4957, A2 => n1298, ZN => n4959);
   U1947 : XNOR2_X1 port map( A => n1299, B => n1383, ZN => n7055);
   U1948 : XNOR2_X1 port map( A => n1884, B => n7489, ZN => n1561);
   U1949 : XNOR2_X1 port map( A => n1300, B => n5118, ZN => n5119);
   U1950 : MUX2_X2 port map( A => n1890, B => n1889, S => n859, Z => n1888);
   U1951 : OAI21_X1 port map( B1 => n6374, B2 => n250, A => n6341, ZN => n1303)
                           ;
   U1952 : OR2_X1 port map( A1 => n6022, A2 => n892, ZN => n1304);
   U1953 : NAND2_X1 port map( A1 => n6021, A2 => n1304, ZN => n6098);
   U1954 : BUF_X1 port map( A => n8276, Z => n2269);
   U1955 : NAND2_X1 port map( A1 => n4801, A2 => n312, ZN => n4803);
   U1956 : OR2_X1 port map( A1 => n1120, A2 => n6482, ZN => n1306);
   U1957 : NAND2_X1 port map( A1 => n6481, A2 => n1306, ZN => n6483);
   U1958 : XNOR2_X1 port map( A => n1660, B => n7010, ZN => n1307);
   U1959 : XOR2_X1 port map( A => n1561, B => n921, Z => n1308);
   U1960 : OR2_X1 port map( A1 => n2266, A2 => n6846, ZN => n1309);
   U1961 : NAND2_X1 port map( A1 => n1309, A2 => n6788, ZN => n6836);
   U1962 : OR2_X1 port map( A1 => n5553, A2 => n1198, ZN => n1310);
   U1963 : NAND2_X1 port map( A1 => n5552, A2 => n1310, ZN => n5594);
   U1964 : NOR2_X1 port map( A1 => n5588, A2 => n5587, ZN => n1311);
   U1965 : NOR2_X1 port map( A1 => n5586, A2 => n1787, ZN => n1312);
   U1966 : XNOR2_X1 port map( A => n6836, B => n1879, ZN => n1313);
   U1967 : XOR2_X1 port map( A => n5804, B => n1897, Z => n1314);
   U1968 : INV_X1 port map( A => n4891, ZN => n1315);
   U1969 : OR2_X1 port map( A1 => n7453, A2 => n882, ZN => n1316);
   U1970 : OAI22_X1 port map( A1 => n2191, A2 => n17195, B1 => n2229, B2 => 
                           n494, ZN => n4896);
   U1971 : AND2_X1 port map( A1 => n1354, A2 => n1875, ZN => n1319);
   U1972 : INV_X1 port map( A => n577, ZN => n1320);
   U1973 : NAND2_X1 port map( A1 => n5701, A2 => n1321, ZN => n5685);
   U1974 : INV_X1 port map( A => n5134, ZN => n1322);
   U1975 : XNOR2_X1 port map( A => n1335, B => n7014, ZN => n1343);
   U1976 : NAND2_X1 port map( A1 => n1669, A2 => n1670, ZN => n1323);
   U1978 : MUX2_X1 port map( A => n6675, B => n6676, S => n6594, Z => n7027);
   U1979 : INV_X1 port map( A => n913, ZN => n6580);
   U1980 : AND2_X1 port map( A1 => n1699, A2 => n7040, ZN => n1796);
   U1981 : OR2_X1 port map( A1 => n5266, A2 => n5265, ZN => n1327);
   U1982 : NAND2_X1 port map( A1 => n1327, A2 => n5264, ZN => n5769);
   U1983 : OR2_X1 port map( A1 => n5774, A2 => n5773, ZN => n1328);
   U1984 : NAND2_X1 port map( A1 => n5772, A2 => n1328, ZN => n6711);
   U1985 : OR2_X1 port map( A1 => n5848, A2 => n1671, ZN => n1330);
   U1986 : NAND2_X1 port map( A1 => n925, A2 => n1330, ZN => n6045);
   U1987 : OR2_X1 port map( A1 => n7420, A2 => n565, ZN => n1331);
   U1988 : AND2_X1 port map( A1 => n7479, A2 => n7480, ZN => n1905);
   U1989 : OAI21_X1 port map( B1 => n1852, B2 => n1843, A => n6918, ZN => n1333
                           );
   U1990 : OAI21_X1 port map( B1 => n6908, B2 => n1850, A => n6906, ZN => n1334
                           );
   U1991 : MUX2_X1 port map( A => n6676, B => n6675, S => n7771, Z => n1335);
   U1992 : XNOR2_X1 port map( A => n6451, B => n909, ZN => n6449);
   U1993 : MUX2_X2 port map( A => n5793, B => n5794, S => n936, Z => n6754);
   U1994 : XNOR2_X1 port map( A => n725, B => n7393, ZN => n7276);
   U1995 : NAND2_X1 port map( A1 => n7055, A2 => n7647, ZN => n1336);
   U1996 : INV_X1 port map( A => n1347, ZN => n7041);
   U1997 : AND2_X1 port map( A1 => n4959, A2 => n1495, ZN => n1337);
   U1998 : NAND2_X1 port map( A1 => n7029, A2 => n1338, ZN => n7013);
   U1999 : NAND2_X1 port map( A1 => n7053, A2 => n7471, ZN => n1339);
   U2000 : OR2_X1 port map( A1 => n6082, A2 => n6081, ZN => n1340);
   U2001 : NAND2_X1 port map( A1 => n6826, A2 => n6594, ZN => n1341);
   U2002 : XNOR2_X1 port map( A => n5738, B => n1342, ZN => n5739);
   U2003 : XNOR2_X1 port map( A => n929, B => n5734, ZN => n1342);
   U2004 : XNOR2_X1 port map( A => n7029, B => n1343, ZN => n1348);
   U2005 : OR2_X1 port map( A1 => n7000, A2 => n7002, ZN => n1344);
   U2006 : NAND2_X1 port map( A1 => n6999, A2 => n1344, ZN => n7245);
   U2007 : OAI21_X1 port map( B1 => n1586, B2 => n6590, A => n572, ZN => n1345)
                           ;
   U2008 : OR2_X1 port map( A1 => n1732, A2 => n7003, ZN => n1346);
   U2009 : NAND2_X1 port map( A1 => n1346, A2 => n201, ZN => n6999);
   U2010 : MUX2_X2 port map( A => n4769, B => n4768, S => n2250, Z => n4935);
   U2011 : XNOR2_X1 port map( A => n1722, B => n7028, ZN => n1349);
   U2012 : INV_X1 port map( A => n680, ZN => n4596);
   U2013 : NAND2_X1 port map( A1 => n4909, A2 => n4908, ZN => n1353);
   U2014 : AND2_X1 port map( A1 => n2131, A2 => n8208, ZN => n1355);
   U2015 : AND3_X1 port map( A1 => n4568, A2 => n4569, A3 => n1355, ZN => n1550
                           );
   U2016 : XNOR2_X1 port map( A => n1357, B => n5127, ZN => n1356);
   U2017 : XOR2_X1 port map( A => n1043, B => n1801, Z => n1357);
   U2018 : AND2_X1 port map( A1 => n5701, A2 => n5702, ZN => n1359);
   U2019 : NOR2_X1 port map( A1 => n1359, A2 => n5700, ZN => n5703);
   U2020 : XNOR2_X1 port map( A => n1735, B => n4904, ZN => n1360);
   U2021 : OR2_X1 port map( A1 => n6325, A2 => n6326, ZN => n1361);
   U2022 : NAND2_X1 port map( A1 => n1361, A2 => n603, ZN => n6317);
   U2023 : OR2_X1 port map( A1 => n1718, A2 => n6316, ZN => n1362);
   U2024 : NAND2_X1 port map( A1 => n1362, A2 => n6317, ZN => n6297);
   U2025 : OR2_X1 port map( A1 => n5813, A2 => n5815, ZN => n1363);
   U2026 : NAND2_X1 port map( A1 => n5718, A2 => n1363, ZN => n5958);
   U2027 : XNOR2_X1 port map( A => n1735, B => n4904, ZN => n5122);
   U2028 : NAND2_X1 port map( A1 => n1057, A2 => n319, ZN => n4741);
   U2029 : OR2_X1 port map( A1 => n5349, A2 => n5299, ZN => n1364);
   U2030 : NAND2_X1 port map( A1 => n5210, A2 => n1364, ZN => n5344);
   U2031 : OR2_X1 port map( A1 => n5357, A2 => n5296, ZN => n1365);
   U2032 : NAND2_X1 port map( A1 => n5209, A2 => n1365, ZN => n5353);
   U2033 : OR2_X1 port map( A1 => n4973, A2 => n5030, ZN => n1366);
   U2034 : OR2_X1 port map( A1 => n4972, A2 => n5037, ZN => n1367);
   U2035 : NAND3_X1 port map( A1 => n1366, A2 => n1367, A3 => n4971, ZN => 
                           n5022);
   U2036 : MUX2_X2 port map( A => n5011, B => n5010, S => n2249, Z => n5349);
   U2037 : AND2_X1 port map( A1 => n1547, A2 => n1546, ZN => n1368);
   U2038 : XOR2_X1 port map( A => n1371, B => n1864, Z => n1370);
   U2039 : OAI33_X1 port map( A1 => n622, A2 => n5036, A3 => n2249, B1 => n5035
                           , B2 => n5034, B3 => n5033, ZN => n1371);
   U2040 : INV_X1 port map( A => n2129, ZN => n1606);
   U2041 : XOR2_X1 port map( A => n5075, B => n5087, Z => n5088);
   U2042 : AND2_X1 port map( A1 => n6780, A2 => n6779, ZN => n1372);
   U2043 : OR2_X1 port map( A1 => n5760, A2 => n5763, ZN => n1373);
   U2044 : NAND2_X1 port map( A1 => n1373, A2 => n5756, ZN => n5757);
   U2045 : AND2_X1 port map( A1 => n6763, A2 => n322, ZN => n6766);
   U2046 : MUX2_X1 port map( A => DataPath_i_PIPLIN_IN1_9_port, B => 
                           DataPath_i_PIPLIN_A_9_port, S => CU_I_n108, Z => 
                           n1374);
   U2047 : XNOR2_X1 port map( A => n5622, B => n1375, ZN => n5627);
   U2048 : XNOR2_X1 port map( A => n504, B => n5624, ZN => n1375);
   U2049 : XNOR2_X1 port map( A => n560, B => n6880, ZN => n6731);
   U2050 : XNOR2_X1 port map( A => n6731, B => n1376, ZN => n6743);
   U2051 : XNOR2_X1 port map( A => n785, B => n6049, ZN => n6051);
   U2052 : INV_X1 port map( A => n1602, ZN => n4804);
   U2054 : XNOR2_X1 port map( A => n6879, B => n6882, ZN => n6850);
   U2055 : INV_X1 port map( A => n6882, ZN => n6880);
   U2056 : NOR2_X1 port map( A1 => n5796, A2 => n875, ZN => n1377);
   U2057 : NAND2_X1 port map( A1 => n5676, A2 => n1378, ZN => n5669);
   U2058 : OAI221_X1 port map( B1 => n4953, B2 => n5191, C1 => n1579, C2 => 
                           n4952, A => n4951, ZN => n1379);
   U2059 : OAI22_X1 port map( A1 => n6020, A2 => n1646, B1 => n1008, B2 => 
                           n6019, ZN => n6106);
   U2060 : MUX2_X2 port map( A => n6940, B => n6939, S => n2243, Z => n6946);
   U2061 : XNOR2_X1 port map( A => n1380, B => n1152, ZN => n6261);
   U2063 : XNOR2_X1 port map( A => n1381, B => n1261, ZN => n1725);
   U2064 : XNOR2_X1 port map( A => n1193, B => n7025, ZN => n1381);
   U2065 : NAND2_X1 port map( A1 => n5674, A2 => n1382, ZN => n5665);
   U2066 : OAI21_X1 port map( B1 => n7045, B2 => n7044, A => n7043, ZN => n1383
                           );
   U2067 : OR2_X1 port map( A1 => n6652, A2 => n1537, ZN => n1384);
   U2068 : CLKBUF_X1 port map( A => n6635, Z => n1385);
   U2070 : INV_X1 port map( A => n1386, ZN => n1387);
   U2071 : XNOR2_X1 port map( A => n6980, B => n1388, ZN => n1678);
   U2072 : XNOR2_X1 port map( A => n1763, B => n1717, ZN => n1583);
   U2073 : AND2_X1 port map( A1 => n1236, A2 => n5319, ZN => n1390);
   U2074 : MUX2_X2 port map( A => n1392, B => n1393, S => n6495, Z => n1391);
   U2075 : OR2_X1 port map( A1 => n17162, A2 => n6115, ZN => n1394);
   U2076 : NAND2_X1 port map( A1 => n5985, A2 => n1394, ZN => n6104);
   U2077 : XNOR2_X1 port map( A => n6253, B => n1398, ZN => n1395);
   U2078 : NAND2_X1 port map( A1 => n6450, A2 => n1679, ZN => n1396);
   U2079 : OR2_X1 port map( A1 => n6583, A2 => n6634, ZN => n1397);
   U2080 : NAND2_X1 port map( A1 => n6582, A2 => n1397, ZN => n6631);
   U2081 : INV_X1 port map( A => n1131, ZN => n1398);
   U2082 : XNOR2_X1 port map( A => n1484, B => n1399, ZN => n5993);
   U2083 : AND2_X1 port map( A1 => n1105, A2 => n1494, ZN => n1399);
   U2084 : CLKBUF_X1 port map( A => n854, Z => n1401);
   U2085 : NAND2_X1 port map( A1 => n6565, A2 => n6369, ZN => n1402);
   U2086 : NAND2_X1 port map( A1 => n6564, A2 => n1702, ZN => n1403);
   U2087 : NAND2_X1 port map( A1 => n1403, A2 => n1402, ZN => n6576);
   U2088 : NAND2_X1 port map( A1 => n6688, A2 => n7771, ZN => n1404);
   U2089 : NAND2_X1 port map( A1 => n6689, A2 => n6594, ZN => n1405);
   U2090 : NAND2_X1 port map( A1 => n1404, A2 => n1405, ZN => n7006);
   U2091 : OAI21_X1 port map( B1 => n6471, B2 => n6473, A => n203, ZN => n1406)
                           ;
   U2092 : MUX2_X2 port map( A => n6533, B => n6532, S => n1702, Z => n6585);
   U2093 : INV_X1 port map( A => n1758, ZN => n4600);
   U2094 : INV_X1 port map( A => n1542, ZN => n1619);
   U2095 : OR2_X1 port map( A1 => n6403, A2 => n6360, ZN => n1409);
   U2096 : NAND2_X1 port map( A1 => n6359, A2 => n1409, ZN => n6387);
   U2097 : OR2_X1 port map( A1 => n6805, A2 => n6806, ZN => n1410);
   U2098 : OR2_X1 port map( A1 => n7030, A2 => n7014, ZN => n1411);
   U2099 : NAND2_X1 port map( A1 => n1125, A2 => n1411, ZN => n6693);
   U2100 : NAND2_X1 port map( A1 => n7014, A2 => n1412, ZN => n1413);
   U2101 : INV_X1 port map( A => n1576, ZN => n1412);
   U2102 : OAI22_X1 port map( A1 => n2229, A2 => n7244, B1 => n2227, B2 => 
                           n7243, ZN => n7014);
   U2103 : XNOR2_X1 port map( A => n1414, B => n578, ZN => n7061);
   U2104 : XNOR2_X1 port map( A => n7057, B => n7059, ZN => n1414);
   U2105 : XNOR2_X1 port map( A => n1417, B => n6666, ZN => n6676);
   U2106 : XNOR2_X1 port map( A => n6661, B => n6673, ZN => n1417);
   U2107 : INV_X1 port map( A => n882, ZN => n1418);
   U2108 : MUX2_X1 port map( A => n1748, B => n1749, S => n6594, Z => n1419);
   U2109 : MUX2_X1 port map( A => n1748, B => n1749, S => n6594, Z => n1420);
   U2110 : OR2_X1 port map( A1 => n6236, A2 => n6237, ZN => n1421);
   U2111 : NAND2_X1 port map( A1 => n1421, A2 => n6238, ZN => n6226);
   U2112 : NAND2_X1 port map( A1 => n1470, A2 => n1469, ZN => n1763);
   U2113 : NAND2_X1 port map( A1 => n1573, A2 => n1572, ZN => n6132);
   U2114 : AND2_X1 port map( A1 => n1177, A2 => n6994, ZN => n1422);
   U2115 : XNOR2_X1 port map( A => n696, B => n6171, ZN => n1592);
   U2116 : AND2_X1 port map( A1 => n6842, A2 => n1313, ZN => n1513);
   U2117 : NAND2_X1 port map( A1 => n1198, A2 => n1618, ZN => n1425);
   U2118 : NAND2_X1 port map( A1 => n1423, A2 => n1424, ZN => n1426);
   U2119 : NAND2_X1 port map( A1 => n1426, A2 => n1425, ZN => n5605);
   U2120 : INV_X1 port map( A => n613, ZN => n1423);
   U2121 : INV_X1 port map( A => n1618, ZN => n1424);
   U2122 : INV_X1 port map( A => n5599, ZN => n1618);
   U2123 : AND2_X1 port map( A1 => n729, A2 => n4949, ZN => n1427);
   U2124 : NAND2_X1 port map( A1 => n4821, A2 => n316, ZN => n4824);
   U2125 : INV_X1 port map( A => n510, ZN => n1428);
   U2126 : NAND2_X1 port map( A1 => n5438, A2 => n5439, ZN => n1659);
   U2127 : CLKBUF_X1 port map( A => n8255, Z => n1429);
   U2128 : INV_X1 port map( A => n7318, ZN => n8276);
   U2129 : XNOR2_X1 port map( A => n5708, B => n5692, ZN => n5715);
   U2130 : XNOR2_X1 port map( A => n1668, B => n1430, ZN => n5636);
   U2131 : MUX2_X1 port map( A => n2171, B => n2170, S => n2168, Z => n1711);
   U2132 : XNOR2_X1 port map( A => n4960, B => n5091, ZN => n5093);
   U2133 : XOR2_X1 port map( A => n5093, B => n5098, Z => n1824);
   U2134 : XNOR2_X1 port map( A => n4560, B => n8208, ZN => n4565);
   U2135 : XNOR2_X1 port map( A => n1248, B => n1727, ZN => n6294);
   U2136 : INV_X1 port map( A => n5815, ZN => n1431);
   U2137 : XOR2_X1 port map( A => n6095, B => n6100, Z => n1656);
   U2138 : AND2_X1 port map( A1 => n6089, A2 => n2266, ZN => n1432);
   U2139 : AND3_X1 port map( A1 => n1593, A2 => n6066, A3 => n1432, ZN => n6086
                           );
   U2140 : INV_X1 port map( A => n934, ZN => n1433);
   U2141 : XNOR2_X1 port map( A => n1434, B => n5884, ZN => n5885);
   U2142 : XOR2_X1 port map( A => n5879, B => n5827, Z => n1434);
   U2143 : XNOR2_X1 port map( A => n5072, B => n4963, ZN => n5079);
   U2144 : XOR2_X1 port map( A => n5657, B => n5658, Z => n5656);
   U2145 : XNOR2_X1 port map( A => n713, B => n5991, ZN => n5992);
   U2146 : NAND2_X1 port map( A1 => n5960, A2 => n1435, ZN => n1436);
   U2147 : NAND2_X1 port map( A1 => n5961, A2 => n1588, ZN => n1437);
   U2148 : NAND2_X1 port map( A1 => n1437, A2 => n1436, ZN => n8255);
   U2149 : INV_X1 port map( A => n1588, ZN => n1435);
   U2150 : INV_X1 port map( A => n526, ZN => n1438);
   U2151 : INV_X1 port map( A => n2267, ZN => n1588);
   U2152 : CLKBUF_X1 port map( A => n510, Z => n1439);
   U2153 : NAND2_X1 port map( A1 => n563, A2 => n1441, ZN => n1443);
   U2154 : NAND2_X1 port map( A1 => n6189, A2 => n1443, ZN => n6263);
   U2155 : INV_X1 port map( A => n6271, ZN => n1441);
   U2156 : INV_X1 port map( A => n6272, ZN => n1442);
   U2157 : OR2_X1 port map( A1 => n664, A2 => n5548, ZN => n1444);
   U2158 : INV_X1 port map( A => n5987, ZN => n1445);
   U2159 : AND2_X1 port map( A1 => n1669, A2 => n1670, ZN => n1446);
   U2160 : XOR2_X1 port map( A => n1332, B => n1865, Z => n1447);
   U2161 : OR2_X1 port map( A1 => n6840, A2 => n6842, ZN => n7400);
   U2162 : OR2_X1 port map( A1 => n4728, A2 => n4673, ZN => n1448);
   U2163 : NAND2_X1 port map( A1 => n1448, A2 => n4672, ZN => n4674);
   U2164 : INV_X1 port map( A => n1372, ZN => n1449);
   U2165 : OR2_X1 port map( A1 => n4709, A2 => n4684, ZN => n1450);
   U2166 : NAND2_X1 port map( A1 => n1450, A2 => n4683, ZN => n4704);
   U2167 : OR2_X1 port map( A1 => n4715, A2 => n4681, ZN => n1451);
   U2168 : NAND2_X1 port map( A1 => n1451, A2 => n4680, ZN => n4711);
   U2169 : AND2_X1 port map( A1 => n1876, A2 => n6778, ZN => n1452);
   U2170 : AND2_X1 port map( A1 => n1877, A2 => n1210, ZN => n1453);
   U2171 : NOR3_X1 port map( A1 => n1452, A2 => n1453, A3 => n6777, ZN => n6779
                           );
   U2172 : XOR2_X1 port map( A => n517, B => n1798, Z => n1454);
   U2173 : MUX2_X2 port map( A => n5766, B => n5765, S => n2250, Z => n6736);
   U2175 : OR2_X1 port map( A1 => n1084, A2 => n1814, ZN => n1582);
   U2176 : XNOR2_X1 port map( A => n1456, B => n5136, ZN => n5139);
   U2177 : NAND2_X1 port map( A1 => n574, A2 => n315, ZN => n6786);
   U2178 : OR2_X1 port map( A1 => n5827, A2 => n5879, ZN => n1457);
   U2179 : NAND2_X1 port map( A1 => n5826, A2 => n1457, ZN => n5866);
   U2180 : XNOR2_X1 port map( A => n952, B => n5829, ZN => n1667);
   U2181 : AND2_X1 port map( A1 => n5155, A2 => n5154, ZN => n5141);
   U2182 : NAND2_X1 port map( A1 => n6505, A2 => n6515, ZN => n1458);
   U2183 : NAND2_X1 port map( A1 => n1459, A2 => n1458, ZN => n1479);
   U2184 : XNOR2_X1 port map( A => n1460, B => n6674, ZN => n6675);
   U2185 : OR2_X1 port map( A1 => n4955, A2 => n4954, ZN => n1461);
   U2186 : NAND2_X1 port map( A1 => n4916, A2 => n1461, ZN => n5092);
   U2187 : OR2_X1 port map( A1 => n5569, A2 => n471, ZN => n1462);
   U2188 : NAND2_X1 port map( A1 => n5525, A2 => n1462, ZN => n5560);
   U2189 : XNOR2_X1 port map( A => n7469, B => n7470, ZN => n1463);
   U2190 : OR2_X1 port map( A1 => n5562, A2 => n5561, ZN => n1464);
   U2191 : NAND2_X1 port map( A1 => n5527, A2 => n1464, ZN => n5795);
   U2192 : OR2_X1 port map( A1 => n4918, A2 => n1611, ZN => n1465);
   U2193 : NAND2_X1 port map( A1 => n4917, A2 => n1465, ZN => n5067);
   U2194 : MUX2_X2 port map( A => n4796, B => n4795, S => n804, Z => n4954);
   U2195 : MUX2_X2 port map( A => n7468, B => n7467, S => n7712, Z => n7469);
   U2196 : XNOR2_X1 port map( A => n1475, B => n1468, ZN => n6504);
   U2197 : NAND2_X1 port map( A1 => n1765, A2 => n6495, ZN => n1469);
   U2198 : NAND2_X1 port map( A1 => n1764, A2 => n7835, ZN => n1470);
   U2199 : OAI21_X1 port map( B1 => n1744, B2 => n5831, A => n5830, ZN => n1471
                           );
   U2200 : XNOR2_X1 port map( A => n1729, B => n7417, ZN => n1472);
   U2201 : XNOR2_X1 port map( A => n1473, B => n856, ZN => n5678);
   U2202 : XNOR2_X1 port map( A => n600, B => n5824, ZN => n5889);
   U2203 : INV_X1 port map( A => n1513, ZN => n7279);
   U2204 : XNOR2_X1 port map( A => n6235, B => n1474, ZN => n6240);
   U2205 : XNOR2_X1 port map( A => n6234, B => n6233, ZN => n1474);
   U2206 : XNOR2_X1 port map( A => n1182, B => n6590, ZN => n1610);
   U2207 : AOI21_X1 port map( B1 => n7426, B2 => n947, A => n1832, ZN => n6985)
                           ;
   U2208 : OR2_X1 port map( A1 => n6501, A2 => n1094, ZN => n1476);
   U2209 : NAND2_X1 port map( A1 => n6466, A2 => n1476, ZN => n6800);
   U2210 : OR2_X1 port map( A1 => n1718, A2 => n6319, ZN => n1477);
   U2211 : NAND2_X1 port map( A1 => n1477, A2 => n6318, ZN => n6303);
   U2212 : OR2_X1 port map( A1 => n6323, A2 => n6326, ZN => n1478);
   U2213 : NAND2_X1 port map( A1 => n1478, A2 => n6211, ZN => n6318);
   U2214 : OR2_X1 port map( A1 => n6677, A2 => n6681, ZN => n6663);
   U2215 : XOR2_X1 port map( A => n6516, B => n1479, Z => n6517);
   U2216 : INV_X1 port map( A => n8241, ZN => n1480);
   U2218 : OR2_X1 port map( A1 => n5045, A2 => n5046, ZN => n1482);
   U2219 : NAND2_X1 port map( A1 => n5047, A2 => n1482, ZN => n4923);
   U2220 : OR2_X1 port map( A1 => n5829, A2 => n952, ZN => n1483);
   U2221 : XNOR2_X1 port map( A => n5987, B => n5990, ZN => n1484);
   U2222 : NAND3_X1 port map( A1 => n6162, A2 => n6159, A3 => n341, ZN => n6161
                           );
   U2223 : AND2_X1 port map( A1 => n6009, A2 => n1557, ZN => n1485);
   U2224 : XOR2_X1 port map( A => n6037, B => n6049, Z => n6052);
   U2226 : XNOR2_X1 port map( A => n1133, B => n6574, ZN => n6620);
   U2227 : OR2_X1 port map( A1 => n6403, A2 => n6406, ZN => n1486);
   U2228 : NAND2_X1 port map( A1 => n6338, A2 => n1486, ZN => n6379);
   U2229 : OR2_X1 port map( A1 => n6346, A2 => n780, ZN => n1487);
   U2230 : NAND2_X1 port map( A1 => n6334, A2 => n1487, ZN => n6433);
   U2231 : OR2_X1 port map( A1 => n6421, A2 => n6410, ZN => n1489);
   U2232 : CLKBUF_X1 port map( A => n6441, Z => n1490);
   U2233 : CLKBUF_X1 port map( A => n7033, Z => n1491);
   U2234 : NAND2_X1 port map( A1 => n2163, A2 => n5812, ZN => n1493);
   U2235 : NAND2_X2 port map( A1 => n609, A2 => n7109, ZN => n8089);
   U2236 : OR2_X1 port map( A1 => n5868, A2 => n951, ZN => n1494);
   U2237 : NAND2_X1 port map( A1 => n1105, A2 => n1494, ZN => n5988);
   U2238 : OR2_X1 port map( A1 => n5091, A2 => n4960, ZN => n1495);
   U2239 : NAND2_X1 port map( A1 => n4959, A2 => n1495, ZN => n5075);
   U2240 : OR2_X1 port map( A1 => n5052, A2 => n5053, ZN => n1497);
   U2241 : NAND3_X1 port map( A1 => n1496, A2 => n1497, A3 => n4965, ZN => 
                           n5048);
   U2242 : OR2_X1 port map( A1 => n1408, A2 => n7054, ZN => n1498);
   U2243 : NAND2_X1 port map( A1 => n1498, A2 => n1383, ZN => n7046);
   U2244 : AND2_X1 port map( A1 => n6834, A2 => n859, ZN => n6697);
   U2246 : XNOR2_X1 port map( A => n1499, B => n5079, ZN => n5082);
   U2247 : NAND2_X1 port map( A1 => n5074, A2 => n5073, ZN => n1499);
   U2248 : MUX2_X2 port map( A => n5082, B => n5081, S => n2248, Z => n5405);
   U2249 : XNOR2_X1 port map( A => n6041, B => n6040, ZN => n1500);
   U2250 : OR2_X1 port map( A1 => n5818, A2 => n5936, ZN => n1501);
   U2251 : NAND2_X1 port map( A1 => n5817, A2 => n1501, ZN => n5929);
   U2252 : AND2_X1 port map( A1 => n6976, A2 => n1447, ZN => n1502);
   U2253 : XNOR2_X1 port map( A => n1504, B => n1503, ZN => n6798);
   U2254 : XNOR2_X1 port map( A => n6977, B => n6976, ZN => n1504);
   U2255 : XOR2_X1 port map( A => n6836, B => n1879, Z => n6840);
   U2256 : XNOR2_X1 port map( A => n6113, B => n1505, ZN => n6117);
   U2258 : XNOR2_X1 port map( A => n7019, B => n7022, ZN => n1631);
   U2259 : XNOR2_X1 port map( A => n1263, B => n6683, ZN => n1559);
   U2260 : XNOR2_X1 port map( A => n1628, B => n1506, ZN => n6431);
   U2261 : XNOR2_X1 port map( A => n6430, B => n1032, ZN => n1506);
   U2262 : OR2_X1 port map( A1 => n5588, A2 => n896, ZN => n1508);
   U2263 : NAND2_X1 port map( A1 => n5524, A2 => n1508, ZN => n5566);
   U2264 : OR2_X1 port map( A1 => n6041, A2 => n5836, ZN => n1509);
   U2265 : NAND2_X1 port map( A1 => n1509, A2 => n5835, ZN => n6945);
   U2266 : OAI221_X1 port map( B1 => n5841, B2 => n5840, C1 => n5839, C2 => 
                           n6776, A => n5838, ZN => n1510);
   U2267 : XNOR2_X1 port map( A => n6397, B => n1511, ZN => n6398);
   U2268 : XNOR2_X1 port map( A => n1512, B => n1152, ZN => n6260);
   U2269 : XNOR2_X1 port map( A => n6259, B => n6258, ZN => n1512);
   U2270 : XNOR2_X1 port map( A => n776, B => n6176, ZN => n6179);
   U2272 : XNOR2_X1 port map( A => n1389, B => n6237, ZN => n1591);
   U2273 : INV_X1 port map( A => n5897, ZN => n1514);
   U2274 : MUX2_X2 port map( A => n1678, B => n1677, S => n529, Z => n1676);
   U2275 : NAND2_X1 port map( A1 => n6104, A2 => n1515, ZN => n5986);
   U2276 : AND2_X1 port map( A1 => n1551, A2 => n1067, ZN => n1516);
   U2277 : NAND2_X1 port map( A1 => n1617, A2 => n4532, ZN => n1518);
   U2278 : OR2_X2 port map( A1 => n1518, A2 => n1519, ZN => n4522);
   U2279 : OR2_X1 port map( A1 => n4457, A2 => n4456, ZN => n1519);
   U2280 : INV_X1 port map( A => n8045, ZN => n1520);
   U2281 : NAND2_X1 port map( A1 => n7454, A2 => n7771, ZN => n1521);
   U2282 : NAND2_X1 port map( A1 => n7455, A2 => n6594, ZN => n1522);
   U2283 : NAND2_X1 port map( A1 => n1521, A2 => n1522, ZN => n7456);
   U2284 : INV_X1 port map( A => n8045, ZN => n2237);
   U2285 : OR2_X1 port map( A1 => n6151, A2 => n670, ZN => n1523);
   U2286 : NAND2_X1 port map( A1 => n5967, A2 => n1523, ZN => n6143);
   U2287 : NOR2_X1 port map( A1 => n8128, A2 => n8130, ZN => n1524);
   U2288 : NOR2_X1 port map( A1 => n8129, A2 => n8128, ZN => n1525);
   U2289 : NOR2_X1 port map( A1 => n663, A2 => n8130, ZN => n1526);
   U2290 : OR2_X1 port map( A1 => n4790, A2 => n4660, ZN => n1527);
   U2291 : NAND2_X1 port map( A1 => n4793, A2 => n1527, ZN => n4661);
   U2292 : OR2_X1 port map( A1 => n4784, A2 => n4665, ZN => n1528);
   U2293 : NAND2_X1 port map( A1 => n1528, A2 => n4664, ZN => n4779);
   U2294 : OR2_X1 port map( A1 => n4791, A2 => n4662, ZN => n1529);
   U2295 : NAND2_X1 port map( A1 => n4661, A2 => n1529, ZN => n4786);
   U2296 : INV_X1 port map( A => n1170, ZN => n1530);
   U2297 : NAND2_X1 port map( A1 => n5355, A2 => n936, ZN => n1531);
   U2298 : MUX2_X1 port map( A => n5161, B => n5160, S => n2247, Z => n1532);
   U2299 : OR2_X1 port map( A1 => n5928, A2 => n5927, ZN => n1534);
   U2300 : NAND2_X1 port map( A1 => n5929, A2 => n1534, ZN => n5819);
   U2302 : MUX2_X1 port map( A => n265, B => n4303, S => n547, Z => n8045);
   U2303 : XNOR2_X1 port map( A => n5585, B => n1535, ZN => n5591);
   U2304 : XNOR2_X1 port map( A => n896, B => n5588, ZN => n1535);
   U2305 : XNOR2_X1 port map( A => n5908, B => n5909, ZN => n1538);
   U2306 : AND2_X1 port map( A1 => n832, A2 => n4943, ZN => n1539);
   U2307 : INV_X1 port map( A => n7063, ZN => n1541);
   U2308 : MUX2_X1 port map( A => n5161, B => n5160, S => n2247, Z => n8151);
   U2309 : MUX2_X1 port map( A => n1543, B => n1544, S => CU_I_n108, Z => n1542
                           );
   U2310 : AND2_X1 port map( A1 => n4588, A2 => n4587, ZN => n1564);
   U2311 : OR2_X1 port map( A1 => n4790, A2 => n4791, ZN => n1545);
   U2312 : NAND2_X1 port map( A1 => n4792, A2 => n1545, ZN => n4607);
   U2313 : OR2_X1 port map( A1 => n4663, A2 => n4665, ZN => n1546);
   U2314 : OR2_X1 port map( A1 => n4660, A2 => n4662, ZN => n1547);
   U2315 : NAND2_X1 port map( A1 => n4607, A2 => n1547, ZN => n4785);
   U2316 : XOR2_X1 port map( A => n6249, B => n6254, Z => n6257);
   U2317 : INV_X2 port map( A => n2237, ZN => n2236);
   U2318 : OAI221_X1 port map( B1 => n1863, B2 => n310, C1 => n1863, C2 => 
                           n7297, A => n6897, ZN => n6911);
   U2319 : NAND2_X1 port map( A1 => n7064, A2 => n7581, ZN => n1548);
   U2320 : OAI21_X1 port map( B1 => n4565, B2 => n554, A => n4564, ZN => n1549)
                           ;
   U2321 : NAND2_X1 port map( A1 => n6568, A2 => n1551, ZN => n6630);
   U2322 : OR2_X1 port map( A1 => n5818, A2 => n5943, ZN => n1553);
   U2323 : NAND2_X1 port map( A1 => n5720, A2 => n1553, ZN => n5926);
   U2324 : OR2_X1 port map( A1 => n670, A2 => n6160, ZN => n1554);
   U2325 : NAND2_X1 port map( A1 => n6007, A2 => n1554, ZN => n6144);
   U2326 : OR2_X1 port map( A1 => n6436, A2 => n6354, ZN => n1555);
   U2327 : OR2_X1 port map( A1 => n1888, A2 => n6448, ZN => n1556);
   U2328 : NAND2_X1 port map( A1 => n1163, A2 => n1556, ZN => n6425);
   U2329 : OR2_X1 port map( A1 => n6142, A2 => n17163, ZN => n1557);
   U2330 : NAND2_X1 port map( A1 => n6009, A2 => n1557, ZN => n6011);
   U2331 : XNOR2_X1 port map( A => n6617, B => n1558, ZN => n1868);
   U2332 : XNOR2_X1 port map( A => n1133, B => n6574, ZN => n1558);
   U2333 : XNOR2_X1 port map( A => n482, B => n1559, ZN => n1640);
   U2334 : XNOR2_X1 port map( A => n6407, B => n1560, ZN => n6408);
   U2335 : XNOR2_X1 port map( A => n1660, B => n7010, ZN => n7034);
   U2336 : XNOR2_X1 port map( A => n5266, B => n5265, ZN => n5237);
   U2337 : XNOR2_X1 port map( A => n1561, B => n921, ZN => n7481);
   U2338 : XNOR2_X1 port map( A => n5910, B => n1562, ZN => n5911);
   U2339 : NAND2_X1 port map( A1 => n605, A2 => n5907, ZN => n1562);
   U2340 : XNOR2_X1 port map( A => n1061, B => n6105, ZN => n6111);
   U2341 : XNOR2_X1 port map( A => n1675, B => n1563, ZN => n1665);
   U2342 : NAND2_X1 port map( A1 => n7021, A2 => n7020, ZN => n1563);
   U2343 : CLKBUF_X1 port map( A => n6834, Z => n1565);
   U2344 : INV_X1 port map( A => n4541, ZN => n1566);
   U2345 : OR2_X1 port map( A1 => n5122, A2 => n5145, ZN => n1568);
   U2346 : XOR2_X2 port map( A => n4859, B => n4858, Z => n4904);
   U2347 : XNOR2_X1 port map( A => n1570, B => n5980, ZN => n5981);
   U2348 : XOR2_X1 port map( A => n5979, B => n935, Z => n1570);
   U2349 : NAND2_X1 port map( A1 => n5911, A2 => n1571, ZN => n1572);
   U2350 : NAND2_X1 port map( A1 => n5912, A2 => n1584, ZN => n1573);
   U2351 : INV_X1 port map( A => n1584, ZN => n1571);
   U2352 : OR2_X1 port map( A1 => n6197, A2 => n6221, ZN => n1574);
   U2353 : NAND2_X1 port map( A1 => n6249, A2 => n1574, ZN => n6193);
   U2354 : OR2_X1 port map( A1 => n6205, A2 => n6328, ZN => n1575);
   U2355 : NAND2_X1 port map( A1 => n1575, A2 => n6327, ZN => n6185);
   U2356 : INV_X1 port map( A => n1732, ZN => n7002);
   U2357 : MUX2_X1 port map( A => n6181, B => n6180, S => n2265, Z => n1577);
   U2358 : XNOR2_X1 port map( A => n880, B => n6793, ZN => n6342);
   U2359 : INV_X1 port map( A => n4830, ZN => n1579);
   U2361 : CLKBUF_X1 port map( A => n1577, Z => n1581);
   U2362 : MUX2_X1 port map( A => n6181, B => n6180, S => n2265, Z => n8238);
   U2363 : XNOR2_X1 port map( A => n1582, B => n6794, ZN => n6799);
   U2364 : XNOR2_X1 port map( A => n1583, B => n7451, ZN => n1748);
   U2365 : AND2_X1 port map( A1 => CU_I_n108, A2 => DataPath_i_PIPLIN_A_3_port,
                           ZN => n4450);
   U2366 : XNOR2_X1 port map( A => n1301, B => n7000, ZN => n6817);
   U2367 : XNOR2_X1 port map( A => n619, B => n6363, ZN => n1595);
   U2368 : XNOR2_X1 port map( A => n6509, B => n1585, ZN => n6518);
   U2369 : XNOR2_X1 port map( A => n850, B => n6515, ZN => n1585);
   U2370 : INV_X1 port map( A => n6598, ZN => n1586);
   U2371 : OR2_X1 port map( A1 => n5091, A2 => n5090, ZN => n1587);
   U2372 : NAND2_X1 port map( A1 => n5092, A2 => n1587, ZN => n5085);
   U2373 : XNOR2_X1 port map( A => n6562, B => n1406, ZN => n6565);
   U2374 : XNOR2_X1 port map( A => n868, B => n6215, ZN => n6278);
   U2375 : XNOR2_X1 port map( A => n6278, B => n6285, ZN => n6286);
   U2376 : XNOR2_X1 port map( A => n204, B => n1589, ZN => n1757);
   U2377 : XNOR2_X1 port map( A => n6255, B => n6254, ZN => n6256);
   U2378 : XNOR2_X1 port map( A => n1590, B => n6386, ZN => n6395);
   U2379 : XNOR2_X1 port map( A => n958, B => n6392, ZN => n1590);
   U2380 : XNOR2_X1 port map( A => n6645, B => n718, ZN => n6659);
   U2381 : XNOR2_X1 port map( A => n1682, B => n5805, ZN => n5858);
   U2382 : AND3_X1 port map( A1 => n6053, A2 => n6075, A3 => n6054, ZN => n5994
                           );
   U2383 : XNOR2_X1 port map( A => n6238, B => n1591, ZN => n6239);
   U2384 : XNOR2_X1 port map( A => n1592, B => n6170, ZN => n6174);
   U2385 : NAND2_X1 port map( A1 => n6098, A2 => n6084, ZN => n1593);
   U2386 : INV_X1 port map( A => n783, ZN => n1594);
   U2387 : XNOR2_X1 port map( A => n1595, B => n6393, ZN => n6394);
   U2388 : XNOR2_X1 port map( A => n6011, B => n1596, ZN => n1720);
   U2389 : XNOR2_X1 port map( A => n6748, B => n6853, ZN => n6749);
   U2390 : MUX2_X2 port map( A => n6445, B => n6444, S => n7973, Z => n6469);
   U2391 : XNOR2_X1 port map( A => n5889, B => n1597, ZN => n5891);
   U2392 : NAND2_X1 port map( A1 => n588, A2 => n5872, ZN => n1597);
   U2393 : XNOR2_X1 port map( A => n6135, B => n1598, ZN => n6137);
   U2394 : INV_X1 port map( A => n1415, ZN => n1599);
   U2395 : AND2_X1 port map( A1 => n5386, A2 => n5385, ZN => n1600);
   U2396 : AND2_X1 port map( A1 => n571, A2 => n6084, ZN => n1601);
   U2397 : XNOR2_X1 port map( A => n17251, B => n5920, ZN => n1629);
   U2398 : AND2_X1 port map( A1 => n1839, A2 => n4809, ZN => n1602);
   U2399 : OR2_X1 port map( A1 => n461, A2 => n6136, ZN => n6120);
   U2400 : XNOR2_X1 port map( A => n5560, B => n1603, ZN => n1683);
   U2401 : XNOR2_X1 port map( A => n17183, B => n5809, ZN => n5916);
   U2402 : XNOR2_X1 port map( A => n5976, B => n5916, ZN => n5917);
   U2403 : OR2_X1 port map( A1 => n4624, A2 => n4733, ZN => n4670);
   U2404 : XNOR2_X1 port map( A => n5563, B => n1604, ZN => n5564);
   U2405 : XNOR2_X1 port map( A => n1605, B => n816, ZN => n5404);
   U2406 : XNOR2_X1 port map( A => n17214, B => n5401, ZN => n1605);
   U2407 : AND2_X1 port map( A1 => n5721, A2 => n1714, ZN => n1608);
   U2408 : AND2_X1 port map( A1 => n5721, A2 => n1714, ZN => n1609);
   U2409 : XNOR2_X1 port map( A => n1610, B => n6597, ZN => n6602);
   U2410 : INV_X1 port map( A => n1064, ZN => n1611);
   U2411 : INV_X1 port map( A => n1676, ZN => n7432);
   U2412 : OR2_X1 port map( A1 => n546, A2 => n8188, ZN => n4894);
   U2413 : XNOR2_X1 port map( A => n5399, B => n5402, ZN => n5403);
   U2414 : NAND2_X1 port map( A1 => n632, A2 => n1612, ZN => n1613);
   U2415 : NAND2_X1 port map( A1 => n1613, A2 => n1781, ZN => n6691);
   U2416 : INV_X1 port map( A => n7705, ZN => n1612);
   U2417 : CLKBUF_X1 port map( A => n6636, Z => n1615);
   U2418 : OR2_X1 port map( A1 => n1580, A2 => n6629, ZN => n1616);
   U2419 : NAND2_X1 port map( A1 => n6584, A2 => n1616, ZN => n6624);
   U2420 : INV_X1 port map( A => n1536, ZN => n7012);
   U2421 : XNOR2_X1 port map( A => n6525, B => n6483, ZN => n1653);
   U2422 : INV_X1 port map( A => n1753, ZN => n5818);
   U2423 : INV_X1 port map( A => n1651, ZN => n6623);
   U2424 : INV_X1 port map( A => n1689, ZN => n6583);
   U2425 : XOR2_X1 port map( A => n5042, B => n5028, Z => n5043);
   U2426 : XNOR2_X1 port map( A => n6573, B => n6829, ZN => n6593);
   U2427 : XNOR2_X1 port map( A => n1620, B => n5788, ZN => n5316);
   U2428 : XNOR2_X1 port map( A => n5241, B => n5787, ZN => n1620);
   U2429 : AND2_X1 port map( A1 => n5164, A2 => n1288, ZN => n1621);
   U2430 : AND2_X1 port map( A1 => n6223, A2 => n6222, ZN => n6225);
   U2431 : OR2_X1 port map( A1 => n1389, A2 => n6233, ZN => n1622);
   U2432 : NAND2_X1 port map( A1 => n6226, A2 => n1622, ZN => n6227);
   U2433 : OAI21_X1 port map( B1 => n6920, B2 => n5316, A => n5315, ZN => n5797
                           );
   U2434 : XNOR2_X1 port map( A => n6433, B => n6355, ZN => n6434);
   U2435 : XNOR2_X1 port map( A => n1623, B => n5956, ZN => n2171);
   U2436 : XNOR2_X1 port map( A => n1635, B => n1624, ZN => n6432);
   U2437 : XOR2_X1 port map( A => n1031, B => n6430, Z => n1624);
   U2438 : XNOR2_X1 port map( A => n5921, B => n5820, ZN => n5922);
   U2439 : XNOR2_X1 port map( A => n1625, B => n692, ZN => n6147);
   U2440 : XNOR2_X1 port map( A => n6010, B => n6145, ZN => n1625);
   U2441 : XNOR2_X1 port map( A => n1626, B => n6527, ZN => n6533);
   U2442 : XNOR2_X1 port map( A => n222, B => n6449, ZN => n6454);
   U2443 : XNOR2_X1 port map( A => n1627, B => n1644, ZN => n6230);
   U2444 : XNOR2_X1 port map( A => n1323, B => n6695, ZN => n1627);
   U2445 : XNOR2_X1 port map( A => n6983, B => n6984, ZN => n6803);
   U2446 : XNOR2_X1 port map( A => n6375, B => n980, ZN => n6376);
   U2447 : INV_X1 port map( A => n839, ZN => n7009);
   U2448 : NAND2_X1 port map( A1 => n6427, A2 => n6428, ZN => n1628);
   U2449 : XNOR2_X1 port map( A => n6010, B => n6145, ZN => n1721);
   U2450 : XNOR2_X1 port map( A => n6622, B => n1103, ZN => n6628);
   U2451 : XNOR2_X1 port map( A => n6103, B => n6108, ZN => n6109);
   U2452 : XNOR2_X1 port map( A => n6109, B => n6106, ZN => n6110);
   U2453 : XNOR2_X1 port map( A => n1629, B => n1609, ZN => n5923);
   U2454 : XNOR2_X1 port map( A => n6228, B => n6227, ZN => n6229);
   U2455 : XNOR2_X1 port map( A => n6823, B => n6822, ZN => n6645);
   U2456 : INV_X1 port map( A => n6366, ZN => n6796);
   U2457 : XNOR2_X1 port map( A => n1510, B => n6784, ZN => n6033);
   U2458 : XNOR2_X1 port map( A => n6733, B => n6736, ZN => n5775);
   U2459 : XNOR2_X1 port map( A => n1170, B => n5274, ZN => n5461);
   U2460 : XNOR2_X1 port map( A => n1159, B => n6809, ZN => n6573);
   U2461 : XNOR2_X1 port map( A => n616, B => n6822, ZN => n1761);
   U2462 : INV_X1 port map( A => n1106, ZN => n6032);
   U2463 : XNOR2_X1 port map( A => n585, B => n6994, ZN => n6813);
   U2464 : XNOR2_X1 port map( A => n1632, B => n1631, ZN => n1666);
   U2465 : NAND2_X1 port map( A1 => n7459, A2 => n7460, ZN => n1632);
   U2466 : XNOR2_X1 port map( A => n1030, B => n7487, ZN => n1633);
   U2467 : BUF_X1 port map( A => n5856, Z => n1682);
   U2468 : XNOR2_X1 port map( A => n504, B => n5624, ZN => n5625);
   U2469 : XNOR2_X1 port map( A => n1181, B => n6599, ZN => n6600);
   U2470 : XNOR2_X1 port map( A => n1633, B => n7073, ZN => n7074);
   U2471 : XNOR2_X1 port map( A => n5929, B => n1634, ZN => n5930);
   U2472 : XNOR2_X1 port map( A => n660, B => n5927, ZN => n1634);
   U2473 : NAND2_X1 port map( A1 => n6425, A2 => n6426, ZN => n1635);
   U2474 : OAI22_X2 port map( A1 => n2230, A2 => n7316, B1 => n1242, B2 => 
                           n2227, ZN => n5145);
   U2475 : AND2_X1 port map( A1 => n8199, A2 => n1878, ZN => n1636);
   U2476 : OR2_X1 port map( A1 => n6684, A2 => n1537, ZN => n1637);
   U2477 : OR2_X1 port map( A1 => n566, A2 => n6683, ZN => n1638);
   U2478 : NAND2_X1 port map( A1 => n482, A2 => n1638, ZN => n6667);
   U2479 : OAI21_X1 port map( B1 => n4566, B2 => n4565, A => n4564, ZN => n8199
                           );
   U2480 : XNOR2_X1 port map( A => n6474, B => n6560, ZN => n6562);
   U2481 : XNOR2_X1 port map( A => n991, B => n1874, ZN => n1641);
   U2482 : XNOR2_X1 port map( A => n6520, B => n1643, ZN => n1756);
   U2483 : XNOR2_X1 port map( A => n6519, B => n6522, ZN => n1643);
   U2484 : NOR2_X1 port map( A1 => n1352, A2 => n5955, ZN => n1645);
   U2485 : AND2_X1 port map( A1 => n6018, A2 => n6017, ZN => n1646);
   U2486 : XNOR2_X1 port map( A => n5066, B => n4935, ZN => n5069);
   U2487 : XNOR2_X1 port map( A => n5861, B => n591, ZN => n5862);
   U2488 : INV_X1 port map( A => n1420, ZN => n7464);
   U2489 : XNOR2_X1 port map( A => n778, B => n5289, ZN => n5382);
   U2490 : XNOR2_X1 port map( A => n5633, B => n664, ZN => n5634);
   U2491 : OR2_X1 port map( A1 => n6145, A2 => n17163, ZN => n1648);
   U2492 : NAND2_X1 port map( A1 => n5354, A2 => n2245, ZN => n1649);
   U2493 : NAND2_X1 port map( A1 => n1531, A2 => n890, ZN => n5593);
   U2494 : OAI21_X1 port map( B1 => n214, B2 => n1849, A => n6506, ZN => n1650)
                           ;
   U2495 : MUX2_X2 port map( A => n1652, B => n1653, S => n1702, Z => n1651);
   U2496 : XNOR2_X1 port map( A => n6525, B => n214, ZN => n1652);
   U2497 : XNOR2_X1 port map( A => n1654, B => n5865, ZN => n5870);
   U2498 : XNOR2_X1 port map( A => n951, B => n5868, ZN => n1654);
   U2499 : INV_X1 port map( A => n4570, ZN => n4561);
   U2500 : OR2_X1 port map( A1 => n1836, A2 => n694, ZN => n1658);
   U2501 : XNOR2_X1 port map( A => n942, B => n5707, ZN => n5708);
   U2502 : MUX2_X1 port map( A => n207, B => n436, S => n7771, Z => n1655);
   U2503 : XNOR2_X1 port map( A => n826, B => n1656, ZN => n6101);
   U2504 : OR2_X1 port map( A1 => n706, A2 => n5546, ZN => n1657);
   U2505 : NAND2_X1 port map( A1 => n5545, A2 => n1657, ZN => n5631);
   U2506 : XNOR2_X1 port map( A => n237, B => n1630, ZN => n1675);
   U2507 : XNOR2_X1 port map( A => n6083, B => n1398, ZN => n6197);
   U2508 : XNOR2_X1 port map( A => n1658, B => n5366, ZN => n5372);
   U2509 : XNOR2_X1 port map( A => n1176, B => n1659, ZN => n5448);
   U2510 : XNOR2_X1 port map( A => n1728, B => n695, ZN => n1662);
   U2511 : INV_X1 port map( A => n934, ZN => n5978);
   U2512 : XNOR2_X1 port map( A => n6694, B => n6695, ZN => n6228);
   U2513 : XNOR2_X1 port map( A => n17156, B => n7478, ZN => n1663);
   U2514 : XNOR2_X1 port map( A => n1663, B => n7472, ZN => n7050);
   U2515 : INV_X1 port map( A => n1142, ZN => n7047);
   U2516 : XNOR2_X1 port map( A => n17250, B => n5920, ZN => n5921);
   U2518 : XNOR2_X1 port map( A => n5139, B => n5141, ZN => n5142);
   U2519 : XNOR2_X1 port map( A => n1667, B => n1277, ZN => n5869);
   U2520 : NAND2_X1 port map( A1 => n5629, A2 => n5630, ZN => n1668);
   U2521 : NAND2_X1 port map( A1 => n6034, A2 => n2266, ZN => n1669);
   U2522 : NAND2_X1 port map( A1 => n6035, A2 => n750, ZN => n1670);
   U2523 : NAND2_X1 port map( A1 => n755, A2 => n1670, ZN => n6694);
   U2524 : INV_X1 port map( A => n1655, ZN => n1672);
   U2525 : XNOR2_X1 port map( A => n933, B => n5896, ZN => n5895);
   U2526 : XNOR2_X1 port map( A => n6613, B => n580, ZN => n6614);
   U2527 : XNOR2_X1 port map( A => n1673, B => n7489, ZN => n1871);
   U2528 : XNOR2_X1 port map( A => n1905, B => n1463, ZN => n1673);
   U2529 : XNOR2_X1 port map( A => n6133, B => n6134, ZN => n6138);
   U2530 : XNOR2_X1 port map( A => n6398, B => n1674, ZN => n6402);
   U2531 : NAND2_X1 port map( A1 => n652, A2 => n606, ZN => n1674);
   U2532 : XNOR2_X1 port map( A => n6467, B => n989, ZN => n6494);
   U2533 : XNOR2_X1 port map( A => n6991, B => n6591, ZN => n6592);
   U2534 : MUX2_X2 port map( A => n1823, B => n1824, S => n2248, Z => n1822);
   U2535 : XNOR2_X1 port map( A => n5855, B => n1671, ZN => n6027);
   U2536 : XNOR2_X1 port map( A => n202, B => n599, ZN => n6825);
   U2537 : XNOR2_X1 port map( A => n4910, B => n4938, ZN => n4939);
   U2538 : XNOR2_X1 port map( A => n1472, B => n6973, ZN => n1677);
   U2539 : OR2_X1 port map( A1 => n909, A2 => n6451, ZN => n1679);
   U2540 : NAND2_X1 port map( A1 => n6450, A2 => n1679, ZN => n6427);
   U2541 : OR2_X1 port map( A1 => n5099, A2 => n5100, ZN => n1680);
   U2542 : NAND2_X1 port map( A1 => n1228, A2 => n1680, ZN => n4916);
   U2543 : XNOR2_X1 port map( A => n1683, B => n5561, ZN => n5565);
   U2544 : XOR2_X1 port map( A => n6042, B => n5844, Z => n1686);
   U2545 : OR2_X1 port map( A1 => n6237, A2 => n1389, ZN => n1687);
   U2546 : OR2_X1 port map( A1 => n6114, A2 => n6019, ZN => n1688);
   U2547 : NAND2_X1 port map( A1 => n6113, A2 => n1688, ZN => n5985);
   U2548 : XNOR2_X1 port map( A => n6541, B => n6542, ZN => n1690);
   U2549 : XNOR2_X1 port map( A => n6550, B => n6549, ZN => n1691);
   U2551 : AND2_X1 port map( A1 => n6609, A2 => n6610, ZN => n1692);
   U2552 : XNOR2_X1 port map( A => n862, B => n6982, ZN => n1698);
   U2553 : AND2_X1 port map( A1 => n1226, A2 => n339, ZN => n1694);
   U2554 : AND2_X1 port map( A1 => n1810, A2 => n6059, ZN => n1695);
   U2555 : NOR3_X1 port map( A1 => n6058, A2 => n1695, A3 => n1694, ZN => n6063
                           );
   U2556 : INV_X1 port map( A => n1723, ZN => n7044);
   U2557 : OR2_X1 port map( A1 => n7024, A2 => n7005, ZN => n1696);
   U2558 : NAND2_X1 port map( A1 => n1696, A2 => n1260, ZN => n7020);
   U2559 : NOR2_X1 port map( A1 => n2162, A2 => n1352, ZN => n1697);
   U2560 : OR2_X1 port map( A1 => n6288, A2 => n6292, ZN => n6275);
   U2561 : XNOR2_X1 port map( A => n6492, B => n618, ZN => n6493);
   U2562 : XNOR2_X1 port map( A => n947, B => n1698, ZN => n1752);
   U2563 : MUX2_X2 port map( A => n6463, B => n6462, S => n7973, Z => n6524);
   U2564 : XNOR2_X1 port map( A => n5631, B => n5634, ZN => n5635);
   U2565 : MUX2_X2 port map( A => n1700, B => n1701, S => n4436, Z => n1699);
   U2566 : XNOR2_X1 port map( A => n1307, B => n1491, ZN => n1700);
   U2567 : OR2_X1 port map( A1 => n5948, A2 => n5955, ZN => n5933);
   U2568 : MUX2_X2 port map( A => n5071, B => n5070, S => n2248, Z => n5499);
   U2569 : OR2_X1 port map( A1 => n5859, A2 => n5860, ZN => n1703);
   U2570 : OR2_X1 port map( A1 => n4777, A2 => n4668, ZN => n1704);
   U2571 : NAND2_X1 port map( A1 => n1706, A2 => n5930, ZN => n1707);
   U2572 : NAND2_X1 port map( A1 => n5931, A2 => n2168, ZN => n1708);
   U2573 : NAND2_X1 port map( A1 => n1708, A2 => n1707, ZN => n5998);
   U2574 : INV_X1 port map( A => n2168, ZN => n1706);
   U2575 : CLKBUF_X1 port map( A => n1827, Z => n1709);
   U2576 : CLKBUF_X1 port map( A => n17187, Z => n1710);
   U2577 : INV_X1 port map( A => n6654, ZN => n1712);
   U2578 : MUX2_X1 port map( A => n6453, B => n6454, S => n529, Z => n1713);
   U2579 : OR2_X1 port map( A1 => n5927, A2 => n5924, ZN => n1714);
   U2580 : INV_X1 port map( A => n6002, ZN => n1715);
   U2581 : XNOR2_X1 port map( A => n6810, B => n6812, ZN => n6591);
   U2582 : XNOR2_X1 port map( A => n5610, B => n1778, ZN => n5616);
   U2583 : XNOR2_X1 port map( A => n5883, B => n5889, ZN => n5890);
   U2584 : XNOR2_X1 port map( A => n1576, B => n7031, ZN => n1722);
   U2585 : XNOR2_X1 port map( A => n5324, B => n5328, ZN => n5325);
   U2586 : XNOR2_X1 port map( A => n1750, B => n6990, ZN => n6808);
   U2587 : MUX2_X2 port map( A => n4693, B => n4692, S => n2250, Z => n5235);
   U2588 : XNOR2_X1 port map( A => n5593, B => n5521, ZN => n5595);
   U2589 : XNOR2_X1 port map( A => n6199, B => n974, ZN => n6218);
   U2590 : XNOR2_X1 port map( A => n1693, B => n7474, ZN => n7048);
   U2591 : INV_X1 port map( A => n7477, ZN => n7476);
   U2592 : XNOR2_X1 port map( A => n6526, B => n6530, ZN => n6531);
   U2593 : INV_X1 port map( A => n565, ZN => n7418);
   U2594 : XNOR2_X1 port map( A => n5987, B => n5990, ZN => n5991);
   U2595 : XNOR2_X1 port map( A => n1400, B => n6802, ZN => n6467);
   U2596 : XNOR2_X1 port map( A => n1193, B => n7025, ZN => n7026);
   U2597 : XNOR2_X1 port map( A => n897, B => n6374, ZN => n6375);
   U2598 : NAND2_X1 port map( A1 => n6187, A2 => n6289, ZN => n1727);
   U2600 : XNOR2_X1 port map( A => n6548, B => n6534, ZN => n6549);
   U2601 : XNOR2_X1 port map( A => n6626, B => n6623, ZN => n6627);
   U2602 : XNOR2_X1 port map( A => n6680, B => n6681, ZN => n1728);
   U2603 : XNOR2_X1 port map( A => n5790, B => n5791, ZN => n5310);
   U2604 : XNOR2_X1 port map( A => n6970, B => n6969, ZN => n1729);
   U2605 : XNOR2_X1 port map( A => n1353, B => n4904, ZN => n4942);
   U2606 : MUX2_X2 port map( A => n5992, B => n5993, S => n1731, Z => n6023);
   U2607 : XNOR2_X1 port map( A => n6808, B => n6807, ZN => n1733);
   U2608 : XNOR2_X1 port map( A => n6813, B => n6814, ZN => n1734);
   U2609 : OR2_X2 port map( A1 => n4522, A2 => n4458, ZN => n4518);
   U2610 : XNOR2_X1 port map( A => n5046, B => n4969, ZN => n5049);
   U2611 : NAND2_X1 port map( A1 => n4903, A2 => n4908, ZN => n1735);
   U2612 : XNOR2_X1 port map( A => n5145, B => n1360, ZN => n5159);
   U2613 : XNOR2_X1 port map( A => n1773, B => n1295, ZN => n5454);
   U2614 : XNOR2_X1 port map( A => n5695, B => n1736, ZN => n5705);
   U2616 : OR2_X1 port map( A1 => n4783, A2 => n4663, ZN => n1737);
   U2617 : NAND2_X1 port map( A1 => n4786, A2 => n1737, ZN => n4664);
   U2618 : OR2_X1 port map( A1 => n4776, A2 => n4666, ZN => n1738);
   U2619 : OR2_X1 port map( A1 => n5528, A2 => n5549, ZN => n1739);
   U2620 : NAND2_X1 port map( A1 => n5610, A2 => n1739, ZN => n5520);
   U2621 : OR2_X1 port map( A1 => n868, A2 => n6215, ZN => n1740);
   U2622 : NAND2_X1 port map( A1 => n6214, A2 => n1740, ZN => n6265);
   U2623 : XNOR2_X1 port map( A => n1741, B => n5926, ZN => n5931);
   U2624 : XNOR2_X1 port map( A => n5925, B => n5924, ZN => n1741);
   U2625 : XNOR2_X1 port map( A => n6531, B => n6528, ZN => n6532);
   U2626 : INV_X1 port map( A => n4614, ZN => n1742);
   U2627 : NAND3_X1 port map( A1 => n4610, A2 => n4734, A3 => n320, ZN => n4611
                           );
   U2628 : OAI221_X1 port map( B1 => n8039, B2 => n8089, C1 => n8038, C2 => 
                           n8037, A => n8036, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n170);
   U2629 : OAI221_X1 port map( B1 => n7998, B2 => n8089, C1 => 
                           DataPath_ALUhw_SHIFTER_HW_n411, C2 => n7997, A => 
                           n7996, ZN => DataPath_ALUhw_SHIFTER_HW_n147);
   U2630 : XNOR2_X1 port map( A => n717, B => n6684, ZN => n6687);
   U2631 : INV_X1 port map( A => n5989, ZN => n1744);
   U2632 : XNOR2_X1 port map( A => n5708, B => n5713, ZN => n5714);
   U2633 : MUX2_X2 port map( A => n5715, B => n5714, S => n2243, Z => n8269);
   U2634 : MUX2_X2 port map( A => n6287, B => n6286, S => n8229, Z => n6410);
   U2635 : MUX2_X2 port map( A => n5051, B => n5050, S => n2248, Z => n5386);
   U2636 : INV_X1 port map( A => n1132, ZN => n6616);
   U2637 : INV_X1 port map( A => n1177, ZN => n6993);
   U2638 : XNOR2_X1 port map( A => n1012, B => n5625, ZN => n5626);
   U2639 : MUX2_X2 port map( A => n5557, B => n5556, S => n2243, Z => n6041);
   U2640 : XNOR2_X1 port map( A => n6803, B => n6833, ZN => n1751);
   U2641 : OAI21_X1 port map( B1 => n4582, B2 => n4581, A => n4854, ZN => n4883
                           );
   U2642 : XNOR2_X1 port map( A => n5667, B => n5668, ZN => n1754);
   U2643 : XNOR2_X1 port map( A => n6501, B => n643, ZN => n6502);
   U2644 : XNOR2_X1 port map( A => n6499, B => n6502, ZN => n6503);
   U2645 : XNOR2_X1 port map( A => n469, B => n6600, ZN => n6601);
   U2646 : XNOR2_X1 port map( A => n6097, B => n738, ZN => n6102);
   U2647 : XNOR2_X1 port map( A => n1003, B => n6267, ZN => n6268);
   U2648 : XNOR2_X1 port map( A => n6624, B => n6625, ZN => n6626);
   U2650 : XNOR2_X1 port map( A => n6981, B => n1759, ZN => n6987);
   U2651 : XNOR2_X1 port map( A => n1676, B => n7430, ZN => n1759);
   U2652 : XNOR2_X1 port map( A => n1037, B => n6246, ZN => n6247);
   U2653 : XNOR2_X1 port map( A => n5026, B => n5042, ZN => n5044);
   U2654 : XNOR2_X1 port map( A => n1400, B => n6806, ZN => n6492);
   U2655 : MUX2_X1 port map( A => DataPath_i_PIPLIN_B_2_port, B => 
                           DataPath_i_PIPLIN_IN2_2_port, S => i_S2, Z => n1760)
                           ;
   U2656 : XNOR2_X1 port map( A => n1761, B => n626, ZN => n6658);
   U2657 : XNOR2_X1 port map( A => n1762, B => n6985, ZN => n6986);
   U2658 : XNOR2_X1 port map( A => n7433, B => n1676, ZN => n1762);
   U2659 : XNOR2_X1 port map( A => n6997, B => n6996, ZN => n1764);
   U2660 : XNOR2_X1 port map( A => n6988, B => n6989, ZN => n1765);
   U2661 : XNOR2_X1 port map( A => n4528, B => n2262, ZN => n4581);
   U2662 : XNOR2_X1 port map( A => n5079, B => n5080, ZN => n5081);
   U2663 : XNOR2_X1 port map( A => n1766, B => n5589, ZN => n5590);
   U2664 : XNOR2_X1 port map( A => n7004, B => n1767, ZN => n7018);
   U2665 : XNOR2_X1 port map( A => n1419, B => n1726, ZN => n1767);
   U2666 : XOR2_X2 port map( A => n7865, B => n1702, Z => n7256);
   U2667 : NAND2_X2 port map( A1 => n6370, A2 => n7265, ZN => n7266);
   U2668 : XOR2_X2 port map( A => n7933, B => n7973, Z => n7265);
   U2669 : NAND2_X2 port map( A1 => n6232, A2 => n7272, ZN => n7274);
   U2670 : XOR2_X2 port map( A => n8215, B => n8229, Z => n7272);
   U2671 : BUF_X2 port map( A => n7296, Z => n2184);
   U2672 : INV_X2 port map( A => n2263, ZN => n2260);
   U2673 : MUX2_X2 port map( A => n5089, B => n5088, S => n2248, Z => n5422);
   U2674 : XNOR2_X1 port map( A => n1768, B => n5482, ZN => n5494);
   U2675 : XNOR2_X1 port map( A => n552, B => n5490, ZN => n1768);
   U2676 : INV_X2 port map( A => n1899, ZN => n2220);
   U2677 : INV_X2 port map( A => n1898, ZN => n2217);
   U2678 : INV_X2 port map( A => n1898, ZN => n2218);
   U2679 : CLKBUF_X3 port map( A => n8135, Z => n2243);
   U2680 : XOR2_X1 port map( A => n4570, B => n2155, Z => n4439);
   U2681 : CLKBUF_X3 port map( A => n7290, Z => n2185);
   U2682 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n600, B2 => 
                           n8019, C1 => n8018, C2 => n8037, A => n8017, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n156);
   U2683 : NAND3_X1 port map( A1 => n1907, A2 => n17175, A3 => n2260, ZN => 
                           n1769);
   U2684 : INV_X2 port map( A => n1935, ZN => n2213);
   U2685 : INV_X2 port map( A => n1934, ZN => n2215);
   U2687 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_14_port, A2 => n8325, ZN 
                           => n1770);
   U2688 : AND2_X1 port map( A1 => DataPath_i_ALU_OUT_13_port, A2 => n8325, ZN 
                           => n1771);
   U2689 : INV_X1 port map( A => n3707, ZN => n3638);
   U2690 : INV_X1 port map( A => n3706, ZN => n3633);
   U2691 : INV_X1 port map( A => n3706, ZN => n3634);
   U2692 : INV_X1 port map( A => n3707, ZN => n3637);
   U2693 : INV_X1 port map( A => n3707, ZN => n3636);
   U2694 : INV_X1 port map( A => n3704, ZN => n3631);
   U2695 : INV_X1 port map( A => n3708, ZN => n3639);
   U2696 : INV_X1 port map( A => n3708, ZN => n3640);
   U2697 : INV_X1 port map( A => n3708, ZN => n3641);
   U2698 : BUF_X1 port map( A => n3709, Z => n3706);
   U2699 : BUF_X1 port map( A => n3709, Z => n3708);
   U2700 : BUF_X1 port map( A => n3709, Z => n3707);
   U2701 : BUF_X1 port map( A => n3710, Z => n3704);
   U2702 : BUF_X1 port map( A => n3710, Z => n3705);
   U2703 : BUF_X1 port map( A => n3728, Z => n3651);
   U2704 : BUF_X1 port map( A => n3730, Z => n3644);
   U2705 : BUF_X1 port map( A => n3727, Z => n3653);
   U2706 : BUF_X1 port map( A => n3730, Z => n3645);
   U2707 : BUF_X1 port map( A => n3729, Z => n3648);
   U2708 : BUF_X1 port map( A => n3729, Z => n3646);
   U2709 : BUF_X1 port map( A => n3728, Z => n3649);
   U2710 : BUF_X1 port map( A => n3729, Z => n3647);
   U2711 : BUF_X1 port map( A => n3728, Z => n3650);
   U2712 : BUF_X1 port map( A => n3727, Z => n3652);
   U2713 : BUF_X1 port map( A => n3730, Z => n3643);
   U2714 : BUF_X1 port map( A => n3718, Z => n3680);
   U2715 : BUF_X1 port map( A => n3712, Z => n3699);
   U2716 : BUF_X1 port map( A => n3722, Z => n3668);
   U2717 : BUF_X1 port map( A => n3727, Z => n3654);
   U2718 : BUF_X1 port map( A => n3714, Z => n3693);
   U2719 : BUF_X1 port map( A => n3716, Z => n3687);
   U2720 : BUF_X1 port map( A => n3720, Z => n3675);
   U2721 : BUF_X1 port map( A => n3711, Z => n3700);
   U2722 : BUF_X1 port map( A => n3718, Z => n3681);
   U2723 : BUF_X1 port map( A => n3722, Z => n3669);
   U2724 : BUF_X1 port map( A => n3713, Z => n3694);
   U2725 : BUF_X1 port map( A => n3715, Z => n3689);
   U2726 : BUF_X1 port map( A => n3719, Z => n3677);
   U2727 : BUF_X1 port map( A => n3717, Z => n3683);
   U2728 : BUF_X1 port map( A => n3726, Z => n3656);
   U2729 : BUF_X1 port map( A => n3721, Z => n3671);
   U2730 : BUF_X1 port map( A => n3713, Z => n3696);
   U2731 : BUF_X1 port map( A => n3711, Z => n3702);
   U2732 : BUF_X1 port map( A => n3723, Z => n3665);
   U2733 : BUF_X1 port map( A => n3725, Z => n3660);
   U2734 : BUF_X1 port map( A => n3715, Z => n3690);
   U2735 : BUF_X1 port map( A => n3719, Z => n3678);
   U2736 : BUF_X1 port map( A => n3717, Z => n3684);
   U2737 : BUF_X1 port map( A => n3710, Z => n3703);
   U2738 : BUF_X1 port map( A => n3721, Z => n3672);
   U2739 : BUF_X1 port map( A => n3726, Z => n3657);
   U2740 : BUF_X1 port map( A => n3712, Z => n3697);
   U2741 : BUF_X1 port map( A => n3724, Z => n3663);
   U2742 : BUF_X1 port map( A => n3723, Z => n3666);
   U2743 : BUF_X1 port map( A => n3724, Z => n3661);
   U2744 : BUF_X1 port map( A => n3718, Z => n3679);
   U2745 : BUF_X1 port map( A => n3716, Z => n3686);
   U2746 : BUF_X1 port map( A => n3720, Z => n3674);
   U2747 : BUF_X1 port map( A => n3725, Z => n3659);
   U2748 : BUF_X1 port map( A => n3725, Z => n3658);
   U2749 : BUF_X1 port map( A => n3711, Z => n3701);
   U2750 : BUF_X1 port map( A => n3713, Z => n3695);
   U2751 : BUF_X1 port map( A => n3715, Z => n3688);
   U2752 : BUF_X1 port map( A => n3717, Z => n3682);
   U2753 : BUF_X1 port map( A => n3719, Z => n3676);
   U2754 : BUF_X1 port map( A => n3721, Z => n3670);
   U2755 : BUF_X1 port map( A => n3723, Z => n3664);
   U2756 : BUF_X1 port map( A => n3712, Z => n3698);
   U2757 : BUF_X1 port map( A => n3714, Z => n3691);
   U2758 : BUF_X1 port map( A => n3716, Z => n3685);
   U2759 : BUF_X1 port map( A => n3726, Z => n3655);
   U2760 : BUF_X1 port map( A => n3714, Z => n3692);
   U2761 : BUF_X1 port map( A => n3720, Z => n3673);
   U2762 : BUF_X1 port map( A => n3722, Z => n3667);
   U2763 : BUF_X1 port map( A => n3724, Z => n3662);
   U2764 : BUF_X1 port map( A => DataPath_WRF_CUhw_n113, Z => n3259);
   U2765 : BUF_X1 port map( A => DataPath_WRF_CUhw_n113, Z => n3260);
   U2766 : BUF_X1 port map( A => DataPath_WRF_CUhw_n113, Z => n3261);
   U2767 : INV_X1 port map( A => n5485, ZN => n5486);
   U2768 : AOI21_X1 port map( B1 => n5935, B2 => n5934, A => n1645, ZN => n5938
                           );
   U2769 : AND2_X1 port map( A1 => n5736, A2 => n5737, ZN => n5738);
   U2770 : AND2_X1 port map( A1 => n5450, A2 => n5449, ZN => n5451);
   U2771 : AND2_X1 port map( A1 => n5899, A2 => n5898, ZN => n5900);
   U2772 : AND2_X1 port map( A1 => n5441, A2 => n5442, ZN => n1773);
   U2773 : NAND2_X1 port map( A1 => n5653, A2 => n5654, ZN => n5655);
   U2774 : AND2_X1 port map( A1 => n4837, A2 => n4848, ZN => n1774);
   U2775 : AND2_X1 port map( A1 => n5903, A2 => n5904, ZN => n5905);
   U2776 : NAND2_X1 port map( A1 => n5939, A2 => n5953, ZN => n5942);
   U2777 : INV_X1 port map( A => n3371, ZN => n3301);
   U2778 : INV_X1 port map( A => n3370, ZN => n3297);
   U2779 : INV_X1 port map( A => n3370, ZN => n3298);
   U2780 : INV_X1 port map( A => n3371, ZN => n3300);
   U2781 : INV_X1 port map( A => n3371, ZN => n3302);
   U2782 : INV_X1 port map( A => n3370, ZN => n3296);
   U2783 : INV_X1 port map( A => n3483, ZN => n3414);
   U2784 : INV_X1 port map( A => n3482, ZN => n3410);
   U2785 : INV_X1 port map( A => n3483, ZN => n3413);
   U2786 : INV_X1 port map( A => n3483, ZN => n3412);
   U2787 : INV_X1 port map( A => n3595, ZN => n3526);
   U2788 : INV_X1 port map( A => n3594, ZN => n3522);
   U2789 : INV_X1 port map( A => n3595, ZN => n3525);
   U2790 : INV_X1 port map( A => n3595, ZN => n3524);
   U2791 : INV_X1 port map( A => n3819, ZN => n3749);
   U2792 : INV_X1 port map( A => n3818, ZN => n3744);
   U2793 : INV_X1 port map( A => n3818, ZN => n3745);
   U2794 : INV_X1 port map( A => n3819, ZN => n3750);
   U2795 : INV_X1 port map( A => n3818, ZN => n3743);
   U2796 : INV_X1 port map( A => n3819, ZN => n3748);
   U2797 : INV_X1 port map( A => n3819, ZN => n3747);
   U2798 : INV_X1 port map( A => n3480, ZN => n3407);
   U2799 : INV_X1 port map( A => n3481, ZN => n3408);
   U2800 : INV_X1 port map( A => n3592, ZN => n3519);
   U2801 : INV_X1 port map( A => n3593, ZN => n3520);
   U2802 : INV_X1 port map( A => n3484, ZN => n3415);
   U2803 : INV_X1 port map( A => n3596, ZN => n3527);
   U2804 : INV_X1 port map( A => n3820, ZN => n3751);
   U2805 : INV_X1 port map( A => n3372, ZN => n3303);
   U2806 : INV_X1 port map( A => n3372, ZN => n3304);
   U2807 : INV_X1 port map( A => n3372, ZN => n3305);
   U2808 : INV_X1 port map( A => n3484, ZN => n3416);
   U2809 : INV_X1 port map( A => n3484, ZN => n3417);
   U2810 : INV_X1 port map( A => n3596, ZN => n3528);
   U2811 : INV_X1 port map( A => n3596, ZN => n3529);
   U2812 : INV_X1 port map( A => n3820, ZN => n3752);
   U2813 : INV_X1 port map( A => n3820, ZN => n3753);
   U2814 : BUF_X1 port map( A => n3620, Z => n3710);
   U2815 : BUF_X1 port map( A => n3620, Z => n3709);
   U2816 : BUF_X1 port map( A => n14260, Z => n2486);
   U2817 : BUF_X1 port map( A => n14260, Z => n2487);
   U2818 : BUF_X1 port map( A => n14260, Z => n2488);
   U2819 : BUF_X1 port map( A => n3731, Z => n3642);
   U2820 : BUF_X1 port map( A => n3627, Z => n3731);
   U2821 : BUF_X1 port map( A => n3626, Z => n3729);
   U2822 : BUF_X1 port map( A => n3626, Z => n3728);
   U2823 : BUF_X1 port map( A => n3626, Z => n3727);
   U2824 : BUF_X1 port map( A => n3623, Z => n3718);
   U2825 : BUF_X1 port map( A => n3625, Z => n3725);
   U2826 : BUF_X1 port map( A => n3620, Z => n3711);
   U2827 : BUF_X1 port map( A => n3621, Z => n3713);
   U2828 : BUF_X1 port map( A => n3622, Z => n3715);
   U2829 : BUF_X1 port map( A => n3622, Z => n3717);
   U2830 : BUF_X1 port map( A => n3623, Z => n3719);
   U2831 : BUF_X1 port map( A => n3624, Z => n3721);
   U2832 : BUF_X1 port map( A => n3624, Z => n3723);
   U2833 : BUF_X1 port map( A => n3621, Z => n3712);
   U2834 : BUF_X1 port map( A => n3622, Z => n3716);
   U2835 : BUF_X1 port map( A => n3625, Z => n3726);
   U2836 : BUF_X1 port map( A => n3621, Z => n3714);
   U2837 : BUF_X1 port map( A => n3623, Z => n3720);
   U2838 : BUF_X1 port map( A => n3624, Z => n3722);
   U2839 : BUF_X1 port map( A => n3625, Z => n3724);
   U2840 : BUF_X1 port map( A => n3627, Z => n3730);
   U2841 : NAND2_X1 port map( A1 => n3258, A2 => n4264, ZN => 
                           DataPath_WRF_CUhw_n113);
   U2842 : XNOR2_X1 port map( A => n6435, B => n6436, ZN => n6437);
   U2843 : XNOR2_X1 port map( A => n1077, B => n6625, ZN => n6622);
   U2844 : XNOR2_X1 port map( A => n620, B => n5909, ZN => n5910);
   U2845 : XNOR2_X1 port map( A => n1043, B => n1801, ZN => n4945);
   U2846 : BUF_X2 port map( A => n7312, Z => n2221);
   U2847 : CLKBUF_X1 port map( A => n7312, Z => n2222);
   U2848 : AND2_X1 port map( A1 => n5665, A2 => n5666, ZN => n5667);
   U2849 : BUF_X2 port map( A => n7303, Z => n2180);
   U2850 : NAND2_X1 port map( A1 => n5271, A2 => n5490, ZN => n5278);
   U2851 : INV_X1 port map( A => n5476, ZN => n5271);
   U2852 : AND2_X1 port map( A1 => n5406, A2 => n5407, ZN => n5410);
   U2853 : XNOR2_X1 port map( A => n4829, B => n4828, ZN => n1777);
   U2854 : BUF_X2 port map( A => n7303, Z => n2181);
   U2855 : CLKBUF_X3 port map( A => n7296, Z => n2183);
   U2856 : INV_X1 port map( A => n5955, ZN => n2162);
   U2857 : XNOR2_X1 port map( A => n975, B => n5608, ZN => n1778);
   U2858 : NAND2_X1 port map( A1 => n6118, A2 => n6016, ZN => n6015);
   U2859 : INV_X1 port map( A => n6023, ZN => n6198);
   U2861 : AND2_X1 port map( A1 => n7803, A2 => n6648, ZN => n1782);
   U2862 : INV_X1 port map( A => n6136, ZN => n2156);
   U2863 : AOI21_X1 port map( B1 => n5942, B2 => n5941, A => n1697, ZN => n5945
                           );
   U2864 : AND2_X1 port map( A1 => n1177, A2 => n6990, ZN => n1786);
   U2865 : AND2_X1 port map( A1 => n5592, A2 => n1647, ZN => n1787);
   U2866 : AND2_X1 port map( A1 => n6177, A2 => n6157, ZN => n1788);
   U2867 : AND2_X1 port map( A1 => n6841, A2 => n6840, ZN => n1792);
   U2868 : AND2_X1 port map( A1 => n825, A2 => n7460, ZN => n7015);
   U2869 : AND2_X1 port map( A1 => n6141, A2 => n1134, ZN => n1793);
   U2870 : AND2_X1 port map( A1 => n5821, A2 => n5920, ZN => n1794);
   U2871 : OR2_X1 port map( A1 => n6152, A2 => n6164, ZN => n6153);
   U2872 : XNOR2_X1 port map( A => n742, B => n1856, ZN => n7972);
   U2873 : NOR2_X2 port map( A1 => n8583, A2 => n8584, ZN => 
                           DataPath_RF_internal_inloc_data_0_0_port);
   U2874 : INV_X1 port map( A => n13107, ZN => n11611);
   U2875 : NOR2_X2 port map( A1 => n8581, A2 => n8582, ZN => 
                           DataPath_RF_internal_inloc_data_1_31_port);
   U2876 : INV_X1 port map( A => n13339, ZN => n12579);
   U2877 : NOR2_X2 port map( A1 => n8579, A2 => n8580, ZN => 
                           DataPath_RF_internal_inloc_data_1_30_port);
   U2878 : INV_X1 port map( A => n13340, ZN => n12539);
   U2879 : NOR2_X2 port map( A1 => n8577, A2 => n8578, ZN => 
                           DataPath_RF_internal_inloc_data_1_29_port);
   U2880 : INV_X1 port map( A => n13342, ZN => n12459);
   U2881 : NOR2_X2 port map( A1 => n8575, A2 => n8576, ZN => 
                           DataPath_RF_internal_inloc_data_1_28_port);
   U2882 : INV_X1 port map( A => n13247, ZN => n12416);
   U2883 : NOR2_X2 port map( A1 => n8573, A2 => n8574, ZN => 
                           DataPath_RF_internal_inloc_data_1_27_port);
   U2884 : INV_X1 port map( A => n13344, ZN => n12379);
   U2885 : NOR2_X2 port map( A1 => n8571, A2 => n8572, ZN => 
                           DataPath_RF_internal_inloc_data_1_26_port);
   U2886 : INV_X1 port map( A => n13345, ZN => n12339);
   U2887 : NOR2_X2 port map( A1 => n8523, A2 => n8524, ZN => 
                           DataPath_RF_internal_inloc_data_1_2_port);
   U2888 : INV_X1 port map( A => n13341, ZN => n12499);
   U2889 : NOR2_X2 port map( A1 => n8517, A2 => n8518, ZN => 
                           DataPath_RF_internal_inloc_data_2_31_port);
   U2890 : INV_X1 port map( A => n13595, ZN => n12587);
   U2891 : NOR2_X2 port map( A1 => n8515, A2 => n8516, ZN => 
                           DataPath_RF_internal_inloc_data_2_30_port);
   U2892 : INV_X1 port map( A => n13596, ZN => n12547);
   U2893 : NOR2_X2 port map( A1 => n8513, A2 => n8514, ZN => 
                           DataPath_RF_internal_inloc_data_2_29_port);
   U2894 : INV_X1 port map( A => n13598, ZN => n12467);
   U2895 : NOR2_X2 port map( A1 => n8511, A2 => n8512, ZN => 
                           DataPath_RF_internal_inloc_data_2_28_port);
   U2896 : INV_X1 port map( A => n13503, ZN => n12424);
   U2897 : NOR2_X2 port map( A1 => n8509, A2 => n8510, ZN => 
                           DataPath_RF_internal_inloc_data_2_27_port);
   U2898 : INV_X1 port map( A => n13600, ZN => n12387);
   U2899 : NOR2_X2 port map( A1 => n8507, A2 => n8508, ZN => 
                           DataPath_RF_internal_inloc_data_2_26_port);
   U2900 : INV_X1 port map( A => n13601, ZN => n12347);
   U2901 : NOR2_X2 port map( A1 => n8459, A2 => n8460, ZN => 
                           DataPath_RF_internal_inloc_data_2_2_port);
   U2902 : INV_X1 port map( A => n13597, ZN => n12507);
   U2903 : NOR2_X2 port map( A1 => n8447, A2 => n8448, ZN => 
                           DataPath_RF_internal_inloc_data_3_28_port);
   U2904 : INV_X1 port map( A => n13759, ZN => n12432);
   U2905 : NOR2_X2 port map( A1 => n8419, A2 => n8420, ZN => 
                           DataPath_RF_internal_inloc_data_3_14_port);
   U2906 : INV_X1 port map( A => n13870, ZN => n11835);
   U2907 : NOR2_X2 port map( A1 => n8417, A2 => n8418, ZN => 
                           DataPath_RF_internal_inloc_data_3_13_port);
   U2908 : INV_X1 port map( A => n13871, ZN => n11795);
   U2909 : NOR2_X2 port map( A1 => n8415, A2 => n8416, ZN => 
                           DataPath_RF_internal_inloc_data_3_12_port);
   U2910 : INV_X1 port map( A => n13872, ZN => n11755);
   U2911 : NOR2_X2 port map( A1 => n8413, A2 => n8414, ZN => 
                           DataPath_RF_internal_inloc_data_3_11_port);
   U2912 : INV_X1 port map( A => n13873, ZN => n11715);
   U2913 : NOR2_X2 port map( A1 => n8411, A2 => n8412, ZN => 
                           DataPath_RF_internal_inloc_data_3_10_port);
   U2914 : INV_X1 port map( A => n13874, ZN => n11675);
   U2915 : NOR2_X2 port map( A1 => n8409, A2 => n8410, ZN => 
                           DataPath_RF_internal_inloc_data_3_9_port);
   U2916 : INV_X1 port map( A => n13844, ZN => n12875);
   U2917 : NOR2_X2 port map( A1 => n8407, A2 => n8408, ZN => 
                           DataPath_RF_internal_inloc_data_3_8_port);
   U2918 : INV_X1 port map( A => n13845, ZN => n12835);
   U2919 : NOR2_X2 port map( A1 => n8405, A2 => n8406, ZN => 
                           DataPath_RF_internal_inloc_data_3_7_port);
   U2920 : INV_X1 port map( A => n13846, ZN => n12795);
   U2921 : NOR2_X2 port map( A1 => n8403, A2 => n8404, ZN => 
                           DataPath_RF_internal_inloc_data_3_6_port);
   U2922 : INV_X1 port map( A => n13847, ZN => n12755);
   U2923 : NOR2_X2 port map( A1 => n8401, A2 => n8402, ZN => 
                           DataPath_RF_internal_inloc_data_3_5_port);
   U2924 : INV_X1 port map( A => n13848, ZN => n12715);
   U2925 : NOR2_X2 port map( A1 => n8399, A2 => n8400, ZN => 
                           DataPath_RF_internal_inloc_data_3_4_port);
   U2926 : INV_X1 port map( A => n13849, ZN => n12675);
   U2927 : NOR2_X2 port map( A1 => n8397, A2 => n8398, ZN => 
                           DataPath_RF_internal_inloc_data_3_3_port);
   U2928 : INV_X1 port map( A => n13850, ZN => n12635);
   U2929 : NOR2_X2 port map( A1 => n8391, A2 => n8392, ZN => 
                           DataPath_RF_internal_inloc_data_3_0_port);
   U2930 : INV_X1 port map( A => n13875, ZN => n11635);
   U2931 : NOR2_X2 port map( A1 => n8383, A2 => n8384, ZN => 
                           DataPath_RF_internal_inloc_data_4_28_port);
   U2932 : INV_X1 port map( A => n14015, ZN => n12440);
   U2933 : NOR2_X2 port map( A1 => n8355, A2 => n8356, ZN => 
                           DataPath_RF_internal_inloc_data_4_14_port);
   U2934 : INV_X1 port map( A => n14126, ZN => n11843);
   U2935 : NOR2_X2 port map( A1 => n8353, A2 => n8354, ZN => 
                           DataPath_RF_internal_inloc_data_4_13_port);
   U2936 : INV_X1 port map( A => n14127, ZN => n11803);
   U2937 : NOR2_X2 port map( A1 => n8351, A2 => n8352, ZN => 
                           DataPath_RF_internal_inloc_data_4_12_port);
   U2938 : INV_X1 port map( A => n14128, ZN => n11763);
   U2939 : NOR2_X2 port map( A1 => n8349, A2 => n8350, ZN => 
                           DataPath_RF_internal_inloc_data_4_11_port);
   U2940 : INV_X1 port map( A => n14129, ZN => n11723);
   U2941 : NOR2_X2 port map( A1 => n8347, A2 => n8348, ZN => 
                           DataPath_RF_internal_inloc_data_4_10_port);
   U2942 : INV_X1 port map( A => n14130, ZN => n11683);
   U2943 : NOR2_X2 port map( A1 => n8345, A2 => n8346, ZN => 
                           DataPath_RF_internal_inloc_data_4_9_port);
   U2944 : INV_X1 port map( A => n14100, ZN => n12883);
   U2945 : NOR2_X2 port map( A1 => n8343, A2 => n8344, ZN => 
                           DataPath_RF_internal_inloc_data_4_8_port);
   U2946 : INV_X1 port map( A => n14101, ZN => n12843);
   U2947 : NOR2_X2 port map( A1 => n8341, A2 => n8342, ZN => 
                           DataPath_RF_internal_inloc_data_4_7_port);
   U2948 : INV_X1 port map( A => n14102, ZN => n12803);
   U2949 : NOR2_X2 port map( A1 => n8339, A2 => n8340, ZN => 
                           DataPath_RF_internal_inloc_data_4_6_port);
   U2950 : INV_X1 port map( A => n14103, ZN => n12763);
   U2951 : NOR2_X2 port map( A1 => n8337, A2 => n8338, ZN => 
                           DataPath_RF_internal_inloc_data_4_5_port);
   U2952 : INV_X1 port map( A => n14104, ZN => n12723);
   U2953 : NOR2_X2 port map( A1 => n8335, A2 => n8336, ZN => 
                           DataPath_RF_internal_inloc_data_4_4_port);
   U2954 : INV_X1 port map( A => n14105, ZN => n12683);
   U2955 : NOR2_X2 port map( A1 => n8333, A2 => n8334, ZN => 
                           DataPath_RF_internal_inloc_data_4_3_port);
   U2956 : INV_X1 port map( A => n14106, ZN => n12643);
   U2957 : NOR2_X2 port map( A1 => n8327, A2 => n8328, ZN => 
                           DataPath_RF_internal_inloc_data_4_0_port);
   U2958 : INV_X1 port map( A => n14131, ZN => n11643);
   U2959 : INV_X1 port map( A => n8025, ZN => n8305);
   U2960 : INV_X1 port map( A => n8030, ZN => n8306);
   U2961 : OAI22_X1 port map( A1 => n8289, A2 => n1769, B1 => n8286, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n533);
   U2962 : OAI22_X1 port map( A1 => n8292, A2 => n2984, B1 => n8291, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n148);
   U2963 : OAI22_X1 port map( A1 => n8286, A2 => n2984, B1 => n8289, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n500);
   U2964 : OAI22_X1 port map( A1 => n8290, A2 => n1769, B1 => n8289, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n520);
   U2965 : OAI22_X1 port map( A1 => n8290, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8289, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n180);
   U2966 : NOR2_X2 port map( A1 => n8645, A2 => n8646, ZN => 
                           DataPath_RF_internal_inloc_data_0_31_port);
   U2967 : INV_X1 port map( A => n13115, ZN => n12572);
   U2968 : NOR2_X2 port map( A1 => n8643, A2 => n8644, ZN => 
                           DataPath_RF_internal_inloc_data_0_30_port);
   U2969 : INV_X1 port map( A => n13116, ZN => n12532);
   U2970 : NOR2_X2 port map( A1 => n8641, A2 => n8642, ZN => 
                           DataPath_RF_internal_inloc_data_0_29_port);
   U2971 : INV_X1 port map( A => n13118, ZN => n12452);
   U2972 : NOR2_X2 port map( A1 => n8639, A2 => n8640, ZN => 
                           DataPath_RF_internal_inloc_data_0_28_port);
   U2973 : INV_X1 port map( A => n13119, ZN => n12412);
   U2974 : NOR2_X2 port map( A1 => n8637, A2 => n8638, ZN => 
                           DataPath_RF_internal_inloc_data_0_27_port);
   U2975 : INV_X1 port map( A => n13120, ZN => n12372);
   U2976 : NOR2_X2 port map( A1 => n8635, A2 => n8636, ZN => 
                           DataPath_RF_internal_inloc_data_0_26_port);
   U2977 : INV_X1 port map( A => n13121, ZN => n12332);
   U2978 : NOR2_X2 port map( A1 => n8633, A2 => n8634, ZN => 
                           DataPath_RF_internal_inloc_data_0_25_port);
   U2979 : INV_X1 port map( A => n13122, ZN => n12292);
   U2980 : NOR2_X2 port map( A1 => n8631, A2 => n8632, ZN => 
                           DataPath_RF_internal_inloc_data_0_24_port);
   U2981 : INV_X1 port map( A => n13123, ZN => n12252);
   U2982 : NOR2_X2 port map( A1 => n8629, A2 => n8630, ZN => 
                           DataPath_RF_internal_inloc_data_0_23_port);
   U2983 : INV_X1 port map( A => n13124, ZN => n12212);
   U2984 : NOR2_X2 port map( A1 => n8627, A2 => n8628, ZN => 
                           DataPath_RF_internal_inloc_data_0_22_port);
   U2985 : INV_X1 port map( A => n13125, ZN => n12172);
   U2986 : NOR2_X2 port map( A1 => n8625, A2 => n8626, ZN => 
                           DataPath_RF_internal_inloc_data_0_21_port);
   U2987 : INV_X1 port map( A => n13126, ZN => n12132);
   U2988 : NOR2_X2 port map( A1 => n8623, A2 => n8624, ZN => 
                           DataPath_RF_internal_inloc_data_0_20_port);
   U2989 : INV_X1 port map( A => n13127, ZN => n12092);
   U2990 : NOR2_X2 port map( A1 => n8621, A2 => n8622, ZN => 
                           DataPath_RF_internal_inloc_data_0_19_port);
   U2991 : INV_X1 port map( A => n13129, ZN => n12012);
   U2992 : NOR2_X2 port map( A1 => n8619, A2 => n8620, ZN => 
                           DataPath_RF_internal_inloc_data_0_18_port);
   U2993 : INV_X1 port map( A => n13130, ZN => n11972);
   U2994 : NOR2_X2 port map( A1 => n8617, A2 => n8618, ZN => 
                           DataPath_RF_internal_inloc_data_0_17_port);
   U2995 : INV_X1 port map( A => n13131, ZN => n11932);
   U2996 : NOR2_X2 port map( A1 => n8615, A2 => n8616, ZN => 
                           DataPath_RF_internal_inloc_data_0_16_port);
   U2997 : INV_X1 port map( A => n13132, ZN => n11892);
   U2998 : NOR2_X2 port map( A1 => n8613, A2 => n8614, ZN => 
                           DataPath_RF_internal_inloc_data_0_15_port);
   U2999 : INV_X1 port map( A => n13133, ZN => n11852);
   U3000 : NOR2_X2 port map( A1 => n8611, A2 => n8612, ZN => 
                           DataPath_RF_internal_inloc_data_0_14_port);
   U3001 : INV_X1 port map( A => n13134, ZN => n11812);
   U3002 : NOR2_X2 port map( A1 => n8609, A2 => n8610, ZN => 
                           DataPath_RF_internal_inloc_data_0_13_port);
   U3003 : INV_X1 port map( A => n13135, ZN => n11772);
   U3004 : NOR2_X2 port map( A1 => n8607, A2 => n8608, ZN => 
                           DataPath_RF_internal_inloc_data_0_12_port);
   U3005 : INV_X1 port map( A => n13136, ZN => n11732);
   U3006 : NOR2_X2 port map( A1 => n8605, A2 => n8606, ZN => 
                           DataPath_RF_internal_inloc_data_0_11_port);
   U3007 : INV_X1 port map( A => n13137, ZN => n11692);
   U3008 : NOR2_X2 port map( A1 => n8603, A2 => n8604, ZN => 
                           DataPath_RF_internal_inloc_data_0_10_port);
   U3009 : INV_X1 port map( A => n13138, ZN => n11652);
   U3010 : NOR2_X2 port map( A1 => n8601, A2 => n8602, ZN => 
                           DataPath_RF_internal_inloc_data_0_9_port);
   U3011 : INV_X1 port map( A => n13108, ZN => n12852);
   U3012 : NOR2_X2 port map( A1 => n8599, A2 => n8600, ZN => 
                           DataPath_RF_internal_inloc_data_0_8_port);
   U3013 : INV_X1 port map( A => n13109, ZN => n12812);
   U3014 : NOR2_X2 port map( A1 => n8597, A2 => n8598, ZN => 
                           DataPath_RF_internal_inloc_data_0_7_port);
   U3015 : INV_X1 port map( A => n13110, ZN => n12772);
   U3016 : NOR2_X2 port map( A1 => n8595, A2 => n8596, ZN => 
                           DataPath_RF_internal_inloc_data_0_6_port);
   U3017 : INV_X1 port map( A => n13111, ZN => n12732);
   U3018 : NOR2_X2 port map( A1 => n8593, A2 => n8594, ZN => 
                           DataPath_RF_internal_inloc_data_0_5_port);
   U3019 : INV_X1 port map( A => n13112, ZN => n12692);
   U3020 : NOR2_X2 port map( A1 => n8591, A2 => n8592, ZN => 
                           DataPath_RF_internal_inloc_data_0_4_port);
   U3021 : INV_X1 port map( A => n13113, ZN => n12652);
   U3022 : NOR2_X2 port map( A1 => n8589, A2 => n8590, ZN => 
                           DataPath_RF_internal_inloc_data_0_3_port);
   U3023 : INV_X1 port map( A => n13114, ZN => n12612);
   U3024 : NOR2_X2 port map( A1 => n8587, A2 => n8588, ZN => 
                           DataPath_RF_internal_inloc_data_0_2_port);
   U3025 : INV_X1 port map( A => n13117, ZN => n12492);
   U3026 : NOR2_X2 port map( A1 => n8585, A2 => n8586, ZN => 
                           DataPath_RF_internal_inloc_data_0_1_port);
   U3027 : INV_X1 port map( A => n13128, ZN => n12052);
   U3028 : NOR2_X2 port map( A1 => n8569, A2 => n8570, ZN => 
                           DataPath_RF_internal_inloc_data_1_25_port);
   U3029 : INV_X1 port map( A => n13346, ZN => n12299);
   U3030 : NOR2_X2 port map( A1 => n8567, A2 => n8568, ZN => 
                           DataPath_RF_internal_inloc_data_1_24_port);
   U3031 : INV_X1 port map( A => n13347, ZN => n12259);
   U3032 : NOR2_X2 port map( A1 => n8565, A2 => n8566, ZN => 
                           DataPath_RF_internal_inloc_data_1_23_port);
   U3033 : INV_X1 port map( A => n13348, ZN => n12219);
   U3034 : NOR2_X2 port map( A1 => n8563, A2 => n8564, ZN => 
                           DataPath_RF_internal_inloc_data_1_22_port);
   U3035 : INV_X1 port map( A => n13349, ZN => n12179);
   U3036 : NOR2_X2 port map( A1 => n8561, A2 => n8562, ZN => 
                           DataPath_RF_internal_inloc_data_1_21_port);
   U3037 : INV_X1 port map( A => n13350, ZN => n12139);
   U3038 : NOR2_X2 port map( A1 => n8559, A2 => n8560, ZN => 
                           DataPath_RF_internal_inloc_data_1_20_port);
   U3039 : INV_X1 port map( A => n13351, ZN => n12099);
   U3040 : NOR2_X2 port map( A1 => n8557, A2 => n8558, ZN => 
                           DataPath_RF_internal_inloc_data_1_19_port);
   U3041 : INV_X1 port map( A => n13353, ZN => n12019);
   U3042 : NOR2_X2 port map( A1 => n8555, A2 => n8556, ZN => 
                           DataPath_RF_internal_inloc_data_1_18_port);
   U3043 : INV_X1 port map( A => n13354, ZN => n11979);
   U3044 : NOR2_X2 port map( A1 => n8553, A2 => n8554, ZN => 
                           DataPath_RF_internal_inloc_data_1_17_port);
   U3045 : INV_X1 port map( A => n13355, ZN => n11939);
   U3046 : NOR2_X2 port map( A1 => n8551, A2 => n8552, ZN => 
                           DataPath_RF_internal_inloc_data_1_16_port);
   U3047 : INV_X1 port map( A => n13356, ZN => n11899);
   U3048 : NOR2_X2 port map( A1 => n8549, A2 => n8550, ZN => 
                           DataPath_RF_internal_inloc_data_1_15_port);
   U3049 : INV_X1 port map( A => n13389, ZN => n11860);
   U3050 : NOR2_X2 port map( A1 => n8547, A2 => n8548, ZN => 
                           DataPath_RF_internal_inloc_data_1_14_port);
   U3051 : INV_X1 port map( A => n13358, ZN => n11819);
   U3052 : NOR2_X2 port map( A1 => n8545, A2 => n8546, ZN => 
                           DataPath_RF_internal_inloc_data_1_13_port);
   U3053 : INV_X1 port map( A => n13359, ZN => n11779);
   U3054 : NOR2_X2 port map( A1 => n8543, A2 => n8544, ZN => 
                           DataPath_RF_internal_inloc_data_1_12_port);
   U3055 : INV_X1 port map( A => n13360, ZN => n11739);
   U3056 : NOR2_X2 port map( A1 => n8541, A2 => n8542, ZN => 
                           DataPath_RF_internal_inloc_data_1_11_port);
   U3057 : INV_X1 port map( A => n13361, ZN => n11699);
   U3058 : NOR2_X2 port map( A1 => n8539, A2 => n8540, ZN => 
                           DataPath_RF_internal_inloc_data_1_10_port);
   U3059 : INV_X1 port map( A => n13362, ZN => n11659);
   U3060 : NOR2_X2 port map( A1 => n8537, A2 => n8538, ZN => 
                           DataPath_RF_internal_inloc_data_1_9_port);
   U3061 : INV_X1 port map( A => n13332, ZN => n12859);
   U3062 : NOR2_X2 port map( A1 => n8535, A2 => n8536, ZN => 
                           DataPath_RF_internal_inloc_data_1_8_port);
   U3063 : INV_X1 port map( A => n13333, ZN => n12819);
   U3064 : NOR2_X2 port map( A1 => n8533, A2 => n8534, ZN => 
                           DataPath_RF_internal_inloc_data_1_7_port);
   U3065 : INV_X1 port map( A => n13334, ZN => n12779);
   U3066 : NOR2_X2 port map( A1 => n8531, A2 => n8532, ZN => 
                           DataPath_RF_internal_inloc_data_1_6_port);
   U3067 : INV_X1 port map( A => n13335, ZN => n12739);
   U3068 : NOR2_X2 port map( A1 => n8529, A2 => n8530, ZN => 
                           DataPath_RF_internal_inloc_data_1_5_port);
   U3069 : INV_X1 port map( A => n13336, ZN => n12699);
   U3070 : NOR2_X2 port map( A1 => n8527, A2 => n8528, ZN => 
                           DataPath_RF_internal_inloc_data_1_4_port);
   U3071 : INV_X1 port map( A => n13337, ZN => n12659);
   U3072 : NOR2_X2 port map( A1 => n8525, A2 => n8526, ZN => 
                           DataPath_RF_internal_inloc_data_1_3_port);
   U3073 : INV_X1 port map( A => n13338, ZN => n12619);
   U3074 : NOR2_X2 port map( A1 => n8521, A2 => n8522, ZN => 
                           DataPath_RF_internal_inloc_data_1_1_port);
   U3075 : INV_X1 port map( A => n13352, ZN => n12059);
   U3076 : NOR2_X2 port map( A1 => n8519, A2 => n8520, ZN => 
                           DataPath_RF_internal_inloc_data_1_0_port);
   U3077 : INV_X1 port map( A => n13363, ZN => n11619);
   U3078 : NOR2_X2 port map( A1 => n8505, A2 => n8506, ZN => 
                           DataPath_RF_internal_inloc_data_2_25_port);
   U3079 : INV_X1 port map( A => n13602, ZN => n12307);
   U3080 : NOR2_X2 port map( A1 => n8503, A2 => n8504, ZN => 
                           DataPath_RF_internal_inloc_data_2_24_port);
   U3081 : INV_X1 port map( A => n13603, ZN => n12267);
   U3082 : NOR2_X2 port map( A1 => n8501, A2 => n8502, ZN => 
                           DataPath_RF_internal_inloc_data_2_23_port);
   U3083 : INV_X1 port map( A => n13604, ZN => n12227);
   U3084 : NOR2_X2 port map( A1 => n8499, A2 => n8500, ZN => 
                           DataPath_RF_internal_inloc_data_2_22_port);
   U3085 : INV_X1 port map( A => n13605, ZN => n12187);
   U3086 : NOR2_X2 port map( A1 => n8497, A2 => n8498, ZN => 
                           DataPath_RF_internal_inloc_data_2_21_port);
   U3087 : INV_X1 port map( A => n13606, ZN => n12147);
   U3088 : NOR2_X2 port map( A1 => n8495, A2 => n8496, ZN => 
                           DataPath_RF_internal_inloc_data_2_20_port);
   U3089 : INV_X1 port map( A => n13607, ZN => n12107);
   U3090 : NOR2_X2 port map( A1 => n8493, A2 => n8494, ZN => 
                           DataPath_RF_internal_inloc_data_2_19_port);
   U3091 : INV_X1 port map( A => n13609, ZN => n12027);
   U3092 : NOR2_X2 port map( A1 => n8491, A2 => n8492, ZN => 
                           DataPath_RF_internal_inloc_data_2_18_port);
   U3093 : INV_X1 port map( A => n13610, ZN => n11987);
   U3094 : NOR2_X2 port map( A1 => n8489, A2 => n8490, ZN => 
                           DataPath_RF_internal_inloc_data_2_17_port);
   U3095 : INV_X1 port map( A => n13611, ZN => n11947);
   U3096 : NOR2_X2 port map( A1 => n8487, A2 => n8488, ZN => 
                           DataPath_RF_internal_inloc_data_2_16_port);
   U3097 : INV_X1 port map( A => n13612, ZN => n11907);
   U3098 : NOR2_X2 port map( A1 => n8485, A2 => n8486, ZN => 
                           DataPath_RF_internal_inloc_data_2_15_port);
   U3099 : INV_X1 port map( A => n13645, ZN => n11868);
   U3100 : NOR2_X2 port map( A1 => n8483, A2 => n8484, ZN => 
                           DataPath_RF_internal_inloc_data_2_14_port);
   U3101 : INV_X1 port map( A => n13614, ZN => n11827);
   U3102 : NOR2_X2 port map( A1 => n8481, A2 => n8482, ZN => 
                           DataPath_RF_internal_inloc_data_2_13_port);
   U3103 : INV_X1 port map( A => n13615, ZN => n11787);
   U3104 : NOR2_X2 port map( A1 => n8479, A2 => n8480, ZN => 
                           DataPath_RF_internal_inloc_data_2_12_port);
   U3105 : INV_X1 port map( A => n13616, ZN => n11747);
   U3106 : NOR2_X2 port map( A1 => n8477, A2 => n8478, ZN => 
                           DataPath_RF_internal_inloc_data_2_11_port);
   U3107 : INV_X1 port map( A => n13617, ZN => n11707);
   U3108 : NOR2_X2 port map( A1 => n8475, A2 => n8476, ZN => 
                           DataPath_RF_internal_inloc_data_2_10_port);
   U3109 : INV_X1 port map( A => n13618, ZN => n11667);
   U3110 : NOR2_X2 port map( A1 => n8473, A2 => n8474, ZN => 
                           DataPath_RF_internal_inloc_data_2_9_port);
   U3111 : INV_X1 port map( A => n13588, ZN => n12867);
   U3112 : NOR2_X2 port map( A1 => n8471, A2 => n8472, ZN => 
                           DataPath_RF_internal_inloc_data_2_8_port);
   U3113 : INV_X1 port map( A => n13589, ZN => n12827);
   U3114 : NOR2_X2 port map( A1 => n8469, A2 => n8470, ZN => 
                           DataPath_RF_internal_inloc_data_2_7_port);
   U3115 : INV_X1 port map( A => n13590, ZN => n12787);
   U3116 : NOR2_X2 port map( A1 => n8467, A2 => n8468, ZN => 
                           DataPath_RF_internal_inloc_data_2_6_port);
   U3117 : INV_X1 port map( A => n13591, ZN => n12747);
   U3118 : NOR2_X2 port map( A1 => n8465, A2 => n8466, ZN => 
                           DataPath_RF_internal_inloc_data_2_5_port);
   U3119 : INV_X1 port map( A => n13592, ZN => n12707);
   U3120 : NOR2_X2 port map( A1 => n8463, A2 => n8464, ZN => 
                           DataPath_RF_internal_inloc_data_2_4_port);
   U3121 : INV_X1 port map( A => n13593, ZN => n12667);
   U3122 : NOR2_X2 port map( A1 => n8461, A2 => n8462, ZN => 
                           DataPath_RF_internal_inloc_data_2_3_port);
   U3123 : INV_X1 port map( A => n13594, ZN => n12627);
   U3124 : NOR2_X2 port map( A1 => n8457, A2 => n8458, ZN => 
                           DataPath_RF_internal_inloc_data_2_1_port);
   U3125 : INV_X1 port map( A => n13608, ZN => n12067);
   U3126 : NOR2_X2 port map( A1 => n8455, A2 => n8456, ZN => 
                           DataPath_RF_internal_inloc_data_2_0_port);
   U3127 : INV_X1 port map( A => n13619, ZN => n11627);
   U3128 : NOR2_X2 port map( A1 => n8453, A2 => n8454, ZN => 
                           DataPath_RF_internal_inloc_data_3_31_port);
   U3129 : INV_X1 port map( A => n13851, ZN => n12595);
   U3130 : NOR2_X2 port map( A1 => n8451, A2 => n8452, ZN => 
                           DataPath_RF_internal_inloc_data_3_30_port);
   U3131 : INV_X1 port map( A => n13852, ZN => n12555);
   U3132 : NOR2_X2 port map( A1 => n8449, A2 => n8450, ZN => 
                           DataPath_RF_internal_inloc_data_3_29_port);
   U3133 : INV_X1 port map( A => n13854, ZN => n12475);
   U3134 : NOR2_X2 port map( A1 => n8445, A2 => n8446, ZN => 
                           DataPath_RF_internal_inloc_data_3_27_port);
   U3135 : INV_X1 port map( A => n13856, ZN => n12395);
   U3136 : NOR2_X2 port map( A1 => n8443, A2 => n8444, ZN => 
                           DataPath_RF_internal_inloc_data_3_26_port);
   U3137 : INV_X1 port map( A => n13857, ZN => n12355);
   U3138 : NOR2_X2 port map( A1 => n8441, A2 => n8442, ZN => 
                           DataPath_RF_internal_inloc_data_3_25_port);
   U3139 : INV_X1 port map( A => n13858, ZN => n12315);
   U3140 : NOR2_X2 port map( A1 => n8439, A2 => n8440, ZN => 
                           DataPath_RF_internal_inloc_data_3_24_port);
   U3141 : INV_X1 port map( A => n13859, ZN => n12275);
   U3142 : NOR2_X2 port map( A1 => n8437, A2 => n8438, ZN => 
                           DataPath_RF_internal_inloc_data_3_23_port);
   U3143 : INV_X1 port map( A => n13860, ZN => n12235);
   U3144 : NOR2_X2 port map( A1 => n8435, A2 => n8436, ZN => 
                           DataPath_RF_internal_inloc_data_3_22_port);
   U3145 : INV_X1 port map( A => n13861, ZN => n12195);
   U3146 : NOR2_X2 port map( A1 => n8433, A2 => n8434, ZN => 
                           DataPath_RF_internal_inloc_data_3_21_port);
   U3147 : INV_X1 port map( A => n13862, ZN => n12155);
   U3148 : NOR2_X2 port map( A1 => n8431, A2 => n8432, ZN => 
                           DataPath_RF_internal_inloc_data_3_20_port);
   U3149 : INV_X1 port map( A => n13863, ZN => n12115);
   U3150 : NOR2_X2 port map( A1 => n8429, A2 => n8430, ZN => 
                           DataPath_RF_internal_inloc_data_3_19_port);
   U3151 : INV_X1 port map( A => n13865, ZN => n12035);
   U3152 : NOR2_X2 port map( A1 => n8427, A2 => n8428, ZN => 
                           DataPath_RF_internal_inloc_data_3_18_port);
   U3153 : INV_X1 port map( A => n13866, ZN => n11995);
   U3154 : NOR2_X2 port map( A1 => n8425, A2 => n8426, ZN => 
                           DataPath_RF_internal_inloc_data_3_17_port);
   U3155 : INV_X1 port map( A => n13867, ZN => n11955);
   U3156 : NOR2_X2 port map( A1 => n8423, A2 => n8424, ZN => 
                           DataPath_RF_internal_inloc_data_3_16_port);
   U3157 : INV_X1 port map( A => n13868, ZN => n11915);
   U3158 : NOR2_X2 port map( A1 => n8421, A2 => n8422, ZN => 
                           DataPath_RF_internal_inloc_data_3_15_port);
   U3159 : INV_X1 port map( A => n13901, ZN => n11876);
   U3160 : NOR2_X2 port map( A1 => n8395, A2 => n8396, ZN => 
                           DataPath_RF_internal_inloc_data_3_2_port);
   U3161 : INV_X1 port map( A => n13853, ZN => n12515);
   U3162 : NOR2_X2 port map( A1 => n8393, A2 => n8394, ZN => 
                           DataPath_RF_internal_inloc_data_3_1_port);
   U3163 : INV_X1 port map( A => n13864, ZN => n12075);
   U3164 : NOR2_X2 port map( A1 => n8389, A2 => n8390, ZN => 
                           DataPath_RF_internal_inloc_data_4_31_port);
   U3165 : INV_X1 port map( A => n14107, ZN => n12603);
   U3166 : NOR2_X2 port map( A1 => n8387, A2 => n8388, ZN => 
                           DataPath_RF_internal_inloc_data_4_30_port);
   U3167 : INV_X1 port map( A => n14108, ZN => n12563);
   U3168 : NOR2_X2 port map( A1 => n8385, A2 => n8386, ZN => 
                           DataPath_RF_internal_inloc_data_4_29_port);
   U3169 : INV_X1 port map( A => n14110, ZN => n12483);
   U3170 : NOR2_X2 port map( A1 => n8381, A2 => n8382, ZN => 
                           DataPath_RF_internal_inloc_data_4_27_port);
   U3171 : INV_X1 port map( A => n14112, ZN => n12403);
   U3172 : NOR2_X2 port map( A1 => n8379, A2 => n8380, ZN => 
                           DataPath_RF_internal_inloc_data_4_26_port);
   U3173 : INV_X1 port map( A => n14113, ZN => n12363);
   U3174 : NOR2_X2 port map( A1 => n8377, A2 => n8378, ZN => 
                           DataPath_RF_internal_inloc_data_4_25_port);
   U3175 : INV_X1 port map( A => n14114, ZN => n12323);
   U3176 : NOR2_X2 port map( A1 => n8375, A2 => n8376, ZN => 
                           DataPath_RF_internal_inloc_data_4_24_port);
   U3177 : INV_X1 port map( A => n14115, ZN => n12283);
   U3178 : NOR2_X2 port map( A1 => n8373, A2 => n8374, ZN => 
                           DataPath_RF_internal_inloc_data_4_23_port);
   U3179 : INV_X1 port map( A => n14116, ZN => n12243);
   U3180 : NOR2_X2 port map( A1 => n8371, A2 => n8372, ZN => 
                           DataPath_RF_internal_inloc_data_4_22_port);
   U3181 : INV_X1 port map( A => n14117, ZN => n12203);
   U3182 : NOR2_X2 port map( A1 => n8369, A2 => n8370, ZN => 
                           DataPath_RF_internal_inloc_data_4_21_port);
   U3183 : INV_X1 port map( A => n14118, ZN => n12163);
   U3184 : NOR2_X2 port map( A1 => n8367, A2 => n8368, ZN => 
                           DataPath_RF_internal_inloc_data_4_20_port);
   U3185 : INV_X1 port map( A => n14119, ZN => n12123);
   U3186 : NOR2_X2 port map( A1 => n8365, A2 => n8366, ZN => 
                           DataPath_RF_internal_inloc_data_4_19_port);
   U3187 : INV_X1 port map( A => n14121, ZN => n12043);
   U3188 : NOR2_X2 port map( A1 => n8363, A2 => n8364, ZN => 
                           DataPath_RF_internal_inloc_data_4_18_port);
   U3189 : INV_X1 port map( A => n14122, ZN => n12003);
   U3190 : NOR2_X2 port map( A1 => n8361, A2 => n8362, ZN => 
                           DataPath_RF_internal_inloc_data_4_17_port);
   U3191 : INV_X1 port map( A => n14123, ZN => n11963);
   U3192 : NOR2_X2 port map( A1 => n8359, A2 => n8360, ZN => 
                           DataPath_RF_internal_inloc_data_4_16_port);
   U3193 : INV_X1 port map( A => n14124, ZN => n11923);
   U3194 : NOR2_X2 port map( A1 => n8357, A2 => n8358, ZN => 
                           DataPath_RF_internal_inloc_data_4_15_port);
   U3195 : INV_X1 port map( A => n14157, ZN => n11884);
   U3196 : NOR2_X2 port map( A1 => n8331, A2 => n8332, ZN => 
                           DataPath_RF_internal_inloc_data_4_2_port);
   U3197 : INV_X1 port map( A => n14109, ZN => n12523);
   U3198 : NOR2_X2 port map( A1 => n8329, A2 => n8330, ZN => 
                           DataPath_RF_internal_inloc_data_4_1_port);
   U3199 : INV_X1 port map( A => n14120, ZN => n12083);
   U3200 : OAI22_X1 port map( A1 => n8283, A2 => n2984, B1 => n8284, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n198);
   U3201 : OAI22_X1 port map( A1 => n8297, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8296, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n487);
   U3202 : OAI22_X1 port map( A1 => n8298, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8297, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n472);
   U3203 : OAI22_X1 port map( A1 => n8282, A2 => n2984, B1 => n8283, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n206);
   U3204 : OAI22_X1 port map( A1 => n520, A2 => n2984, B1 => n8293, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n450);
   U3205 : OAI22_X1 port map( A1 => n8284, A2 => n2984, B1 => n8285, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n189);
   U3206 : OAI22_X1 port map( A1 => n11494, A2 => n2984, B1 => n8282, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n216);
   U3207 : OAI22_X1 port map( A1 => n8283, A2 => n1769, B1 => n8282, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n267);
   U3208 : OAI22_X1 port map( A1 => n8293, A2 => n2984, B1 => n8294, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n437);
   U3209 : OAI22_X1 port map( A1 => n11490, A2 => n2984, B1 => n520, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n460);
   U3210 : OAI22_X1 port map( A1 => n11496, A2 => n2984, B1 => n11495, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n410);
   U3211 : BUF_X1 port map( A => n14362, Z => n2504);
   U3212 : BUF_X1 port map( A => n14362, Z => n2505);
   U3213 : BUF_X1 port map( A => n14396, Z => n2510);
   U3214 : BUF_X1 port map( A => n14396, Z => n2511);
   U3215 : BUF_X1 port map( A => n14430, Z => n2516);
   U3216 : BUF_X1 port map( A => n14430, Z => n2517);
   U3217 : BUF_X1 port map( A => n14464, Z => n2522);
   U3218 : BUF_X1 port map( A => n14464, Z => n2523);
   U3219 : BUF_X1 port map( A => n14498, Z => n2528);
   U3220 : BUF_X1 port map( A => n14498, Z => n2529);
   U3221 : BUF_X1 port map( A => n14532, Z => n2534);
   U3222 : BUF_X1 port map( A => n14532, Z => n2535);
   U3223 : BUF_X1 port map( A => n14566, Z => n2540);
   U3224 : BUF_X1 port map( A => n14566, Z => n2541);
   U3225 : BUF_X1 port map( A => n14600, Z => n2546);
   U3226 : BUF_X1 port map( A => n14600, Z => n2547);
   U3227 : BUF_X1 port map( A => n14634, Z => n2552);
   U3228 : BUF_X1 port map( A => n14634, Z => n2553);
   U3229 : BUF_X1 port map( A => n14668, Z => n2558);
   U3230 : BUF_X1 port map( A => n14668, Z => n2559);
   U3231 : BUF_X1 port map( A => n14702, Z => n2564);
   U3232 : BUF_X1 port map( A => n14702, Z => n2565);
   U3233 : BUF_X1 port map( A => n14736, Z => n2570);
   U3234 : BUF_X1 port map( A => n14736, Z => n2571);
   U3235 : BUF_X1 port map( A => n14770, Z => n2576);
   U3236 : BUF_X1 port map( A => n14770, Z => n2577);
   U3237 : BUF_X1 port map( A => n14804, Z => n2582);
   U3238 : BUF_X1 port map( A => n14804, Z => n2583);
   U3239 : BUF_X1 port map( A => n14838, Z => n2588);
   U3240 : BUF_X1 port map( A => n14838, Z => n2589);
   U3241 : BUF_X1 port map( A => n14872, Z => n2594);
   U3242 : BUF_X1 port map( A => n14872, Z => n2595);
   U3243 : BUF_X1 port map( A => n14906, Z => n2600);
   U3244 : BUF_X1 port map( A => n14906, Z => n2601);
   U3245 : BUF_X1 port map( A => n14940, Z => n2606);
   U3246 : BUF_X1 port map( A => n14940, Z => n2607);
   U3247 : BUF_X1 port map( A => n14974, Z => n2612);
   U3248 : BUF_X1 port map( A => n14974, Z => n2613);
   U3249 : BUF_X1 port map( A => n15008, Z => n2618);
   U3250 : BUF_X1 port map( A => n15008, Z => n2619);
   U3251 : BUF_X1 port map( A => n15042, Z => n2624);
   U3252 : BUF_X1 port map( A => n15042, Z => n2625);
   U3253 : BUF_X1 port map( A => n15076, Z => n2630);
   U3254 : BUF_X1 port map( A => n15076, Z => n2631);
   U3255 : BUF_X1 port map( A => n15110, Z => n2636);
   U3256 : BUF_X1 port map( A => n15110, Z => n2637);
   U3257 : BUF_X1 port map( A => n15144, Z => n2642);
   U3258 : BUF_X1 port map( A => n15144, Z => n2643);
   U3259 : BUF_X1 port map( A => n15178, Z => n2648);
   U3260 : BUF_X1 port map( A => n15178, Z => n2649);
   U3261 : BUF_X1 port map( A => n15212, Z => n2654);
   U3262 : BUF_X1 port map( A => n15212, Z => n2655);
   U3263 : BUF_X1 port map( A => n15246, Z => n2660);
   U3264 : BUF_X1 port map( A => n15246, Z => n2661);
   U3265 : BUF_X1 port map( A => n15280, Z => n2666);
   U3266 : BUF_X1 port map( A => n15280, Z => n2667);
   U3267 : BUF_X1 port map( A => n15314, Z => n2672);
   U3268 : BUF_X1 port map( A => n15314, Z => n2673);
   U3269 : BUF_X1 port map( A => n15348, Z => n2678);
   U3270 : BUF_X1 port map( A => n15348, Z => n2679);
   U3271 : BUF_X1 port map( A => n15382, Z => n2684);
   U3272 : BUF_X1 port map( A => n15382, Z => n2685);
   U3273 : BUF_X1 port map( A => n15416, Z => n2690);
   U3274 : BUF_X1 port map( A => n15416, Z => n2691);
   U3275 : BUF_X1 port map( A => n15450, Z => n2696);
   U3276 : BUF_X1 port map( A => n15450, Z => n2697);
   U3277 : BUF_X1 port map( A => n15484, Z => n2702);
   U3278 : BUF_X1 port map( A => n15484, Z => n2703);
   U3279 : BUF_X1 port map( A => n15518, Z => n2708);
   U3280 : BUF_X1 port map( A => n15518, Z => n2709);
   U3281 : BUF_X1 port map( A => n15552, Z => n2714);
   U3282 : BUF_X1 port map( A => n15552, Z => n2715);
   U3283 : BUF_X1 port map( A => n15586, Z => n2720);
   U3284 : BUF_X1 port map( A => n15586, Z => n2721);
   U3285 : BUF_X1 port map( A => n15620, Z => n2726);
   U3286 : BUF_X1 port map( A => n15620, Z => n2727);
   U3287 : BUF_X1 port map( A => n15654, Z => n2732);
   U3288 : BUF_X1 port map( A => n15654, Z => n2733);
   U3289 : BUF_X1 port map( A => n15688, Z => n2738);
   U3290 : BUF_X1 port map( A => n15688, Z => n2739);
   U3291 : BUF_X1 port map( A => n15722, Z => n2744);
   U3292 : BUF_X1 port map( A => n15722, Z => n2745);
   U3293 : BUF_X1 port map( A => n15756, Z => n2750);
   U3294 : BUF_X1 port map( A => n15756, Z => n2751);
   U3295 : BUF_X1 port map( A => n15790, Z => n2756);
   U3296 : BUF_X1 port map( A => n15790, Z => n2757);
   U3297 : BUF_X1 port map( A => n15824, Z => n2762);
   U3298 : BUF_X1 port map( A => n15824, Z => n2763);
   U3299 : BUF_X1 port map( A => n15858, Z => n2768);
   U3300 : BUF_X1 port map( A => n15858, Z => n2769);
   U3301 : BUF_X1 port map( A => n15892, Z => n2774);
   U3302 : BUF_X1 port map( A => n15892, Z => n2775);
   U3303 : BUF_X1 port map( A => n15926, Z => n2780);
   U3304 : BUF_X1 port map( A => n15926, Z => n2781);
   U3305 : BUF_X1 port map( A => n15960, Z => n2786);
   U3306 : BUF_X1 port map( A => n15960, Z => n2787);
   U3307 : BUF_X1 port map( A => n15994, Z => n2792);
   U3308 : BUF_X1 port map( A => n15994, Z => n2793);
   U3309 : BUF_X1 port map( A => n16028, Z => n2798);
   U3310 : BUF_X1 port map( A => n16028, Z => n2799);
   U3311 : BUF_X1 port map( A => n16062, Z => n2804);
   U3312 : BUF_X1 port map( A => n16062, Z => n2805);
   U3313 : BUF_X1 port map( A => n16096, Z => n2810);
   U3314 : BUF_X1 port map( A => n16096, Z => n2811);
   U3315 : BUF_X1 port map( A => n16130, Z => n2816);
   U3316 : BUF_X1 port map( A => n16130, Z => n2817);
   U3317 : BUF_X1 port map( A => n16164, Z => n2822);
   U3318 : BUF_X1 port map( A => n16164, Z => n2823);
   U3319 : BUF_X1 port map( A => n16198, Z => n2828);
   U3320 : BUF_X1 port map( A => n16198, Z => n2829);
   U3321 : BUF_X1 port map( A => n16232, Z => n2834);
   U3322 : BUF_X1 port map( A => n16232, Z => n2835);
   U3323 : BUF_X1 port map( A => n16266, Z => n2840);
   U3324 : BUF_X1 port map( A => n16266, Z => n2841);
   U3325 : BUF_X1 port map( A => n16300, Z => n2846);
   U3326 : BUF_X1 port map( A => n16300, Z => n2847);
   U3327 : BUF_X1 port map( A => n16334, Z => n2852);
   U3328 : BUF_X1 port map( A => n16334, Z => n2853);
   U3329 : BUF_X1 port map( A => n16368, Z => n2858);
   U3330 : BUF_X1 port map( A => n16368, Z => n2859);
   U3331 : BUF_X1 port map( A => n16402, Z => n2864);
   U3332 : BUF_X1 port map( A => n16402, Z => n2865);
   U3333 : BUF_X1 port map( A => n16436, Z => n2870);
   U3334 : BUF_X1 port map( A => n16436, Z => n2871);
   U3335 : BUF_X1 port map( A => n16470, Z => n2876);
   U3336 : BUF_X1 port map( A => n16470, Z => n2877);
   U3337 : BUF_X1 port map( A => n16504, Z => n2882);
   U3338 : BUF_X1 port map( A => n16504, Z => n2883);
   U3339 : BUF_X1 port map( A => n16538, Z => n2888);
   U3340 : BUF_X1 port map( A => n16538, Z => n2889);
   U3341 : BUF_X1 port map( A => n16572, Z => n2894);
   U3342 : BUF_X1 port map( A => n16572, Z => n2895);
   U3343 : BUF_X1 port map( A => n16606, Z => n2900);
   U3344 : BUF_X1 port map( A => n16606, Z => n2901);
   U3345 : BUF_X1 port map( A => n16640, Z => n2906);
   U3346 : BUF_X1 port map( A => n16640, Z => n2907);
   U3347 : BUF_X1 port map( A => n16674, Z => n2912);
   U3348 : BUF_X1 port map( A => n16674, Z => n2913);
   U3349 : BUF_X1 port map( A => n16708, Z => n2918);
   U3350 : BUF_X1 port map( A => n16708, Z => n2919);
   U3351 : BUF_X1 port map( A => n16742, Z => n2924);
   U3352 : BUF_X1 port map( A => n16742, Z => n2925);
   U3353 : BUF_X1 port map( A => n16776, Z => n2930);
   U3354 : BUF_X1 port map( A => n16776, Z => n2931);
   U3355 : BUF_X1 port map( A => n16810, Z => n2936);
   U3356 : BUF_X1 port map( A => n16810, Z => n2937);
   U3357 : BUF_X1 port map( A => n16844, Z => n2942);
   U3358 : BUF_X1 port map( A => n16844, Z => n2943);
   U3359 : BUF_X1 port map( A => n16878, Z => n2948);
   U3360 : BUF_X1 port map( A => n16878, Z => n2949);
   U3361 : BUF_X1 port map( A => n16912, Z => n2954);
   U3362 : BUF_X1 port map( A => n16912, Z => n2955);
   U3363 : BUF_X1 port map( A => n16946, Z => n2960);
   U3364 : BUF_X1 port map( A => n16946, Z => n2961);
   U3365 : BUF_X1 port map( A => n16980, Z => n2966);
   U3366 : BUF_X1 port map( A => n16980, Z => n2967);
   U3367 : BUF_X1 port map( A => n17014, Z => n2972);
   U3368 : BUF_X1 port map( A => n17014, Z => n2973);
   U3369 : BUF_X1 port map( A => n17048, Z => n2978);
   U3370 : BUF_X1 port map( A => n17048, Z => n2979);
   U3371 : OAI22_X1 port map( A1 => n8294, A2 => n2984, B1 => n8295, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n424);
   U3372 : OAI22_X1 port map( A1 => n8295, A2 => n2984, B1 => n8296, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n397);
   U3373 : OAI22_X1 port map( A1 => n8297, A2 => n1769, B1 => n8296, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n430);
   U3374 : OAI22_X1 port map( A1 => n8296, A2 => n1769, B1 => n8295, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n443);
   U3375 : OAI22_X1 port map( A1 => n8296, A2 => n2984, B1 => n8297, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n385);
   U3376 : OAI22_X1 port map( A1 => n8302, A2 => n1769, B1 => n8301, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n378);
   U3377 : OAI22_X1 port map( A1 => n8301, A2 => n1769, B1 => n8298, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n390);
   U3378 : OAI22_X1 port map( A1 => n8317, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8308, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n289);
   U3379 : OAI22_X1 port map( A1 => n8308, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8318, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n303);
   U3380 : OAI22_X1 port map( A1 => n8318, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8313, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n317);
   U3381 : BUF_X1 port map( A => n14362, Z => n2506);
   U3382 : BUF_X1 port map( A => n14396, Z => n2512);
   U3383 : BUF_X1 port map( A => n14430, Z => n2518);
   U3384 : BUF_X1 port map( A => n14464, Z => n2524);
   U3385 : BUF_X1 port map( A => n14498, Z => n2530);
   U3386 : BUF_X1 port map( A => n14532, Z => n2536);
   U3387 : BUF_X1 port map( A => n14566, Z => n2542);
   U3388 : BUF_X1 port map( A => n14600, Z => n2548);
   U3389 : BUF_X1 port map( A => n14634, Z => n2554);
   U3390 : BUF_X1 port map( A => n14668, Z => n2560);
   U3391 : BUF_X1 port map( A => n14702, Z => n2566);
   U3392 : BUF_X1 port map( A => n14736, Z => n2572);
   U3393 : BUF_X1 port map( A => n14770, Z => n2578);
   U3394 : BUF_X1 port map( A => n14804, Z => n2584);
   U3395 : BUF_X1 port map( A => n14838, Z => n2590);
   U3396 : BUF_X1 port map( A => n14872, Z => n2596);
   U3397 : BUF_X1 port map( A => n14906, Z => n2602);
   U3398 : BUF_X1 port map( A => n14940, Z => n2608);
   U3399 : BUF_X1 port map( A => n14974, Z => n2614);
   U3400 : BUF_X1 port map( A => n15008, Z => n2620);
   U3401 : BUF_X1 port map( A => n15042, Z => n2626);
   U3402 : BUF_X1 port map( A => n15076, Z => n2632);
   U3403 : BUF_X1 port map( A => n15110, Z => n2638);
   U3404 : BUF_X1 port map( A => n15144, Z => n2644);
   U3405 : BUF_X1 port map( A => n15178, Z => n2650);
   U3406 : BUF_X1 port map( A => n15212, Z => n2656);
   U3407 : BUF_X1 port map( A => n15246, Z => n2662);
   U3408 : BUF_X1 port map( A => n15280, Z => n2668);
   U3409 : BUF_X1 port map( A => n15314, Z => n2674);
   U3410 : BUF_X1 port map( A => n15348, Z => n2680);
   U3411 : BUF_X1 port map( A => n15382, Z => n2686);
   U3412 : BUF_X1 port map( A => n15416, Z => n2692);
   U3413 : BUF_X1 port map( A => n15450, Z => n2698);
   U3414 : BUF_X1 port map( A => n15484, Z => n2704);
   U3415 : BUF_X1 port map( A => n15518, Z => n2710);
   U3416 : BUF_X1 port map( A => n15552, Z => n2716);
   U3417 : BUF_X1 port map( A => n15586, Z => n2722);
   U3418 : BUF_X1 port map( A => n15620, Z => n2728);
   U3419 : BUF_X1 port map( A => n15654, Z => n2734);
   U3420 : BUF_X1 port map( A => n15688, Z => n2740);
   U3421 : BUF_X1 port map( A => n15722, Z => n2746);
   U3422 : BUF_X1 port map( A => n15756, Z => n2752);
   U3423 : BUF_X1 port map( A => n15790, Z => n2758);
   U3424 : BUF_X1 port map( A => n15824, Z => n2764);
   U3425 : BUF_X1 port map( A => n15858, Z => n2770);
   U3426 : BUF_X1 port map( A => n15892, Z => n2776);
   U3427 : BUF_X1 port map( A => n15926, Z => n2782);
   U3428 : BUF_X1 port map( A => n15960, Z => n2788);
   U3429 : BUF_X1 port map( A => n15994, Z => n2794);
   U3430 : BUF_X1 port map( A => n16028, Z => n2800);
   U3431 : BUF_X1 port map( A => n16062, Z => n2806);
   U3432 : BUF_X1 port map( A => n16096, Z => n2812);
   U3433 : BUF_X1 port map( A => n16130, Z => n2818);
   U3434 : BUF_X1 port map( A => n16164, Z => n2824);
   U3435 : BUF_X1 port map( A => n16198, Z => n2830);
   U3436 : BUF_X1 port map( A => n16232, Z => n2836);
   U3437 : BUF_X1 port map( A => n16266, Z => n2842);
   U3438 : BUF_X1 port map( A => n16300, Z => n2848);
   U3439 : BUF_X1 port map( A => n16334, Z => n2854);
   U3440 : BUF_X1 port map( A => n16368, Z => n2860);
   U3441 : BUF_X1 port map( A => n16402, Z => n2866);
   U3442 : BUF_X1 port map( A => n16436, Z => n2872);
   U3443 : BUF_X1 port map( A => n16470, Z => n2878);
   U3444 : BUF_X1 port map( A => n16504, Z => n2884);
   U3445 : BUF_X1 port map( A => n16538, Z => n2890);
   U3446 : BUF_X1 port map( A => n16572, Z => n2896);
   U3447 : BUF_X1 port map( A => n16606, Z => n2902);
   U3448 : BUF_X1 port map( A => n16640, Z => n2908);
   U3449 : BUF_X1 port map( A => n16674, Z => n2914);
   U3450 : BUF_X1 port map( A => n16708, Z => n2920);
   U3451 : BUF_X1 port map( A => n16742, Z => n2926);
   U3452 : BUF_X1 port map( A => n16776, Z => n2932);
   U3453 : BUF_X1 port map( A => n16810, Z => n2938);
   U3454 : BUF_X1 port map( A => n16844, Z => n2944);
   U3455 : BUF_X1 port map( A => n16878, Z => n2950);
   U3456 : BUF_X1 port map( A => n16912, Z => n2956);
   U3457 : BUF_X1 port map( A => n16946, Z => n2962);
   U3458 : BUF_X1 port map( A => n16980, Z => n2968);
   U3459 : BUF_X1 port map( A => n17014, Z => n2974);
   U3460 : BUF_X1 port map( A => n17048, Z => n2980);
   U3461 : XNOR2_X1 port map( A => n4271, B => n2146, ZN => n1797);
   U3462 : BUF_X1 port map( A => n3373, Z => n3371);
   U3463 : BUF_X1 port map( A => n3373, Z => n3372);
   U3464 : BUF_X1 port map( A => n3373, Z => n3370);
   U3465 : BUF_X1 port map( A => n3485, Z => n3482);
   U3466 : BUF_X1 port map( A => n3485, Z => n3484);
   U3467 : BUF_X1 port map( A => n3485, Z => n3483);
   U3468 : BUF_X1 port map( A => n3597, Z => n3594);
   U3469 : BUF_X1 port map( A => n3597, Z => n3596);
   U3470 : BUF_X1 port map( A => n3597, Z => n3595);
   U3471 : BUF_X1 port map( A => n3821, Z => n3818);
   U3472 : BUF_X1 port map( A => n3821, Z => n3820);
   U3473 : BUF_X1 port map( A => n3821, Z => n3819);
   U3474 : BUF_X1 port map( A => n3374, Z => n3368);
   U3475 : BUF_X1 port map( A => n3374, Z => n3369);
   U3476 : BUF_X1 port map( A => n3486, Z => n3480);
   U3477 : BUF_X1 port map( A => n3486, Z => n3481);
   U3478 : BUF_X1 port map( A => n3598, Z => n3592);
   U3479 : BUF_X1 port map( A => n3598, Z => n3593);
   U3480 : BUF_X1 port map( A => n3822, Z => n3816);
   U3481 : BUF_X1 port map( A => n3822, Z => n3817);
   U3482 : AND2_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_28_port, A2
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_26_port,
                           ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_28_port);
   U3483 : AND2_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_26_port, A2
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_25_port,
                           ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_26_port);
   U3484 : AND2_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_24_port, A2
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_20_port,
                           ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_3_24_port);
   U3485 : BUF_X1 port map( A => n3630, Z => n3620);
   U3486 : NOR2_X1 port map( A1 => n2491, A2 => n4182, ZN => n14260);
   U3487 : BUF_X1 port map( A => n14294, Z => n2492);
   U3488 : BUF_X1 port map( A => n14294, Z => n2493);
   U3489 : BUF_X1 port map( A => n14328, Z => n2498);
   U3490 : BUF_X1 port map( A => n14328, Z => n2499);
   U3491 : BUF_X1 port map( A => n14294, Z => n2494);
   U3492 : BUF_X1 port map( A => n14328, Z => n2500);
   U3493 : BUF_X1 port map( A => n3392, Z => n3315);
   U3494 : BUF_X1 port map( A => n3394, Z => n3308);
   U3495 : BUF_X1 port map( A => n3391, Z => n3317);
   U3496 : BUF_X1 port map( A => n3394, Z => n3309);
   U3497 : BUF_X1 port map( A => n3393, Z => n3312);
   U3498 : BUF_X1 port map( A => n3393, Z => n3310);
   U3499 : BUF_X1 port map( A => n3392, Z => n3313);
   U3500 : BUF_X1 port map( A => n3393, Z => n3311);
   U3501 : BUF_X1 port map( A => n3392, Z => n3314);
   U3502 : BUF_X1 port map( A => n3391, Z => n3316);
   U3503 : BUF_X1 port map( A => n3394, Z => n3307);
   U3504 : BUF_X1 port map( A => n3504, Z => n3427);
   U3505 : BUF_X1 port map( A => n3506, Z => n3420);
   U3506 : BUF_X1 port map( A => n3503, Z => n3429);
   U3507 : BUF_X1 port map( A => n3506, Z => n3421);
   U3508 : BUF_X1 port map( A => n3505, Z => n3424);
   U3509 : BUF_X1 port map( A => n3505, Z => n3422);
   U3510 : BUF_X1 port map( A => n3504, Z => n3425);
   U3511 : BUF_X1 port map( A => n3505, Z => n3423);
   U3512 : BUF_X1 port map( A => n3504, Z => n3426);
   U3513 : BUF_X1 port map( A => n3503, Z => n3428);
   U3514 : BUF_X1 port map( A => n3506, Z => n3419);
   U3515 : BUF_X1 port map( A => n3616, Z => n3539);
   U3516 : BUF_X1 port map( A => n3618, Z => n3532);
   U3517 : BUF_X1 port map( A => n3615, Z => n3541);
   U3518 : BUF_X1 port map( A => n3618, Z => n3533);
   U3519 : BUF_X1 port map( A => n3617, Z => n3536);
   U3520 : BUF_X1 port map( A => n3617, Z => n3534);
   U3521 : BUF_X1 port map( A => n3616, Z => n3537);
   U3522 : BUF_X1 port map( A => n3617, Z => n3535);
   U3523 : BUF_X1 port map( A => n3616, Z => n3538);
   U3524 : BUF_X1 port map( A => n3615, Z => n3540);
   U3525 : BUF_X1 port map( A => n3618, Z => n3531);
   U3526 : BUF_X1 port map( A => n3840, Z => n3763);
   U3527 : BUF_X1 port map( A => n3842, Z => n3756);
   U3528 : BUF_X1 port map( A => n3839, Z => n3765);
   U3529 : BUF_X1 port map( A => n3842, Z => n3757);
   U3530 : BUF_X1 port map( A => n3841, Z => n3760);
   U3531 : BUF_X1 port map( A => n3841, Z => n3758);
   U3532 : BUF_X1 port map( A => n3840, Z => n3761);
   U3533 : BUF_X1 port map( A => n3841, Z => n3759);
   U3534 : BUF_X1 port map( A => n3840, Z => n3762);
   U3535 : BUF_X1 port map( A => n3839, Z => n3764);
   U3536 : BUF_X1 port map( A => n3842, Z => n3755);
   U3537 : BUF_X1 port map( A => n3382, Z => n3344);
   U3538 : BUF_X1 port map( A => n3376, Z => n3363);
   U3539 : BUF_X1 port map( A => n3386, Z => n3332);
   U3540 : BUF_X1 port map( A => n3391, Z => n3318);
   U3541 : BUF_X1 port map( A => n3378, Z => n3357);
   U3542 : BUF_X1 port map( A => n3380, Z => n3351);
   U3543 : BUF_X1 port map( A => n3384, Z => n3339);
   U3544 : BUF_X1 port map( A => n3375, Z => n3364);
   U3545 : BUF_X1 port map( A => n3382, Z => n3345);
   U3546 : BUF_X1 port map( A => n3386, Z => n3333);
   U3547 : BUF_X1 port map( A => n3377, Z => n3358);
   U3548 : BUF_X1 port map( A => n3379, Z => n3353);
   U3549 : BUF_X1 port map( A => n3383, Z => n3341);
   U3550 : BUF_X1 port map( A => n3381, Z => n3347);
   U3551 : BUF_X1 port map( A => n3385, Z => n3335);
   U3552 : BUF_X1 port map( A => n3390, Z => n3320);
   U3553 : BUF_X1 port map( A => n3377, Z => n3360);
   U3554 : BUF_X1 port map( A => n3375, Z => n3366);
   U3555 : BUF_X1 port map( A => n3387, Z => n3329);
   U3556 : BUF_X1 port map( A => n3389, Z => n3324);
   U3557 : BUF_X1 port map( A => n3379, Z => n3354);
   U3558 : BUF_X1 port map( A => n3383, Z => n3342);
   U3559 : BUF_X1 port map( A => n3381, Z => n3348);
   U3560 : BUF_X1 port map( A => n3374, Z => n3367);
   U3561 : BUF_X1 port map( A => n3385, Z => n3336);
   U3562 : BUF_X1 port map( A => n3390, Z => n3321);
   U3563 : BUF_X1 port map( A => n3376, Z => n3361);
   U3564 : BUF_X1 port map( A => n3388, Z => n3327);
   U3565 : BUF_X1 port map( A => n3387, Z => n3330);
   U3566 : BUF_X1 port map( A => n3388, Z => n3325);
   U3567 : BUF_X1 port map( A => n3382, Z => n3343);
   U3568 : BUF_X1 port map( A => n3380, Z => n3350);
   U3569 : BUF_X1 port map( A => n3384, Z => n3338);
   U3570 : BUF_X1 port map( A => n3389, Z => n3323);
   U3571 : BUF_X1 port map( A => n3389, Z => n3322);
   U3572 : BUF_X1 port map( A => n3375, Z => n3365);
   U3573 : BUF_X1 port map( A => n3377, Z => n3359);
   U3574 : BUF_X1 port map( A => n3379, Z => n3352);
   U3575 : BUF_X1 port map( A => n3381, Z => n3346);
   U3576 : BUF_X1 port map( A => n3383, Z => n3340);
   U3577 : BUF_X1 port map( A => n3385, Z => n3334);
   U3578 : BUF_X1 port map( A => n3387, Z => n3328);
   U3579 : BUF_X1 port map( A => n3378, Z => n3356);
   U3580 : BUF_X1 port map( A => n3384, Z => n3337);
   U3581 : BUF_X1 port map( A => n3386, Z => n3331);
   U3582 : BUF_X1 port map( A => n3388, Z => n3326);
   U3583 : BUF_X1 port map( A => n3376, Z => n3362);
   U3584 : BUF_X1 port map( A => n3378, Z => n3355);
   U3585 : BUF_X1 port map( A => n3380, Z => n3349);
   U3586 : BUF_X1 port map( A => n3390, Z => n3319);
   U3587 : BUF_X1 port map( A => n3494, Z => n3456);
   U3588 : BUF_X1 port map( A => n3488, Z => n3475);
   U3589 : BUF_X1 port map( A => n3498, Z => n3444);
   U3590 : BUF_X1 port map( A => n3503, Z => n3430);
   U3591 : BUF_X1 port map( A => n3490, Z => n3469);
   U3592 : BUF_X1 port map( A => n3492, Z => n3463);
   U3593 : BUF_X1 port map( A => n3496, Z => n3451);
   U3594 : BUF_X1 port map( A => n3487, Z => n3476);
   U3595 : BUF_X1 port map( A => n3494, Z => n3457);
   U3596 : BUF_X1 port map( A => n3498, Z => n3445);
   U3597 : BUF_X1 port map( A => n3489, Z => n3470);
   U3598 : BUF_X1 port map( A => n3491, Z => n3465);
   U3599 : BUF_X1 port map( A => n3495, Z => n3453);
   U3600 : BUF_X1 port map( A => n3493, Z => n3459);
   U3601 : BUF_X1 port map( A => n3502, Z => n3432);
   U3602 : BUF_X1 port map( A => n3497, Z => n3447);
   U3603 : BUF_X1 port map( A => n3489, Z => n3472);
   U3604 : BUF_X1 port map( A => n3487, Z => n3478);
   U3605 : BUF_X1 port map( A => n3499, Z => n3441);
   U3606 : BUF_X1 port map( A => n3501, Z => n3436);
   U3607 : BUF_X1 port map( A => n3491, Z => n3466);
   U3608 : BUF_X1 port map( A => n3495, Z => n3454);
   U3609 : BUF_X1 port map( A => n3493, Z => n3460);
   U3610 : BUF_X1 port map( A => n3486, Z => n3479);
   U3611 : BUF_X1 port map( A => n3497, Z => n3448);
   U3612 : BUF_X1 port map( A => n3502, Z => n3433);
   U3613 : BUF_X1 port map( A => n3488, Z => n3473);
   U3614 : BUF_X1 port map( A => n3500, Z => n3439);
   U3615 : BUF_X1 port map( A => n3499, Z => n3442);
   U3616 : BUF_X1 port map( A => n3500, Z => n3437);
   U3617 : BUF_X1 port map( A => n3494, Z => n3455);
   U3618 : BUF_X1 port map( A => n3492, Z => n3462);
   U3619 : BUF_X1 port map( A => n3496, Z => n3450);
   U3620 : BUF_X1 port map( A => n3501, Z => n3435);
   U3621 : BUF_X1 port map( A => n3501, Z => n3434);
   U3622 : BUF_X1 port map( A => n3487, Z => n3477);
   U3623 : BUF_X1 port map( A => n3489, Z => n3471);
   U3624 : BUF_X1 port map( A => n3491, Z => n3464);
   U3625 : BUF_X1 port map( A => n3493, Z => n3458);
   U3626 : BUF_X1 port map( A => n3495, Z => n3452);
   U3627 : BUF_X1 port map( A => n3497, Z => n3446);
   U3628 : BUF_X1 port map( A => n3499, Z => n3440);
   U3629 : BUF_X1 port map( A => n3488, Z => n3474);
   U3630 : BUF_X1 port map( A => n3490, Z => n3467);
   U3631 : BUF_X1 port map( A => n3492, Z => n3461);
   U3632 : BUF_X1 port map( A => n3502, Z => n3431);
   U3633 : BUF_X1 port map( A => n3490, Z => n3468);
   U3634 : BUF_X1 port map( A => n3496, Z => n3449);
   U3635 : BUF_X1 port map( A => n3498, Z => n3443);
   U3636 : BUF_X1 port map( A => n3500, Z => n3438);
   U3637 : BUF_X1 port map( A => n3606, Z => n3568);
   U3638 : BUF_X1 port map( A => n3600, Z => n3587);
   U3639 : BUF_X1 port map( A => n3610, Z => n3556);
   U3640 : BUF_X1 port map( A => n3615, Z => n3542);
   U3641 : BUF_X1 port map( A => n3602, Z => n3581);
   U3642 : BUF_X1 port map( A => n3604, Z => n3575);
   U3643 : BUF_X1 port map( A => n3608, Z => n3563);
   U3644 : BUF_X1 port map( A => n3599, Z => n3588);
   U3645 : BUF_X1 port map( A => n3606, Z => n3569);
   U3646 : BUF_X1 port map( A => n3610, Z => n3557);
   U3647 : BUF_X1 port map( A => n3601, Z => n3582);
   U3648 : BUF_X1 port map( A => n3603, Z => n3577);
   U3649 : BUF_X1 port map( A => n3607, Z => n3565);
   U3650 : BUF_X1 port map( A => n3605, Z => n3571);
   U3651 : BUF_X1 port map( A => n3614, Z => n3544);
   U3652 : BUF_X1 port map( A => n3609, Z => n3559);
   U3653 : BUF_X1 port map( A => n3601, Z => n3584);
   U3654 : BUF_X1 port map( A => n3599, Z => n3590);
   U3655 : BUF_X1 port map( A => n3611, Z => n3553);
   U3656 : BUF_X1 port map( A => n3613, Z => n3548);
   U3657 : BUF_X1 port map( A => n3603, Z => n3578);
   U3658 : BUF_X1 port map( A => n3607, Z => n3566);
   U3659 : BUF_X1 port map( A => n3605, Z => n3572);
   U3660 : BUF_X1 port map( A => n3598, Z => n3591);
   U3661 : BUF_X1 port map( A => n3609, Z => n3560);
   U3662 : BUF_X1 port map( A => n3614, Z => n3545);
   U3663 : BUF_X1 port map( A => n3600, Z => n3585);
   U3664 : BUF_X1 port map( A => n3612, Z => n3551);
   U3665 : BUF_X1 port map( A => n3611, Z => n3554);
   U3666 : BUF_X1 port map( A => n3612, Z => n3549);
   U3667 : BUF_X1 port map( A => n3606, Z => n3567);
   U3668 : BUF_X1 port map( A => n3604, Z => n3574);
   U3669 : BUF_X1 port map( A => n3608, Z => n3562);
   U3670 : BUF_X1 port map( A => n3613, Z => n3547);
   U3671 : BUF_X1 port map( A => n3613, Z => n3546);
   U3672 : BUF_X1 port map( A => n3599, Z => n3589);
   U3673 : BUF_X1 port map( A => n3601, Z => n3583);
   U3674 : BUF_X1 port map( A => n3603, Z => n3576);
   U3675 : BUF_X1 port map( A => n3605, Z => n3570);
   U3676 : BUF_X1 port map( A => n3607, Z => n3564);
   U3677 : BUF_X1 port map( A => n3609, Z => n3558);
   U3678 : BUF_X1 port map( A => n3611, Z => n3552);
   U3679 : BUF_X1 port map( A => n3600, Z => n3586);
   U3680 : BUF_X1 port map( A => n3602, Z => n3579);
   U3681 : BUF_X1 port map( A => n3604, Z => n3573);
   U3682 : BUF_X1 port map( A => n3614, Z => n3543);
   U3683 : BUF_X1 port map( A => n3602, Z => n3580);
   U3684 : BUF_X1 port map( A => n3608, Z => n3561);
   U3685 : BUF_X1 port map( A => n3610, Z => n3555);
   U3686 : BUF_X1 port map( A => n3612, Z => n3550);
   U3687 : BUF_X1 port map( A => n3830, Z => n3792);
   U3688 : BUF_X1 port map( A => n3824, Z => n3811);
   U3689 : BUF_X1 port map( A => n3834, Z => n3780);
   U3690 : BUF_X1 port map( A => n3839, Z => n3766);
   U3691 : BUF_X1 port map( A => n3826, Z => n3805);
   U3692 : BUF_X1 port map( A => n3828, Z => n3799);
   U3693 : BUF_X1 port map( A => n3832, Z => n3787);
   U3694 : BUF_X1 port map( A => n3823, Z => n3812);
   U3695 : BUF_X1 port map( A => n3830, Z => n3793);
   U3696 : BUF_X1 port map( A => n3834, Z => n3781);
   U3697 : BUF_X1 port map( A => n3825, Z => n3806);
   U3698 : BUF_X1 port map( A => n3827, Z => n3801);
   U3699 : BUF_X1 port map( A => n3831, Z => n3789);
   U3700 : BUF_X1 port map( A => n3829, Z => n3795);
   U3701 : BUF_X1 port map( A => n3838, Z => n3768);
   U3702 : BUF_X1 port map( A => n3833, Z => n3783);
   U3703 : BUF_X1 port map( A => n3825, Z => n3808);
   U3704 : BUF_X1 port map( A => n3823, Z => n3814);
   U3705 : BUF_X1 port map( A => n3835, Z => n3777);
   U3706 : BUF_X1 port map( A => n3837, Z => n3772);
   U3707 : BUF_X1 port map( A => n3827, Z => n3802);
   U3708 : BUF_X1 port map( A => n3831, Z => n3790);
   U3709 : BUF_X1 port map( A => n3829, Z => n3796);
   U3710 : BUF_X1 port map( A => n3822, Z => n3815);
   U3711 : BUF_X1 port map( A => n3833, Z => n3784);
   U3712 : BUF_X1 port map( A => n3838, Z => n3769);
   U3713 : BUF_X1 port map( A => n3824, Z => n3809);
   U3714 : BUF_X1 port map( A => n3836, Z => n3775);
   U3715 : BUF_X1 port map( A => n3835, Z => n3778);
   U3716 : BUF_X1 port map( A => n3836, Z => n3773);
   U3717 : BUF_X1 port map( A => n3830, Z => n3791);
   U3718 : BUF_X1 port map( A => n3828, Z => n3798);
   U3719 : BUF_X1 port map( A => n3832, Z => n3786);
   U3720 : BUF_X1 port map( A => n3837, Z => n3771);
   U3721 : BUF_X1 port map( A => n3837, Z => n3770);
   U3722 : BUF_X1 port map( A => n3823, Z => n3813);
   U3723 : BUF_X1 port map( A => n3825, Z => n3807);
   U3724 : BUF_X1 port map( A => n3827, Z => n3800);
   U3725 : BUF_X1 port map( A => n3829, Z => n3794);
   U3726 : BUF_X1 port map( A => n3831, Z => n3788);
   U3727 : BUF_X1 port map( A => n3833, Z => n3782);
   U3728 : BUF_X1 port map( A => n3835, Z => n3776);
   U3729 : BUF_X1 port map( A => n3824, Z => n3810);
   U3730 : BUF_X1 port map( A => n3826, Z => n3803);
   U3731 : BUF_X1 port map( A => n3828, Z => n3797);
   U3732 : BUF_X1 port map( A => n3838, Z => n3767);
   U3733 : BUF_X1 port map( A => n3826, Z => n3804);
   U3734 : BUF_X1 port map( A => n3832, Z => n3785);
   U3735 : BUF_X1 port map( A => n3834, Z => n3779);
   U3736 : BUF_X1 port map( A => n3836, Z => n3774);
   U3737 : BUF_X1 port map( A => n3628, Z => n3626);
   U3738 : BUF_X1 port map( A => n3629, Z => n3622);
   U3739 : BUF_X1 port map( A => n3629, Z => n3623);
   U3740 : BUF_X1 port map( A => n3629, Z => n3624);
   U3741 : BUF_X1 port map( A => n3628, Z => n3625);
   U3742 : BUF_X1 port map( A => n3630, Z => n3621);
   U3743 : BUF_X1 port map( A => n3628, Z => n3627);
   U3744 : INV_X1 port map( A => n4221, ZN => n4266);
   U3745 : INV_X1 port map( A => n4220, ZN => n4259);
   U3746 : INV_X1 port map( A => n4220, ZN => n4258);
   U3747 : INV_X1 port map( A => n4220, ZN => n4264);
   U3748 : INV_X1 port map( A => n4220, ZN => n4263);
   U3749 : INV_X1 port map( A => n4220, ZN => n4261);
   U3750 : INV_X1 port map( A => n4220, ZN => n4262);
   U3751 : INV_X1 port map( A => n4218, ZN => n4260);
   U3752 : INV_X1 port map( A => n4219, ZN => n4265);
   U3753 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n22, Z => n3012);
   U3754 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n24, Z => n3018);
   U3755 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n26, Z => n3024);
   U3756 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n28, Z => n3030);
   U3757 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n10, Z => n2988);
   U3758 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n12, Z => n2994);
   U3759 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n14, Z => n3000);
   U3760 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n16, Z => n3006);
   U3761 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n22, Z => n3013);
   U3762 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n24, Z => n3019);
   U3763 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n26, Z => n3025);
   U3764 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n28, Z => n3031);
   U3765 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n10, Z => n2989);
   U3766 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n12, Z => n2995);
   U3767 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n14, Z => n3001);
   U3768 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n16, Z => n3007);
   U3769 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n23, Z => n3015);
   U3770 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n25, Z => n3021);
   U3771 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n27, Z => n3027);
   U3772 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n29, Z => n3033);
   U3773 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n11, Z => n2991);
   U3774 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n13, Z => n2997);
   U3775 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n15, Z => n3003);
   U3776 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n17, Z => n3009);
   U3777 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n23, Z => n3016);
   U3778 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n25, Z => n3022);
   U3779 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n27, Z => n3028);
   U3780 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n29, Z => n3034);
   U3781 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n11, Z => n2992);
   U3782 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n13, Z => n2998);
   U3783 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n15, Z => n3004);
   U3784 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n17, Z => n3010);
   U3785 : BUF_X1 port map( A => DataPath_WRF_CUhw_n112, Z => n3258);
   U3786 : BUF_X1 port map( A => DataPath_WRF_CUhw_n112, Z => n3257);
   U3787 : BUF_X1 port map( A => DataPath_WRF_CUhw_n112, Z => n3256);
   U3788 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n22, Z => n3014);
   U3789 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n24, Z => n3020);
   U3790 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n26, Z => n3026);
   U3791 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n28, Z => n3032);
   U3792 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n10, Z => n2990);
   U3793 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n12, Z => n2996);
   U3794 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n14, Z => n3002);
   U3795 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n16, Z => n3008);
   U3796 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n23, Z => n3017);
   U3797 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n25, Z => n3023);
   U3798 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n27, Z => n3029);
   U3799 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n29, Z => n3035);
   U3800 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n11, Z => n2993);
   U3801 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n13, Z => n2999);
   U3802 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n15, Z => n3005);
   U3803 : BUF_X1 port map( A => DataPath_RF_RDPORT_SPILL_n17, Z => n3011);
   U3804 : XNOR2_X1 port map( A => n6904, B => n1798, ZN => n6761);
   U3805 : XNOR2_X1 port map( A => n6947, B => n6921, ZN => n1798);
   U3806 : INV_X1 port map( A => n2263, ZN => n2261);
   U3808 : XNOR2_X1 port map( A => n5436, B => n5437, ZN => n5445);
   U3809 : XNOR2_X1 port map( A => n5052, B => n5053, ZN => n5058);
   U3810 : XNOR2_X1 port map( A => n4757, B => n4756, ZN => n4762);
   U3811 : XNOR2_X1 port map( A => n5365, B => n5364, ZN => n5366);
   U3812 : XNOR2_X1 port map( A => n725, B => n1799, ZN => n6963);
   U3813 : XNOR2_X1 port map( A => n7404, B => n7391, ZN => n1799);
   U3814 : INV_X1 port map( A => n1873, ZN => n2188);
   U3815 : XNOR2_X1 port map( A => n968, B => n5795, ZN => n5557);
   U3816 : XNOR2_X1 port map( A => n7577, B => n7576, ZN => n1800);
   U3817 : XNOR2_X1 port map( A => n4849, B => n4850, ZN => n1801);
   U3818 : XNOR2_X1 port map( A => n5461, B => n5459, ZN => n5463);
   U3819 : OAI21_X1 port map( B1 => n1550, B2 => n1870, A => n4641, ZN => n8188
                           );
   U3820 : XNOR2_X1 port map( A => n6850, B => n6849, ZN => n1804);
   U3821 : XNOR2_X1 port map( A => n6852, B => n6851, ZN => n1805);
   U3822 : XNOR2_X1 port map( A => n1173, B => n6198, ZN => n1806);
   U3823 : XNOR2_X1 port map( A => n5394, B => n5390, ZN => n5395);
   U3824 : XNOR2_X1 port map( A => n454, B => n7305, ZN => n7306);
   U3826 : XNOR2_X1 port map( A => n7276, B => n589, ZN => n7278);
   U3827 : XNOR2_X1 port map( A => n5724, B => n5725, ZN => n5726);
   U3828 : BUF_X2 port map( A => n2151, Z => n2145);
   U3829 : CLKBUF_X1 port map( A => n2150, Z => n2144);
   U3830 : AND2_X1 port map( A1 => n5652, A2 => n5658, ZN => n1807);
   U3831 : XNOR2_X1 port map( A => n5570, B => n5569, ZN => n1809);
   U3832 : OAI21_X1 port map( B1 => n17230, B2 => n1825, A => n4889, ZN => 
                           n4890);
   U3833 : INV_X1 port map( A => n17195, ZN => n2146);
   U3834 : NOR2_X1 port map( A1 => n1292, A2 => n7507, ZN => n7510);
   U3835 : AND2_X1 port map( A1 => n6251, A2 => n6079, ZN => n1810);
   U3836 : AND2_X1 port map( A1 => n6811, A2 => n6809, ZN => n1811);
   U3837 : AND2_X1 port map( A1 => n5859, A2 => n5805, ZN => n1812);
   U3838 : XNOR2_X1 port map( A => n17151, B => n5101, ZN => n5104);
   U3839 : XNOR2_X1 port map( A => n4946, B => n1817, ZN => n1813);
   U3840 : AND2_X1 port map( A1 => n440, A2 => n6793, ZN => n1814);
   U3841 : AND2_X1 port map( A1 => n6805, A2 => n6802, ZN => n1815);
   U3842 : AND2_X1 port map( A1 => n5859, A2 => n5860, ZN => n1816);
   U3843 : XNOR2_X1 port map( A => n4841, B => n4842, ZN => n1817);
   U3844 : XNOR2_X1 port map( A => n17209, B => n7641, ZN => n1818);
   U3845 : XNOR2_X1 port map( A => n629, B => n7705, ZN => n1819);
   U3846 : XNOR2_X1 port map( A => n1822, B => n5431, ZN => n1820);
   U3847 : XNOR2_X1 port map( A => n833, B => n5186, ZN => n1821);
   U3848 : XNOR2_X1 port map( A => n5649, B => n558, ZN => n5650);
   U3849 : NAND2_X1 port map( A1 => n5157, A2 => n5156, ZN => n5158);
   U3850 : AND2_X1 port map( A1 => n4642, A2 => n8187, ZN => n1825);
   U3851 : XNOR2_X1 port map( A => n5370, B => n5366, ZN => n5371);
   U3852 : XNOR2_X1 port map( A => n5175, B => n5169, ZN => n5176);
   U3853 : INV_X1 port map( A => n6024, ZN => n6251);
   U3854 : AND2_X1 port map( A1 => n1655, A2 => n7022, ZN => n1828);
   U3855 : AND2_X1 port map( A1 => n6977, A2 => n6978, ZN => n1831);
   U3856 : AND2_X1 port map( A1 => n6984, A2 => n1415, ZN => n1832);
   U3857 : AND2_X1 port map( A1 => n4549, A2 => n4548, ZN => n1833);
   U3858 : AND2_X1 port map( A1 => n698, A2 => n5919, ZN => n1834);
   U3859 : AND2_X1 port map( A1 => n5294, A2 => n5364, ZN => n1835);
   U3860 : AND2_X1 port map( A1 => n1370, A2 => n5292, ZN => n1836);
   U3861 : AND2_X1 port map( A1 => n5297, A2 => n5296, ZN => n1837);
   U3862 : AND2_X1 port map( A1 => n4841, A2 => n4842, ZN => n1839);
   U3863 : AND2_X1 port map( A1 => n975, A2 => n5549, ZN => n1840);
   U3864 : AND2_X1 port map( A1 => n6944, A2 => n981, ZN => n1841);
   U3865 : AND2_X1 port map( A1 => n5787, A2 => n5790, ZN => n1842);
   U3866 : AND2_X1 port map( A1 => n6694, A2 => n6696, ZN => n1844);
   U3867 : AND2_X1 port map( A1 => n5572, A2 => n5569, ZN => n1845);
   U3868 : AND2_X1 port map( A1 => n6695, A2 => n1323, ZN => n1846);
   U3869 : AND2_X1 port map( A1 => n6524, A2 => n6484, ZN => n1847);
   U3870 : AND2_X1 port map( A1 => n1134, A2 => n6012, ZN => n1848);
   U3871 : AND2_X1 port map( A1 => n6524, A2 => n6523, ZN => n1849);
   U3872 : NAND2_X1 port map( A1 => n483, A2 => n8198, ZN => n4893);
   U3873 : NAND2_X1 port map( A1 => n7546, A2 => n7547, ZN => n7509);
   U3874 : AND2_X1 port map( A1 => n4640, A2 => n4875, ZN => n1851);
   U3875 : INV_X1 port map( A => n2172, ZN => n6473);
   U3876 : XNOR2_X1 port map( A => n913, B => n7828, ZN => n1853);
   U3877 : XNOR2_X1 port map( A => n7764, B => n1391, ZN => n1854);
   U3878 : INV_X1 port map( A => n2267, ZN => n2168);
   U3879 : INV_X1 port map( A => n3902, ZN => n3900);
   U3880 : NOR2_X1 port map( A1 => n4156, A2 => n3900, ZN => 
                           DataPath_WRF_CUhw_N26_port);
   U3881 : BUF_X1 port map( A => n7989, Z => n2273);
   U3882 : OR2_X1 port map( A1 => n3901, A2 => n4155, ZN => n1855);
   U3883 : XNOR2_X1 port map( A => n765, B => n7964, ZN => n1856);
   U3884 : XNOR2_X1 port map( A => n17166, B => n7895, ZN => n1857);
   U3885 : AND2_X1 port map( A1 => n5845, A2 => n2268, ZN => n1858);
   U3886 : XNOR2_X1 port map( A => n8132, B => n1217, ZN => n8134);
   U3887 : INV_X1 port map( A => n8031, ZN => n8307);
   U3888 : INV_X1 port map( A => n8032, ZN => n8312);
   U3889 : NAND2_X1 port map( A1 => n7747, A2 => n1861, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n181);
   U3890 : INV_X1 port map( A => n4127, ZN => n4118);
   U3891 : NAND2_X1 port map( A1 => n7747, A2 => n7746, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n182);
   U3892 : AOI21_X1 port map( B1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_12_port, B2
                           => n11511, A => n11518, ZN => n12928);
   U3893 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, A => 
                           DataPath_ALUhw_SHIFTER_HW_n173, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n167);
   U3894 : OAI22_X1 port map( A1 => n8287, A2 => n1769, B1 => n8291, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n173);
   U3895 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n445, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n432, A => 
                           DataPath_ALUhw_SHIFTER_HW_n513, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n512);
   U3896 : OAI22_X1 port map( A1 => n8288, A2 => n2984, B1 => n8286, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n513);
   U3897 : AOI221_X1 port map( B1 => n8305, B2 => n521, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n432, A => 
                           DataPath_ALUhw_SHIFTER_HW_n495, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n484);
   U3898 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n405, ZN => n8296);
   U3899 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n432, ZN => n8295);
   U3900 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n405, A => 
                           DataPath_ALUhw_SHIFTER_HW_n482, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n469);
   U3901 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, C1 => n8309, C2 => 
                           n523, A => DataPath_ALUhw_SHIFTER_HW_n217, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n214);
   U3902 : OAI22_X1 port map( A1 => n8284, A2 => n1769, B1 => n8283, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n217);
   U3903 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n392, ZN => n8297);
   U3904 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n211, C1 => n8315, C2 => 
                           n523, A => DataPath_ALUhw_SHIFTER_HW_n268, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n263);
   U3905 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n219, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, A => 
                           DataPath_ALUhw_SHIFTER_HW_n418, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n407);
   U3906 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n269, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n201, A => 
                           DataPath_ALUhw_SHIFTER_HW_n606, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n583);
   U3907 : OAI22_X1 port map( A1 => n8295, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8296, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n481);
   U3908 : OAI22_X1 port map( A1 => n8294, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8295, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n494);
   U3909 : AOI221_X1 port map( B1 => n8311, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, C1 => n8310, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, A => 
                           DataPath_ALUhw_SHIFTER_HW_n507, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n498);
   U3910 : OAI22_X1 port map( A1 => n8293, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8294, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n507);
   U3911 : AOI221_X1 port map( B1 => n8311, B2 => n523, C1 => n8310, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, A => 
                           DataPath_ALUhw_SHIFTER_HW_n190, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n187);
   U3912 : OAI22_X1 port map( A1 => n8287, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8288, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n190);
   U3913 : AOI221_X1 port map( B1 => n8311, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, C1 => n8310, C2 => 
                           n523, A => DataPath_ALUhw_SHIFTER_HW_n199, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n196);
   U3914 : OAI22_X1 port map( A1 => n8291, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8287, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n199);
   U3915 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n380, ZN => n8298);
   U3916 : AOI221_X1 port map( B1 => n8300, B2 => n521, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, A => 
                           DataPath_ALUhw_SHIFTER_HW_n539, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n538);
   U3917 : OAI22_X1 port map( A1 => n8291, A2 => n2984, B1 => n8287, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n539);
   U3918 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, A => 
                           DataPath_ALUhw_SHIFTER_HW_n153, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n144);
   U3919 : OAI22_X1 port map( A1 => n8288, A2 => n1769, B1 => n8287, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n153);
   U3920 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n392, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n405, A => 
                           DataPath_ALUhw_SHIFTER_HW_n466, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n458);
   U3921 : OAI22_X1 port map( A1 => n8294, A2 => n1769, B1 => n8293, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n466);
   U3922 : OAI22_X1 port map( A1 => n8308, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8317, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n260);
   U3923 : OAI22_X1 port map( A1 => n8313, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8318, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n296);
   U3924 : OAI22_X1 port map( A1 => n8319, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8313, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n310);
   U3925 : OAI22_X1 port map( A1 => n8320, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8319, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n324);
   U3926 : OAI22_X1 port map( A1 => n11491, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n191, B1 => n8320, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n192, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n338);
   U3927 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n445, A => 
                           DataPath_ALUhw_SHIFTER_HW_n526, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n525);
   U3928 : OAI22_X1 port map( A1 => n8287, A2 => n2984, B1 => n8288, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n526);
   U3929 : OAI22_X1 port map( A1 => n8286, A2 => n1769, B1 => n8288, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n551);
   U3930 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, A => 
                           DataPath_ALUhw_SHIFTER_HW_n183, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n177);
   U3931 : OAI22_X1 port map( A1 => n8291, A2 => n1769, B1 => n8292, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n183);
   U3932 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, A => 
                           DataPath_ALUhw_SHIFTER_HW_n207, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n204);
   U3933 : OAI22_X1 port map( A1 => n8285, A2 => n1769, B1 => n8284, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n207);
   U3934 : OAI22_X1 port map( A1 => n8295, A2 => n1769, B1 => n8294, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n453);
   U3935 : OAI22_X1 port map( A1 => n11495, A2 => n2984, B1 => n11494, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n266);
   U3936 : OAI22_X1 port map( A1 => n8282, A2 => n1769, B1 => n11494, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n417);
   U3937 : OAI22_X1 port map( A1 => n11494, A2 => n1769, B1 => n11495, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n603);
   U3938 : NOR2_X1 port map( A1 => n2509, A2 => n4180, ZN => n14362);
   U3939 : NOR2_X1 port map( A1 => n2515, A2 => n4179, ZN => n14396);
   U3940 : NOR2_X1 port map( A1 => n2521, A2 => n4179, ZN => n14430);
   U3941 : NOR2_X1 port map( A1 => n2527, A2 => n4178, ZN => n14464);
   U3942 : NOR2_X1 port map( A1 => n2533, A2 => n4178, ZN => n14498);
   U3943 : NOR2_X1 port map( A1 => n2539, A2 => n4177, ZN => n14532);
   U3944 : NOR2_X1 port map( A1 => n2545, A2 => n4177, ZN => n14566);
   U3945 : NOR2_X1 port map( A1 => n2551, A2 => n4176, ZN => n14600);
   U3946 : NOR2_X1 port map( A1 => n2557, A2 => n4176, ZN => n14634);
   U3947 : NOR2_X1 port map( A1 => n2563, A2 => n4175, ZN => n14668);
   U3948 : NOR2_X1 port map( A1 => n2569, A2 => n4175, ZN => n14702);
   U3949 : NOR2_X1 port map( A1 => n2575, A2 => n4174, ZN => n14736);
   U3950 : NOR2_X1 port map( A1 => n2581, A2 => n4174, ZN => n14770);
   U3951 : NOR2_X1 port map( A1 => n2587, A2 => n4173, ZN => n14804);
   U3952 : NOR2_X1 port map( A1 => n2593, A2 => n4173, ZN => n14838);
   U3953 : NOR2_X1 port map( A1 => n2599, A2 => n4172, ZN => n14872);
   U3954 : NOR2_X1 port map( A1 => n2605, A2 => n4171, ZN => n14906);
   U3955 : NOR2_X1 port map( A1 => n2611, A2 => n4171, ZN => n14940);
   U3956 : NOR2_X1 port map( A1 => n2617, A2 => n4170, ZN => n14974);
   U3957 : NOR2_X1 port map( A1 => n2623, A2 => n4170, ZN => n15008);
   U3958 : NOR2_X1 port map( A1 => n2629, A2 => n4169, ZN => n15042);
   U3959 : NOR2_X1 port map( A1 => n2635, A2 => n4169, ZN => n15076);
   U3960 : NOR2_X1 port map( A1 => n2641, A2 => n4168, ZN => n15110);
   U3961 : NOR2_X1 port map( A1 => n2647, A2 => n4168, ZN => n15144);
   U3962 : NOR2_X1 port map( A1 => n2653, A2 => n4167, ZN => n15178);
   U3963 : NOR2_X1 port map( A1 => n2659, A2 => n4167, ZN => n15212);
   U3964 : NOR2_X1 port map( A1 => n2665, A2 => n4166, ZN => n15246);
   U3965 : NOR2_X1 port map( A1 => n2671, A2 => n4166, ZN => n15280);
   U3966 : NOR2_X1 port map( A1 => n2677, A2 => n4165, ZN => n15314);
   U3967 : NOR2_X1 port map( A1 => n2683, A2 => n4165, ZN => n15348);
   U3968 : NOR2_X1 port map( A1 => n2689, A2 => n4164, ZN => n15382);
   U3969 : NOR2_X1 port map( A1 => n2695, A2 => n4164, ZN => n15416);
   U3970 : NOR2_X1 port map( A1 => n2701, A2 => n4163, ZN => n15450);
   U3971 : NOR2_X1 port map( A1 => n2707, A2 => n4163, ZN => n15484);
   U3972 : NOR2_X1 port map( A1 => n2713, A2 => n4162, ZN => n15518);
   U3973 : NOR2_X1 port map( A1 => n2719, A2 => n4162, ZN => n15552);
   U3974 : NOR2_X1 port map( A1 => n2725, A2 => n4161, ZN => n15586);
   U3975 : NOR2_X1 port map( A1 => n2731, A2 => n4161, ZN => n15620);
   U3976 : NOR2_X1 port map( A1 => n2737, A2 => n4160, ZN => n15654);
   U3977 : NOR2_X1 port map( A1 => n2743, A2 => n4160, ZN => n15688);
   U3978 : NOR2_X1 port map( A1 => n2749, A2 => n4159, ZN => n15722);
   U3979 : NOR2_X1 port map( A1 => n2755, A2 => n4159, ZN => n15756);
   U3980 : NOR2_X1 port map( A1 => n2761, A2 => n4158, ZN => n15790);
   U3981 : NOR2_X1 port map( A1 => n2767, A2 => n4158, ZN => n15824);
   U3982 : NOR2_X1 port map( A1 => n2773, A2 => n4157, ZN => n15858);
   U3983 : NOR2_X1 port map( A1 => n2779, A2 => n4202, ZN => n15892);
   U3984 : NOR2_X1 port map( A1 => n2785, A2 => n4201, ZN => n15926);
   U3985 : NOR2_X1 port map( A1 => n2791, A2 => n4201, ZN => n15960);
   U3986 : NOR2_X1 port map( A1 => n2797, A2 => n4200, ZN => n15994);
   U3987 : NOR2_X1 port map( A1 => n2803, A2 => n4200, ZN => n16028);
   U3988 : NOR2_X1 port map( A1 => n2809, A2 => n4199, ZN => n16062);
   U3989 : NOR2_X1 port map( A1 => n2815, A2 => n4199, ZN => n16096);
   U3990 : NOR2_X1 port map( A1 => n2821, A2 => n4198, ZN => n16130);
   U3991 : NOR2_X1 port map( A1 => n2827, A2 => n4198, ZN => n16164);
   U3992 : NOR2_X1 port map( A1 => n2833, A2 => n4197, ZN => n16198);
   U3993 : NOR2_X1 port map( A1 => n2839, A2 => n4197, ZN => n16232);
   U3994 : NOR2_X1 port map( A1 => n2845, A2 => n4196, ZN => n16266);
   U3995 : NOR2_X1 port map( A1 => n2851, A2 => n4196, ZN => n16300);
   U3996 : NOR2_X1 port map( A1 => n2857, A2 => n4195, ZN => n16334);
   U3997 : NOR2_X1 port map( A1 => n2863, A2 => n4195, ZN => n16368);
   U3998 : NOR2_X1 port map( A1 => n2869, A2 => n4194, ZN => n16402);
   U3999 : NOR2_X1 port map( A1 => n2875, A2 => n4194, ZN => n16436);
   U4000 : NOR2_X1 port map( A1 => n2881, A2 => n4193, ZN => n16470);
   U4001 : NOR2_X1 port map( A1 => n2887, A2 => n4192, ZN => n16504);
   U4002 : NOR2_X1 port map( A1 => n2893, A2 => n4192, ZN => n16538);
   U4003 : NOR2_X1 port map( A1 => n2899, A2 => n4191, ZN => n16572);
   U4004 : NOR2_X1 port map( A1 => n2905, A2 => n4191, ZN => n16606);
   U4005 : NOR2_X1 port map( A1 => n2911, A2 => n4190, ZN => n16640);
   U4006 : NOR2_X1 port map( A1 => n2917, A2 => n4190, ZN => n16674);
   U4007 : NOR2_X1 port map( A1 => n2923, A2 => n4189, ZN => n16708);
   U4008 : NOR2_X1 port map( A1 => n2929, A2 => n4189, ZN => n16742);
   U4009 : NOR2_X1 port map( A1 => n2935, A2 => n4188, ZN => n16776);
   U4010 : NOR2_X1 port map( A1 => n2941, A2 => n4188, ZN => n16810);
   U4011 : NOR2_X1 port map( A1 => n2947, A2 => n4187, ZN => n16844);
   U4012 : NOR2_X1 port map( A1 => n2953, A2 => n4187, ZN => n16878);
   U4013 : NOR2_X1 port map( A1 => n2959, A2 => n4186, ZN => n16912);
   U4014 : NOR2_X1 port map( A1 => n2965, A2 => n4186, ZN => n16946);
   U4015 : NOR2_X1 port map( A1 => n2971, A2 => n4185, ZN => n16980);
   U4016 : NOR2_X1 port map( A1 => n2977, A2 => n4185, ZN => n17014);
   U4017 : NOR2_X1 port map( A1 => n2983, A2 => n4184, ZN => n17048);
   U4018 : AOI21_X1 port map( B1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_3_16_port, B2
                           => n11511, A => n11517, ZN => n12929);
   U4019 : AND2_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_16_port, A2
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_12_port,
                           ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_3_16_port);
   U4020 : INV_X1 port map( A => n12923, ZN => n11517);
   U4021 : AOI21_X1 port map( B1 => n11518, B2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_16_port, A 
                           => n11520, ZN => n12923);
   U4022 : INV_X1 port map( A => n4117, ZN => n4108);
   U4023 : BUF_X1 port map( A => n7989, Z => n2274);
   U4024 : OAI22_X1 port map( A1 => n8298, A2 => n2984, B1 => n8301, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n360);
   U4025 : OAI22_X1 port map( A1 => n8298, A2 => n1769, B1 => n8297, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n403);
   U4026 : OAI22_X1 port map( A1 => n8319, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8320, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n345);
   U4027 : OAI22_X1 port map( A1 => n8297, A2 => n2984, B1 => n8298, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n150, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n373);
   U4028 : OAI22_X1 port map( A1 => n8303, A2 => n1769, B1 => n8302, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n367);
   U4029 : OAI22_X1 port map( A1 => n11493, A2 => n1769, B1 => n8303, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n155, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n354);
   U4030 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_2_port
                           , A2 => n11511, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_2_port
                           , B2 => n12927, ZN => n12896);
   U4031 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_1_port
                           , A2 => n11511, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_1_port
                           , B2 => n12927, ZN => n12897);
   U4032 : AOI22_X1 port map( A1 => n2429, A2 => n3299, B1 => n4006, B2 => 
                           n3322, ZN => n13132);
   U4033 : AOI22_X1 port map( A1 => n2351, A2 => n3413, B1 => n3934, B2 => 
                           n3462, ZN => n13247);
   U4034 : AOI22_X1 port map( A1 => n2429, A2 => n3410, B1 => n4006, B2 => 
                           n3434, ZN => n13356);
   U4035 : AOI22_X1 port map( A1 => n2436, A2 => n3413, B1 => n4013, B2 => 
                           n3441, ZN => n13389);
   U4036 : AOI22_X1 port map( A1 => n2441, A2 => n3408, B1 => n4018, B2 => 
                           n3433, ZN => n13358);
   U4037 : AOI22_X1 port map( A1 => n2447, A2 => n3411, B1 => n4024, B2 => 
                           n3436, ZN => n13359);
   U4038 : AOI22_X1 port map( A1 => n2453, A2 => n3410, B1 => n4030, B2 => 
                           n3433, ZN => n13360);
   U4039 : AOI22_X1 port map( A1 => n2459, A2 => n3414, B1 => n4036, B2 => 
                           n3433, ZN => n13361);
   U4040 : AOI22_X1 port map( A1 => n2465, A2 => n3407, B1 => n4042, B2 => 
                           n3437, ZN => n13362);
   U4041 : AOI22_X1 port map( A1 => n2471, A2 => n3409, B1 => n4102, B2 => 
                           n3438, ZN => n13363);
   U4042 : AOI22_X1 port map( A1 => n2352, A2 => n3525, B1 => n3935, B2 => 
                           n3574, ZN => n13503);
   U4043 : AOI22_X1 port map( A1 => n2430, A2 => n3522, B1 => n4007, B2 => 
                           n3546, ZN => n13612);
   U4044 : AOI22_X1 port map( A1 => n2436, A2 => n3525, B1 => n4013, B2 => 
                           n3553, ZN => n13645);
   U4045 : AOI22_X1 port map( A1 => n2442, A2 => n3519, B1 => n4019, B2 => 
                           n3545, ZN => n13614);
   U4046 : AOI22_X1 port map( A1 => n2448, A2 => n3523, B1 => n4025, B2 => 
                           n3548, ZN => n13615);
   U4047 : AOI22_X1 port map( A1 => n2454, A2 => n3522, B1 => n4031, B2 => 
                           n3545, ZN => n13616);
   U4048 : AOI22_X1 port map( A1 => n2460, A2 => n3526, B1 => n4037, B2 => 
                           n3545, ZN => n13617);
   U4049 : AOI22_X1 port map( A1 => n2466, A2 => n3520, B1 => n4043, B2 => 
                           n3549, ZN => n13618);
   U4050 : AOI22_X1 port map( A1 => n2472, A2 => n3521, B1 => n4103, B2 => 
                           n3550, ZN => n13619);
   U4051 : AOI22_X1 port map( A1 => n2353, A2 => n3634, B1 => n3936, B2 => 
                           n3686, ZN => n13759);
   U4052 : AOI22_X1 port map( A1 => n2431, A2 => n3633, B1 => n4008, B2 => 
                           n3658, ZN => n13868);
   U4053 : AOI22_X1 port map( A1 => n2437, A2 => n3637, B1 => n4014, B2 => 
                           n3665, ZN => n13901);
   U4054 : AOI22_X1 port map( A1 => n2443, A2 => n3634, B1 => n4020, B2 => 
                           n3657, ZN => n13870);
   U4055 : AOI22_X1 port map( A1 => n2449, A2 => n3635, B1 => n4026, B2 => 
                           n3660, ZN => n13871);
   U4056 : AOI22_X1 port map( A1 => n2455, A2 => n3633, B1 => n4032, B2 => 
                           n3657, ZN => n13872);
   U4057 : AOI22_X1 port map( A1 => n2461, A2 => n3638, B1 => n4038, B2 => 
                           n3657, ZN => n13873);
   U4058 : AOI22_X1 port map( A1 => n2467, A2 => n3634, B1 => n4044, B2 => 
                           n3661, ZN => n13874);
   U4059 : AOI22_X1 port map( A1 => n2473, A2 => n3632, B1 => n4104, B2 => 
                           n3662, ZN => n13875);
   U4060 : AOI22_X1 port map( A1 => n2353, A2 => n3744, B1 => n3936, B2 => 
                           n3798, ZN => n14015);
   U4061 : AOI22_X1 port map( A1 => n2431, A2 => n3746, B1 => n4008, B2 => 
                           n3770, ZN => n14124);
   U4062 : AOI22_X1 port map( A1 => n2438, A2 => n3748, B1 => n4015, B2 => 
                           n3777, ZN => n14157);
   U4063 : AOI22_X1 port map( A1 => n2443, A2 => n3747, B1 => n4020, B2 => 
                           n3769, ZN => n14126);
   U4064 : AOI22_X1 port map( A1 => n2449, A2 => n3747, B1 => n4026, B2 => 
                           n3772, ZN => n14127);
   U4065 : AOI22_X1 port map( A1 => n2455, A2 => n3747, B1 => n4032, B2 => 
                           n3769, ZN => n14128);
   U4066 : AOI22_X1 port map( A1 => n2461, A2 => n3747, B1 => n4038, B2 => 
                           n3769, ZN => n14129);
   U4067 : AOI22_X1 port map( A1 => n2467, A2 => n3747, B1 => n4044, B2 => 
                           n3773, ZN => n14130);
   U4068 : AOI22_X1 port map( A1 => n2473, A2 => n3747, B1 => n4104, B2 => 
                           n3774, ZN => n14131);
   U4069 : AOI22_X1 port map( A1 => n2435, A2 => n3295, B1 => n4012, B2 => 
                           n3320, ZN => n13133);
   U4070 : AOI22_X1 port map( A1 => n2441, A2 => n3301, B1 => n4018, B2 => 
                           n3321, ZN => n13134);
   U4071 : AOI22_X1 port map( A1 => n2447, A2 => n3300, B1 => n4024, B2 => 
                           n3324, ZN => n13135);
   U4072 : AOI22_X1 port map( A1 => n2453, A2 => n3295, B1 => n4030, B2 => 
                           n3321, ZN => n13136);
   U4073 : AOI22_X1 port map( A1 => n2459, A2 => n3305, B1 => n4036, B2 => 
                           n3321, ZN => n13137);
   U4074 : AOI22_X1 port map( A1 => n2465, A2 => n3303, B1 => n4042, B2 => 
                           n3325, ZN => n13138);
   U4075 : AOI22_X1 port map( A1 => n2327, A2 => n3303, B1 => n3916, B2 => 
                           n3320, ZN => n13115);
   U4076 : AOI22_X1 port map( A1 => n2333, A2 => n3304, B1 => n3922, B2 => 
                           n3318, ZN => n13116);
   U4077 : AOI22_X1 port map( A1 => n2345, A2 => n3295, B1 => n3928, B2 => 
                           n3318, ZN => n13118);
   U4078 : AOI22_X1 port map( A1 => n2351, A2 => n3304, B1 => n3934, B2 => 
                           n3318, ZN => n13119);
   U4079 : AOI22_X1 port map( A1 => n2357, A2 => n3305, B1 => n3940, B2 => 
                           n3322, ZN => n13120);
   U4080 : AOI22_X1 port map( A1 => n2363, A2 => n3302, B1 => n3946, B2 => 
                           n3318, ZN => n13121);
   U4081 : AOI22_X1 port map( A1 => n2369, A2 => n3301, B1 => n3952, B2 => 
                           n3324, ZN => n13122);
   U4082 : AOI22_X1 port map( A1 => n2375, A2 => n3303, B1 => n3958, B2 => 
                           n3323, ZN => n13123);
   U4083 : AOI22_X1 port map( A1 => n2381, A2 => n3299, B1 => n3964, B2 => 
                           n3324, ZN => n13124);
   U4084 : AOI22_X1 port map( A1 => n2387, A2 => n3297, B1 => n3970, B2 => 
                           n3319, ZN => n13125);
   U4085 : AOI22_X1 port map( A1 => n2393, A2 => n3298, B1 => n3976, B2 => 
                           n3323, ZN => n13126);
   U4086 : AOI22_X1 port map( A1 => n2399, A2 => n3296, B1 => n3982, B2 => 
                           n3319, ZN => n13127);
   U4087 : AOI22_X1 port map( A1 => n2411, A2 => n3299, B1 => n3988, B2 => 
                           n3321, ZN => n13129);
   U4088 : AOI22_X1 port map( A1 => n2417, A2 => n3300, B1 => n3994, B2 => 
                           n3320, ZN => n13130);
   U4089 : AOI22_X1 port map( A1 => n2423, A2 => n3302, B1 => n4000, B2 => 
                           n3320, ZN => n13131);
   U4090 : AOI22_X1 port map( A1 => n2339, A2 => n3303, B1 => n4090, B2 => 
                           n3322, ZN => n13117);
   U4091 : AOI22_X1 port map( A1 => n2405, A2 => n3301, B1 => n4096, B2 => 
                           n3319, ZN => n13128);
   U4092 : AOI22_X1 port map( A1 => n2471, A2 => n3295, B1 => n4102, B2 => 
                           n3319, ZN => n13107);
   U4093 : AOI22_X1 port map( A1 => n2327, A2 => n3408, B1 => n3916, B2 => 
                           n3432, ZN => n13339);
   U4094 : AOI22_X1 port map( A1 => n2333, A2 => n3408, B1 => n3922, B2 => 
                           n3430, ZN => n13340);
   U4095 : AOI22_X1 port map( A1 => n2345, A2 => n3408, B1 => n3928, B2 => 
                           n3430, ZN => n13342);
   U4096 : AOI22_X1 port map( A1 => n2357, A2 => n3408, B1 => n3940, B2 => 
                           n3434, ZN => n13344);
   U4097 : AOI22_X1 port map( A1 => n2363, A2 => n3407, B1 => n3946, B2 => 
                           n3430, ZN => n13345);
   U4098 : AOI22_X1 port map( A1 => n2369, A2 => n3407, B1 => n3952, B2 => 
                           n3436, ZN => n13346);
   U4099 : AOI22_X1 port map( A1 => n2375, A2 => n3407, B1 => n3958, B2 => 
                           n3435, ZN => n13347);
   U4100 : AOI22_X1 port map( A1 => n2381, A2 => n3407, B1 => n3964, B2 => 
                           n3436, ZN => n13348);
   U4101 : AOI22_X1 port map( A1 => n2387, A2 => n3407, B1 => n3970, B2 => 
                           n3431, ZN => n13349);
   U4102 : AOI22_X1 port map( A1 => n2393, A2 => n3407, B1 => n3976, B2 => 
                           n3435, ZN => n13350);
   U4103 : AOI22_X1 port map( A1 => n2399, A2 => n3407, B1 => n3982, B2 => 
                           n3431, ZN => n13351);
   U4104 : AOI22_X1 port map( A1 => n2411, A2 => n3407, B1 => n3988, B2 => 
                           n3433, ZN => n13353);
   U4105 : AOI22_X1 port map( A1 => n2417, A2 => n3407, B1 => n3994, B2 => 
                           n3432, ZN => n13354);
   U4106 : AOI22_X1 port map( A1 => n2423, A2 => n3407, B1 => n4000, B2 => 
                           n3432, ZN => n13355);
   U4107 : AOI22_X1 port map( A1 => n2339, A2 => n3408, B1 => n4090, B2 => 
                           n3434, ZN => n13341);
   U4108 : AOI22_X1 port map( A1 => n2405, A2 => n3407, B1 => n4096, B2 => 
                           n3431, ZN => n13352);
   U4109 : AOI22_X1 port map( A1 => n2328, A2 => n3520, B1 => n3917, B2 => 
                           n3544, ZN => n13595);
   U4110 : AOI22_X1 port map( A1 => n2334, A2 => n3520, B1 => n3923, B2 => 
                           n3542, ZN => n13596);
   U4111 : AOI22_X1 port map( A1 => n2346, A2 => n3520, B1 => n3929, B2 => 
                           n3542, ZN => n13598);
   U4112 : AOI22_X1 port map( A1 => n2358, A2 => n3520, B1 => n3941, B2 => 
                           n3546, ZN => n13600);
   U4113 : AOI22_X1 port map( A1 => n2364, A2 => n3519, B1 => n3947, B2 => 
                           n3542, ZN => n13601);
   U4114 : AOI22_X1 port map( A1 => n2370, A2 => n3519, B1 => n3953, B2 => 
                           n3548, ZN => n13602);
   U4115 : AOI22_X1 port map( A1 => n2376, A2 => n3519, B1 => n3959, B2 => 
                           n3547, ZN => n13603);
   U4116 : AOI22_X1 port map( A1 => n2382, A2 => n3519, B1 => n3965, B2 => 
                           n3548, ZN => n13604);
   U4117 : AOI22_X1 port map( A1 => n2388, A2 => n3519, B1 => n3971, B2 => 
                           n3543, ZN => n13605);
   U4118 : AOI22_X1 port map( A1 => n2394, A2 => n3519, B1 => n3977, B2 => 
                           n3547, ZN => n13606);
   U4119 : AOI22_X1 port map( A1 => n2400, A2 => n3519, B1 => n3983, B2 => 
                           n3543, ZN => n13607);
   U4120 : AOI22_X1 port map( A1 => n2412, A2 => n3519, B1 => n3989, B2 => 
                           n3545, ZN => n13609);
   U4121 : AOI22_X1 port map( A1 => n2418, A2 => n3519, B1 => n3995, B2 => 
                           n3544, ZN => n13610);
   U4122 : AOI22_X1 port map( A1 => n2424, A2 => n3519, B1 => n4001, B2 => 
                           n3544, ZN => n13611);
   U4123 : AOI22_X1 port map( A1 => n2340, A2 => n3520, B1 => n4091, B2 => 
                           n3546, ZN => n13597);
   U4124 : AOI22_X1 port map( A1 => n2406, A2 => n3519, B1 => n4097, B2 => 
                           n3543, ZN => n13608);
   U4125 : AOI22_X1 port map( A1 => n2329, A2 => n3641, B1 => n3918, B2 => 
                           n3656, ZN => n13851);
   U4126 : AOI22_X1 port map( A1 => n2335, A2 => n3640, B1 => n3924, B2 => 
                           n3654, ZN => n13852);
   U4127 : AOI22_X1 port map( A1 => n2347, A2 => n3639, B1 => n3930, B2 => 
                           n3654, ZN => n13854);
   U4128 : AOI22_X1 port map( A1 => n2359, A2 => n3631, B1 => n3942, B2 => 
                           n3658, ZN => n13856);
   U4129 : AOI22_X1 port map( A1 => n2365, A2 => n3631, B1 => n3948, B2 => 
                           n3654, ZN => n13857);
   U4130 : AOI22_X1 port map( A1 => n2371, A2 => n3631, B1 => n3954, B2 => 
                           n3660, ZN => n13858);
   U4131 : AOI22_X1 port map( A1 => n2377, A2 => n3631, B1 => n3960, B2 => 
                           n3659, ZN => n13859);
   U4132 : AOI22_X1 port map( A1 => n2383, A2 => n3631, B1 => n3966, B2 => 
                           n3660, ZN => n13860);
   U4133 : AOI22_X1 port map( A1 => n2389, A2 => n3631, B1 => n3972, B2 => 
                           n3655, ZN => n13861);
   U4134 : AOI22_X1 port map( A1 => n2395, A2 => n3631, B1 => n3978, B2 => 
                           n3659, ZN => n13862);
   U4135 : AOI22_X1 port map( A1 => n2401, A2 => n3631, B1 => n3984, B2 => 
                           n3655, ZN => n13863);
   U4136 : AOI22_X1 port map( A1 => n2413, A2 => n3631, B1 => n3990, B2 => 
                           n3657, ZN => n13865);
   U4137 : AOI22_X1 port map( A1 => n2419, A2 => n3631, B1 => n3996, B2 => 
                           n3656, ZN => n13866);
   U4138 : AOI22_X1 port map( A1 => n2425, A2 => n3631, B1 => n4002, B2 => 
                           n3656, ZN => n13867);
   U4139 : AOI22_X1 port map( A1 => n2341, A2 => n3641, B1 => n4092, B2 => 
                           n3658, ZN => n13853);
   U4140 : AOI22_X1 port map( A1 => n2407, A2 => n3631, B1 => n4098, B2 => 
                           n3655, ZN => n13864);
   U4141 : AOI22_X1 port map( A1 => n2329, A2 => n3749, B1 => n3918, B2 => 
                           n3768, ZN => n14107);
   U4142 : AOI22_X1 port map( A1 => n2335, A2 => n3750, B1 => n3924, B2 => 
                           n3766, ZN => n14108);
   U4143 : AOI22_X1 port map( A1 => n2347, A2 => n3747, B1 => n3930, B2 => 
                           n3766, ZN => n14110);
   U4144 : AOI22_X1 port map( A1 => n2359, A2 => n3752, B1 => n3942, B2 => 
                           n3770, ZN => n14112);
   U4145 : AOI22_X1 port map( A1 => n2365, A2 => n3746, B1 => n3948, B2 => 
                           n3766, ZN => n14113);
   U4146 : AOI22_X1 port map( A1 => n2371, A2 => n3748, B1 => n3954, B2 => 
                           n3772, ZN => n14114);
   U4147 : AOI22_X1 port map( A1 => n2377, A2 => n3749, B1 => n3960, B2 => 
                           n3771, ZN => n14115);
   U4148 : AOI22_X1 port map( A1 => n2383, A2 => n3750, B1 => n3966, B2 => 
                           n3772, ZN => n14116);
   U4149 : AOI22_X1 port map( A1 => n2389, A2 => n3747, B1 => n3972, B2 => 
                           n3767, ZN => n14117);
   U4150 : AOI22_X1 port map( A1 => n2395, A2 => n3743, B1 => n3978, B2 => 
                           n3771, ZN => n14118);
   U4151 : AOI22_X1 port map( A1 => n2401, A2 => n3753, B1 => n3984, B2 => 
                           n3767, ZN => n14119);
   U4152 : AOI22_X1 port map( A1 => n2413, A2 => n3751, B1 => n3990, B2 => 
                           n3769, ZN => n14121);
   U4153 : AOI22_X1 port map( A1 => n2419, A2 => n3753, B1 => n3996, B2 => 
                           n3768, ZN => n14122);
   U4154 : AOI22_X1 port map( A1 => n2425, A2 => n3752, B1 => n4002, B2 => 
                           n3768, ZN => n14123);
   U4155 : AOI22_X1 port map( A1 => n2341, A2 => n3744, B1 => n4092, B2 => 
                           n3770, ZN => n14109);
   U4156 : AOI22_X1 port map( A1 => n2407, A2 => n3743, B1 => n4098, B2 => 
                           n3767, ZN => n14120);
   U4157 : AOI22_X1 port map( A1 => n11511, A2 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_3_port
                           , B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_3_port
                           , B2 => n12927, ZN => n12895);
   U4158 : AOI22_X1 port map( A1 => n3369, A2 => n4048, B1 => n2288, B2 => 
                           n3304, ZN => n13108);
   U4159 : AOI22_X1 port map( A1 => n4054, A2 => n3306, B1 => n2294, B2 => 
                           n3305, ZN => n13109);
   U4160 : AOI22_X1 port map( A1 => n4060, A2 => n3306, B1 => n2300, B2 => 
                           n3304, ZN => n13110);
   U4161 : AOI22_X1 port map( A1 => n4066, A2 => n3307, B1 => n2306, B2 => 
                           n3305, ZN => n13111);
   U4162 : AOI22_X1 port map( A1 => n4072, A2 => n3307, B1 => n2312, B2 => 
                           n3305, ZN => n13112);
   U4163 : AOI22_X1 port map( A1 => n4078, A2 => n3307, B1 => n2318, B2 => 
                           n3305, ZN => n13113);
   U4164 : AOI22_X1 port map( A1 => n4084, A2 => n3307, B1 => n2324, B2 => 
                           n3305, ZN => n13114);
   U4165 : AOI22_X1 port map( A1 => n3481, A2 => n4048, B1 => n2288, B2 => 
                           n3417, ZN => n13332);
   U4166 : AOI22_X1 port map( A1 => n4054, A2 => n3418, B1 => n2294, B2 => 
                           n3417, ZN => n13333);
   U4167 : AOI22_X1 port map( A1 => n4060, A2 => n3418, B1 => n2300, B2 => 
                           n3417, ZN => n13334);
   U4168 : AOI22_X1 port map( A1 => n4066, A2 => n3419, B1 => n2306, B2 => 
                           n3417, ZN => n13335);
   U4169 : AOI22_X1 port map( A1 => n4072, A2 => n3419, B1 => n2312, B2 => 
                           n3417, ZN => n13336);
   U4170 : AOI22_X1 port map( A1 => n4078, A2 => n3419, B1 => n2318, B2 => 
                           n3417, ZN => n13337);
   U4171 : AOI22_X1 port map( A1 => n4084, A2 => n3419, B1 => n2324, B2 => 
                           n3417, ZN => n13338);
   U4172 : AOI22_X1 port map( A1 => n3593, A2 => n4049, B1 => n2287, B2 => 
                           n3529, ZN => n13588);
   U4173 : AOI22_X1 port map( A1 => n4055, A2 => n3530, B1 => n2293, B2 => 
                           n3529, ZN => n13589);
   U4174 : AOI22_X1 port map( A1 => n4061, A2 => n3530, B1 => n2299, B2 => 
                           n3529, ZN => n13590);
   U4175 : AOI22_X1 port map( A1 => n4067, A2 => n3531, B1 => n2305, B2 => 
                           n3529, ZN => n13591);
   U4176 : AOI22_X1 port map( A1 => n4073, A2 => n3531, B1 => n2311, B2 => 
                           n3529, ZN => n13592);
   U4177 : AOI22_X1 port map( A1 => n4079, A2 => n3531, B1 => n2317, B2 => 
                           n3529, ZN => n13593);
   U4178 : AOI22_X1 port map( A1 => n4085, A2 => n3531, B1 => n2323, B2 => 
                           n3529, ZN => n13594);
   U4179 : AOI22_X1 port map( A1 => n3705, A2 => n4050, B1 => n2286, B2 => 
                           n3640, ZN => n13844);
   U4180 : AOI22_X1 port map( A1 => n4056, A2 => n3642, B1 => n2292, B2 => 
                           n3641, ZN => n13845);
   U4181 : AOI22_X1 port map( A1 => n4062, A2 => n3642, B1 => n2298, B2 => 
                           n3631, ZN => n13846);
   U4182 : AOI22_X1 port map( A1 => n4068, A2 => n3643, B1 => n2304, B2 => 
                           n3639, ZN => n13847);
   U4183 : AOI22_X1 port map( A1 => n4074, A2 => n3643, B1 => n2310, B2 => 
                           n3631, ZN => n13848);
   U4184 : AOI22_X1 port map( A1 => n4080, A2 => n3643, B1 => n2316, B2 => 
                           n3631, ZN => n13849);
   U4185 : AOI22_X1 port map( A1 => n4086, A2 => n3643, B1 => n2322, B2 => 
                           n3640, ZN => n13850);
   U4186 : AOI22_X1 port map( A1 => n3817, A2 => n4050, B1 => n2286, B2 => 
                           n3753, ZN => n14100);
   U4187 : AOI22_X1 port map( A1 => n4056, A2 => n3754, B1 => n2292, B2 => 
                           n3753, ZN => n14101);
   U4188 : AOI22_X1 port map( A1 => n4062, A2 => n3754, B1 => n2298, B2 => 
                           n3753, ZN => n14102);
   U4189 : AOI22_X1 port map( A1 => n4068, A2 => n3755, B1 => n2304, B2 => 
                           n3753, ZN => n14103);
   U4190 : AOI22_X1 port map( A1 => n4074, A2 => n3755, B1 => n2310, B2 => 
                           n3753, ZN => n14104);
   U4191 : AOI22_X1 port map( A1 => n4080, A2 => n3755, B1 => n2316, B2 => 
                           n3753, ZN => n14105);
   U4192 : AOI22_X1 port map( A1 => n4086, A2 => n3755, B1 => n2322, B2 => 
                           n3753, ZN => n14106);
   U4193 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_2_port
                           , A2 => n11506, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_2_port
                           , B2 => n12928, ZN => n12899);
   U4194 : AOI22_X1 port map( A1 => n11506, A2 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_3_port
                           , B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_3_port
                           , B2 => n12928, ZN => n12898);
   U4195 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n509, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n510, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n511, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n512, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_108_port);
   U4196 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n445, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n509);
   U4197 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, C1 => n8309, C2 => 
                           n521, A => DataPath_ALUhw_SHIFTER_HW_n520, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n511);
   U4198 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n496, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n497, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n498, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n499, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_109_port);
   U4199 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n432, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n496);
   U4200 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n432, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n405, A => 
                           DataPath_ALUhw_SHIFTER_HW_n500, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n499);
   U4201 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n445, A => 
                           DataPath_ALUhw_SHIFTER_HW_n508, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n497);
   U4202 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n185, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n186, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n187, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n188, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_102_port);
   U4203 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, C1 => n8312, C2 => 
                           n523, ZN => DataPath_ALUhw_SHIFTER_HW_n185);
   U4204 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, A => 
                           DataPath_ALUhw_SHIFTER_HW_n189, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n188);
   U4205 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, A => 
                           DataPath_ALUhw_SHIFTER_HW_n193, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n186);
   U4206 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n175, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n176, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n177, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n178, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_103_port);
   U4207 : AOI222_X1 port map( A1 => n8306, A2 => n523, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n175);
   U4208 : AOI221_X1 port map( B1 => n8304, B2 => n523, C1 => n260, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, A => 
                           DataPath_ALUhw_SHIFTER_HW_n180, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n178);
   U4209 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, A => 
                           DataPath_ALUhw_SHIFTER_HW_n184, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n176);
   U4210 : AOI21_X1 port map( B1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_4_28_port, B2
                           => n8326, A => n11523, ZN => n12932);
   U4211 : AND2_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_28_port, A2
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_3_24_port,
                           ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_4_28_port);
   U4212 : INV_X1 port map( A => n12925, ZN => n11523);
   U4213 : AOI21_X1 port map( B1 => n11524, B2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_28_port, A 
                           => n11531, ZN => n12925);
   U4214 : AOI21_X1 port map( B1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_3_24_port, B2
                           => n8326, A => n11524, ZN => n12931);
   U4215 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n142, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n143, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n144, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n145, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_105_port);
   U4216 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n164, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n142);
   U4217 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, A => 
                           DataPath_ALUhw_SHIFTER_HW_n157, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n143);
   U4218 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, C1 => n8299, C2 => 
                           n521, A => DataPath_ALUhw_SHIFTER_HW_n148, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n145);
   U4219 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n522, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n523, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n524, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n525, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_107_port);
   U4220 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n522);
   U4221 : AOI221_X1 port map( B1 => n8314, B2 => n521, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, A => 
                           DataPath_ALUhw_SHIFTER_HW_n533, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n524);
   U4222 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n212, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n213, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n214, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n215, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_99_port);
   U4223 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n219, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n211, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n212);
   U4224 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n164, A => 
                           DataPath_ALUhw_SHIFTER_HW_n216, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n215);
   U4225 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n202, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n203, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n204, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n205, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_100_port);
   U4226 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n211, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n164, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n201, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n202);
   U4227 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n164, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, A => 
                           DataPath_ALUhw_SHIFTER_HW_n206, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n205);
   U4228 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n269, ZN => n11494);
   U4229 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n535, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n536, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n537, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n538, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_106_port);
   U4230 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n164, B1 => n8307, B2 => 
                           n521, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n535);
   U4231 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, A => 
                           DataPath_ALUhw_SHIFTER_HW_n552, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n536);
   U4232 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, A => 
                           DataPath_ALUhw_SHIFTER_HW_n551, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n537);
   U4233 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n456, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n457, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n458, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n459, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_112_port);
   U4234 : AOI222_X1 port map( A1 => n8306, A2 => n521, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n380, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n456);
   U4235 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n380, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n344, A => 
                           DataPath_ALUhw_SHIFTER_HW_n460, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n459);
   U4236 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n445, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n392, A => 
                           DataPath_ALUhw_SHIFTER_HW_n467, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n457);
   U4237 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n165, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n166, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n167, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n168, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_104_port);
   U4238 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n165);
   U4239 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, A => n11489, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n168);
   U4240 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n164, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, A => 
                           DataPath_ALUhw_SHIFTER_HW_n174, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n166);
   U4241 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n483, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n484, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n485, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n486, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_110_port);
   U4242 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n405, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n483);
   U4243 : AOI221_X1 port map( B1 => n8304, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, C1 => n260, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, A => 
                           DataPath_ALUhw_SHIFTER_HW_n487, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n486);
   U4244 : AOI221_X1 port map( B1 => n8311, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, C1 => n8310, C2 => 
                           n521, A => DataPath_ALUhw_SHIFTER_HW_n494, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n485);
   U4245 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n468, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n469, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n470, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n471, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_111_port);
   U4246 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n392, C1 => n8312, C2 => 
                           n521, ZN => DataPath_ALUhw_SHIFTER_HW_n468);
   U4247 : AOI221_X1 port map( B1 => n8304, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n146, C1 => n260, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, A => 
                           DataPath_ALUhw_SHIFTER_HW_n472, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n471);
   U4248 : AOI221_X1 port map( B1 => n8311, B2 => n521, C1 => n8310, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, A => 
                           DataPath_ALUhw_SHIFTER_HW_n481, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n470);
   U4249 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n194, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n195, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n196, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n197, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_101_port);
   U4250 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n201, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n194);
   U4251 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n156, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n172, A => 
                           DataPath_ALUhw_SHIFTER_HW_n198, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n197);
   U4252 : AOI221_X1 port map( B1 => n8305, B2 => n523, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n164, A => 
                           DataPath_ALUhw_SHIFTER_HW_n200, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n195);
   U4253 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n262, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n263, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n264, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n265, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_98_port);
   U4254 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n269, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n219, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n262);
   U4255 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, A => 
                           DataPath_ALUhw_SHIFTER_HW_n266, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n265);
   U4256 : AOI221_X1 port map( B1 => n8314, B2 => n523, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, A => 
                           DataPath_ALUhw_SHIFTER_HW_n267, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n264);
   U4257 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n406, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n407, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n408, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n409, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_97_port);
   U4258 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n419, B1 => n8307, B2 => 
                           n523, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n269, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n406);
   U4259 : AOI221_X1 port map( B1 => n8300, B2 => n523, C1 => n8299, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, A => 
                           DataPath_ALUhw_SHIFTER_HW_n410, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n409);
   U4260 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n201, A => 
                           DataPath_ALUhw_SHIFTER_HW_n417, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n408);
   U4261 : AOI21_X1 port map( B1 => n8324, B2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_26_port, A 
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_26_port,
                           ZN => n12915);
   U4262 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n419, ZN => n11495);
   U4263 : BUF_X1 port map( A => n2281, Z => n2276);
   U4264 : BUF_X1 port map( A => n2281, Z => n2277);
   U4265 : BUF_X1 port map( A => n2280, Z => n2278);
   U4266 : AND2_X1 port map( A1 => n1861, A2 => n2130, ZN => n1859);
   U4267 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n588, ZN => n11496);
   U4268 : BUF_X1 port map( A => n7989, Z => n2275);
   U4269 : XNOR2_X1 port map( A => n4270, B => n2154, ZN => n1860);
   U4270 : BUF_X1 port map( A => n7970, Z => n2187);
   U4271 : INV_X1 port map( A => n12892, ZN => n11515);
   U4272 : AOI22_X1 port map( A1 => n11516, A2 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_3_port
                           , B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_3_port
                           , B2 => n12926, ZN => n12892);
   U4273 : AND2_X1 port map( A1 => n364, A2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_27_port, ZN
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_28_port)
                           ;
   U4274 : AND2_X1 port map( A1 => n375, A2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_22_port, ZN
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_24_port)
                           ;
   U4275 : AND2_X1 port map( A1 => n373, A2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_10_port, ZN
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_12_port)
                           ;
   U4276 : AND2_X1 port map( A1 => n376, A2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_18_port, ZN
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_20_port)
                           ;
   U4277 : BUF_X1 port map( A => n2280, Z => n2279);
   U4278 : AND2_X1 port map( A1 => n830, A2 => n2264, ZN => n1861);
   U4279 : INV_X1 port map( A => n12893, ZN => n11514);
   U4280 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_2_port
                           , A2 => n11516, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_2_port
                           , B2 => n12926, ZN => n12893);
   U4281 : INV_X1 port map( A => n12894, ZN => n11513);
   U4282 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_1_port
                           , A2 => n11516, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_1_port
                           , B2 => n12926, ZN => n12894);
   U4283 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n169, ZN => n11489);
   U4284 : AOI22_X1 port map( A1 => n523, A2 => n260, B1 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, B2 => n8304, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n169);
   U4285 : BUF_X1 port map( A => n3284, Z => n3373);
   U4286 : BUF_X1 port map( A => n3284, Z => n3374);
   U4287 : BUF_X1 port map( A => n3396, Z => n3486);
   U4288 : BUF_X1 port map( A => n3396, Z => n3485);
   U4289 : BUF_X1 port map( A => n3508, Z => n3598);
   U4290 : BUF_X1 port map( A => n3508, Z => n3597);
   U4291 : BUF_X1 port map( A => n3732, Z => n3822);
   U4292 : BUF_X1 port map( A => n3732, Z => n3821);
   U4293 : INV_X1 port map( A => n13090, ZN => n12291);
   U4294 : AOI22_X1 port map( A1 => n2369, A2 => n3295, B1 => n3952, B2 => 
                           n3364, ZN => n13090);
   U4295 : INV_X1 port map( A => n13091, ZN => n12251);
   U4296 : AOI22_X1 port map( A1 => n2375, A2 => n3295, B1 => n3958, B2 => 
                           n3364, ZN => n13091);
   U4297 : INV_X1 port map( A => n13092, ZN => n12211);
   U4298 : AOI22_X1 port map( A1 => n2381, A2 => n3295, B1 => n3964, B2 => 
                           n3364, ZN => n13092);
   U4299 : INV_X1 port map( A => n13093, ZN => n12171);
   U4300 : AOI22_X1 port map( A1 => n2387, A2 => n3295, B1 => n3970, B2 => 
                           n3364, ZN => n13093);
   U4301 : INV_X1 port map( A => n13094, ZN => n12131);
   U4302 : AOI22_X1 port map( A1 => n2393, A2 => n3295, B1 => n3976, B2 => 
                           n3365, ZN => n13094);
   U4303 : INV_X1 port map( A => n13095, ZN => n12091);
   U4304 : AOI22_X1 port map( A1 => n2399, A2 => n3295, B1 => n3982, B2 => 
                           n3365, ZN => n13095);
   U4305 : INV_X1 port map( A => n13097, ZN => n12011);
   U4306 : AOI22_X1 port map( A1 => n2411, A2 => n3295, B1 => n3988, B2 => 
                           n3365, ZN => n13097);
   U4307 : INV_X1 port map( A => n13098, ZN => n11971);
   U4308 : AOI22_X1 port map( A1 => n2417, A2 => n3295, B1 => n3994, B2 => 
                           n3366, ZN => n13098);
   U4309 : INV_X1 port map( A => n13099, ZN => n11931);
   U4310 : AOI22_X1 port map( A1 => n2423, A2 => n3295, B1 => n4000, B2 => 
                           n3366, ZN => n13099);
   U4311 : INV_X1 port map( A => n13100, ZN => n11891);
   U4312 : AOI22_X1 port map( A1 => n2429, A2 => n3295, B1 => n4006, B2 => 
                           n3366, ZN => n13100);
   U4313 : INV_X1 port map( A => n13101, ZN => n11851);
   U4314 : AOI22_X1 port map( A1 => n2435, A2 => n3295, B1 => n4012, B2 => 
                           n3367, ZN => n13101);
   U4315 : INV_X1 port map( A => n13096, ZN => n12051);
   U4316 : AOI22_X1 port map( A1 => n2405, A2 => n3295, B1 => n4096, B2 => 
                           n3365, ZN => n13096);
   U4317 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n65, ZN => n11647);
   U4318 : AOI22_X1 port map( A1 => n2474, A2 => n3299, B1 => n4105, B2 => 
                           n3356, ZN => DataPath_RF_MUX_SELINPUT_8_n65);
   U4319 : INV_X1 port map( A => n13314, ZN => n12298);
   U4320 : AOI22_X1 port map( A1 => n2369, A2 => n3409, B1 => n3952, B2 => 
                           n3476, ZN => n13314);
   U4321 : INV_X1 port map( A => n13315, ZN => n12258);
   U4322 : AOI22_X1 port map( A1 => n2375, A2 => n3409, B1 => n3958, B2 => 
                           n3476, ZN => n13315);
   U4323 : INV_X1 port map( A => n13316, ZN => n12218);
   U4324 : AOI22_X1 port map( A1 => n2381, A2 => n3409, B1 => n3964, B2 => 
                           n3476, ZN => n13316);
   U4325 : INV_X1 port map( A => n13317, ZN => n12178);
   U4326 : AOI22_X1 port map( A1 => n2387, A2 => n3409, B1 => n3970, B2 => 
                           n3476, ZN => n13317);
   U4327 : INV_X1 port map( A => n13318, ZN => n12138);
   U4328 : AOI22_X1 port map( A1 => n2393, A2 => n3409, B1 => n3976, B2 => 
                           n3477, ZN => n13318);
   U4329 : INV_X1 port map( A => n13319, ZN => n12098);
   U4330 : AOI22_X1 port map( A1 => n2399, A2 => n3409, B1 => n3982, B2 => 
                           n3477, ZN => n13319);
   U4331 : INV_X1 port map( A => n13321, ZN => n12018);
   U4332 : AOI22_X1 port map( A1 => n2411, A2 => n3409, B1 => n3988, B2 => 
                           n3477, ZN => n13321);
   U4333 : INV_X1 port map( A => n13322, ZN => n11978);
   U4334 : AOI22_X1 port map( A1 => n2417, A2 => n3409, B1 => n3994, B2 => 
                           n3478, ZN => n13322);
   U4335 : INV_X1 port map( A => n13323, ZN => n11938);
   U4336 : AOI22_X1 port map( A1 => n2423, A2 => n3409, B1 => n4000, B2 => 
                           n3478, ZN => n13323);
   U4337 : INV_X1 port map( A => n13324, ZN => n11898);
   U4338 : AOI22_X1 port map( A1 => n2429, A2 => n3409, B1 => n4006, B2 => 
                           n3478, ZN => n13324);
   U4339 : INV_X1 port map( A => n13325, ZN => n11858);
   U4340 : AOI22_X1 port map( A1 => n2435, A2 => n3409, B1 => n4012, B2 => 
                           n3479, ZN => n13325);
   U4341 : INV_X1 port map( A => n13320, ZN => n12058);
   U4342 : AOI22_X1 port map( A1 => n2405, A2 => n3409, B1 => n4096, B2 => 
                           n3477, ZN => n13320);
   U4343 : INV_X1 port map( A => n13570, ZN => n12306);
   U4344 : AOI22_X1 port map( A1 => n2370, A2 => n3521, B1 => n3953, B2 => 
                           n3588, ZN => n13570);
   U4345 : INV_X1 port map( A => n13571, ZN => n12266);
   U4346 : AOI22_X1 port map( A1 => n2376, A2 => n3521, B1 => n3959, B2 => 
                           n3588, ZN => n13571);
   U4347 : INV_X1 port map( A => n13572, ZN => n12226);
   U4348 : AOI22_X1 port map( A1 => n2382, A2 => n3521, B1 => n3965, B2 => 
                           n3588, ZN => n13572);
   U4349 : INV_X1 port map( A => n13573, ZN => n12186);
   U4350 : AOI22_X1 port map( A1 => n2388, A2 => n3521, B1 => n3971, B2 => 
                           n3588, ZN => n13573);
   U4351 : INV_X1 port map( A => n13574, ZN => n12146);
   U4352 : AOI22_X1 port map( A1 => n2394, A2 => n3521, B1 => n3977, B2 => 
                           n3589, ZN => n13574);
   U4353 : INV_X1 port map( A => n13575, ZN => n12106);
   U4354 : AOI22_X1 port map( A1 => n2400, A2 => n3521, B1 => n3983, B2 => 
                           n3589, ZN => n13575);
   U4355 : INV_X1 port map( A => n13577, ZN => n12026);
   U4356 : AOI22_X1 port map( A1 => n2412, A2 => n3521, B1 => n3989, B2 => 
                           n3589, ZN => n13577);
   U4357 : INV_X1 port map( A => n13578, ZN => n11986);
   U4358 : AOI22_X1 port map( A1 => n2418, A2 => n3521, B1 => n3995, B2 => 
                           n3590, ZN => n13578);
   U4359 : INV_X1 port map( A => n13579, ZN => n11946);
   U4360 : AOI22_X1 port map( A1 => n2424, A2 => n3521, B1 => n4001, B2 => 
                           n3590, ZN => n13579);
   U4361 : INV_X1 port map( A => n13580, ZN => n11906);
   U4362 : AOI22_X1 port map( A1 => n2430, A2 => n3521, B1 => n4007, B2 => 
                           n3590, ZN => n13580);
   U4363 : INV_X1 port map( A => n13581, ZN => n11866);
   U4364 : AOI22_X1 port map( A1 => n2436, A2 => n3521, B1 => n4013, B2 => 
                           n3591, ZN => n13581);
   U4365 : INV_X1 port map( A => n13576, ZN => n12066);
   U4366 : AOI22_X1 port map( A1 => n2406, A2 => n3521, B1 => n4097, B2 => 
                           n3589, ZN => n13576);
   U4367 : INV_X1 port map( A => n13826, ZN => n12314);
   U4368 : AOI22_X1 port map( A1 => n2371, A2 => n3632, B1 => n3954, B2 => 
                           n3700, ZN => n13826);
   U4369 : INV_X1 port map( A => n13827, ZN => n12274);
   U4370 : AOI22_X1 port map( A1 => n2377, A2 => n3632, B1 => n3960, B2 => 
                           n3700, ZN => n13827);
   U4371 : INV_X1 port map( A => n13828, ZN => n12234);
   U4372 : AOI22_X1 port map( A1 => n2383, A2 => n3632, B1 => n3966, B2 => 
                           n3700, ZN => n13828);
   U4373 : INV_X1 port map( A => n13829, ZN => n12194);
   U4374 : AOI22_X1 port map( A1 => n2389, A2 => n3632, B1 => n3972, B2 => 
                           n3700, ZN => n13829);
   U4375 : INV_X1 port map( A => n13830, ZN => n12154);
   U4376 : AOI22_X1 port map( A1 => n2395, A2 => n3632, B1 => n3978, B2 => 
                           n3701, ZN => n13830);
   U4377 : INV_X1 port map( A => n13831, ZN => n12114);
   U4378 : AOI22_X1 port map( A1 => n2401, A2 => n3632, B1 => n3984, B2 => 
                           n3701, ZN => n13831);
   U4379 : INV_X1 port map( A => n13833, ZN => n12034);
   U4380 : AOI22_X1 port map( A1 => n2413, A2 => n3632, B1 => n3990, B2 => 
                           n3701, ZN => n13833);
   U4381 : INV_X1 port map( A => n13834, ZN => n11994);
   U4382 : AOI22_X1 port map( A1 => n2419, A2 => n3632, B1 => n3996, B2 => 
                           n3702, ZN => n13834);
   U4383 : INV_X1 port map( A => n13835, ZN => n11954);
   U4384 : AOI22_X1 port map( A1 => n2425, A2 => n3632, B1 => n4002, B2 => 
                           n3702, ZN => n13835);
   U4385 : INV_X1 port map( A => n13836, ZN => n11914);
   U4386 : AOI22_X1 port map( A1 => n2431, A2 => n3632, B1 => n4008, B2 => 
                           n3702, ZN => n13836);
   U4387 : INV_X1 port map( A => n13837, ZN => n11874);
   U4388 : AOI22_X1 port map( A1 => n2437, A2 => n3632, B1 => n4014, B2 => 
                           n3703, ZN => n13837);
   U4389 : INV_X1 port map( A => n13832, ZN => n12074);
   U4390 : AOI22_X1 port map( A1 => n2407, A2 => n3632, B1 => n4098, B2 => 
                           n3701, ZN => n13832);
   U4391 : INV_X1 port map( A => n14082, ZN => n12322);
   U4392 : AOI22_X1 port map( A1 => n2371, A2 => n3752, B1 => n3954, B2 => 
                           n3812, ZN => n14082);
   U4393 : INV_X1 port map( A => n14083, ZN => n12282);
   U4394 : AOI22_X1 port map( A1 => n2377, A2 => n3751, B1 => n3960, B2 => 
                           n3812, ZN => n14083);
   U4395 : INV_X1 port map( A => n14084, ZN => n12242);
   U4396 : AOI22_X1 port map( A1 => n2383, A2 => n3743, B1 => n3966, B2 => 
                           n3812, ZN => n14084);
   U4397 : INV_X1 port map( A => n14085, ZN => n12202);
   U4398 : AOI22_X1 port map( A1 => n2389, A2 => n3753, B1 => n3972, B2 => 
                           n3812, ZN => n14085);
   U4399 : INV_X1 port map( A => n14086, ZN => n12162);
   U4400 : AOI22_X1 port map( A1 => n2395, A2 => n3752, B1 => n3978, B2 => 
                           n3813, ZN => n14086);
   U4401 : INV_X1 port map( A => n14087, ZN => n12122);
   U4402 : AOI22_X1 port map( A1 => n2401, A2 => n3751, B1 => n3984, B2 => 
                           n3813, ZN => n14087);
   U4403 : INV_X1 port map( A => n14089, ZN => n12042);
   U4404 : AOI22_X1 port map( A1 => n2413, A2 => n3753, B1 => n3990, B2 => 
                           n3813, ZN => n14089);
   U4405 : INV_X1 port map( A => n14090, ZN => n12002);
   U4406 : AOI22_X1 port map( A1 => n2419, A2 => n3752, B1 => n3996, B2 => 
                           n3814, ZN => n14090);
   U4407 : INV_X1 port map( A => n14091, ZN => n11962);
   U4408 : AOI22_X1 port map( A1 => n2425, A2 => n3751, B1 => n4002, B2 => 
                           n3814, ZN => n14091);
   U4409 : INV_X1 port map( A => n14092, ZN => n11922);
   U4410 : AOI22_X1 port map( A1 => n2431, A2 => n3753, B1 => n4008, B2 => 
                           n3814, ZN => n14092);
   U4411 : INV_X1 port map( A => n14093, ZN => n11882);
   U4412 : AOI22_X1 port map( A1 => n2437, A2 => n3752, B1 => n4014, B2 => 
                           n3815, ZN => n14093);
   U4413 : INV_X1 port map( A => n14088, ZN => n12082);
   U4414 : AOI22_X1 port map( A1 => n2407, A2 => n3751, B1 => n4098, B2 => 
                           n3813, ZN => n14088);
   U4415 : INV_X1 port map( A => n13203, ZN => n11614);
   U4416 : AOI22_X1 port map( A1 => n2471, A2 => n3299, B1 => n4102, B2 => 
                           n3337, ZN => n13203);
   U4417 : INV_X1 port map( A => n13407, ZN => n12421);
   U4418 : AOI22_X1 port map( A1 => n2352, A2 => n3411, B1 => n3935, B2 => 
                           n3444, ZN => n13407);
   U4419 : INV_X1 port map( A => n13663, ZN => n12429);
   U4420 : AOI22_X1 port map( A1 => n2352, A2 => n3523, B1 => n3935, B2 => 
                           n3556, ZN => n13663);
   U4421 : INV_X1 port map( A => n13919, ZN => n12437);
   U4422 : AOI22_X1 port map( A1 => n2353, A2 => n3635, B1 => n3936, B2 => 
                           n3668, ZN => n13919);
   U4423 : INV_X1 port map( A => n14175, ZN => n12445);
   U4424 : AOI22_X1 port map( A1 => n2354, A2 => n3746, B1 => n3937, B2 => 
                           n3780, ZN => n14175);
   U4425 : INV_X1 port map( A => n12988, ZN => n12528);
   U4426 : AOI22_X1 port map( A1 => n2333, A2 => n3299, B1 => n3922, B2 => 
                           n3343, ZN => n12988);
   U4427 : INV_X1 port map( A => n12990, ZN => n12448);
   U4428 : AOI22_X1 port map( A1 => n2345, A2 => n3299, B1 => n3928, B2 => 
                           n3344, ZN => n12990);
   U4429 : INV_X1 port map( A => n12991, ZN => n12408);
   U4430 : AOI22_X1 port map( A1 => n2351, A2 => n3299, B1 => n3934, B2 => 
                           n3344, ZN => n12991);
   U4431 : INV_X1 port map( A => n12992, ZN => n12368);
   U4432 : AOI22_X1 port map( A1 => n2357, A2 => n3299, B1 => n3940, B2 => 
                           n3344, ZN => n12992);
   U4433 : INV_X1 port map( A => n12993, ZN => n12328);
   U4434 : AOI22_X1 port map( A1 => n2363, A2 => n3299, B1 => n3946, B2 => 
                           n3344, ZN => n12993);
   U4435 : INV_X1 port map( A => n12994, ZN => n12288);
   U4436 : AOI22_X1 port map( A1 => n2369, A2 => n3299, B1 => n3952, B2 => 
                           n3345, ZN => n12994);
   U4437 : INV_X1 port map( A => n12995, ZN => n12248);
   U4438 : AOI22_X1 port map( A1 => n2375, A2 => n3299, B1 => n3958, B2 => 
                           n3345, ZN => n12995);
   U4439 : INV_X1 port map( A => n12996, ZN => n12208);
   U4440 : AOI22_X1 port map( A1 => n2381, A2 => n3299, B1 => n3964, B2 => 
                           n3345, ZN => n12996);
   U4441 : INV_X1 port map( A => n12997, ZN => n12168);
   U4442 : AOI22_X1 port map( A1 => n2387, A2 => n3299, B1 => n3970, B2 => 
                           n3345, ZN => n12997);
   U4443 : INV_X1 port map( A => n12989, ZN => n12488);
   U4444 : AOI22_X1 port map( A1 => n2339, A2 => n3299, B1 => n4090, B2 => 
                           n3343, ZN => n12989);
   U4445 : INV_X1 port map( A => n13212, ZN => n12535);
   U4446 : AOI22_X1 port map( A1 => n2333, A2 => n3411, B1 => n3922, B2 => 
                           n3455, ZN => n13212);
   U4447 : INV_X1 port map( A => n13214, ZN => n12455);
   U4448 : AOI22_X1 port map( A1 => n2345, A2 => n3411, B1 => n3928, B2 => 
                           n3456, ZN => n13214);
   U4449 : INV_X1 port map( A => n13215, ZN => n12415);
   U4450 : AOI22_X1 port map( A1 => n2351, A2 => n3411, B1 => n3934, B2 => 
                           n3456, ZN => n13215);
   U4451 : INV_X1 port map( A => n13216, ZN => n12375);
   U4452 : AOI22_X1 port map( A1 => n2357, A2 => n3411, B1 => n3940, B2 => 
                           n3456, ZN => n13216);
   U4453 : INV_X1 port map( A => n13217, ZN => n12335);
   U4454 : AOI22_X1 port map( A1 => n2363, A2 => n3411, B1 => n3946, B2 => 
                           n3456, ZN => n13217);
   U4455 : INV_X1 port map( A => n13218, ZN => n12295);
   U4456 : AOI22_X1 port map( A1 => n2369, A2 => n3411, B1 => n3952, B2 => 
                           n3457, ZN => n13218);
   U4457 : INV_X1 port map( A => n13219, ZN => n12255);
   U4458 : AOI22_X1 port map( A1 => n2375, A2 => n3411, B1 => n3958, B2 => 
                           n3457, ZN => n13219);
   U4459 : INV_X1 port map( A => n13220, ZN => n12215);
   U4460 : AOI22_X1 port map( A1 => n2381, A2 => n3411, B1 => n3964, B2 => 
                           n3457, ZN => n13220);
   U4461 : INV_X1 port map( A => n13221, ZN => n12175);
   U4462 : AOI22_X1 port map( A1 => n2387, A2 => n3411, B1 => n3970, B2 => 
                           n3457, ZN => n13221);
   U4463 : INV_X1 port map( A => n13357, ZN => n11859);
   U4464 : AOI22_X1 port map( A1 => n2435, A2 => n3411, B1 => n4012, B2 => 
                           n3432, ZN => n13357);
   U4465 : INV_X1 port map( A => n13213, ZN => n12495);
   U4466 : AOI22_X1 port map( A1 => n2339, A2 => n3411, B1 => n4090, B2 => 
                           n3455, ZN => n13213);
   U4467 : INV_X1 port map( A => n13468, ZN => n12543);
   U4468 : AOI22_X1 port map( A1 => n2334, A2 => n3523, B1 => n3923, B2 => 
                           n3567, ZN => n13468);
   U4469 : INV_X1 port map( A => n13470, ZN => n12463);
   U4470 : AOI22_X1 port map( A1 => n2346, A2 => n3523, B1 => n3929, B2 => 
                           n3568, ZN => n13470);
   U4471 : INV_X1 port map( A => n13471, ZN => n12423);
   U4472 : AOI22_X1 port map( A1 => n2352, A2 => n3523, B1 => n3935, B2 => 
                           n3568, ZN => n13471);
   U4473 : INV_X1 port map( A => n13472, ZN => n12383);
   U4474 : AOI22_X1 port map( A1 => n2358, A2 => n3523, B1 => n3941, B2 => 
                           n3568, ZN => n13472);
   U4475 : INV_X1 port map( A => n13473, ZN => n12343);
   U4476 : AOI22_X1 port map( A1 => n2364, A2 => n3523, B1 => n3947, B2 => 
                           n3568, ZN => n13473);
   U4477 : INV_X1 port map( A => n13474, ZN => n12303);
   U4478 : AOI22_X1 port map( A1 => n2370, A2 => n3523, B1 => n3953, B2 => 
                           n3569, ZN => n13474);
   U4479 : INV_X1 port map( A => n13475, ZN => n12263);
   U4480 : AOI22_X1 port map( A1 => n2376, A2 => n3523, B1 => n3959, B2 => 
                           n3569, ZN => n13475);
   U4481 : INV_X1 port map( A => n13476, ZN => n12223);
   U4482 : AOI22_X1 port map( A1 => n2382, A2 => n3523, B1 => n3965, B2 => 
                           n3569, ZN => n13476);
   U4483 : INV_X1 port map( A => n13477, ZN => n12183);
   U4484 : AOI22_X1 port map( A1 => n2388, A2 => n3523, B1 => n3971, B2 => 
                           n3569, ZN => n13477);
   U4485 : INV_X1 port map( A => n13613, ZN => n11867);
   U4486 : AOI22_X1 port map( A1 => n2436, A2 => n3523, B1 => n4013, B2 => 
                           n3544, ZN => n13613);
   U4487 : INV_X1 port map( A => n13469, ZN => n12503);
   U4488 : AOI22_X1 port map( A1 => n2340, A2 => n3523, B1 => n4091, B2 => 
                           n3567, ZN => n13469);
   U4489 : INV_X1 port map( A => n13724, ZN => n12551);
   U4490 : AOI22_X1 port map( A1 => n2334, A2 => n3635, B1 => n3923, B2 => 
                           n3679, ZN => n13724);
   U4491 : INV_X1 port map( A => n13726, ZN => n12471);
   U4492 : AOI22_X1 port map( A1 => n2346, A2 => n3635, B1 => n3929, B2 => 
                           n3680, ZN => n13726);
   U4493 : INV_X1 port map( A => n13727, ZN => n12431);
   U4494 : AOI22_X1 port map( A1 => n2352, A2 => n3635, B1 => n3935, B2 => 
                           n3680, ZN => n13727);
   U4495 : INV_X1 port map( A => n13728, ZN => n12391);
   U4496 : AOI22_X1 port map( A1 => n2358, A2 => n3635, B1 => n3941, B2 => 
                           n3680, ZN => n13728);
   U4497 : INV_X1 port map( A => n13729, ZN => n12351);
   U4498 : AOI22_X1 port map( A1 => n2364, A2 => n3635, B1 => n3947, B2 => 
                           n3680, ZN => n13729);
   U4499 : INV_X1 port map( A => n13730, ZN => n12311);
   U4500 : AOI22_X1 port map( A1 => n2370, A2 => n3635, B1 => n3953, B2 => 
                           n3681, ZN => n13730);
   U4501 : INV_X1 port map( A => n13731, ZN => n12271);
   U4502 : AOI22_X1 port map( A1 => n2376, A2 => n3635, B1 => n3959, B2 => 
                           n3681, ZN => n13731);
   U4503 : INV_X1 port map( A => n13732, ZN => n12231);
   U4504 : AOI22_X1 port map( A1 => n2382, A2 => n3635, B1 => n3965, B2 => 
                           n3681, ZN => n13732);
   U4505 : INV_X1 port map( A => n13733, ZN => n12191);
   U4506 : AOI22_X1 port map( A1 => n2388, A2 => n3635, B1 => n3971, B2 => 
                           n3681, ZN => n13733);
   U4507 : INV_X1 port map( A => n13869, ZN => n11875);
   U4508 : AOI22_X1 port map( A1 => n2437, A2 => n3635, B1 => n4014, B2 => 
                           n3656, ZN => n13869);
   U4509 : INV_X1 port map( A => n13725, ZN => n12511);
   U4510 : AOI22_X1 port map( A1 => n2340, A2 => n3635, B1 => n4091, B2 => 
                           n3679, ZN => n13725);
   U4511 : INV_X1 port map( A => n13980, ZN => n12559);
   U4512 : AOI22_X1 port map( A1 => n2335, A2 => n3746, B1 => n3924, B2 => 
                           n3791, ZN => n13980);
   U4513 : INV_X1 port map( A => n13982, ZN => n12479);
   U4514 : AOI22_X1 port map( A1 => n2347, A2 => n3746, B1 => n3930, B2 => 
                           n3792, ZN => n13982);
   U4515 : INV_X1 port map( A => n13983, ZN => n12439);
   U4516 : AOI22_X1 port map( A1 => n2353, A2 => n3746, B1 => n3936, B2 => 
                           n3792, ZN => n13983);
   U4517 : INV_X1 port map( A => n13984, ZN => n12399);
   U4518 : AOI22_X1 port map( A1 => n2359, A2 => n3746, B1 => n3942, B2 => 
                           n3792, ZN => n13984);
   U4519 : INV_X1 port map( A => n13985, ZN => n12359);
   U4520 : AOI22_X1 port map( A1 => n2365, A2 => n3746, B1 => n3948, B2 => 
                           n3792, ZN => n13985);
   U4521 : INV_X1 port map( A => n13986, ZN => n12319);
   U4522 : AOI22_X1 port map( A1 => n2371, A2 => n3746, B1 => n3954, B2 => 
                           n3793, ZN => n13986);
   U4523 : INV_X1 port map( A => n13987, ZN => n12279);
   U4524 : AOI22_X1 port map( A1 => n2377, A2 => n3746, B1 => n3960, B2 => 
                           n3793, ZN => n13987);
   U4525 : INV_X1 port map( A => n13988, ZN => n12239);
   U4526 : AOI22_X1 port map( A1 => n2383, A2 => n3746, B1 => n3966, B2 => 
                           n3793, ZN => n13988);
   U4527 : INV_X1 port map( A => n13989, ZN => n12199);
   U4528 : AOI22_X1 port map( A1 => n2389, A2 => n3746, B1 => n3972, B2 => 
                           n3793, ZN => n13989);
   U4529 : INV_X1 port map( A => n14125, ZN => n11883);
   U4530 : AOI22_X1 port map( A1 => n2437, A2 => n3746, B1 => n4014, B2 => 
                           n3768, ZN => n14125);
   U4531 : INV_X1 port map( A => n13981, ZN => n12519);
   U4532 : AOI22_X1 port map( A1 => n2341, A2 => n3746, B1 => n4092, B2 => 
                           n3791, ZN => n13981);
   U4533 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n34, ZN => n12887);
   U4534 : AOI22_X1 port map( A1 => n3369, A2 => n4051, B1 => n2287, B2 => 
                           n3302, ZN => DataPath_RF_MUX_SELINPUT_8_n34);
   U4535 : INV_X1 port map( A => n13076, ZN => n12851);
   U4536 : AOI22_X1 port map( A1 => n3368, A2 => n4048, B1 => n2288, B2 => 
                           n3304, ZN => n13076);
   U4537 : INV_X1 port map( A => n13077, ZN => n12811);
   U4538 : AOI22_X1 port map( A1 => n4054, A2 => n3311, B1 => n2294, B2 => 
                           n3305, ZN => n13077);
   U4539 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n35, ZN => n12847);
   U4540 : AOI22_X1 port map( A1 => n4057, A2 => n3312, B1 => n2293, B2 => 
                           n3304, ZN => DataPath_RF_MUX_SELINPUT_8_n35);
   U4541 : INV_X1 port map( A => n13078, ZN => n12771);
   U4542 : AOI22_X1 port map( A1 => n4060, A2 => n3313, B1 => n2300, B2 => 
                           n3304, ZN => n13078);
   U4543 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n36, ZN => n12807);
   U4544 : AOI22_X1 port map( A1 => n4063, A2 => n3306, B1 => n2299, B2 => 
                           n3295, ZN => DataPath_RF_MUX_SELINPUT_8_n36);
   U4545 : INV_X1 port map( A => n13079, ZN => n12731);
   U4546 : AOI22_X1 port map( A1 => n4066, A2 => n3313, B1 => n2306, B2 => 
                           n3304, ZN => n13079);
   U4547 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n37, ZN => n12767);
   U4548 : AOI22_X1 port map( A1 => n4069, A2 => n3312, B1 => n2305, B2 => 
                           n3303, ZN => DataPath_RF_MUX_SELINPUT_8_n37);
   U4549 : INV_X1 port map( A => n13080, ZN => n12691);
   U4550 : AOI22_X1 port map( A1 => n4072, A2 => n3310, B1 => n2312, B2 => 
                           n3305, ZN => n13080);
   U4551 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n38, ZN => n12727);
   U4552 : AOI22_X1 port map( A1 => n4075, A2 => n3312, B1 => n2311, B2 => 
                           n3305, ZN => DataPath_RF_MUX_SELINPUT_8_n38);
   U4553 : INV_X1 port map( A => n13081, ZN => n12651);
   U4554 : AOI22_X1 port map( A1 => n4078, A2 => n3308, B1 => n2318, B2 => 
                           n3305, ZN => n13081);
   U4555 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n39, ZN => n12687);
   U4556 : AOI22_X1 port map( A1 => n4081, A2 => n3309, B1 => n2317, B2 => 
                           n3303, ZN => DataPath_RF_MUX_SELINPUT_8_n39);
   U4557 : INV_X1 port map( A => n13082, ZN => n12611);
   U4558 : AOI22_X1 port map( A1 => n4084, A2 => n3310, B1 => n2324, B2 => 
                           n3305, ZN => n13082);
   U4559 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n40, ZN => n12647);
   U4560 : AOI22_X1 port map( A1 => n4087, A2 => n3311, B1 => n2323, B2 => 
                           n3303, ZN => DataPath_RF_MUX_SELINPUT_8_n40);
   U4561 : INV_X1 port map( A => n13300, ZN => n12858);
   U4562 : AOI22_X1 port map( A1 => n3480, A2 => n4048, B1 => n2288, B2 => 
                           n3417, ZN => n13300);
   U4563 : INV_X1 port map( A => n13428, ZN => n12862);
   U4564 : AOI22_X1 port map( A1 => n3481, A2 => n4049, B1 => n2287, B2 => 
                           n3416, ZN => n13428);
   U4565 : INV_X1 port map( A => n13301, ZN => n12818);
   U4566 : AOI22_X1 port map( A1 => n4054, A2 => n3423, B1 => n2294, B2 => 
                           n3416, ZN => n13301);
   U4567 : INV_X1 port map( A => n13429, ZN => n12822);
   U4568 : AOI22_X1 port map( A1 => n4055, A2 => n3424, B1 => n2293, B2 => 
                           n3416, ZN => n13429);
   U4569 : INV_X1 port map( A => n13302, ZN => n12778);
   U4570 : AOI22_X1 port map( A1 => n4060, A2 => n3425, B1 => n2300, B2 => 
                           n3416, ZN => n13302);
   U4571 : INV_X1 port map( A => n13430, ZN => n12782);
   U4572 : AOI22_X1 port map( A1 => n4061, A2 => n3418, B1 => n2299, B2 => 
                           n3416, ZN => n13430);
   U4573 : INV_X1 port map( A => n13303, ZN => n12738);
   U4574 : AOI22_X1 port map( A1 => n4066, A2 => n3425, B1 => n2306, B2 => 
                           n3415, ZN => n13303);
   U4575 : INV_X1 port map( A => n13431, ZN => n12742);
   U4576 : AOI22_X1 port map( A1 => n4067, A2 => n3424, B1 => n2305, B2 => 
                           n3416, ZN => n13431);
   U4577 : INV_X1 port map( A => n13304, ZN => n12698);
   U4578 : AOI22_X1 port map( A1 => n4072, A2 => n3422, B1 => n2312, B2 => 
                           n3407, ZN => n13304);
   U4579 : INV_X1 port map( A => n13432, ZN => n12702);
   U4580 : AOI22_X1 port map( A1 => n4073, A2 => n3424, B1 => n2311, B2 => 
                           n3416, ZN => n13432);
   U4581 : INV_X1 port map( A => n13305, ZN => n12658);
   U4582 : AOI22_X1 port map( A1 => n4078, A2 => n3420, B1 => n2318, B2 => 
                           n3408, ZN => n13305);
   U4583 : INV_X1 port map( A => n13433, ZN => n12662);
   U4584 : AOI22_X1 port map( A1 => n4079, A2 => n3421, B1 => n2317, B2 => 
                           n3417, ZN => n13433);
   U4585 : INV_X1 port map( A => n13306, ZN => n12618);
   U4586 : AOI22_X1 port map( A1 => n4084, A2 => n3422, B1 => n2324, B2 => 
                           n3417, ZN => n13306);
   U4587 : INV_X1 port map( A => n13434, ZN => n12622);
   U4588 : AOI22_X1 port map( A1 => n4085, A2 => n3423, B1 => n2323, B2 => 
                           n3415, ZN => n13434);
   U4589 : INV_X1 port map( A => n13556, ZN => n12866);
   U4590 : AOI22_X1 port map( A1 => n3592, A2 => n4049, B1 => n2287, B2 => 
                           n3529, ZN => n13556);
   U4591 : INV_X1 port map( A => n13684, ZN => n12870);
   U4592 : AOI22_X1 port map( A1 => n3593, A2 => n4049, B1 => n2287, B2 => 
                           n3528, ZN => n13684);
   U4593 : INV_X1 port map( A => n13557, ZN => n12826);
   U4594 : AOI22_X1 port map( A1 => n4055, A2 => n3535, B1 => n2293, B2 => 
                           n3528, ZN => n13557);
   U4595 : INV_X1 port map( A => n13685, ZN => n12830);
   U4596 : AOI22_X1 port map( A1 => n4055, A2 => n3536, B1 => n2293, B2 => 
                           n3528, ZN => n13685);
   U4597 : INV_X1 port map( A => n13558, ZN => n12786);
   U4598 : AOI22_X1 port map( A1 => n4061, A2 => n3537, B1 => n2299, B2 => 
                           n3528, ZN => n13558);
   U4599 : INV_X1 port map( A => n13686, ZN => n12790);
   U4600 : AOI22_X1 port map( A1 => n4061, A2 => n3530, B1 => n2299, B2 => 
                           n3528, ZN => n13686);
   U4601 : INV_X1 port map( A => n13559, ZN => n12746);
   U4602 : AOI22_X1 port map( A1 => n4067, A2 => n3537, B1 => n2305, B2 => 
                           n3527, ZN => n13559);
   U4603 : INV_X1 port map( A => n13687, ZN => n12750);
   U4604 : AOI22_X1 port map( A1 => n4067, A2 => n3536, B1 => n2305, B2 => 
                           n3528, ZN => n13687);
   U4605 : INV_X1 port map( A => n13560, ZN => n12706);
   U4606 : AOI22_X1 port map( A1 => n4073, A2 => n3534, B1 => n2311, B2 => 
                           n3520, ZN => n13560);
   U4607 : INV_X1 port map( A => n13688, ZN => n12710);
   U4608 : AOI22_X1 port map( A1 => n4073, A2 => n3536, B1 => n2311, B2 => 
                           n3528, ZN => n13688);
   U4609 : INV_X1 port map( A => n13561, ZN => n12666);
   U4610 : AOI22_X1 port map( A1 => n4079, A2 => n3532, B1 => n2317, B2 => 
                           n3519, ZN => n13561);
   U4611 : INV_X1 port map( A => n13689, ZN => n12670);
   U4612 : AOI22_X1 port map( A1 => n4079, A2 => n3533, B1 => n2317, B2 => 
                           n3529, ZN => n13689);
   U4613 : INV_X1 port map( A => n13562, ZN => n12626);
   U4614 : AOI22_X1 port map( A1 => n4085, A2 => n3534, B1 => n2323, B2 => 
                           n3529, ZN => n13562);
   U4615 : INV_X1 port map( A => n13690, ZN => n12630);
   U4616 : AOI22_X1 port map( A1 => n4085, A2 => n3535, B1 => n2323, B2 => 
                           n3527, ZN => n13690);
   U4617 : INV_X1 port map( A => n13812, ZN => n12874);
   U4618 : AOI22_X1 port map( A1 => n3704, A2 => n4050, B1 => n2286, B2 => 
                           n3641, ZN => n13812);
   U4619 : INV_X1 port map( A => n13940, ZN => n12878);
   U4620 : AOI22_X1 port map( A1 => n3705, A2 => n4050, B1 => n2286, B2 => 
                           n3640, ZN => n13940);
   U4621 : INV_X1 port map( A => n13813, ZN => n12834);
   U4622 : AOI22_X1 port map( A1 => n4056, A2 => n3647, B1 => n2292, B2 => 
                           n3641, ZN => n13813);
   U4623 : INV_X1 port map( A => n13941, ZN => n12838);
   U4624 : AOI22_X1 port map( A1 => n4056, A2 => n3648, B1 => n2292, B2 => 
                           n3640, ZN => n13941);
   U4625 : INV_X1 port map( A => n13814, ZN => n12794);
   U4626 : AOI22_X1 port map( A1 => n4062, A2 => n3649, B1 => n2298, B2 => 
                           n3641, ZN => n13814);
   U4627 : INV_X1 port map( A => n13942, ZN => n12798);
   U4628 : AOI22_X1 port map( A1 => n4062, A2 => n3642, B1 => n2298, B2 => 
                           n3640, ZN => n13942);
   U4629 : INV_X1 port map( A => n13815, ZN => n12754);
   U4630 : AOI22_X1 port map( A1 => n4068, A2 => n3649, B1 => n2304, B2 => 
                           n3641, ZN => n13815);
   U4631 : INV_X1 port map( A => n13943, ZN => n12758);
   U4632 : AOI22_X1 port map( A1 => n4068, A2 => n3648, B1 => n2304, B2 => 
                           n3640, ZN => n13943);
   U4633 : INV_X1 port map( A => n13816, ZN => n12714);
   U4634 : AOI22_X1 port map( A1 => n4074, A2 => n3646, B1 => n2310, B2 => 
                           n3641, ZN => n13816);
   U4635 : INV_X1 port map( A => n13944, ZN => n12718);
   U4636 : AOI22_X1 port map( A1 => n4074, A2 => n3648, B1 => n2310, B2 => 
                           n3640, ZN => n13944);
   U4637 : INV_X1 port map( A => n13817, ZN => n12674);
   U4638 : AOI22_X1 port map( A1 => n4080, A2 => n3644, B1 => n2316, B2 => 
                           n3641, ZN => n13817);
   U4639 : INV_X1 port map( A => n13945, ZN => n12678);
   U4640 : AOI22_X1 port map( A1 => n4080, A2 => n3645, B1 => n2316, B2 => 
                           n3631, ZN => n13945);
   U4641 : INV_X1 port map( A => n13818, ZN => n12634);
   U4642 : AOI22_X1 port map( A1 => n4086, A2 => n3646, B1 => n2322, B2 => 
                           n3641, ZN => n13818);
   U4643 : INV_X1 port map( A => n13946, ZN => n12638);
   U4644 : AOI22_X1 port map( A1 => n4086, A2 => n3647, B1 => n2322, B2 => 
                           n3631, ZN => n13946);
   U4645 : INV_X1 port map( A => n14068, ZN => n12882);
   U4646 : AOI22_X1 port map( A1 => n3816, A2 => n4050, B1 => n2286, B2 => 
                           n3748, ZN => n14068);
   U4647 : INV_X1 port map( A => n14196, ZN => n12886);
   U4648 : AOI22_X1 port map( A1 => n3817, A2 => n4051, B1 => n2285, B2 => 
                           n3744, ZN => n14196);
   U4649 : INV_X1 port map( A => n14069, ZN => n12842);
   U4650 : AOI22_X1 port map( A1 => n4056, A2 => n3759, B1 => n2292, B2 => 
                           n3744, ZN => n14069);
   U4651 : INV_X1 port map( A => n14197, ZN => n12846);
   U4652 : AOI22_X1 port map( A1 => n4057, A2 => n3760, B1 => n2291, B2 => 
                           n3745, ZN => n14197);
   U4653 : INV_X1 port map( A => n14070, ZN => n12802);
   U4654 : AOI22_X1 port map( A1 => n4062, A2 => n3761, B1 => n2298, B2 => 
                           n3745, ZN => n14070);
   U4655 : INV_X1 port map( A => n14198, ZN => n12806);
   U4656 : AOI22_X1 port map( A1 => n4063, A2 => n3754, B1 => n2297, B2 => 
                           n3747, ZN => n14198);
   U4657 : INV_X1 port map( A => n14071, ZN => n12762);
   U4658 : AOI22_X1 port map( A1 => n4068, A2 => n3761, B1 => n2304, B2 => 
                           n3749, ZN => n14071);
   U4659 : INV_X1 port map( A => n14199, ZN => n12766);
   U4660 : AOI22_X1 port map( A1 => n4069, A2 => n3760, B1 => n2303, B2 => 
                           n3748, ZN => n14199);
   U4661 : INV_X1 port map( A => n14072, ZN => n12722);
   U4662 : AOI22_X1 port map( A1 => n4074, A2 => n3758, B1 => n2310, B2 => 
                           n3748, ZN => n14072);
   U4663 : INV_X1 port map( A => n14200, ZN => n12726);
   U4664 : AOI22_X1 port map( A1 => n4075, A2 => n3760, B1 => n2309, B2 => 
                           n3749, ZN => n14200);
   U4665 : INV_X1 port map( A => n14073, ZN => n12682);
   U4666 : AOI22_X1 port map( A1 => n4080, A2 => n3756, B1 => n2316, B2 => 
                           n3750, ZN => n14073);
   U4667 : INV_X1 port map( A => n14201, ZN => n12686);
   U4668 : AOI22_X1 port map( A1 => n4081, A2 => n3757, B1 => n2315, B2 => 
                           n3752, ZN => n14201);
   U4669 : INV_X1 port map( A => n14074, ZN => n12642);
   U4670 : AOI22_X1 port map( A1 => n4086, A2 => n3758, B1 => n2322, B2 => 
                           n3747, ZN => n14074);
   U4671 : INV_X1 port map( A => n14202, ZN => n12646);
   U4672 : AOI22_X1 port map( A1 => n4087, A2 => n3759, B1 => n2321, B2 => 
                           n3752, ZN => n14202);
   U4673 : INV_X1 port map( A => n13044, ZN => n12850);
   U4674 : AOI22_X1 port map( A1 => n3368, A2 => n4048, B1 => n2288, B2 => 
                           n3304, ZN => n13044);
   U4675 : INV_X1 port map( A => n13172, ZN => n12854);
   U4676 : AOI22_X1 port map( A1 => n3368, A2 => n4048, B1 => n2288, B2 => 
                           n3305, ZN => n13172);
   U4677 : INV_X1 port map( A => n13045, ZN => n12810);
   U4678 : AOI22_X1 port map( A1 => n4054, A2 => n3317, B1 => n2294, B2 => 
                           n3295, ZN => n13045);
   U4679 : INV_X1 port map( A => n13173, ZN => n12814);
   U4680 : AOI22_X1 port map( A1 => n4054, A2 => n3316, B1 => n2294, B2 => 
                           n3305, ZN => n13173);
   U4681 : INV_X1 port map( A => n13046, ZN => n12770);
   U4682 : AOI22_X1 port map( A1 => n4060, A2 => n3317, B1 => n2300, B2 => 
                           n3304, ZN => n13046);
   U4683 : INV_X1 port map( A => n13174, ZN => n12774);
   U4684 : AOI22_X1 port map( A1 => n4060, A2 => n3308, B1 => n2300, B2 => 
                           n3305, ZN => n13174);
   U4685 : INV_X1 port map( A => n13047, ZN => n12730);
   U4686 : AOI22_X1 port map( A1 => n4066, A2 => n3314, B1 => n2306, B2 => 
                           n3303, ZN => n13047);
   U4687 : INV_X1 port map( A => n13175, ZN => n12734);
   U4688 : AOI22_X1 port map( A1 => n4066, A2 => n3314, B1 => n2306, B2 => 
                           n3304, ZN => n13175);
   U4689 : INV_X1 port map( A => n13048, ZN => n12690);
   U4690 : AOI22_X1 port map( A1 => n4072, A2 => n3317, B1 => n2312, B2 => 
                           n3304, ZN => n13048);
   U4691 : INV_X1 port map( A => n13176, ZN => n12694);
   U4692 : AOI22_X1 port map( A1 => n4072, A2 => n3316, B1 => n2312, B2 => 
                           n3304, ZN => n13176);
   U4693 : INV_X1 port map( A => n13049, ZN => n12650);
   U4694 : AOI22_X1 port map( A1 => n4078, A2 => n3317, B1 => n2318, B2 => 
                           n3305, ZN => n13049);
   U4695 : INV_X1 port map( A => n13177, ZN => n12654);
   U4696 : AOI22_X1 port map( A1 => n4078, A2 => n3309, B1 => n2318, B2 => 
                           n3304, ZN => n13177);
   U4697 : INV_X1 port map( A => n13050, ZN => n12610);
   U4698 : AOI22_X1 port map( A1 => n4084, A2 => n3314, B1 => n2324, B2 => 
                           n3304, ZN => n13050);
   U4699 : INV_X1 port map( A => n13178, ZN => n12614);
   U4700 : AOI22_X1 port map( A1 => n4084, A2 => n3314, B1 => n2324, B2 => 
                           n3304, ZN => n13178);
   U4701 : INV_X1 port map( A => n13268, ZN => n12857);
   U4702 : AOI22_X1 port map( A1 => n3480, A2 => n4048, B1 => n2288, B2 => 
                           n3416, ZN => n13268);
   U4703 : INV_X1 port map( A => n13396, ZN => n12861);
   U4704 : AOI22_X1 port map( A1 => n3480, A2 => n4049, B1 => n2287, B2 => 
                           n3417, ZN => n13396);
   U4705 : INV_X1 port map( A => n13269, ZN => n12817);
   U4706 : AOI22_X1 port map( A1 => n4054, A2 => n3429, B1 => n2294, B2 => 
                           n3416, ZN => n13269);
   U4707 : INV_X1 port map( A => n13397, ZN => n12821);
   U4708 : AOI22_X1 port map( A1 => n4055, A2 => n3428, B1 => n2293, B2 => 
                           n3417, ZN => n13397);
   U4709 : INV_X1 port map( A => n13270, ZN => n12777);
   U4710 : AOI22_X1 port map( A1 => n4060, A2 => n3429, B1 => n2300, B2 => 
                           n3416, ZN => n13270);
   U4711 : INV_X1 port map( A => n13398, ZN => n12781);
   U4712 : AOI22_X1 port map( A1 => n4061, A2 => n3420, B1 => n2299, B2 => 
                           n3416, ZN => n13398);
   U4713 : INV_X1 port map( A => n13271, ZN => n12737);
   U4714 : AOI22_X1 port map( A1 => n4066, A2 => n3426, B1 => n2306, B2 => 
                           n3416, ZN => n13271);
   U4715 : INV_X1 port map( A => n13399, ZN => n12741);
   U4716 : AOI22_X1 port map( A1 => n4067, A2 => n3426, B1 => n2305, B2 => 
                           n3417, ZN => n13399);
   U4717 : INV_X1 port map( A => n13272, ZN => n12697);
   U4718 : AOI22_X1 port map( A1 => n4072, A2 => n3429, B1 => n2312, B2 => 
                           n3416, ZN => n13272);
   U4719 : INV_X1 port map( A => n13400, ZN => n12701);
   U4720 : AOI22_X1 port map( A1 => n4073, A2 => n3428, B1 => n2311, B2 => 
                           n3415, ZN => n13400);
   U4721 : INV_X1 port map( A => n13273, ZN => n12657);
   U4722 : AOI22_X1 port map( A1 => n4078, A2 => n3429, B1 => n2318, B2 => 
                           n3416, ZN => n13273);
   U4723 : INV_X1 port map( A => n13401, ZN => n12661);
   U4724 : AOI22_X1 port map( A1 => n4079, A2 => n3421, B1 => n2317, B2 => 
                           n3407, ZN => n13401);
   U4725 : INV_X1 port map( A => n13274, ZN => n12617);
   U4726 : AOI22_X1 port map( A1 => n4084, A2 => n3426, B1 => n2324, B2 => 
                           n3416, ZN => n13274);
   U4727 : INV_X1 port map( A => n13402, ZN => n12621);
   U4728 : AOI22_X1 port map( A1 => n4085, A2 => n3426, B1 => n2323, B2 => 
                           n3408, ZN => n13402);
   U4729 : INV_X1 port map( A => n13524, ZN => n12865);
   U4730 : AOI22_X1 port map( A1 => n3592, A2 => n4049, B1 => n2287, B2 => 
                           n3528, ZN => n13524);
   U4731 : INV_X1 port map( A => n13652, ZN => n12869);
   U4732 : AOI22_X1 port map( A1 => n3592, A2 => n4049, B1 => n2287, B2 => 
                           n3529, ZN => n13652);
   U4733 : INV_X1 port map( A => n13525, ZN => n12825);
   U4734 : AOI22_X1 port map( A1 => n4055, A2 => n3541, B1 => n2293, B2 => 
                           n3528, ZN => n13525);
   U4735 : INV_X1 port map( A => n13653, ZN => n12829);
   U4736 : AOI22_X1 port map( A1 => n4055, A2 => n3540, B1 => n2293, B2 => 
                           n3529, ZN => n13653);
   U4737 : INV_X1 port map( A => n13526, ZN => n12785);
   U4738 : AOI22_X1 port map( A1 => n4061, A2 => n3541, B1 => n2299, B2 => 
                           n3528, ZN => n13526);
   U4739 : INV_X1 port map( A => n13654, ZN => n12789);
   U4740 : AOI22_X1 port map( A1 => n4061, A2 => n3532, B1 => n2299, B2 => 
                           n3528, ZN => n13654);
   U4741 : INV_X1 port map( A => n13527, ZN => n12745);
   U4742 : AOI22_X1 port map( A1 => n4067, A2 => n3538, B1 => n2305, B2 => 
                           n3528, ZN => n13527);
   U4743 : INV_X1 port map( A => n13655, ZN => n12749);
   U4744 : AOI22_X1 port map( A1 => n4067, A2 => n3538, B1 => n2305, B2 => 
                           n3529, ZN => n13655);
   U4745 : INV_X1 port map( A => n13528, ZN => n12705);
   U4746 : AOI22_X1 port map( A1 => n4073, A2 => n3541, B1 => n2311, B2 => 
                           n3528, ZN => n13528);
   U4747 : INV_X1 port map( A => n13656, ZN => n12709);
   U4748 : AOI22_X1 port map( A1 => n4073, A2 => n3540, B1 => n2311, B2 => 
                           n3527, ZN => n13656);
   U4749 : INV_X1 port map( A => n13529, ZN => n12665);
   U4750 : AOI22_X1 port map( A1 => n4079, A2 => n3541, B1 => n2317, B2 => 
                           n3528, ZN => n13529);
   U4751 : INV_X1 port map( A => n13657, ZN => n12669);
   U4752 : AOI22_X1 port map( A1 => n4079, A2 => n3533, B1 => n2317, B2 => 
                           n3520, ZN => n13657);
   U4753 : INV_X1 port map( A => n13530, ZN => n12625);
   U4754 : AOI22_X1 port map( A1 => n4085, A2 => n3538, B1 => n2323, B2 => 
                           n3528, ZN => n13530);
   U4755 : INV_X1 port map( A => n13658, ZN => n12629);
   U4756 : AOI22_X1 port map( A1 => n4085, A2 => n3538, B1 => n2323, B2 => 
                           n3519, ZN => n13658);
   U4757 : INV_X1 port map( A => n13780, ZN => n12873);
   U4758 : AOI22_X1 port map( A1 => n3704, A2 => n4050, B1 => n2286, B2 => 
                           n3640, ZN => n13780);
   U4759 : INV_X1 port map( A => n13908, ZN => n12877);
   U4760 : AOI22_X1 port map( A1 => n3704, A2 => n4050, B1 => n2286, B2 => 
                           n3638, ZN => n13908);
   U4761 : INV_X1 port map( A => n13781, ZN => n12833);
   U4762 : AOI22_X1 port map( A1 => n4056, A2 => n3653, B1 => n2292, B2 => 
                           n3640, ZN => n13781);
   U4763 : INV_X1 port map( A => n13909, ZN => n12837);
   U4764 : AOI22_X1 port map( A1 => n4056, A2 => n3652, B1 => n2292, B2 => 
                           n3636, ZN => n13909);
   U4765 : INV_X1 port map( A => n13782, ZN => n12793);
   U4766 : AOI22_X1 port map( A1 => n4062, A2 => n3653, B1 => n2298, B2 => 
                           n3640, ZN => n13782);
   U4767 : INV_X1 port map( A => n13910, ZN => n12797);
   U4768 : AOI22_X1 port map( A1 => n4062, A2 => n3644, B1 => n2298, B2 => 
                           n3641, ZN => n13910);
   U4769 : INV_X1 port map( A => n13783, ZN => n12753);
   U4770 : AOI22_X1 port map( A1 => n4068, A2 => n3650, B1 => n2304, B2 => 
                           n3640, ZN => n13783);
   U4771 : INV_X1 port map( A => n13911, ZN => n12757);
   U4772 : AOI22_X1 port map( A1 => n4068, A2 => n3650, B1 => n2304, B2 => 
                           n3635, ZN => n13911);
   U4773 : INV_X1 port map( A => n13784, ZN => n12713);
   U4774 : AOI22_X1 port map( A1 => n4074, A2 => n3653, B1 => n2310, B2 => 
                           n3640, ZN => n13784);
   U4775 : INV_X1 port map( A => n13912, ZN => n12717);
   U4776 : AOI22_X1 port map( A1 => n4074, A2 => n3652, B1 => n2310, B2 => 
                           n3641, ZN => n13912);
   U4777 : INV_X1 port map( A => n13785, ZN => n12673);
   U4778 : AOI22_X1 port map( A1 => n4080, A2 => n3653, B1 => n2316, B2 => 
                           n3640, ZN => n13785);
   U4779 : INV_X1 port map( A => n13913, ZN => n12677);
   U4780 : AOI22_X1 port map( A1 => n4080, A2 => n3645, B1 => n2316, B2 => 
                           n3641, ZN => n13913);
   U4781 : INV_X1 port map( A => n13786, ZN => n12633);
   U4782 : AOI22_X1 port map( A1 => n4086, A2 => n3650, B1 => n2322, B2 => 
                           n3641, ZN => n13786);
   U4783 : INV_X1 port map( A => n13914, ZN => n12637);
   U4784 : AOI22_X1 port map( A1 => n4086, A2 => n3650, B1 => n2322, B2 => 
                           n3641, ZN => n13914);
   U4785 : INV_X1 port map( A => n14036, ZN => n12881);
   U4786 : AOI22_X1 port map( A1 => n3816, A2 => n4050, B1 => n2286, B2 => 
                           n3747, ZN => n14036);
   U4787 : INV_X1 port map( A => n14164, ZN => n12885);
   U4788 : AOI22_X1 port map( A1 => n3816, A2 => n4051, B1 => n2285, B2 => 
                           n3753, ZN => n14164);
   U4789 : INV_X1 port map( A => n14037, ZN => n12841);
   U4790 : AOI22_X1 port map( A1 => n4056, A2 => n3765, B1 => n2292, B2 => 
                           n3748, ZN => n14037);
   U4791 : INV_X1 port map( A => n14165, ZN => n12845);
   U4792 : AOI22_X1 port map( A1 => n4057, A2 => n3764, B1 => n2291, B2 => 
                           n3753, ZN => n14165);
   U4793 : INV_X1 port map( A => n14038, ZN => n12801);
   U4794 : AOI22_X1 port map( A1 => n4062, A2 => n3765, B1 => n2298, B2 => 
                           n3749, ZN => n14038);
   U4795 : INV_X1 port map( A => n14166, ZN => n12805);
   U4796 : AOI22_X1 port map( A1 => n4063, A2 => n3756, B1 => n2297, B2 => 
                           n3746, ZN => n14166);
   U4797 : INV_X1 port map( A => n14039, ZN => n12761);
   U4798 : AOI22_X1 port map( A1 => n4068, A2 => n3762, B1 => n2304, B2 => 
                           n3750, ZN => n14039);
   U4799 : INV_X1 port map( A => n14167, ZN => n12765);
   U4800 : AOI22_X1 port map( A1 => n4069, A2 => n3762, B1 => n2303, B2 => 
                           n3753, ZN => n14167);
   U4801 : INV_X1 port map( A => n14040, ZN => n12721);
   U4802 : AOI22_X1 port map( A1 => n4074, A2 => n3765, B1 => n2310, B2 => 
                           n3746, ZN => n14040);
   U4803 : INV_X1 port map( A => n14168, ZN => n12725);
   U4804 : AOI22_X1 port map( A1 => n4075, A2 => n3764, B1 => n2309, B2 => 
                           n3746, ZN => n14168);
   U4805 : INV_X1 port map( A => n14041, ZN => n12681);
   U4806 : AOI22_X1 port map( A1 => n4080, A2 => n3765, B1 => n2316, B2 => 
                           n3746, ZN => n14041);
   U4807 : INV_X1 port map( A => n14169, ZN => n12685);
   U4808 : AOI22_X1 port map( A1 => n4081, A2 => n3757, B1 => n2315, B2 => 
                           n3744, ZN => n14169);
   U4809 : INV_X1 port map( A => n14042, ZN => n12641);
   U4810 : AOI22_X1 port map( A1 => n4086, A2 => n3762, B1 => n2322, B2 => 
                           n3747, ZN => n14042);
   U4811 : INV_X1 port map( A => n14170, ZN => n12645);
   U4812 : AOI22_X1 port map( A1 => n4087, A2 => n3762, B1 => n2321, B2 => 
                           n3745, ZN => n14170);
   U4813 : INV_X1 port map( A => n13364, ZN => n12860);
   U4814 : AOI22_X1 port map( A1 => n3480, A2 => n4049, B1 => n2288, B2 => 
                           n3415, ZN => n13364);
   U4815 : INV_X1 port map( A => n13620, ZN => n12868);
   U4816 : AOI22_X1 port map( A1 => n3592, A2 => n4049, B1 => n2287, B2 => 
                           n3527, ZN => n13620);
   U4817 : INV_X1 port map( A => n13876, ZN => n12876);
   U4818 : AOI22_X1 port map( A1 => n3704, A2 => n4050, B1 => n2286, B2 => 
                           n3639, ZN => n13876);
   U4819 : INV_X1 port map( A => n14132, ZN => n12884);
   U4820 : AOI22_X1 port map( A1 => n3816, A2 => n4051, B1 => n2285, B2 => 
                           n3751, ZN => n14132);
   U4821 : INV_X1 port map( A => n13012, ZN => n12849);
   U4822 : AOI22_X1 port map( A1 => n3369, A2 => n4048, B1 => n2288, B2 => 
                           n3303, ZN => n13012);
   U4823 : INV_X1 port map( A => n13140, ZN => n12853);
   U4824 : AOI22_X1 port map( A1 => n3368, A2 => n4048, B1 => n2288, B2 => 
                           n3303, ZN => n13140);
   U4825 : INV_X1 port map( A => n13013, ZN => n12809);
   U4826 : AOI22_X1 port map( A1 => n4054, A2 => n3315, B1 => n2294, B2 => 
                           n3303, ZN => n13013);
   U4827 : INV_X1 port map( A => n13141, ZN => n12813);
   U4828 : AOI22_X1 port map( A1 => n4054, A2 => n3309, B1 => n2294, B2 => 
                           n3304, ZN => n13141);
   U4829 : INV_X1 port map( A => n13014, ZN => n12769);
   U4830 : AOI22_X1 port map( A1 => n4060, A2 => n3308, B1 => n2300, B2 => 
                           n3303, ZN => n13014);
   U4831 : INV_X1 port map( A => n13015, ZN => n12729);
   U4832 : AOI22_X1 port map( A1 => n4066, A2 => n3313, B1 => n2306, B2 => 
                           n3303, ZN => n13015);
   U4833 : INV_X1 port map( A => n13016, ZN => n12689);
   U4834 : AOI22_X1 port map( A1 => n4072, A2 => n3315, B1 => n2312, B2 => 
                           n3303, ZN => n13016);
   U4835 : INV_X1 port map( A => n13017, ZN => n12649);
   U4836 : AOI22_X1 port map( A1 => n4078, A2 => n3316, B1 => n2318, B2 => 
                           n3303, ZN => n13017);
   U4837 : INV_X1 port map( A => n13145, ZN => n12653);
   U4838 : AOI22_X1 port map( A1 => n4078, A2 => n3312, B1 => n2318, B2 => 
                           n3305, ZN => n13145);
   U4839 : INV_X1 port map( A => n13018, ZN => n12609);
   U4840 : AOI22_X1 port map( A1 => n4084, A2 => n3313, B1 => n2324, B2 => 
                           n3303, ZN => n13018);
   U4841 : INV_X1 port map( A => n13236, ZN => n12856);
   U4842 : AOI22_X1 port map( A1 => n3481, A2 => n4048, B1 => n2288, B2 => 
                           n3407, ZN => n13236);
   U4843 : INV_X1 port map( A => n13237, ZN => n12816);
   U4844 : AOI22_X1 port map( A1 => n4054, A2 => n3427, B1 => n2294, B2 => 
                           n3408, ZN => n13237);
   U4845 : INV_X1 port map( A => n13238, ZN => n12776);
   U4846 : AOI22_X1 port map( A1 => n4060, A2 => n3420, B1 => n2300, B2 => 
                           n3417, ZN => n13238);
   U4847 : INV_X1 port map( A => n13239, ZN => n12736);
   U4848 : AOI22_X1 port map( A1 => n4066, A2 => n3425, B1 => n2306, B2 => 
                           n3415, ZN => n13239);
   U4849 : INV_X1 port map( A => n13240, ZN => n12696);
   U4850 : AOI22_X1 port map( A1 => n4072, A2 => n3427, B1 => n2312, B2 => 
                           n3416, ZN => n13240);
   U4851 : INV_X1 port map( A => n13241, ZN => n12656);
   U4852 : AOI22_X1 port map( A1 => n4078, A2 => n3428, B1 => n2318, B2 => 
                           n3407, ZN => n13241);
   U4853 : INV_X1 port map( A => n13369, ZN => n12660);
   U4854 : AOI22_X1 port map( A1 => n4079, A2 => n3424, B1 => n2318, B2 => 
                           n3417, ZN => n13369);
   U4855 : INV_X1 port map( A => n13242, ZN => n12616);
   U4856 : AOI22_X1 port map( A1 => n4084, A2 => n3425, B1 => n2324, B2 => 
                           n3408, ZN => n13242);
   U4857 : INV_X1 port map( A => n13370, ZN => n12620);
   U4858 : AOI22_X1 port map( A1 => n4085, A2 => n3428, B1 => n2324, B2 => 
                           n3417, ZN => n13370);
   U4859 : INV_X1 port map( A => n13492, ZN => n12864);
   U4860 : AOI22_X1 port map( A1 => n3593, A2 => n4049, B1 => n2287, B2 => 
                           n3520, ZN => n13492);
   U4861 : INV_X1 port map( A => n13493, ZN => n12824);
   U4862 : AOI22_X1 port map( A1 => n4055, A2 => n3539, B1 => n2293, B2 => 
                           n3519, ZN => n13493);
   U4863 : INV_X1 port map( A => n13494, ZN => n12784);
   U4864 : AOI22_X1 port map( A1 => n4061, A2 => n3532, B1 => n2299, B2 => 
                           n3529, ZN => n13494);
   U4865 : INV_X1 port map( A => n13495, ZN => n12744);
   U4866 : AOI22_X1 port map( A1 => n4067, A2 => n3537, B1 => n2305, B2 => 
                           n3527, ZN => n13495);
   U4867 : INV_X1 port map( A => n13496, ZN => n12704);
   U4868 : AOI22_X1 port map( A1 => n4073, A2 => n3539, B1 => n2311, B2 => 
                           n3528, ZN => n13496);
   U4869 : INV_X1 port map( A => n13497, ZN => n12664);
   U4870 : AOI22_X1 port map( A1 => n4079, A2 => n3540, B1 => n2317, B2 => 
                           n3520, ZN => n13497);
   U4871 : INV_X1 port map( A => n13625, ZN => n12668);
   U4872 : AOI22_X1 port map( A1 => n4079, A2 => n3536, B1 => n2317, B2 => 
                           n3529, ZN => n13625);
   U4873 : INV_X1 port map( A => n13498, ZN => n12624);
   U4874 : AOI22_X1 port map( A1 => n4085, A2 => n3537, B1 => n2323, B2 => 
                           n3519, ZN => n13498);
   U4875 : INV_X1 port map( A => n13626, ZN => n12628);
   U4876 : AOI22_X1 port map( A1 => n4085, A2 => n3540, B1 => n2323, B2 => 
                           n3529, ZN => n13626);
   U4877 : INV_X1 port map( A => n13748, ZN => n12872);
   U4878 : AOI22_X1 port map( A1 => n3705, A2 => n4050, B1 => n2286, B2 => 
                           n3640, ZN => n13748);
   U4879 : INV_X1 port map( A => n13749, ZN => n12832);
   U4880 : AOI22_X1 port map( A1 => n4056, A2 => n3651, B1 => n2292, B2 => 
                           n3639, ZN => n13749);
   U4881 : INV_X1 port map( A => n13750, ZN => n12792);
   U4882 : AOI22_X1 port map( A1 => n4062, A2 => n3644, B1 => n2298, B2 => 
                           n3631, ZN => n13750);
   U4883 : INV_X1 port map( A => n13751, ZN => n12752);
   U4884 : AOI22_X1 port map( A1 => n4068, A2 => n3649, B1 => n2304, B2 => 
                           n3639, ZN => n13751);
   U4885 : INV_X1 port map( A => n13752, ZN => n12712);
   U4886 : AOI22_X1 port map( A1 => n4074, A2 => n3651, B1 => n2310, B2 => 
                           n3641, ZN => n13752);
   U4887 : INV_X1 port map( A => n13753, ZN => n12672);
   U4888 : AOI22_X1 port map( A1 => n4080, A2 => n3652, B1 => n2316, B2 => 
                           n3640, ZN => n13753);
   U4889 : INV_X1 port map( A => n13881, ZN => n12676);
   U4890 : AOI22_X1 port map( A1 => n4080, A2 => n3648, B1 => n2316, B2 => 
                           n3631, ZN => n13881);
   U4891 : INV_X1 port map( A => n13754, ZN => n12632);
   U4892 : AOI22_X1 port map( A1 => n4086, A2 => n3649, B1 => n2322, B2 => 
                           n3639, ZN => n13754);
   U4893 : INV_X1 port map( A => n13882, ZN => n12636);
   U4894 : AOI22_X1 port map( A1 => n4086, A2 => n3652, B1 => n2322, B2 => 
                           n3641, ZN => n13882);
   U4895 : INV_X1 port map( A => n14004, ZN => n12880);
   U4896 : AOI22_X1 port map( A1 => n3817, A2 => n4050, B1 => n2286, B2 => 
                           n3752, ZN => n14004);
   U4897 : INV_X1 port map( A => n14005, ZN => n12840);
   U4898 : AOI22_X1 port map( A1 => n4056, A2 => n3763, B1 => n2292, B2 => 
                           n3752, ZN => n14005);
   U4899 : INV_X1 port map( A => n14006, ZN => n12800);
   U4900 : AOI22_X1 port map( A1 => n4062, A2 => n3756, B1 => n2298, B2 => 
                           n3752, ZN => n14006);
   U4901 : INV_X1 port map( A => n14007, ZN => n12760);
   U4902 : AOI22_X1 port map( A1 => n4068, A2 => n3761, B1 => n2304, B2 => 
                           n3752, ZN => n14007);
   U4903 : INV_X1 port map( A => n14008, ZN => n12720);
   U4904 : AOI22_X1 port map( A1 => n4074, A2 => n3763, B1 => n2310, B2 => 
                           n3752, ZN => n14008);
   U4905 : INV_X1 port map( A => n14009, ZN => n12680);
   U4906 : AOI22_X1 port map( A1 => n4080, A2 => n3764, B1 => n2316, B2 => 
                           n3752, ZN => n14009);
   U4907 : INV_X1 port map( A => n14137, ZN => n12684);
   U4908 : AOI22_X1 port map( A1 => n4081, A2 => n3760, B1 => n2315, B2 => 
                           n3753, ZN => n14137);
   U4909 : INV_X1 port map( A => n14010, ZN => n12640);
   U4910 : AOI22_X1 port map( A1 => n4086, A2 => n3761, B1 => n2322, B2 => 
                           n3752, ZN => n14010);
   U4911 : INV_X1 port map( A => n14138, ZN => n12644);
   U4912 : AOI22_X1 port map( A1 => n4087, A2 => n3764, B1 => n2321, B2 => 
                           n3753, ZN => n14138);
   U4913 : INV_X1 port map( A => n13365, ZN => n12820);
   U4914 : AOI22_X1 port map( A1 => n4055, A2 => n3421, B1 => n2294, B2 => 
                           n3415, ZN => n13365);
   U4915 : INV_X1 port map( A => n13366, ZN => n12780);
   U4916 : AOI22_X1 port map( A1 => n4061, A2 => n3423, B1 => n2300, B2 => 
                           n3407, ZN => n13366);
   U4917 : INV_X1 port map( A => n13367, ZN => n12740);
   U4918 : AOI22_X1 port map( A1 => n4067, A2 => n3427, B1 => n2306, B2 => 
                           n3408, ZN => n13367);
   U4919 : INV_X1 port map( A => n13368, ZN => n12700);
   U4920 : AOI22_X1 port map( A1 => n4073, A2 => n3427, B1 => n2312, B2 => 
                           n3417, ZN => n13368);
   U4921 : INV_X1 port map( A => n13621, ZN => n12828);
   U4922 : AOI22_X1 port map( A1 => n4055, A2 => n3533, B1 => n2293, B2 => 
                           n3527, ZN => n13621);
   U4923 : INV_X1 port map( A => n13622, ZN => n12788);
   U4924 : AOI22_X1 port map( A1 => n4061, A2 => n3535, B1 => n2299, B2 => 
                           n3520, ZN => n13622);
   U4925 : INV_X1 port map( A => n13623, ZN => n12748);
   U4926 : AOI22_X1 port map( A1 => n4067, A2 => n3539, B1 => n2305, B2 => 
                           n3519, ZN => n13623);
   U4927 : INV_X1 port map( A => n13624, ZN => n12708);
   U4928 : AOI22_X1 port map( A1 => n4073, A2 => n3539, B1 => n2311, B2 => 
                           n3529, ZN => n13624);
   U4929 : INV_X1 port map( A => n13877, ZN => n12836);
   U4930 : AOI22_X1 port map( A1 => n4056, A2 => n3645, B1 => n2292, B2 => 
                           n3633, ZN => n13877);
   U4931 : INV_X1 port map( A => n13878, ZN => n12796);
   U4932 : AOI22_X1 port map( A1 => n4062, A2 => n3647, B1 => n2298, B2 => 
                           n3634, ZN => n13878);
   U4933 : INV_X1 port map( A => n13879, ZN => n12756);
   U4934 : AOI22_X1 port map( A1 => n4068, A2 => n3651, B1 => n2304, B2 => 
                           n3632, ZN => n13879);
   U4935 : INV_X1 port map( A => n13880, ZN => n12716);
   U4936 : AOI22_X1 port map( A1 => n4074, A2 => n3651, B1 => n2310, B2 => 
                           n3637, ZN => n13880);
   U4937 : INV_X1 port map( A => n14133, ZN => n12844);
   U4938 : AOI22_X1 port map( A1 => n4057, A2 => n3757, B1 => n2291, B2 => 
                           n3749, ZN => n14133);
   U4939 : INV_X1 port map( A => n14134, ZN => n12804);
   U4940 : AOI22_X1 port map( A1 => n4063, A2 => n3759, B1 => n2297, B2 => 
                           n3750, ZN => n14134);
   U4941 : INV_X1 port map( A => n14135, ZN => n12764);
   U4942 : AOI22_X1 port map( A1 => n4069, A2 => n3763, B1 => n2303, B2 => 
                           n3749, ZN => n14135);
   U4943 : INV_X1 port map( A => n14136, ZN => n12724);
   U4944 : AOI22_X1 port map( A1 => n4075, A2 => n3763, B1 => n2309, B2 => 
                           n3748, ZN => n14136);
   U4945 : INV_X1 port map( A => n13142, ZN => n12773);
   U4946 : AOI22_X1 port map( A1 => n4060, A2 => n3311, B1 => n2300, B2 => 
                           n3301, ZN => n13142);
   U4947 : INV_X1 port map( A => n13143, ZN => n12733);
   U4948 : AOI22_X1 port map( A1 => n4066, A2 => n3315, B1 => n2306, B2 => 
                           n3300, ZN => n13143);
   U4949 : INV_X1 port map( A => n13144, ZN => n12693);
   U4950 : AOI22_X1 port map( A1 => n4072, A2 => n3315, B1 => n2312, B2 => 
                           n3301, ZN => n13144);
   U4951 : INV_X1 port map( A => n13146, ZN => n12613);
   U4952 : AOI22_X1 port map( A1 => n4084, A2 => n3316, B1 => n2324, B2 => 
                           n3301, ZN => n13146);
   U4953 : INV_X1 port map( A => n12981, ZN => n12808);
   U4954 : AOI22_X1 port map( A1 => n4054, A2 => n3310, B1 => n2291, B2 => 
                           n3297, ZN => n12981);
   U4955 : INV_X1 port map( A => n12983, ZN => n12728);
   U4956 : AOI22_X1 port map( A1 => n4066, A2 => n3310, B1 => n2303, B2 => 
                           n3298, ZN => n12983);
   U4957 : INV_X1 port map( A => n12986, ZN => n12608);
   U4958 : AOI22_X1 port map( A1 => n4084, A2 => n3306, B1 => n2321, B2 => 
                           n3296, ZN => n12986);
   U4959 : INV_X1 port map( A => n13206, ZN => n12775);
   U4960 : AOI22_X1 port map( A1 => n4060, A2 => n3420, B1 => n2300, B2 => 
                           n3415, ZN => n13206);
   U4961 : INV_X1 port map( A => n13207, ZN => n12735);
   U4962 : AOI22_X1 port map( A1 => n4066, A2 => n3422, B1 => n2306, B2 => 
                           n3415, ZN => n13207);
   U4963 : INV_X1 port map( A => n13208, ZN => n12695);
   U4964 : AOI22_X1 port map( A1 => n4072, A2 => n3423, B1 => n2312, B2 => 
                           n3415, ZN => n13208);
   U4965 : INV_X1 port map( A => n13462, ZN => n12783);
   U4966 : AOI22_X1 port map( A1 => n4061, A2 => n3532, B1 => n2299, B2 => 
                           n3527, ZN => n13462);
   U4967 : INV_X1 port map( A => n13463, ZN => n12743);
   U4968 : AOI22_X1 port map( A1 => n4067, A2 => n3534, B1 => n2305, B2 => 
                           n3527, ZN => n13463);
   U4969 : INV_X1 port map( A => n13464, ZN => n12703);
   U4970 : AOI22_X1 port map( A1 => n4073, A2 => n3535, B1 => n2311, B2 => 
                           n3527, ZN => n13464);
   U4971 : INV_X1 port map( A => n13718, ZN => n12791);
   U4972 : AOI22_X1 port map( A1 => n4061, A2 => n3644, B1 => n2299, B2 => 
                           n3639, ZN => n13718);
   U4973 : INV_X1 port map( A => n13719, ZN => n12751);
   U4974 : AOI22_X1 port map( A1 => n4067, A2 => n3646, B1 => n2305, B2 => 
                           n3639, ZN => n13719);
   U4975 : INV_X1 port map( A => n13720, ZN => n12711);
   U4976 : AOI22_X1 port map( A1 => n4073, A2 => n3647, B1 => n2311, B2 => 
                           n3639, ZN => n13720);
   U4977 : INV_X1 port map( A => n13974, ZN => n12799);
   U4978 : AOI22_X1 port map( A1 => n4062, A2 => n3756, B1 => n2298, B2 => 
                           n3751, ZN => n13974);
   U4979 : INV_X1 port map( A => n13975, ZN => n12759);
   U4980 : AOI22_X1 port map( A1 => n4068, A2 => n3758, B1 => n2304, B2 => 
                           n3751, ZN => n13975);
   U4981 : INV_X1 port map( A => n13976, ZN => n12719);
   U4982 : AOI22_X1 port map( A1 => n4074, A2 => n3759, B1 => n2310, B2 => 
                           n3751, ZN => n13976);
   U4983 : INV_X1 port map( A => n12980, ZN => n12848);
   U4984 : AOI22_X1 port map( A1 => n3369, A2 => n4048, B1 => n2285, B2 => 
                           n3295, ZN => n12980);
   U4985 : INV_X1 port map( A => n12982, ZN => n12768);
   U4986 : AOI22_X1 port map( A1 => n4060, A2 => n3308, B1 => n2297, B2 => 
                           n3303, ZN => n12982);
   U4987 : INV_X1 port map( A => n12984, ZN => n12688);
   U4988 : AOI22_X1 port map( A1 => n4072, A2 => n3311, B1 => n2309, B2 => 
                           n3303, ZN => n12984);
   U4989 : INV_X1 port map( A => n12985, ZN => n12648);
   U4990 : AOI22_X1 port map( A1 => n4078, A2 => n3309, B1 => n2315, B2 => 
                           n3303, ZN => n12985);
   U4991 : INV_X1 port map( A => n13204, ZN => n12855);
   U4992 : AOI22_X1 port map( A1 => n3481, A2 => n4048, B1 => n2288, B2 => 
                           n3416, ZN => n13204);
   U4993 : INV_X1 port map( A => n13205, ZN => n12815);
   U4994 : AOI22_X1 port map( A1 => n4054, A2 => n3422, B1 => n2294, B2 => 
                           n3407, ZN => n13205);
   U4995 : INV_X1 port map( A => n13209, ZN => n12655);
   U4996 : AOI22_X1 port map( A1 => n4078, A2 => n3421, B1 => n2318, B2 => 
                           n3408, ZN => n13209);
   U4997 : INV_X1 port map( A => n13210, ZN => n12615);
   U4998 : AOI22_X1 port map( A1 => n4084, A2 => n3418, B1 => n2324, B2 => 
                           n3417, ZN => n13210);
   U4999 : INV_X1 port map( A => n13460, ZN => n12863);
   U5000 : AOI22_X1 port map( A1 => n3593, A2 => n4049, B1 => n2287, B2 => 
                           n3528, ZN => n13460);
   U5001 : INV_X1 port map( A => n13461, ZN => n12823);
   U5002 : AOI22_X1 port map( A1 => n4055, A2 => n3534, B1 => n2293, B2 => 
                           n3520, ZN => n13461);
   U5003 : INV_X1 port map( A => n13465, ZN => n12663);
   U5004 : AOI22_X1 port map( A1 => n4079, A2 => n3533, B1 => n2317, B2 => 
                           n3519, ZN => n13465);
   U5005 : INV_X1 port map( A => n13466, ZN => n12623);
   U5006 : AOI22_X1 port map( A1 => n4085, A2 => n3530, B1 => n2323, B2 => 
                           n3529, ZN => n13466);
   U5007 : INV_X1 port map( A => n13716, ZN => n12871);
   U5008 : AOI22_X1 port map( A1 => n3705, A2 => n4049, B1 => n2287, B2 => 
                           n3640, ZN => n13716);
   U5009 : INV_X1 port map( A => n13717, ZN => n12831);
   U5010 : AOI22_X1 port map( A1 => n4055, A2 => n3646, B1 => n2293, B2 => 
                           n3641, ZN => n13717);
   U5011 : INV_X1 port map( A => n13721, ZN => n12671);
   U5012 : AOI22_X1 port map( A1 => n4079, A2 => n3645, B1 => n2317, B2 => 
                           n3640, ZN => n13721);
   U5013 : INV_X1 port map( A => n13722, ZN => n12631);
   U5014 : AOI22_X1 port map( A1 => n4085, A2 => n3642, B1 => n2323, B2 => 
                           n3639, ZN => n13722);
   U5015 : INV_X1 port map( A => n13972, ZN => n12879);
   U5016 : AOI22_X1 port map( A1 => n3817, A2 => n4050, B1 => n2286, B2 => 
                           n3750, ZN => n13972);
   U5017 : INV_X1 port map( A => n13973, ZN => n12839);
   U5018 : AOI22_X1 port map( A1 => n4056, A2 => n3758, B1 => n2292, B2 => 
                           n3752, ZN => n13973);
   U5019 : INV_X1 port map( A => n13977, ZN => n12679);
   U5020 : AOI22_X1 port map( A1 => n4080, A2 => n3757, B1 => n2316, B2 => 
                           n3752, ZN => n13977);
   U5021 : INV_X1 port map( A => n13978, ZN => n12639);
   U5022 : AOI22_X1 port map( A1 => n4086, A2 => n3754, B1 => n2322, B2 => 
                           n3752, ZN => n13978);
   U5023 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_3_0_port, Z => 
                           n3630);
   U5024 : INV_X1 port map( A => n13083, ZN => n12571);
   U5025 : AOI22_X1 port map( A1 => n2327, A2 => n3297, B1 => n3916, B2 => 
                           n3362, ZN => n13083);
   U5026 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n41, ZN => n12607);
   U5027 : AOI22_X1 port map( A1 => n2330, A2 => n3297, B1 => n3919, B2 => 
                           n3337, ZN => DataPath_RF_MUX_SELINPUT_8_n41);
   U5028 : INV_X1 port map( A => n13084, ZN => n12531);
   U5029 : AOI22_X1 port map( A1 => n2333, A2 => n3298, B1 => n3922, B2 => 
                           n3362, ZN => n13084);
   U5030 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n42, ZN => n12567);
   U5031 : AOI22_X1 port map( A1 => n2336, A2 => n3298, B1 => n3925, B2 => 
                           n3337, ZN => DataPath_RF_MUX_SELINPUT_8_n42);
   U5032 : INV_X1 port map( A => n13086, ZN => n12451);
   U5033 : AOI22_X1 port map( A1 => n2345, A2 => n3296, B1 => n3928, B2 => 
                           n3363, ZN => n13086);
   U5034 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n44, ZN => n12487);
   U5035 : AOI22_X1 port map( A1 => n2348, A2 => n3301, B1 => n3931, B2 => 
                           n3338, ZN => DataPath_RF_MUX_SELINPUT_8_n44);
   U5036 : INV_X1 port map( A => n13087, ZN => n12411);
   U5037 : AOI22_X1 port map( A1 => n2351, A2 => n3300, B1 => n3934, B2 => 
                           n3363, ZN => n13087);
   U5038 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n45, ZN => n12447);
   U5039 : AOI22_X1 port map( A1 => n2354, A2 => n3301, B1 => n3937, B2 => 
                           n3338, ZN => DataPath_RF_MUX_SELINPUT_8_n45);
   U5040 : INV_X1 port map( A => n13088, ZN => n12371);
   U5041 : AOI22_X1 port map( A1 => n2357, A2 => n3302, B1 => n3940, B2 => 
                           n3363, ZN => n13088);
   U5042 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n46, ZN => n12407);
   U5043 : AOI22_X1 port map( A1 => n2360, A2 => n3301, B1 => n3943, B2 => 
                           n3338, ZN => DataPath_RF_MUX_SELINPUT_8_n46);
   U5044 : INV_X1 port map( A => n13089, ZN => n12331);
   U5045 : AOI22_X1 port map( A1 => n2363, A2 => n3301, B1 => n3946, B2 => 
                           n3363, ZN => n13089);
   U5046 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n47, ZN => n12367);
   U5047 : AOI22_X1 port map( A1 => n2366, A2 => n3301, B1 => n3949, B2 => 
                           n3339, ZN => DataPath_RF_MUX_SELINPUT_8_n47);
   U5048 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n48, ZN => n12327);
   U5049 : AOI22_X1 port map( A1 => n2372, A2 => n3301, B1 => n3955, B2 => 
                           n3339, ZN => DataPath_RF_MUX_SELINPUT_8_n48);
   U5050 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n49, ZN => n12287);
   U5051 : AOI22_X1 port map( A1 => n2378, A2 => n3301, B1 => n3961, B2 => 
                           n3339, ZN => DataPath_RF_MUX_SELINPUT_8_n49);
   U5052 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n50, ZN => n12247);
   U5053 : AOI22_X1 port map( A1 => n2384, A2 => n3301, B1 => n3967, B2 => 
                           n3339, ZN => DataPath_RF_MUX_SELINPUT_8_n50);
   U5054 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n51, ZN => n12207);
   U5055 : AOI22_X1 port map( A1 => n2390, A2 => n3301, B1 => n3973, B2 => 
                           n3340, ZN => DataPath_RF_MUX_SELINPUT_8_n51);
   U5056 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n52, ZN => n12167);
   U5057 : AOI22_X1 port map( A1 => n2396, A2 => n3301, B1 => n3979, B2 => 
                           n3340, ZN => DataPath_RF_MUX_SELINPUT_8_n52);
   U5058 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n53, ZN => n12127);
   U5059 : AOI22_X1 port map( A1 => n2402, A2 => n3301, B1 => n3985, B2 => 
                           n3340, ZN => DataPath_RF_MUX_SELINPUT_8_n53);
   U5060 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n55, ZN => n12047);
   U5061 : AOI22_X1 port map( A1 => n2414, A2 => n3302, B1 => n3991, B2 => 
                           n3341, ZN => DataPath_RF_MUX_SELINPUT_8_n55);
   U5062 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n56, ZN => n12007);
   U5063 : AOI22_X1 port map( A1 => n2420, A2 => n3299, B1 => n3997, B2 => 
                           n3341, ZN => DataPath_RF_MUX_SELINPUT_8_n56);
   U5064 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n57, ZN => n11967);
   U5065 : AOI22_X1 port map( A1 => n2426, A2 => n3300, B1 => n4003, B2 => 
                           n3341, ZN => DataPath_RF_MUX_SELINPUT_8_n57);
   U5066 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n58, ZN => n11927);
   U5067 : AOI22_X1 port map( A1 => n2432, A2 => n3302, B1 => n4009, B2 => 
                           n3341, ZN => DataPath_RF_MUX_SELINPUT_8_n58);
   U5068 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n59, ZN => n11887);
   U5069 : AOI22_X1 port map( A1 => n2438, A2 => n3301, B1 => n4015, B2 => 
                           n3342, ZN => DataPath_RF_MUX_SELINPUT_8_n59);
   U5070 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n60, ZN => n11847);
   U5071 : AOI22_X1 port map( A1 => n2444, A2 => n3297, B1 => n4021, B2 => 
                           n3342, ZN => DataPath_RF_MUX_SELINPUT_8_n60);
   U5072 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n61, ZN => n11807);
   U5073 : AOI22_X1 port map( A1 => n2450, A2 => n3298, B1 => n4027, B2 => 
                           n3342, ZN => DataPath_RF_MUX_SELINPUT_8_n61);
   U5074 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n62, ZN => n11767);
   U5075 : AOI22_X1 port map( A1 => n2456, A2 => n3296, B1 => n4033, B2 => 
                           n3342, ZN => DataPath_RF_MUX_SELINPUT_8_n62);
   U5076 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n63, ZN => n11727);
   U5077 : AOI22_X1 port map( A1 => n2462, A2 => n3299, B1 => n4039, B2 => 
                           n3343, ZN => DataPath_RF_MUX_SELINPUT_8_n63);
   U5078 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n64, ZN => n11687);
   U5079 : AOI22_X1 port map( A1 => n2468, A2 => n3300, B1 => n4045, B2 => 
                           n3322, ZN => DataPath_RF_MUX_SELINPUT_8_n64);
   U5080 : INV_X1 port map( A => n13085, ZN => n12491);
   U5081 : AOI22_X1 port map( A1 => n2339, A2 => n3302, B1 => n4090, B2 => 
                           n3362, ZN => n13085);
   U5082 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n43, ZN => n12527);
   U5083 : AOI22_X1 port map( A1 => n2342, A2 => n3296, B1 => n4093, B2 => 
                           n3338, ZN => DataPath_RF_MUX_SELINPUT_8_n43);
   U5084 : INV_X1 port map( A => DataPath_RF_MUX_SELINPUT_8_n54, ZN => n12087);
   U5085 : AOI22_X1 port map( A1 => n2408, A2 => n3302, B1 => n4099, B2 => 
                           n3340, ZN => DataPath_RF_MUX_SELINPUT_8_n54);
   U5086 : INV_X1 port map( A => n13307, ZN => n12578);
   U5087 : AOI22_X1 port map( A1 => n2327, A2 => n3409, B1 => n3916, B2 => 
                           n3474, ZN => n13307);
   U5088 : INV_X1 port map( A => n13308, ZN => n12538);
   U5089 : AOI22_X1 port map( A1 => n2333, A2 => n3410, B1 => n3922, B2 => 
                           n3474, ZN => n13308);
   U5090 : INV_X1 port map( A => n13310, ZN => n12458);
   U5091 : AOI22_X1 port map( A1 => n2345, A2 => n3410, B1 => n3928, B2 => 
                           n3475, ZN => n13310);
   U5092 : INV_X1 port map( A => n13438, ZN => n12462);
   U5093 : AOI22_X1 port map( A1 => n2346, A2 => n3412, B1 => n3929, B2 => 
                           n3450, ZN => n13438);
   U5094 : INV_X1 port map( A => n13439, ZN => n12422);
   U5095 : AOI22_X1 port map( A1 => n2352, A2 => n3411, B1 => n3935, B2 => 
                           n3450, ZN => n13439);
   U5096 : INV_X1 port map( A => n13311, ZN => n12418);
   U5097 : AOI22_X1 port map( A1 => n2351, A2 => n3409, B1 => n3934, B2 => 
                           n3475, ZN => n13311);
   U5098 : INV_X1 port map( A => n13312, ZN => n12378);
   U5099 : AOI22_X1 port map( A1 => n2357, A2 => n3410, B1 => n3940, B2 => 
                           n3475, ZN => n13312);
   U5100 : INV_X1 port map( A => n13313, ZN => n12338);
   U5101 : AOI22_X1 port map( A1 => n2363, A2 => n3414, B1 => n3946, B2 => 
                           n3475, ZN => n13313);
   U5102 : INV_X1 port map( A => n13442, ZN => n12302);
   U5103 : AOI22_X1 port map( A1 => n2370, A2 => n3410, B1 => n3953, B2 => 
                           n3451, ZN => n13442);
   U5104 : INV_X1 port map( A => n13444, ZN => n12222);
   U5105 : AOI22_X1 port map( A1 => n2382, A2 => n3416, B1 => n3965, B2 => 
                           n3451, ZN => n13444);
   U5106 : INV_X1 port map( A => n13445, ZN => n12182);
   U5107 : AOI22_X1 port map( A1 => n2388, A2 => n3411, B1 => n3971, B2 => 
                           n3452, ZN => n13445);
   U5108 : INV_X1 port map( A => n13446, ZN => n12142);
   U5109 : AOI22_X1 port map( A1 => n2394, A2 => n3414, B1 => n3977, B2 => 
                           n3452, ZN => n13446);
   U5110 : INV_X1 port map( A => n13447, ZN => n12102);
   U5111 : AOI22_X1 port map( A1 => n2400, A2 => n3414, B1 => n3983, B2 => 
                           n3452, ZN => n13447);
   U5112 : INV_X1 port map( A => n13449, ZN => n12022);
   U5113 : AOI22_X1 port map( A1 => n2412, A2 => n3413, B1 => n3989, B2 => 
                           n3453, ZN => n13449);
   U5114 : INV_X1 port map( A => n13450, ZN => n11982);
   U5115 : AOI22_X1 port map( A1 => n2418, A2 => n3413, B1 => n3995, B2 => 
                           n3453, ZN => n13450);
   U5116 : INV_X1 port map( A => n13451, ZN => n11942);
   U5117 : AOI22_X1 port map( A1 => n2424, A2 => n3413, B1 => n4001, B2 => 
                           n3453, ZN => n13451);
   U5118 : INV_X1 port map( A => n13452, ZN => n11902);
   U5119 : AOI22_X1 port map( A1 => n2430, A2 => n3412, B1 => n4007, B2 => 
                           n3453, ZN => n13452);
   U5120 : INV_X1 port map( A => n13453, ZN => n11862);
   U5121 : AOI22_X1 port map( A1 => n2436, A2 => n3411, B1 => n4013, B2 => 
                           n3454, ZN => n13453);
   U5122 : INV_X1 port map( A => n13454, ZN => n11822);
   U5123 : AOI22_X1 port map( A1 => n2442, A2 => n3412, B1 => n4019, B2 => 
                           n3454, ZN => n13454);
   U5124 : INV_X1 port map( A => n13455, ZN => n11782);
   U5125 : AOI22_X1 port map( A1 => n2448, A2 => n3412, B1 => n4025, B2 => 
                           n3454, ZN => n13455);
   U5126 : INV_X1 port map( A => n13456, ZN => n11742);
   U5127 : AOI22_X1 port map( A1 => n2454, A2 => n3412, B1 => n4031, B2 => 
                           n3454, ZN => n13456);
   U5128 : INV_X1 port map( A => n13457, ZN => n11702);
   U5129 : AOI22_X1 port map( A1 => n2460, A2 => n3412, B1 => n4037, B2 => 
                           n3455, ZN => n13457);
   U5130 : INV_X1 port map( A => n13458, ZN => n11662);
   U5131 : AOI22_X1 port map( A1 => n2466, A2 => n3412, B1 => n4043, B2 => 
                           n3434, ZN => n13458);
   U5132 : INV_X1 port map( A => n13309, ZN => n12498);
   U5133 : AOI22_X1 port map( A1 => n2339, A2 => n3414, B1 => n4090, B2 => 
                           n3474, ZN => n13309);
   U5134 : INV_X1 port map( A => n13437, ZN => n12502);
   U5135 : AOI22_X1 port map( A1 => n2340, A2 => n3416, B1 => n4091, B2 => 
                           n3450, ZN => n13437);
   U5136 : INV_X1 port map( A => n13448, ZN => n12062);
   U5137 : AOI22_X1 port map( A1 => n2406, A2 => n3411, B1 => n4097, B2 => 
                           n3452, ZN => n13448);
   U5138 : INV_X1 port map( A => n13459, ZN => n11622);
   U5139 : AOI22_X1 port map( A1 => n2472, A2 => n3412, B1 => n4103, B2 => 
                           n3468, ZN => n13459);
   U5140 : INV_X1 port map( A => n13563, ZN => n12586);
   U5141 : AOI22_X1 port map( A1 => n2328, A2 => n3521, B1 => n3917, B2 => 
                           n3586, ZN => n13563);
   U5142 : INV_X1 port map( A => n13564, ZN => n12546);
   U5143 : AOI22_X1 port map( A1 => n2334, A2 => n3522, B1 => n3923, B2 => 
                           n3586, ZN => n13564);
   U5144 : INV_X1 port map( A => n13566, ZN => n12466);
   U5145 : AOI22_X1 port map( A1 => n2346, A2 => n3522, B1 => n3929, B2 => 
                           n3587, ZN => n13566);
   U5146 : INV_X1 port map( A => n13694, ZN => n12470);
   U5147 : AOI22_X1 port map( A1 => n2346, A2 => n3524, B1 => n3929, B2 => 
                           n3562, ZN => n13694);
   U5148 : INV_X1 port map( A => n13695, ZN => n12430);
   U5149 : AOI22_X1 port map( A1 => n2352, A2 => n3523, B1 => n3935, B2 => 
                           n3562, ZN => n13695);
   U5150 : INV_X1 port map( A => n13567, ZN => n12426);
   U5151 : AOI22_X1 port map( A1 => n2352, A2 => n3521, B1 => n3935, B2 => 
                           n3587, ZN => n13567);
   U5152 : INV_X1 port map( A => n13568, ZN => n12386);
   U5153 : AOI22_X1 port map( A1 => n2358, A2 => n3522, B1 => n3941, B2 => 
                           n3587, ZN => n13568);
   U5154 : INV_X1 port map( A => n13569, ZN => n12346);
   U5155 : AOI22_X1 port map( A1 => n2364, A2 => n3526, B1 => n3947, B2 => 
                           n3587, ZN => n13569);
   U5156 : INV_X1 port map( A => n13698, ZN => n12310);
   U5157 : AOI22_X1 port map( A1 => n2370, A2 => n3522, B1 => n3953, B2 => 
                           n3563, ZN => n13698);
   U5158 : INV_X1 port map( A => n13700, ZN => n12230);
   U5159 : AOI22_X1 port map( A1 => n2382, A2 => n3528, B1 => n3965, B2 => 
                           n3563, ZN => n13700);
   U5160 : INV_X1 port map( A => n13701, ZN => n12190);
   U5161 : AOI22_X1 port map( A1 => n2388, A2 => n3523, B1 => n3971, B2 => 
                           n3564, ZN => n13701);
   U5162 : INV_X1 port map( A => n13702, ZN => n12150);
   U5163 : AOI22_X1 port map( A1 => n2394, A2 => n3526, B1 => n3977, B2 => 
                           n3564, ZN => n13702);
   U5164 : INV_X1 port map( A => n13703, ZN => n12110);
   U5165 : AOI22_X1 port map( A1 => n2400, A2 => n3526, B1 => n3983, B2 => 
                           n3564, ZN => n13703);
   U5166 : INV_X1 port map( A => n13705, ZN => n12030);
   U5167 : AOI22_X1 port map( A1 => n2412, A2 => n3525, B1 => n3989, B2 => 
                           n3565, ZN => n13705);
   U5168 : INV_X1 port map( A => n13706, ZN => n11990);
   U5169 : AOI22_X1 port map( A1 => n2418, A2 => n3525, B1 => n3995, B2 => 
                           n3565, ZN => n13706);
   U5170 : INV_X1 port map( A => n13707, ZN => n11950);
   U5171 : AOI22_X1 port map( A1 => n2424, A2 => n3525, B1 => n4001, B2 => 
                           n3565, ZN => n13707);
   U5172 : INV_X1 port map( A => n13708, ZN => n11910);
   U5173 : AOI22_X1 port map( A1 => n2430, A2 => n3524, B1 => n4007, B2 => 
                           n3565, ZN => n13708);
   U5174 : INV_X1 port map( A => n13709, ZN => n11870);
   U5175 : AOI22_X1 port map( A1 => n2436, A2 => n3523, B1 => n4013, B2 => 
                           n3566, ZN => n13709);
   U5176 : INV_X1 port map( A => n13710, ZN => n11830);
   U5177 : AOI22_X1 port map( A1 => n2442, A2 => n3524, B1 => n4019, B2 => 
                           n3566, ZN => n13710);
   U5178 : INV_X1 port map( A => n13711, ZN => n11790);
   U5179 : AOI22_X1 port map( A1 => n2448, A2 => n3524, B1 => n4025, B2 => 
                           n3566, ZN => n13711);
   U5180 : INV_X1 port map( A => n13712, ZN => n11750);
   U5181 : AOI22_X1 port map( A1 => n2454, A2 => n3524, B1 => n4031, B2 => 
                           n3566, ZN => n13712);
   U5182 : INV_X1 port map( A => n13713, ZN => n11710);
   U5183 : AOI22_X1 port map( A1 => n2460, A2 => n3524, B1 => n4037, B2 => 
                           n3567, ZN => n13713);
   U5184 : INV_X1 port map( A => n13714, ZN => n11670);
   U5185 : AOI22_X1 port map( A1 => n2466, A2 => n3524, B1 => n4043, B2 => 
                           n3546, ZN => n13714);
   U5186 : INV_X1 port map( A => n13565, ZN => n12506);
   U5187 : AOI22_X1 port map( A1 => n2340, A2 => n3526, B1 => n4091, B2 => 
                           n3586, ZN => n13565);
   U5188 : INV_X1 port map( A => n13693, ZN => n12510);
   U5189 : AOI22_X1 port map( A1 => n2340, A2 => n3529, B1 => n4091, B2 => 
                           n3562, ZN => n13693);
   U5190 : INV_X1 port map( A => n13704, ZN => n12070);
   U5191 : AOI22_X1 port map( A1 => n2406, A2 => n3523, B1 => n4097, B2 => 
                           n3564, ZN => n13704);
   U5192 : INV_X1 port map( A => n13715, ZN => n11630);
   U5193 : AOI22_X1 port map( A1 => n2472, A2 => n3524, B1 => n4103, B2 => 
                           n3580, ZN => n13715);
   U5194 : INV_X1 port map( A => n13819, ZN => n12594);
   U5195 : AOI22_X1 port map( A1 => n2329, A2 => n3632, B1 => n3918, B2 => 
                           n3698, ZN => n13819);
   U5196 : INV_X1 port map( A => n13820, ZN => n12554);
   U5197 : AOI22_X1 port map( A1 => n2335, A2 => n3633, B1 => n3924, B2 => 
                           n3698, ZN => n13820);
   U5198 : INV_X1 port map( A => n13822, ZN => n12474);
   U5199 : AOI22_X1 port map( A1 => n2347, A2 => n3633, B1 => n3930, B2 => 
                           n3699, ZN => n13822);
   U5200 : INV_X1 port map( A => n13950, ZN => n12478);
   U5201 : AOI22_X1 port map( A1 => n2347, A2 => n3636, B1 => n3930, B2 => 
                           n3674, ZN => n13950);
   U5202 : INV_X1 port map( A => n13951, ZN => n12438);
   U5203 : AOI22_X1 port map( A1 => n2353, A2 => n3635, B1 => n3936, B2 => 
                           n3674, ZN => n13951);
   U5204 : INV_X1 port map( A => n13823, ZN => n12434);
   U5205 : AOI22_X1 port map( A1 => n2353, A2 => n3632, B1 => n3936, B2 => 
                           n3699, ZN => n13823);
   U5206 : INV_X1 port map( A => n13824, ZN => n12394);
   U5207 : AOI22_X1 port map( A1 => n2359, A2 => n3634, B1 => n3942, B2 => 
                           n3699, ZN => n13824);
   U5208 : INV_X1 port map( A => n13825, ZN => n12354);
   U5209 : AOI22_X1 port map( A1 => n2365, A2 => n3638, B1 => n3948, B2 => 
                           n3699, ZN => n13825);
   U5210 : INV_X1 port map( A => n13954, ZN => n12318);
   U5211 : AOI22_X1 port map( A1 => n2371, A2 => n3633, B1 => n3954, B2 => 
                           n3675, ZN => n13954);
   U5212 : INV_X1 port map( A => n13956, ZN => n12238);
   U5213 : AOI22_X1 port map( A1 => n2383, A2 => n3634, B1 => n3966, B2 => 
                           n3675, ZN => n13956);
   U5214 : INV_X1 port map( A => n13957, ZN => n12198);
   U5215 : AOI22_X1 port map( A1 => n2389, A2 => n3635, B1 => n3972, B2 => 
                           n3676, ZN => n13957);
   U5216 : INV_X1 port map( A => n13958, ZN => n12158);
   U5217 : AOI22_X1 port map( A1 => n2395, A2 => n3638, B1 => n3978, B2 => 
                           n3676, ZN => n13958);
   U5218 : INV_X1 port map( A => n13959, ZN => n12118);
   U5219 : AOI22_X1 port map( A1 => n2401, A2 => n3638, B1 => n3984, B2 => 
                           n3676, ZN => n13959);
   U5220 : INV_X1 port map( A => n13961, ZN => n12038);
   U5221 : AOI22_X1 port map( A1 => n2413, A2 => n3637, B1 => n3990, B2 => 
                           n3677, ZN => n13961);
   U5222 : INV_X1 port map( A => n13962, ZN => n11998);
   U5223 : AOI22_X1 port map( A1 => n2419, A2 => n3637, B1 => n3996, B2 => 
                           n3677, ZN => n13962);
   U5224 : INV_X1 port map( A => n13963, ZN => n11958);
   U5225 : AOI22_X1 port map( A1 => n2425, A2 => n3637, B1 => n4002, B2 => 
                           n3677, ZN => n13963);
   U5226 : INV_X1 port map( A => n13964, ZN => n11918);
   U5227 : AOI22_X1 port map( A1 => n2431, A2 => n3636, B1 => n4008, B2 => 
                           n3677, ZN => n13964);
   U5228 : INV_X1 port map( A => n13965, ZN => n11878);
   U5229 : AOI22_X1 port map( A1 => n2437, A2 => n3635, B1 => n4014, B2 => 
                           n3678, ZN => n13965);
   U5230 : INV_X1 port map( A => n13966, ZN => n11838);
   U5231 : AOI22_X1 port map( A1 => n2443, A2 => n3636, B1 => n4020, B2 => 
                           n3678, ZN => n13966);
   U5232 : INV_X1 port map( A => n13967, ZN => n11798);
   U5233 : AOI22_X1 port map( A1 => n2449, A2 => n3636, B1 => n4026, B2 => 
                           n3678, ZN => n13967);
   U5234 : INV_X1 port map( A => n13968, ZN => n11758);
   U5235 : AOI22_X1 port map( A1 => n2455, A2 => n3636, B1 => n4032, B2 => 
                           n3678, ZN => n13968);
   U5236 : INV_X1 port map( A => n13969, ZN => n11718);
   U5237 : AOI22_X1 port map( A1 => n2461, A2 => n3636, B1 => n4038, B2 => 
                           n3679, ZN => n13969);
   U5238 : INV_X1 port map( A => n13970, ZN => n11678);
   U5239 : AOI22_X1 port map( A1 => n2467, A2 => n3636, B1 => n4044, B2 => 
                           n3658, ZN => n13970);
   U5240 : INV_X1 port map( A => n13821, ZN => n12514);
   U5241 : AOI22_X1 port map( A1 => n2341, A2 => n3638, B1 => n4092, B2 => 
                           n3698, ZN => n13821);
   U5242 : INV_X1 port map( A => n13949, ZN => n12518);
   U5243 : AOI22_X1 port map( A1 => n2341, A2 => n3634, B1 => n4092, B2 => 
                           n3674, ZN => n13949);
   U5244 : INV_X1 port map( A => n13960, ZN => n12078);
   U5245 : AOI22_X1 port map( A1 => n2407, A2 => n3635, B1 => n4098, B2 => 
                           n3676, ZN => n13960);
   U5246 : INV_X1 port map( A => n13971, ZN => n11638);
   U5247 : AOI22_X1 port map( A1 => n2473, A2 => n3636, B1 => n4104, B2 => 
                           n3692, ZN => n13971);
   U5248 : INV_X1 port map( A => n14075, ZN => n12602);
   U5249 : AOI22_X1 port map( A1 => n2329, A2 => n3744, B1 => n3918, B2 => 
                           n3810, ZN => n14075);
   U5250 : INV_X1 port map( A => n14076, ZN => n12562);
   U5251 : AOI22_X1 port map( A1 => n2335, A2 => n3745, B1 => n3924, B2 => 
                           n3810, ZN => n14076);
   U5252 : INV_X1 port map( A => n14078, ZN => n12482);
   U5253 : AOI22_X1 port map( A1 => n2347, A2 => n3749, B1 => n3930, B2 => 
                           n3811, ZN => n14078);
   U5254 : INV_X1 port map( A => n14206, ZN => n12486);
   U5255 : AOI22_X1 port map( A1 => n2348, A2 => n3750, B1 => n3931, B2 => 
                           n3786, ZN => n14206);
   U5256 : INV_X1 port map( A => n14207, ZN => n12446);
   U5257 : AOI22_X1 port map( A1 => n2354, A2 => n3750, B1 => n3937, B2 => 
                           n3786, ZN => n14207);
   U5258 : INV_X1 port map( A => n14079, ZN => n12442);
   U5259 : AOI22_X1 port map( A1 => n2353, A2 => n3750, B1 => n3936, B2 => 
                           n3811, ZN => n14079);
   U5260 : INV_X1 port map( A => n14080, ZN => n12402);
   U5261 : AOI22_X1 port map( A1 => n2359, A2 => n3748, B1 => n3942, B2 => 
                           n3811, ZN => n14080);
   U5262 : INV_X1 port map( A => n14081, ZN => n12362);
   U5263 : AOI22_X1 port map( A1 => n2365, A2 => n3744, B1 => n3948, B2 => 
                           n3811, ZN => n14081);
   U5264 : INV_X1 port map( A => n14210, ZN => n12326);
   U5265 : AOI22_X1 port map( A1 => n2372, A2 => n3750, B1 => n3955, B2 => 
                           n3787, ZN => n14210);
   U5266 : INV_X1 port map( A => n14212, ZN => n12246);
   U5267 : AOI22_X1 port map( A1 => n2384, A2 => n3750, B1 => n3967, B2 => 
                           n3787, ZN => n14212);
   U5268 : INV_X1 port map( A => n14213, ZN => n12206);
   U5269 : AOI22_X1 port map( A1 => n2390, A2 => n3752, B1 => n3973, B2 => 
                           n3788, ZN => n14213);
   U5270 : INV_X1 port map( A => n14214, ZN => n12166);
   U5271 : AOI22_X1 port map( A1 => n2396, A2 => n3749, B1 => n3979, B2 => 
                           n3788, ZN => n14214);
   U5272 : INV_X1 port map( A => n14215, ZN => n12126);
   U5273 : AOI22_X1 port map( A1 => n2402, A2 => n3743, B1 => n3985, B2 => 
                           n3788, ZN => n14215);
   U5274 : INV_X1 port map( A => n14217, ZN => n12046);
   U5275 : AOI22_X1 port map( A1 => n2414, A2 => n3744, B1 => n3991, B2 => 
                           n3789, ZN => n14217);
   U5276 : INV_X1 port map( A => n14218, ZN => n12006);
   U5277 : AOI22_X1 port map( A1 => n2420, A2 => n3750, B1 => n3997, B2 => 
                           n3789, ZN => n14218);
   U5278 : INV_X1 port map( A => n14219, ZN => n11966);
   U5279 : AOI22_X1 port map( A1 => n2426, A2 => n3745, B1 => n4003, B2 => 
                           n3789, ZN => n14219);
   U5280 : INV_X1 port map( A => n14220, ZN => n11926);
   U5281 : AOI22_X1 port map( A1 => n2432, A2 => n3751, B1 => n4009, B2 => 
                           n3789, ZN => n14220);
   U5282 : INV_X1 port map( A => n14221, ZN => n11886);
   U5283 : AOI22_X1 port map( A1 => n2438, A2 => n3747, B1 => n4015, B2 => 
                           n3790, ZN => n14221);
   U5284 : INV_X1 port map( A => n14222, ZN => n11846);
   U5285 : AOI22_X1 port map( A1 => n2444, A2 => n3748, B1 => n4021, B2 => 
                           n3790, ZN => n14222);
   U5286 : INV_X1 port map( A => n14223, ZN => n11806);
   U5287 : AOI22_X1 port map( A1 => n2450, A2 => n3748, B1 => n4027, B2 => 
                           n3790, ZN => n14223);
   U5288 : INV_X1 port map( A => n14224, ZN => n11766);
   U5289 : AOI22_X1 port map( A1 => n2456, A2 => n3748, B1 => n4033, B2 => 
                           n3790, ZN => n14224);
   U5290 : INV_X1 port map( A => n14225, ZN => n11726);
   U5291 : AOI22_X1 port map( A1 => n2462, A2 => n3747, B1 => n4039, B2 => 
                           n3791, ZN => n14225);
   U5292 : INV_X1 port map( A => n14226, ZN => n11686);
   U5293 : AOI22_X1 port map( A1 => n2468, A2 => n3748, B1 => n4045, B2 => 
                           n3770, ZN => n14226);
   U5294 : INV_X1 port map( A => n14077, ZN => n12522);
   U5295 : AOI22_X1 port map( A1 => n2341, A2 => n3745, B1 => n4092, B2 => 
                           n3810, ZN => n14077);
   U5296 : INV_X1 port map( A => n14205, ZN => n12526);
   U5297 : AOI22_X1 port map( A1 => n2342, A2 => n3750, B1 => n4093, B2 => 
                           n3786, ZN => n14205);
   U5298 : INV_X1 port map( A => n14216, ZN => n12086);
   U5299 : AOI22_X1 port map( A1 => n2408, A2 => n3743, B1 => n4099, B2 => 
                           n3788, ZN => n14216);
   U5300 : INV_X1 port map( A => n14227, ZN => n11646);
   U5301 : AOI22_X1 port map( A1 => n2474, A2 => n3748, B1 => n4105, B2 => 
                           n3804, ZN => n14227);
   U5302 : INV_X1 port map( A => n13102, ZN => n11811);
   U5303 : AOI22_X1 port map( A1 => n2441, A2 => n3305, B1 => n4018, B2 => 
                           n3366, ZN => n13102);
   U5304 : INV_X1 port map( A => n13103, ZN => n11771);
   U5305 : AOI22_X1 port map( A1 => n2447, A2 => n3303, B1 => n4024, B2 => 
                           n3367, ZN => n13103);
   U5306 : INV_X1 port map( A => n13104, ZN => n11731);
   U5307 : AOI22_X1 port map( A1 => n2453, A2 => n3304, B1 => n4030, B2 => 
                           n3367, ZN => n13104);
   U5308 : INV_X1 port map( A => n13105, ZN => n11691);
   U5309 : AOI22_X1 port map( A1 => n2459, A2 => n3295, B1 => n4036, B2 => 
                           n3367, ZN => n13105);
   U5310 : INV_X1 port map( A => n13106, ZN => n11651);
   U5311 : AOI22_X1 port map( A1 => n2465, A2 => n3305, B1 => n4042, B2 => 
                           n3327, ZN => n13106);
   U5312 : INV_X1 port map( A => n13326, ZN => n11818);
   U5313 : AOI22_X1 port map( A1 => n2441, A2 => n3408, B1 => n4018, B2 => 
                           n3478, ZN => n13326);
   U5314 : INV_X1 port map( A => n13327, ZN => n11778);
   U5315 : AOI22_X1 port map( A1 => n2447, A2 => n3408, B1 => n4024, B2 => 
                           n3479, ZN => n13327);
   U5316 : INV_X1 port map( A => n13328, ZN => n11738);
   U5317 : AOI22_X1 port map( A1 => n2453, A2 => n3408, B1 => n4030, B2 => 
                           n3479, ZN => n13328);
   U5318 : INV_X1 port map( A => n13329, ZN => n11698);
   U5319 : AOI22_X1 port map( A1 => n2459, A2 => n3408, B1 => n4036, B2 => 
                           n3479, ZN => n13329);
   U5320 : INV_X1 port map( A => n13330, ZN => n11658);
   U5321 : AOI22_X1 port map( A1 => n2465, A2 => n3408, B1 => n4042, B2 => 
                           n3439, ZN => n13330);
   U5322 : INV_X1 port map( A => n13331, ZN => n11618);
   U5323 : AOI22_X1 port map( A1 => n2471, A2 => n3408, B1 => n4102, B2 => 
                           n3431, ZN => n13331);
   U5324 : INV_X1 port map( A => n13582, ZN => n11826);
   U5325 : AOI22_X1 port map( A1 => n2442, A2 => n3520, B1 => n4019, B2 => 
                           n3590, ZN => n13582);
   U5326 : INV_X1 port map( A => n13583, ZN => n11786);
   U5327 : AOI22_X1 port map( A1 => n2448, A2 => n3520, B1 => n4025, B2 => 
                           n3591, ZN => n13583);
   U5328 : INV_X1 port map( A => n13584, ZN => n11746);
   U5329 : AOI22_X1 port map( A1 => n2454, A2 => n3520, B1 => n4031, B2 => 
                           n3591, ZN => n13584);
   U5330 : INV_X1 port map( A => n13585, ZN => n11706);
   U5331 : AOI22_X1 port map( A1 => n2460, A2 => n3520, B1 => n4037, B2 => 
                           n3591, ZN => n13585);
   U5332 : INV_X1 port map( A => n13586, ZN => n11666);
   U5333 : AOI22_X1 port map( A1 => n2466, A2 => n3520, B1 => n4043, B2 => 
                           n3551, ZN => n13586);
   U5334 : INV_X1 port map( A => n13587, ZN => n11626);
   U5335 : AOI22_X1 port map( A1 => n2472, A2 => n3520, B1 => n4103, B2 => 
                           n3543, ZN => n13587);
   U5336 : INV_X1 port map( A => n13838, ZN => n11834);
   U5337 : AOI22_X1 port map( A1 => n2443, A2 => n3640, B1 => n4020, B2 => 
                           n3702, ZN => n13838);
   U5338 : INV_X1 port map( A => n13839, ZN => n11794);
   U5339 : AOI22_X1 port map( A1 => n2449, A2 => n3639, B1 => n4026, B2 => 
                           n3703, ZN => n13839);
   U5340 : INV_X1 port map( A => n13840, ZN => n11754);
   U5341 : AOI22_X1 port map( A1 => n2455, A2 => n3631, B1 => n4032, B2 => 
                           n3703, ZN => n13840);
   U5342 : INV_X1 port map( A => n13841, ZN => n11714);
   U5343 : AOI22_X1 port map( A1 => n2461, A2 => n3641, B1 => n4038, B2 => 
                           n3703, ZN => n13841);
   U5344 : INV_X1 port map( A => n13842, ZN => n11674);
   U5345 : AOI22_X1 port map( A1 => n2467, A2 => n3640, B1 => n4044, B2 => 
                           n3663, ZN => n13842);
   U5346 : INV_X1 port map( A => n13843, ZN => n11634);
   U5347 : AOI22_X1 port map( A1 => n2473, A2 => n3639, B1 => n4104, B2 => 
                           n3655, ZN => n13843);
   U5348 : INV_X1 port map( A => n14094, ZN => n11842);
   U5349 : AOI22_X1 port map( A1 => n2443, A2 => n3743, B1 => n4020, B2 => 
                           n3814, ZN => n14094);
   U5350 : INV_X1 port map( A => n14095, ZN => n11802);
   U5351 : AOI22_X1 port map( A1 => n2449, A2 => n3743, B1 => n4026, B2 => 
                           n3815, ZN => n14095);
   U5352 : INV_X1 port map( A => n14096, ZN => n11762);
   U5353 : AOI22_X1 port map( A1 => n2455, A2 => n3744, B1 => n4032, B2 => 
                           n3815, ZN => n14096);
   U5354 : INV_X1 port map( A => n14097, ZN => n11722);
   U5355 : AOI22_X1 port map( A1 => n2461, A2 => n3745, B1 => n4038, B2 => 
                           n3815, ZN => n14097);
   U5356 : INV_X1 port map( A => n14098, ZN => n11682);
   U5357 : AOI22_X1 port map( A1 => n2467, A2 => n3751, B1 => n4044, B2 => 
                           n3775, ZN => n14098);
   U5358 : INV_X1 port map( A => n14099, ZN => n11642);
   U5359 : AOI22_X1 port map( A1 => n2473, A2 => n3746, B1 => n4104, B2 => 
                           n3767, ZN => n14099);
   U5360 : INV_X1 port map( A => n13435, ZN => n12582);
   U5361 : AOI22_X1 port map( A1 => n2328, A2 => n3415, B1 => n3917, B2 => 
                           n3449, ZN => n13435);
   U5362 : INV_X1 port map( A => n13436, ZN => n12542);
   U5363 : AOI22_X1 port map( A1 => n2334, A2 => n3415, B1 => n3923, B2 => 
                           n3449, ZN => n13436);
   U5364 : INV_X1 port map( A => n13440, ZN => n12382);
   U5365 : AOI22_X1 port map( A1 => n2358, A2 => n3415, B1 => n3941, B2 => 
                           n3450, ZN => n13440);
   U5366 : INV_X1 port map( A => n13441, ZN => n12342);
   U5367 : AOI22_X1 port map( A1 => n2364, A2 => n3415, B1 => n3947, B2 => 
                           n3451, ZN => n13441);
   U5368 : INV_X1 port map( A => n13443, ZN => n12262);
   U5369 : AOI22_X1 port map( A1 => n2376, A2 => n3415, B1 => n3959, B2 => 
                           n3451, ZN => n13443);
   U5370 : INV_X1 port map( A => n13691, ZN => n12590);
   U5371 : AOI22_X1 port map( A1 => n2328, A2 => n3527, B1 => n3917, B2 => 
                           n3561, ZN => n13691);
   U5372 : INV_X1 port map( A => n13692, ZN => n12550);
   U5373 : AOI22_X1 port map( A1 => n2334, A2 => n3527, B1 => n3923, B2 => 
                           n3561, ZN => n13692);
   U5374 : INV_X1 port map( A => n13696, ZN => n12390);
   U5375 : AOI22_X1 port map( A1 => n2358, A2 => n3527, B1 => n3941, B2 => 
                           n3562, ZN => n13696);
   U5376 : INV_X1 port map( A => n13697, ZN => n12350);
   U5377 : AOI22_X1 port map( A1 => n2364, A2 => n3527, B1 => n3947, B2 => 
                           n3563, ZN => n13697);
   U5378 : INV_X1 port map( A => n13699, ZN => n12270);
   U5379 : AOI22_X1 port map( A1 => n2376, A2 => n3527, B1 => n3959, B2 => 
                           n3563, ZN => n13699);
   U5380 : INV_X1 port map( A => n13947, ZN => n12598);
   U5381 : AOI22_X1 port map( A1 => n2329, A2 => n3639, B1 => n3918, B2 => 
                           n3673, ZN => n13947);
   U5382 : INV_X1 port map( A => n13948, ZN => n12558);
   U5383 : AOI22_X1 port map( A1 => n2335, A2 => n3639, B1 => n3924, B2 => 
                           n3673, ZN => n13948);
   U5384 : INV_X1 port map( A => n13952, ZN => n12398);
   U5385 : AOI22_X1 port map( A1 => n2359, A2 => n3639, B1 => n3942, B2 => 
                           n3674, ZN => n13952);
   U5386 : INV_X1 port map( A => n13953, ZN => n12358);
   U5387 : AOI22_X1 port map( A1 => n2365, A2 => n3639, B1 => n3948, B2 => 
                           n3675, ZN => n13953);
   U5388 : INV_X1 port map( A => n13955, ZN => n12278);
   U5389 : AOI22_X1 port map( A1 => n2377, A2 => n3639, B1 => n3960, B2 => 
                           n3675, ZN => n13955);
   U5390 : INV_X1 port map( A => n14203, ZN => n12606);
   U5391 : AOI22_X1 port map( A1 => n2330, A2 => n3751, B1 => n3919, B2 => 
                           n3785, ZN => n14203);
   U5392 : INV_X1 port map( A => n14204, ZN => n12566);
   U5393 : AOI22_X1 port map( A1 => n2336, A2 => n3751, B1 => n3925, B2 => 
                           n3785, ZN => n14204);
   U5394 : INV_X1 port map( A => n14208, ZN => n12406);
   U5395 : AOI22_X1 port map( A1 => n2360, A2 => n3751, B1 => n3943, B2 => 
                           n3786, ZN => n14208);
   U5396 : INV_X1 port map( A => n14209, ZN => n12366);
   U5397 : AOI22_X1 port map( A1 => n2366, A2 => n3751, B1 => n3949, B2 => 
                           n3787, ZN => n14209);
   U5398 : INV_X1 port map( A => n14211, ZN => n12286);
   U5399 : AOI22_X1 port map( A1 => n2378, A2 => n3751, B1 => n3961, B2 => 
                           n3787, ZN => n14211);
   U5400 : INV_X1 port map( A => n13051, ZN => n12570);
   U5401 : AOI22_X1 port map( A1 => n2327, A2 => n3296, B1 => n3916, B2 => 
                           n3355, ZN => n13051);
   U5402 : INV_X1 port map( A => n13179, ZN => n12574);
   U5403 : AOI22_X1 port map( A1 => n2327, A2 => n3301, B1 => n3916, B2 => 
                           n3331, ZN => n13179);
   U5404 : INV_X1 port map( A => n13052, ZN => n12530);
   U5405 : AOI22_X1 port map( A1 => n2333, A2 => n3296, B1 => n3922, B2 => 
                           n3356, ZN => n13052);
   U5406 : INV_X1 port map( A => n13180, ZN => n12534);
   U5407 : AOI22_X1 port map( A1 => n2333, A2 => n3301, B1 => n3922, B2 => 
                           n3331, ZN => n13180);
   U5408 : INV_X1 port map( A => n13054, ZN => n12450);
   U5409 : AOI22_X1 port map( A1 => n2345, A2 => n3296, B1 => n3928, B2 => 
                           n3356, ZN => n13054);
   U5410 : INV_X1 port map( A => n13182, ZN => n12454);
   U5411 : AOI22_X1 port map( A1 => n2345, A2 => n3300, B1 => n3928, B2 => 
                           n3332, ZN => n13182);
   U5412 : INV_X1 port map( A => n13055, ZN => n12410);
   U5413 : AOI22_X1 port map( A1 => n2351, A2 => n3296, B1 => n3934, B2 => 
                           n3357, ZN => n13055);
   U5414 : INV_X1 port map( A => n13183, ZN => n12414);
   U5415 : AOI22_X1 port map( A1 => n2351, A2 => n3300, B1 => n3934, B2 => 
                           n3332, ZN => n13183);
   U5416 : INV_X1 port map( A => n13056, ZN => n12370);
   U5417 : AOI22_X1 port map( A1 => n2357, A2 => n3296, B1 => n3940, B2 => 
                           n3357, ZN => n13056);
   U5418 : INV_X1 port map( A => n13184, ZN => n12374);
   U5419 : AOI22_X1 port map( A1 => n2357, A2 => n3300, B1 => n3940, B2 => 
                           n3332, ZN => n13184);
   U5420 : INV_X1 port map( A => n13057, ZN => n12330);
   U5421 : AOI22_X1 port map( A1 => n2363, A2 => n3296, B1 => n3946, B2 => 
                           n3357, ZN => n13057);
   U5422 : INV_X1 port map( A => n13185, ZN => n12334);
   U5423 : AOI22_X1 port map( A1 => n2363, A2 => n3300, B1 => n3946, B2 => 
                           n3332, ZN => n13185);
   U5424 : INV_X1 port map( A => n13058, ZN => n12290);
   U5425 : AOI22_X1 port map( A1 => n2369, A2 => n3296, B1 => n3952, B2 => 
                           n3357, ZN => n13058);
   U5426 : INV_X1 port map( A => n13186, ZN => n12294);
   U5427 : AOI22_X1 port map( A1 => n2369, A2 => n3300, B1 => n3952, B2 => 
                           n3333, ZN => n13186);
   U5428 : INV_X1 port map( A => n13059, ZN => n12250);
   U5429 : AOI22_X1 port map( A1 => n2375, A2 => n3296, B1 => n3958, B2 => 
                           n3358, ZN => n13059);
   U5430 : INV_X1 port map( A => n13187, ZN => n12254);
   U5431 : AOI22_X1 port map( A1 => n2375, A2 => n3300, B1 => n3958, B2 => 
                           n3333, ZN => n13187);
   U5432 : INV_X1 port map( A => n13060, ZN => n12210);
   U5433 : AOI22_X1 port map( A1 => n2381, A2 => n3297, B1 => n3964, B2 => 
                           n3358, ZN => n13060);
   U5434 : INV_X1 port map( A => n13188, ZN => n12214);
   U5435 : AOI22_X1 port map( A1 => n2381, A2 => n3300, B1 => n3964, B2 => 
                           n3333, ZN => n13188);
   U5436 : INV_X1 port map( A => n13061, ZN => n12170);
   U5437 : AOI22_X1 port map( A1 => n2387, A2 => n3298, B1 => n3970, B2 => 
                           n3358, ZN => n13061);
   U5438 : INV_X1 port map( A => n13189, ZN => n12174);
   U5439 : AOI22_X1 port map( A1 => n2387, A2 => n3300, B1 => n3970, B2 => 
                           n3333, ZN => n13189);
   U5440 : INV_X1 port map( A => n13062, ZN => n12130);
   U5441 : AOI22_X1 port map( A1 => n2393, A2 => n3296, B1 => n3976, B2 => 
                           n3358, ZN => n13062);
   U5442 : INV_X1 port map( A => n13190, ZN => n12134);
   U5443 : AOI22_X1 port map( A1 => n2393, A2 => n3300, B1 => n3976, B2 => 
                           n3334, ZN => n13190);
   U5444 : INV_X1 port map( A => n13063, ZN => n12090);
   U5445 : AOI22_X1 port map( A1 => n2399, A2 => n3300, B1 => n3982, B2 => 
                           n3359, ZN => n13063);
   U5446 : INV_X1 port map( A => n13191, ZN => n12094);
   U5447 : AOI22_X1 port map( A1 => n2399, A2 => n3300, B1 => n3982, B2 => 
                           n3334, ZN => n13191);
   U5448 : INV_X1 port map( A => n13065, ZN => n12010);
   U5449 : AOI22_X1 port map( A1 => n2411, A2 => n3302, B1 => n3988, B2 => 
                           n3359, ZN => n13065);
   U5450 : INV_X1 port map( A => n13193, ZN => n12014);
   U5451 : AOI22_X1 port map( A1 => n2411, A2 => n3300, B1 => n3988, B2 => 
                           n3334, ZN => n13193);
   U5452 : INV_X1 port map( A => n13066, ZN => n11970);
   U5453 : AOI22_X1 port map( A1 => n2417, A2 => n3301, B1 => n3994, B2 => 
                           n3359, ZN => n13066);
   U5454 : INV_X1 port map( A => n13194, ZN => n11974);
   U5455 : AOI22_X1 port map( A1 => n2417, A2 => n3299, B1 => n3994, B2 => 
                           n3335, ZN => n13194);
   U5456 : INV_X1 port map( A => n13067, ZN => n11930);
   U5457 : AOI22_X1 port map( A1 => n2423, A2 => n3299, B1 => n4000, B2 => 
                           n3360, ZN => n13067);
   U5458 : INV_X1 port map( A => n13195, ZN => n11934);
   U5459 : AOI22_X1 port map( A1 => n2423, A2 => n3302, B1 => n4000, B2 => 
                           n3335, ZN => n13195);
   U5460 : INV_X1 port map( A => n13068, ZN => n11890);
   U5461 : AOI22_X1 port map( A1 => n2429, A2 => n3300, B1 => n4006, B2 => 
                           n3360, ZN => n13068);
   U5462 : INV_X1 port map( A => n13196, ZN => n11894);
   U5463 : AOI22_X1 port map( A1 => n2429, A2 => n3301, B1 => n4006, B2 => 
                           n3335, ZN => n13196);
   U5464 : INV_X1 port map( A => n13069, ZN => n11850);
   U5465 : AOI22_X1 port map( A1 => n2435, A2 => n3297, B1 => n4012, B2 => 
                           n3360, ZN => n13069);
   U5466 : INV_X1 port map( A => n13197, ZN => n11854);
   U5467 : AOI22_X1 port map( A1 => n2435, A2 => n3297, B1 => n4012, B2 => 
                           n3335, ZN => n13197);
   U5468 : INV_X1 port map( A => n13070, ZN => n11810);
   U5469 : AOI22_X1 port map( A1 => n2441, A2 => n3298, B1 => n4018, B2 => 
                           n3360, ZN => n13070);
   U5470 : INV_X1 port map( A => n13198, ZN => n11814);
   U5471 : AOI22_X1 port map( A1 => n2441, A2 => n3298, B1 => n4018, B2 => 
                           n3336, ZN => n13198);
   U5472 : INV_X1 port map( A => n13071, ZN => n11770);
   U5473 : AOI22_X1 port map( A1 => n2447, A2 => n3299, B1 => n4024, B2 => 
                           n3361, ZN => n13071);
   U5474 : INV_X1 port map( A => n13199, ZN => n11774);
   U5475 : AOI22_X1 port map( A1 => n2447, A2 => n3296, B1 => n4024, B2 => 
                           n3336, ZN => n13199);
   U5476 : INV_X1 port map( A => n13072, ZN => n11730);
   U5477 : AOI22_X1 port map( A1 => n2453, A2 => n3297, B1 => n4030, B2 => 
                           n3361, ZN => n13072);
   U5478 : INV_X1 port map( A => n13200, ZN => n11734);
   U5479 : AOI22_X1 port map( A1 => n2453, A2 => n3301, B1 => n4030, B2 => 
                           n3336, ZN => n13200);
   U5480 : INV_X1 port map( A => n13073, ZN => n11690);
   U5481 : AOI22_X1 port map( A1 => n2459, A2 => n3298, B1 => n4036, B2 => 
                           n3361, ZN => n13073);
   U5482 : INV_X1 port map( A => n13201, ZN => n11694);
   U5483 : AOI22_X1 port map( A1 => n2459, A2 => n3300, B1 => n4036, B2 => 
                           n3336, ZN => n13201);
   U5484 : INV_X1 port map( A => n13074, ZN => n11650);
   U5485 : AOI22_X1 port map( A1 => n2465, A2 => n3296, B1 => n4042, B2 => 
                           n3361, ZN => n13074);
   U5486 : INV_X1 port map( A => n13202, ZN => n11654);
   U5487 : AOI22_X1 port map( A1 => n2465, A2 => n3299, B1 => n4042, B2 => 
                           n3337, ZN => n13202);
   U5488 : INV_X1 port map( A => n13053, ZN => n12490);
   U5489 : AOI22_X1 port map( A1 => n2339, A2 => n3296, B1 => n4090, B2 => 
                           n3356, ZN => n13053);
   U5490 : INV_X1 port map( A => n13181, ZN => n12494);
   U5491 : AOI22_X1 port map( A1 => n2339, A2 => n3300, B1 => n4090, B2 => 
                           n3331, ZN => n13181);
   U5492 : INV_X1 port map( A => n13064, ZN => n12050);
   U5493 : AOI22_X1 port map( A1 => n2405, A2 => n3296, B1 => n4096, B2 => 
                           n3359, ZN => n13064);
   U5494 : INV_X1 port map( A => n13192, ZN => n12054);
   U5495 : AOI22_X1 port map( A1 => n2405, A2 => n3300, B1 => n4096, B2 => 
                           n3334, ZN => n13192);
   U5496 : INV_X1 port map( A => n13075, ZN => n11610);
   U5497 : AOI22_X1 port map( A1 => n2471, A2 => n3299, B1 => n4102, B2 => 
                           n3362, ZN => n13075);
   U5498 : INV_X1 port map( A => n13275, ZN => n12577);
   U5499 : AOI22_X1 port map( A1 => n2327, A2 => n3409, B1 => n3916, B2 => 
                           n3467, ZN => n13275);
   U5500 : INV_X1 port map( A => n13403, ZN => n12581);
   U5501 : AOI22_X1 port map( A1 => n2328, A2 => n3414, B1 => n3917, B2 => 
                           n3443, ZN => n13403);
   U5502 : INV_X1 port map( A => n13276, ZN => n12537);
   U5503 : AOI22_X1 port map( A1 => n2333, A2 => n3409, B1 => n3922, B2 => 
                           n3468, ZN => n13276);
   U5504 : INV_X1 port map( A => n13404, ZN => n12541);
   U5505 : AOI22_X1 port map( A1 => n2334, A2 => n3414, B1 => n3923, B2 => 
                           n3443, ZN => n13404);
   U5506 : INV_X1 port map( A => n13278, ZN => n12457);
   U5507 : AOI22_X1 port map( A1 => n2345, A2 => n3413, B1 => n3928, B2 => 
                           n3468, ZN => n13278);
   U5508 : INV_X1 port map( A => n13406, ZN => n12461);
   U5509 : AOI22_X1 port map( A1 => n2346, A2 => n3414, B1 => n3929, B2 => 
                           n3444, ZN => n13406);
   U5510 : INV_X1 port map( A => n13279, ZN => n12417);
   U5511 : AOI22_X1 port map( A1 => n2351, A2 => n3412, B1 => n3934, B2 => 
                           n3469, ZN => n13279);
   U5512 : INV_X1 port map( A => n13280, ZN => n12377);
   U5513 : AOI22_X1 port map( A1 => n2357, A2 => n3411, B1 => n3940, B2 => 
                           n3469, ZN => n13280);
   U5514 : INV_X1 port map( A => n13408, ZN => n12381);
   U5515 : AOI22_X1 port map( A1 => n2358, A2 => n3414, B1 => n3941, B2 => 
                           n3444, ZN => n13408);
   U5516 : INV_X1 port map( A => n13281, ZN => n12337);
   U5517 : AOI22_X1 port map( A1 => n2363, A2 => n3414, B1 => n3946, B2 => 
                           n3469, ZN => n13281);
   U5518 : INV_X1 port map( A => n13409, ZN => n12341);
   U5519 : AOI22_X1 port map( A1 => n2364, A2 => n3414, B1 => n3947, B2 => 
                           n3444, ZN => n13409);
   U5520 : INV_X1 port map( A => n13282, ZN => n12297);
   U5521 : AOI22_X1 port map( A1 => n2369, A2 => n3410, B1 => n3952, B2 => 
                           n3469, ZN => n13282);
   U5522 : INV_X1 port map( A => n13410, ZN => n12301);
   U5523 : AOI22_X1 port map( A1 => n2370, A2 => n3414, B1 => n3953, B2 => 
                           n3445, ZN => n13410);
   U5524 : INV_X1 port map( A => n13283, ZN => n12257);
   U5525 : AOI22_X1 port map( A1 => n2375, A2 => n3407, B1 => n3958, B2 => 
                           n3470, ZN => n13283);
   U5526 : INV_X1 port map( A => n13411, ZN => n12261);
   U5527 : AOI22_X1 port map( A1 => n2376, A2 => n3409, B1 => n3959, B2 => 
                           n3445, ZN => n13411);
   U5528 : INV_X1 port map( A => n13284, ZN => n12217);
   U5529 : AOI22_X1 port map( A1 => n2381, A2 => n3410, B1 => n3964, B2 => 
                           n3470, ZN => n13284);
   U5530 : INV_X1 port map( A => n13412, ZN => n12221);
   U5531 : AOI22_X1 port map( A1 => n2382, A2 => n3410, B1 => n3965, B2 => 
                           n3445, ZN => n13412);
   U5532 : INV_X1 port map( A => n13285, ZN => n12177);
   U5533 : AOI22_X1 port map( A1 => n2387, A2 => n3410, B1 => n3970, B2 => 
                           n3470, ZN => n13285);
   U5534 : INV_X1 port map( A => n13413, ZN => n12181);
   U5535 : AOI22_X1 port map( A1 => n2388, A2 => n3414, B1 => n3971, B2 => 
                           n3445, ZN => n13413);
   U5536 : INV_X1 port map( A => n13286, ZN => n12137);
   U5537 : AOI22_X1 port map( A1 => n2393, A2 => n3410, B1 => n3976, B2 => 
                           n3470, ZN => n13286);
   U5538 : INV_X1 port map( A => n13414, ZN => n12141);
   U5539 : AOI22_X1 port map( A1 => n2394, A2 => n3414, B1 => n3977, B2 => 
                           n3446, ZN => n13414);
   U5540 : INV_X1 port map( A => n13287, ZN => n12097);
   U5541 : AOI22_X1 port map( A1 => n2399, A2 => n3410, B1 => n3982, B2 => 
                           n3471, ZN => n13287);
   U5542 : INV_X1 port map( A => n13415, ZN => n12101);
   U5543 : AOI22_X1 port map( A1 => n2400, A2 => n3414, B1 => n3983, B2 => 
                           n3446, ZN => n13415);
   U5544 : INV_X1 port map( A => n13289, ZN => n12017);
   U5545 : AOI22_X1 port map( A1 => n2411, A2 => n3410, B1 => n3988, B2 => 
                           n3471, ZN => n13289);
   U5546 : INV_X1 port map( A => n13417, ZN => n12021);
   U5547 : AOI22_X1 port map( A1 => n2412, A2 => n3413, B1 => n3989, B2 => 
                           n3446, ZN => n13417);
   U5548 : INV_X1 port map( A => n13290, ZN => n11977);
   U5549 : AOI22_X1 port map( A1 => n2417, A2 => n3410, B1 => n3994, B2 => 
                           n3471, ZN => n13290);
   U5550 : INV_X1 port map( A => n13418, ZN => n11981);
   U5551 : AOI22_X1 port map( A1 => n2418, A2 => n3412, B1 => n3995, B2 => 
                           n3447, ZN => n13418);
   U5552 : INV_X1 port map( A => n13291, ZN => n11937);
   U5553 : AOI22_X1 port map( A1 => n2423, A2 => n3410, B1 => n4000, B2 => 
                           n3472, ZN => n13291);
   U5554 : INV_X1 port map( A => n13419, ZN => n11941);
   U5555 : AOI22_X1 port map( A1 => n2424, A2 => n3414, B1 => n4001, B2 => 
                           n3447, ZN => n13419);
   U5556 : INV_X1 port map( A => n13292, ZN => n11897);
   U5557 : AOI22_X1 port map( A1 => n2429, A2 => n3410, B1 => n4006, B2 => 
                           n3472, ZN => n13292);
   U5558 : INV_X1 port map( A => n13420, ZN => n11901);
   U5559 : AOI22_X1 port map( A1 => n2430, A2 => n3411, B1 => n4007, B2 => 
                           n3447, ZN => n13420);
   U5560 : INV_X1 port map( A => n13293, ZN => n11857);
   U5561 : AOI22_X1 port map( A1 => n2435, A2 => n3410, B1 => n4012, B2 => 
                           n3472, ZN => n13293);
   U5562 : INV_X1 port map( A => n13421, ZN => n11861);
   U5563 : AOI22_X1 port map( A1 => n2436, A2 => n3414, B1 => n4013, B2 => 
                           n3447, ZN => n13421);
   U5564 : INV_X1 port map( A => n13294, ZN => n11817);
   U5565 : AOI22_X1 port map( A1 => n2441, A2 => n3410, B1 => n4018, B2 => 
                           n3472, ZN => n13294);
   U5566 : INV_X1 port map( A => n13422, ZN => n11821);
   U5567 : AOI22_X1 port map( A1 => n2442, A2 => n3410, B1 => n4019, B2 => 
                           n3448, ZN => n13422);
   U5568 : INV_X1 port map( A => n13295, ZN => n11777);
   U5569 : AOI22_X1 port map( A1 => n2447, A2 => n3413, B1 => n4024, B2 => 
                           n3473, ZN => n13295);
   U5570 : INV_X1 port map( A => n13423, ZN => n11781);
   U5571 : AOI22_X1 port map( A1 => n2448, A2 => n3414, B1 => n4025, B2 => 
                           n3448, ZN => n13423);
   U5572 : INV_X1 port map( A => n13296, ZN => n11737);
   U5573 : AOI22_X1 port map( A1 => n2453, A2 => n3412, B1 => n4030, B2 => 
                           n3473, ZN => n13296);
   U5574 : INV_X1 port map( A => n13424, ZN => n11741);
   U5575 : AOI22_X1 port map( A1 => n2454, A2 => n3407, B1 => n4031, B2 => 
                           n3448, ZN => n13424);
   U5576 : INV_X1 port map( A => n13297, ZN => n11697);
   U5577 : AOI22_X1 port map( A1 => n2459, A2 => n3413, B1 => n4036, B2 => 
                           n3473, ZN => n13297);
   U5578 : INV_X1 port map( A => n13298, ZN => n11657);
   U5579 : AOI22_X1 port map( A1 => n2465, A2 => n3411, B1 => n4042, B2 => 
                           n3473, ZN => n13298);
   U5580 : INV_X1 port map( A => n13277, ZN => n12497);
   U5581 : AOI22_X1 port map( A1 => n2339, A2 => n3409, B1 => n4090, B2 => 
                           n3468, ZN => n13277);
   U5582 : INV_X1 port map( A => n13405, ZN => n12501);
   U5583 : AOI22_X1 port map( A1 => n2340, A2 => n3414, B1 => n4091, B2 => 
                           n3443, ZN => n13405);
   U5584 : INV_X1 port map( A => n13288, ZN => n12057);
   U5585 : AOI22_X1 port map( A1 => n2405, A2 => n3410, B1 => n4096, B2 => 
                           n3471, ZN => n13288);
   U5586 : INV_X1 port map( A => n13416, ZN => n12061);
   U5587 : AOI22_X1 port map( A1 => n2406, A2 => n3409, B1 => n4097, B2 => 
                           n3446, ZN => n13416);
   U5588 : INV_X1 port map( A => n13299, ZN => n11617);
   U5589 : AOI22_X1 port map( A1 => n2471, A2 => n3410, B1 => n4102, B2 => 
                           n3474, ZN => n13299);
   U5590 : INV_X1 port map( A => n13531, ZN => n12585);
   U5591 : AOI22_X1 port map( A1 => n2328, A2 => n3521, B1 => n3917, B2 => 
                           n3579, ZN => n13531);
   U5592 : INV_X1 port map( A => n13659, ZN => n12589);
   U5593 : AOI22_X1 port map( A1 => n2328, A2 => n3526, B1 => n3917, B2 => 
                           n3555, ZN => n13659);
   U5594 : INV_X1 port map( A => n13532, ZN => n12545);
   U5595 : AOI22_X1 port map( A1 => n2334, A2 => n3521, B1 => n3923, B2 => 
                           n3580, ZN => n13532);
   U5596 : INV_X1 port map( A => n13660, ZN => n12549);
   U5597 : AOI22_X1 port map( A1 => n2334, A2 => n3526, B1 => n3923, B2 => 
                           n3555, ZN => n13660);
   U5598 : INV_X1 port map( A => n13534, ZN => n12465);
   U5599 : AOI22_X1 port map( A1 => n2346, A2 => n3525, B1 => n3929, B2 => 
                           n3580, ZN => n13534);
   U5600 : INV_X1 port map( A => n13662, ZN => n12469);
   U5601 : AOI22_X1 port map( A1 => n2346, A2 => n3526, B1 => n3929, B2 => 
                           n3556, ZN => n13662);
   U5602 : INV_X1 port map( A => n13535, ZN => n12425);
   U5603 : AOI22_X1 port map( A1 => n2352, A2 => n3524, B1 => n3935, B2 => 
                           n3581, ZN => n13535);
   U5604 : INV_X1 port map( A => n13536, ZN => n12385);
   U5605 : AOI22_X1 port map( A1 => n2358, A2 => n3523, B1 => n3941, B2 => 
                           n3581, ZN => n13536);
   U5606 : INV_X1 port map( A => n13664, ZN => n12389);
   U5607 : AOI22_X1 port map( A1 => n2358, A2 => n3526, B1 => n3941, B2 => 
                           n3556, ZN => n13664);
   U5608 : INV_X1 port map( A => n13537, ZN => n12345);
   U5609 : AOI22_X1 port map( A1 => n2364, A2 => n3526, B1 => n3947, B2 => 
                           n3581, ZN => n13537);
   U5610 : INV_X1 port map( A => n13665, ZN => n12349);
   U5611 : AOI22_X1 port map( A1 => n2364, A2 => n3526, B1 => n3947, B2 => 
                           n3556, ZN => n13665);
   U5612 : INV_X1 port map( A => n13538, ZN => n12305);
   U5613 : AOI22_X1 port map( A1 => n2370, A2 => n3522, B1 => n3953, B2 => 
                           n3581, ZN => n13538);
   U5614 : INV_X1 port map( A => n13666, ZN => n12309);
   U5615 : AOI22_X1 port map( A1 => n2370, A2 => n3526, B1 => n3953, B2 => 
                           n3557, ZN => n13666);
   U5616 : INV_X1 port map( A => n13539, ZN => n12265);
   U5617 : AOI22_X1 port map( A1 => n2376, A2 => n3520, B1 => n3959, B2 => 
                           n3582, ZN => n13539);
   U5618 : INV_X1 port map( A => n13667, ZN => n12269);
   U5619 : AOI22_X1 port map( A1 => n2376, A2 => n3521, B1 => n3959, B2 => 
                           n3557, ZN => n13667);
   U5620 : INV_X1 port map( A => n13540, ZN => n12225);
   U5621 : AOI22_X1 port map( A1 => n2382, A2 => n3522, B1 => n3965, B2 => 
                           n3582, ZN => n13540);
   U5622 : INV_X1 port map( A => n13668, ZN => n12229);
   U5623 : AOI22_X1 port map( A1 => n2382, A2 => n3522, B1 => n3965, B2 => 
                           n3557, ZN => n13668);
   U5624 : INV_X1 port map( A => n13541, ZN => n12185);
   U5625 : AOI22_X1 port map( A1 => n2388, A2 => n3522, B1 => n3971, B2 => 
                           n3582, ZN => n13541);
   U5626 : INV_X1 port map( A => n13669, ZN => n12189);
   U5627 : AOI22_X1 port map( A1 => n2388, A2 => n3526, B1 => n3971, B2 => 
                           n3557, ZN => n13669);
   U5628 : INV_X1 port map( A => n13542, ZN => n12145);
   U5629 : AOI22_X1 port map( A1 => n2394, A2 => n3522, B1 => n3977, B2 => 
                           n3582, ZN => n13542);
   U5630 : INV_X1 port map( A => n13670, ZN => n12149);
   U5631 : AOI22_X1 port map( A1 => n2394, A2 => n3526, B1 => n3977, B2 => 
                           n3558, ZN => n13670);
   U5632 : INV_X1 port map( A => n13543, ZN => n12105);
   U5633 : AOI22_X1 port map( A1 => n2400, A2 => n3522, B1 => n3983, B2 => 
                           n3583, ZN => n13543);
   U5634 : INV_X1 port map( A => n13671, ZN => n12109);
   U5635 : AOI22_X1 port map( A1 => n2400, A2 => n3526, B1 => n3983, B2 => 
                           n3558, ZN => n13671);
   U5636 : INV_X1 port map( A => n13545, ZN => n12025);
   U5637 : AOI22_X1 port map( A1 => n2412, A2 => n3522, B1 => n3989, B2 => 
                           n3583, ZN => n13545);
   U5638 : INV_X1 port map( A => n13673, ZN => n12029);
   U5639 : AOI22_X1 port map( A1 => n2412, A2 => n3525, B1 => n3989, B2 => 
                           n3558, ZN => n13673);
   U5640 : INV_X1 port map( A => n13546, ZN => n11985);
   U5641 : AOI22_X1 port map( A1 => n2418, A2 => n3522, B1 => n3995, B2 => 
                           n3583, ZN => n13546);
   U5642 : INV_X1 port map( A => n13674, ZN => n11989);
   U5643 : AOI22_X1 port map( A1 => n2418, A2 => n3524, B1 => n3995, B2 => 
                           n3559, ZN => n13674);
   U5644 : INV_X1 port map( A => n13547, ZN => n11945);
   U5645 : AOI22_X1 port map( A1 => n2424, A2 => n3522, B1 => n4001, B2 => 
                           n3584, ZN => n13547);
   U5646 : INV_X1 port map( A => n13675, ZN => n11949);
   U5647 : AOI22_X1 port map( A1 => n2424, A2 => n3526, B1 => n4001, B2 => 
                           n3559, ZN => n13675);
   U5648 : INV_X1 port map( A => n13548, ZN => n11905);
   U5649 : AOI22_X1 port map( A1 => n2430, A2 => n3522, B1 => n4007, B2 => 
                           n3584, ZN => n13548);
   U5650 : INV_X1 port map( A => n13676, ZN => n11909);
   U5651 : AOI22_X1 port map( A1 => n2430, A2 => n3523, B1 => n4007, B2 => 
                           n3559, ZN => n13676);
   U5652 : INV_X1 port map( A => n13549, ZN => n11865);
   U5653 : AOI22_X1 port map( A1 => n2436, A2 => n3522, B1 => n4013, B2 => 
                           n3584, ZN => n13549);
   U5654 : INV_X1 port map( A => n13677, ZN => n11869);
   U5655 : AOI22_X1 port map( A1 => n2436, A2 => n3526, B1 => n4013, B2 => 
                           n3559, ZN => n13677);
   U5656 : INV_X1 port map( A => n13550, ZN => n11825);
   U5657 : AOI22_X1 port map( A1 => n2442, A2 => n3522, B1 => n4019, B2 => 
                           n3584, ZN => n13550);
   U5658 : INV_X1 port map( A => n13678, ZN => n11829);
   U5659 : AOI22_X1 port map( A1 => n2442, A2 => n3522, B1 => n4019, B2 => 
                           n3560, ZN => n13678);
   U5660 : INV_X1 port map( A => n13551, ZN => n11785);
   U5661 : AOI22_X1 port map( A1 => n2448, A2 => n3525, B1 => n4025, B2 => 
                           n3585, ZN => n13551);
   U5662 : INV_X1 port map( A => n13679, ZN => n11789);
   U5663 : AOI22_X1 port map( A1 => n2448, A2 => n3526, B1 => n4025, B2 => 
                           n3560, ZN => n13679);
   U5664 : INV_X1 port map( A => n13552, ZN => n11745);
   U5665 : AOI22_X1 port map( A1 => n2454, A2 => n3524, B1 => n4031, B2 => 
                           n3585, ZN => n13552);
   U5666 : INV_X1 port map( A => n13680, ZN => n11749);
   U5667 : AOI22_X1 port map( A1 => n2454, A2 => n3520, B1 => n4031, B2 => 
                           n3560, ZN => n13680);
   U5668 : INV_X1 port map( A => n13553, ZN => n11705);
   U5669 : AOI22_X1 port map( A1 => n2460, A2 => n3525, B1 => n4037, B2 => 
                           n3585, ZN => n13553);
   U5670 : INV_X1 port map( A => n13554, ZN => n11665);
   U5671 : AOI22_X1 port map( A1 => n2466, A2 => n3523, B1 => n4043, B2 => 
                           n3585, ZN => n13554);
   U5672 : INV_X1 port map( A => n13533, ZN => n12505);
   U5673 : AOI22_X1 port map( A1 => n2340, A2 => n3521, B1 => n4091, B2 => 
                           n3580, ZN => n13533);
   U5674 : INV_X1 port map( A => n13661, ZN => n12509);
   U5675 : AOI22_X1 port map( A1 => n2340, A2 => n3526, B1 => n4091, B2 => 
                           n3555, ZN => n13661);
   U5676 : INV_X1 port map( A => n13544, ZN => n12065);
   U5677 : AOI22_X1 port map( A1 => n2406, A2 => n3522, B1 => n4097, B2 => 
                           n3583, ZN => n13544);
   U5678 : INV_X1 port map( A => n13672, ZN => n12069);
   U5679 : AOI22_X1 port map( A1 => n2406, A2 => n3521, B1 => n4097, B2 => 
                           n3558, ZN => n13672);
   U5680 : INV_X1 port map( A => n13555, ZN => n11625);
   U5681 : AOI22_X1 port map( A1 => n2472, A2 => n3522, B1 => n4103, B2 => 
                           n3586, ZN => n13555);
   U5682 : INV_X1 port map( A => n13787, ZN => n12593);
   U5683 : AOI22_X1 port map( A1 => n2329, A2 => n3634, B1 => n3918, B2 => 
                           n3691, ZN => n13787);
   U5684 : INV_X1 port map( A => n13915, ZN => n12597);
   U5685 : AOI22_X1 port map( A1 => n2329, A2 => n3638, B1 => n3918, B2 => 
                           n3667, ZN => n13915);
   U5686 : INV_X1 port map( A => n13788, ZN => n12553);
   U5687 : AOI22_X1 port map( A1 => n2335, A2 => n3632, B1 => n3924, B2 => 
                           n3692, ZN => n13788);
   U5688 : INV_X1 port map( A => n13916, ZN => n12557);
   U5689 : AOI22_X1 port map( A1 => n2335, A2 => n3638, B1 => n3924, B2 => 
                           n3667, ZN => n13916);
   U5690 : INV_X1 port map( A => n13790, ZN => n12473);
   U5691 : AOI22_X1 port map( A1 => n2347, A2 => n3637, B1 => n3930, B2 => 
                           n3692, ZN => n13790);
   U5692 : INV_X1 port map( A => n13918, ZN => n12477);
   U5693 : AOI22_X1 port map( A1 => n2347, A2 => n3638, B1 => n3930, B2 => 
                           n3668, ZN => n13918);
   U5694 : INV_X1 port map( A => n13791, ZN => n12433);
   U5695 : AOI22_X1 port map( A1 => n2353, A2 => n3636, B1 => n3936, B2 => 
                           n3693, ZN => n13791);
   U5696 : INV_X1 port map( A => n13792, ZN => n12393);
   U5697 : AOI22_X1 port map( A1 => n2359, A2 => n3635, B1 => n3942, B2 => 
                           n3693, ZN => n13792);
   U5698 : INV_X1 port map( A => n13920, ZN => n12397);
   U5699 : AOI22_X1 port map( A1 => n2359, A2 => n3638, B1 => n3942, B2 => 
                           n3668, ZN => n13920);
   U5700 : INV_X1 port map( A => n13793, ZN => n12353);
   U5701 : AOI22_X1 port map( A1 => n2365, A2 => n3638, B1 => n3948, B2 => 
                           n3693, ZN => n13793);
   U5702 : INV_X1 port map( A => n13921, ZN => n12357);
   U5703 : AOI22_X1 port map( A1 => n2365, A2 => n3638, B1 => n3948, B2 => 
                           n3668, ZN => n13921);
   U5704 : INV_X1 port map( A => n13794, ZN => n12313);
   U5705 : AOI22_X1 port map( A1 => n2371, A2 => n3633, B1 => n3954, B2 => 
                           n3693, ZN => n13794);
   U5706 : INV_X1 port map( A => n13922, ZN => n12317);
   U5707 : AOI22_X1 port map( A1 => n2371, A2 => n3638, B1 => n3954, B2 => 
                           n3669, ZN => n13922);
   U5708 : INV_X1 port map( A => n13795, ZN => n12273);
   U5709 : AOI22_X1 port map( A1 => n2377, A2 => n3634, B1 => n3960, B2 => 
                           n3694, ZN => n13795);
   U5710 : INV_X1 port map( A => n13923, ZN => n12277);
   U5711 : AOI22_X1 port map( A1 => n2377, A2 => n3632, B1 => n3960, B2 => 
                           n3669, ZN => n13923);
   U5712 : INV_X1 port map( A => n13796, ZN => n12233);
   U5713 : AOI22_X1 port map( A1 => n2383, A2 => n3633, B1 => n3966, B2 => 
                           n3694, ZN => n13796);
   U5714 : INV_X1 port map( A => n13924, ZN => n12237);
   U5715 : AOI22_X1 port map( A1 => n2383, A2 => n3633, B1 => n3966, B2 => 
                           n3669, ZN => n13924);
   U5716 : INV_X1 port map( A => n13797, ZN => n12193);
   U5717 : AOI22_X1 port map( A1 => n2389, A2 => n3633, B1 => n3972, B2 => 
                           n3694, ZN => n13797);
   U5718 : INV_X1 port map( A => n13925, ZN => n12197);
   U5719 : AOI22_X1 port map( A1 => n2389, A2 => n3638, B1 => n3972, B2 => 
                           n3669, ZN => n13925);
   U5720 : INV_X1 port map( A => n13798, ZN => n12153);
   U5721 : AOI22_X1 port map( A1 => n2395, A2 => n3633, B1 => n3978, B2 => 
                           n3694, ZN => n13798);
   U5722 : INV_X1 port map( A => n13926, ZN => n12157);
   U5723 : AOI22_X1 port map( A1 => n2395, A2 => n3638, B1 => n3978, B2 => 
                           n3670, ZN => n13926);
   U5724 : INV_X1 port map( A => n13799, ZN => n12113);
   U5725 : AOI22_X1 port map( A1 => n2401, A2 => n3633, B1 => n3984, B2 => 
                           n3695, ZN => n13799);
   U5726 : INV_X1 port map( A => n13927, ZN => n12117);
   U5727 : AOI22_X1 port map( A1 => n2401, A2 => n3638, B1 => n3984, B2 => 
                           n3670, ZN => n13927);
   U5728 : INV_X1 port map( A => n13801, ZN => n12033);
   U5729 : AOI22_X1 port map( A1 => n2413, A2 => n3633, B1 => n3990, B2 => 
                           n3695, ZN => n13801);
   U5730 : INV_X1 port map( A => n13929, ZN => n12037);
   U5731 : AOI22_X1 port map( A1 => n2413, A2 => n3637, B1 => n3990, B2 => 
                           n3670, ZN => n13929);
   U5732 : INV_X1 port map( A => n13802, ZN => n11993);
   U5733 : AOI22_X1 port map( A1 => n2419, A2 => n3633, B1 => n3996, B2 => 
                           n3695, ZN => n13802);
   U5734 : INV_X1 port map( A => n13930, ZN => n11997);
   U5735 : AOI22_X1 port map( A1 => n2419, A2 => n3636, B1 => n3996, B2 => 
                           n3671, ZN => n13930);
   U5736 : INV_X1 port map( A => n13803, ZN => n11953);
   U5737 : AOI22_X1 port map( A1 => n2425, A2 => n3633, B1 => n4002, B2 => 
                           n3696, ZN => n13803);
   U5738 : INV_X1 port map( A => n13931, ZN => n11957);
   U5739 : AOI22_X1 port map( A1 => n2425, A2 => n3638, B1 => n4002, B2 => 
                           n3671, ZN => n13931);
   U5740 : INV_X1 port map( A => n13804, ZN => n11913);
   U5741 : AOI22_X1 port map( A1 => n2431, A2 => n3633, B1 => n4008, B2 => 
                           n3696, ZN => n13804);
   U5742 : INV_X1 port map( A => n13932, ZN => n11917);
   U5743 : AOI22_X1 port map( A1 => n2431, A2 => n3635, B1 => n4008, B2 => 
                           n3671, ZN => n13932);
   U5744 : INV_X1 port map( A => n13805, ZN => n11873);
   U5745 : AOI22_X1 port map( A1 => n2437, A2 => n3633, B1 => n4014, B2 => 
                           n3696, ZN => n13805);
   U5746 : INV_X1 port map( A => n13933, ZN => n11877);
   U5747 : AOI22_X1 port map( A1 => n2437, A2 => n3638, B1 => n4014, B2 => 
                           n3671, ZN => n13933);
   U5748 : INV_X1 port map( A => n13806, ZN => n11833);
   U5749 : AOI22_X1 port map( A1 => n2443, A2 => n3633, B1 => n4020, B2 => 
                           n3696, ZN => n13806);
   U5750 : INV_X1 port map( A => n13934, ZN => n11837);
   U5751 : AOI22_X1 port map( A1 => n2443, A2 => n3633, B1 => n4020, B2 => 
                           n3672, ZN => n13934);
   U5752 : INV_X1 port map( A => n13807, ZN => n11793);
   U5753 : AOI22_X1 port map( A1 => n2449, A2 => n3637, B1 => n4026, B2 => 
                           n3697, ZN => n13807);
   U5754 : INV_X1 port map( A => n13935, ZN => n11797);
   U5755 : AOI22_X1 port map( A1 => n2449, A2 => n3638, B1 => n4026, B2 => 
                           n3672, ZN => n13935);
   U5756 : INV_X1 port map( A => n13808, ZN => n11753);
   U5757 : AOI22_X1 port map( A1 => n2455, A2 => n3636, B1 => n4032, B2 => 
                           n3697, ZN => n13808);
   U5758 : INV_X1 port map( A => n13936, ZN => n11757);
   U5759 : AOI22_X1 port map( A1 => n2455, A2 => n3634, B1 => n4032, B2 => 
                           n3672, ZN => n13936);
   U5760 : INV_X1 port map( A => n13809, ZN => n11713);
   U5761 : AOI22_X1 port map( A1 => n2461, A2 => n3637, B1 => n4038, B2 => 
                           n3697, ZN => n13809);
   U5762 : INV_X1 port map( A => n13810, ZN => n11673);
   U5763 : AOI22_X1 port map( A1 => n2467, A2 => n3635, B1 => n4044, B2 => 
                           n3697, ZN => n13810);
   U5764 : INV_X1 port map( A => n13789, ZN => n12513);
   U5765 : AOI22_X1 port map( A1 => n2341, A2 => n3632, B1 => n4092, B2 => 
                           n3692, ZN => n13789);
   U5766 : INV_X1 port map( A => n13917, ZN => n12517);
   U5767 : AOI22_X1 port map( A1 => n2341, A2 => n3638, B1 => n4092, B2 => 
                           n3667, ZN => n13917);
   U5768 : INV_X1 port map( A => n13800, ZN => n12073);
   U5769 : AOI22_X1 port map( A1 => n2407, A2 => n3633, B1 => n4098, B2 => 
                           n3695, ZN => n13800);
   U5770 : INV_X1 port map( A => n13928, ZN => n12077);
   U5771 : AOI22_X1 port map( A1 => n2407, A2 => n3632, B1 => n4098, B2 => 
                           n3670, ZN => n13928);
   U5772 : INV_X1 port map( A => n13811, ZN => n11633);
   U5773 : AOI22_X1 port map( A1 => n2473, A2 => n3633, B1 => n4104, B2 => 
                           n3698, ZN => n13811);
   U5774 : INV_X1 port map( A => n14043, ZN => n12601);
   U5775 : AOI22_X1 port map( A1 => n2329, A2 => n3743, B1 => n3918, B2 => 
                           n3803, ZN => n14043);
   U5776 : INV_X1 port map( A => n14171, ZN => n12605);
   U5777 : AOI22_X1 port map( A1 => n2330, A2 => n3748, B1 => n3919, B2 => 
                           n3779, ZN => n14171);
   U5778 : INV_X1 port map( A => n14044, ZN => n12561);
   U5779 : AOI22_X1 port map( A1 => n2335, A2 => n3743, B1 => n3924, B2 => 
                           n3804, ZN => n14044);
   U5780 : INV_X1 port map( A => n14172, ZN => n12565);
   U5781 : AOI22_X1 port map( A1 => n2336, A2 => n3749, B1 => n3925, B2 => 
                           n3779, ZN => n14172);
   U5782 : INV_X1 port map( A => n14046, ZN => n12481);
   U5783 : AOI22_X1 port map( A1 => n2347, A2 => n3743, B1 => n3930, B2 => 
                           n3804, ZN => n14046);
   U5784 : INV_X1 port map( A => n14174, ZN => n12485);
   U5785 : AOI22_X1 port map( A1 => n2348, A2 => n3749, B1 => n3931, B2 => 
                           n3780, ZN => n14174);
   U5786 : INV_X1 port map( A => n14047, ZN => n12441);
   U5787 : AOI22_X1 port map( A1 => n2353, A2 => n3743, B1 => n3936, B2 => 
                           n3805, ZN => n14047);
   U5788 : INV_X1 port map( A => n14048, ZN => n12401);
   U5789 : AOI22_X1 port map( A1 => n2359, A2 => n3743, B1 => n3942, B2 => 
                           n3805, ZN => n14048);
   U5790 : INV_X1 port map( A => n14176, ZN => n12405);
   U5791 : AOI22_X1 port map( A1 => n2360, A2 => n3749, B1 => n3943, B2 => 
                           n3780, ZN => n14176);
   U5792 : INV_X1 port map( A => n14049, ZN => n12361);
   U5793 : AOI22_X1 port map( A1 => n2365, A2 => n3743, B1 => n3948, B2 => 
                           n3805, ZN => n14049);
   U5794 : INV_X1 port map( A => n14177, ZN => n12365);
   U5795 : AOI22_X1 port map( A1 => n2366, A2 => n3749, B1 => n3949, B2 => 
                           n3780, ZN => n14177);
   U5796 : INV_X1 port map( A => n14050, ZN => n12321);
   U5797 : AOI22_X1 port map( A1 => n2371, A2 => n3743, B1 => n3954, B2 => 
                           n3805, ZN => n14050);
   U5798 : INV_X1 port map( A => n14178, ZN => n12325);
   U5799 : AOI22_X1 port map( A1 => n2372, A2 => n3749, B1 => n3955, B2 => 
                           n3781, ZN => n14178);
   U5800 : INV_X1 port map( A => n14051, ZN => n12281);
   U5801 : AOI22_X1 port map( A1 => n2377, A2 => n3743, B1 => n3960, B2 => 
                           n3806, ZN => n14051);
   U5802 : INV_X1 port map( A => n14179, ZN => n12285);
   U5803 : AOI22_X1 port map( A1 => n2378, A2 => n3746, B1 => n3961, B2 => 
                           n3781, ZN => n14179);
   U5804 : INV_X1 port map( A => n14052, ZN => n12241);
   U5805 : AOI22_X1 port map( A1 => n2383, A2 => n3744, B1 => n3966, B2 => 
                           n3806, ZN => n14052);
   U5806 : INV_X1 port map( A => n14180, ZN => n12245);
   U5807 : AOI22_X1 port map( A1 => n2384, A2 => n3747, B1 => n3967, B2 => 
                           n3781, ZN => n14180);
   U5808 : INV_X1 port map( A => n14053, ZN => n12201);
   U5809 : AOI22_X1 port map( A1 => n2389, A2 => n3745, B1 => n3972, B2 => 
                           n3806, ZN => n14053);
   U5810 : INV_X1 port map( A => n14181, ZN => n12205);
   U5811 : AOI22_X1 port map( A1 => n2390, A2 => n3749, B1 => n3973, B2 => 
                           n3781, ZN => n14181);
   U5812 : INV_X1 port map( A => n14054, ZN => n12161);
   U5813 : AOI22_X1 port map( A1 => n2395, A2 => n3747, B1 => n3978, B2 => 
                           n3806, ZN => n14054);
   U5814 : INV_X1 port map( A => n14182, ZN => n12165);
   U5815 : AOI22_X1 port map( A1 => n2396, A2 => n3750, B1 => n3979, B2 => 
                           n3782, ZN => n14182);
   U5816 : INV_X1 port map( A => n14055, ZN => n12121);
   U5817 : AOI22_X1 port map( A1 => n2401, A2 => n3746, B1 => n3984, B2 => 
                           n3807, ZN => n14055);
   U5818 : INV_X1 port map( A => n14183, ZN => n12125);
   U5819 : AOI22_X1 port map( A1 => n2402, A2 => n3749, B1 => n3985, B2 => 
                           n3782, ZN => n14183);
   U5820 : INV_X1 port map( A => n14057, ZN => n12041);
   U5821 : AOI22_X1 port map( A1 => n2413, A2 => n3749, B1 => n3990, B2 => 
                           n3807, ZN => n14057);
   U5822 : INV_X1 port map( A => n14185, ZN => n12045);
   U5823 : AOI22_X1 port map( A1 => n2414, A2 => n3750, B1 => n3991, B2 => 
                           n3782, ZN => n14185);
   U5824 : INV_X1 port map( A => n14058, ZN => n12001);
   U5825 : AOI22_X1 port map( A1 => n2419, A2 => n3750, B1 => n3996, B2 => 
                           n3807, ZN => n14058);
   U5826 : INV_X1 port map( A => n14186, ZN => n12005);
   U5827 : AOI22_X1 port map( A1 => n2420, A2 => n3750, B1 => n3997, B2 => 
                           n3783, ZN => n14186);
   U5828 : INV_X1 port map( A => n14059, ZN => n11961);
   U5829 : AOI22_X1 port map( A1 => n2425, A2 => n3748, B1 => n4002, B2 => 
                           n3808, ZN => n14059);
   U5830 : INV_X1 port map( A => n14187, ZN => n11965);
   U5831 : AOI22_X1 port map( A1 => n2426, A2 => n3749, B1 => n4003, B2 => 
                           n3783, ZN => n14187);
   U5832 : INV_X1 port map( A => n14060, ZN => n11921);
   U5833 : AOI22_X1 port map( A1 => n2431, A2 => n3744, B1 => n4008, B2 => 
                           n3808, ZN => n14060);
   U5834 : INV_X1 port map( A => n14188, ZN => n11925);
   U5835 : AOI22_X1 port map( A1 => n2432, A2 => n3750, B1 => n4009, B2 => 
                           n3783, ZN => n14188);
   U5836 : INV_X1 port map( A => n14061, ZN => n11881);
   U5837 : AOI22_X1 port map( A1 => n2437, A2 => n3745, B1 => n4014, B2 => 
                           n3808, ZN => n14061);
   U5838 : INV_X1 port map( A => n14189, ZN => n11885);
   U5839 : AOI22_X1 port map( A1 => n2438, A2 => n3749, B1 => n4015, B2 => 
                           n3783, ZN => n14189);
   U5840 : INV_X1 port map( A => n14062, ZN => n11841);
   U5841 : AOI22_X1 port map( A1 => n2443, A2 => n3749, B1 => n4020, B2 => 
                           n3808, ZN => n14062);
   U5842 : INV_X1 port map( A => n14190, ZN => n11845);
   U5843 : AOI22_X1 port map( A1 => n2444, A2 => n3750, B1 => n4021, B2 => 
                           n3784, ZN => n14190);
   U5844 : INV_X1 port map( A => n14063, ZN => n11801);
   U5845 : AOI22_X1 port map( A1 => n2449, A2 => n3748, B1 => n4026, B2 => 
                           n3809, ZN => n14063);
   U5846 : INV_X1 port map( A => n14191, ZN => n11805);
   U5847 : AOI22_X1 port map( A1 => n2450, A2 => n3749, B1 => n4027, B2 => 
                           n3784, ZN => n14191);
   U5848 : INV_X1 port map( A => n14064, ZN => n11761);
   U5849 : AOI22_X1 port map( A1 => n2455, A2 => n3747, B1 => n4032, B2 => 
                           n3809, ZN => n14064);
   U5850 : INV_X1 port map( A => n14192, ZN => n11765);
   U5851 : AOI22_X1 port map( A1 => n2456, A2 => n3750, B1 => n4033, B2 => 
                           n3784, ZN => n14192);
   U5852 : INV_X1 port map( A => n14065, ZN => n11721);
   U5853 : AOI22_X1 port map( A1 => n2461, A2 => n3746, B1 => n4038, B2 => 
                           n3809, ZN => n14065);
   U5854 : INV_X1 port map( A => n14066, ZN => n11681);
   U5855 : AOI22_X1 port map( A1 => n2467, A2 => n3749, B1 => n4044, B2 => 
                           n3809, ZN => n14066);
   U5856 : INV_X1 port map( A => n14045, ZN => n12521);
   U5857 : AOI22_X1 port map( A1 => n2341, A2 => n3743, B1 => n4092, B2 => 
                           n3804, ZN => n14045);
   U5858 : INV_X1 port map( A => n14173, ZN => n12525);
   U5859 : AOI22_X1 port map( A1 => n2342, A2 => n3749, B1 => n4093, B2 => 
                           n3779, ZN => n14173);
   U5860 : INV_X1 port map( A => n14056, ZN => n12081);
   U5861 : AOI22_X1 port map( A1 => n2407, A2 => n3747, B1 => n4098, B2 => 
                           n3807, ZN => n14056);
   U5862 : INV_X1 port map( A => n14184, ZN => n12085);
   U5863 : AOI22_X1 port map( A1 => n2408, A2 => n3750, B1 => n4099, B2 => 
                           n3782, ZN => n14184);
   U5864 : INV_X1 port map( A => n14067, ZN => n11641);
   U5865 : AOI22_X1 port map( A1 => n2473, A2 => n3750, B1 => n4104, B2 => 
                           n3810, ZN => n14067);
   U5866 : INV_X1 port map( A => n13425, ZN => n11701);
   U5867 : AOI22_X1 port map( A1 => n2460, A2 => n3415, B1 => n4037, B2 => 
                           n3448, ZN => n13425);
   U5868 : INV_X1 port map( A => n13426, ZN => n11661);
   U5869 : AOI22_X1 port map( A1 => n2466, A2 => n3415, B1 => n4043, B2 => 
                           n3449, ZN => n13426);
   U5870 : INV_X1 port map( A => n13427, ZN => n11621);
   U5871 : AOI22_X1 port map( A1 => n2472, A2 => n3415, B1 => n4103, B2 => 
                           n3449, ZN => n13427);
   U5872 : INV_X1 port map( A => n13681, ZN => n11709);
   U5873 : AOI22_X1 port map( A1 => n2460, A2 => n3527, B1 => n4037, B2 => 
                           n3560, ZN => n13681);
   U5874 : INV_X1 port map( A => n13682, ZN => n11669);
   U5875 : AOI22_X1 port map( A1 => n2466, A2 => n3527, B1 => n4043, B2 => 
                           n3561, ZN => n13682);
   U5876 : INV_X1 port map( A => n13683, ZN => n11629);
   U5877 : AOI22_X1 port map( A1 => n2472, A2 => n3527, B1 => n4103, B2 => 
                           n3561, ZN => n13683);
   U5878 : INV_X1 port map( A => n13937, ZN => n11717);
   U5879 : AOI22_X1 port map( A1 => n2461, A2 => n3639, B1 => n4038, B2 => 
                           n3672, ZN => n13937);
   U5880 : INV_X1 port map( A => n13938, ZN => n11677);
   U5881 : AOI22_X1 port map( A1 => n2467, A2 => n3639, B1 => n4044, B2 => 
                           n3673, ZN => n13938);
   U5882 : INV_X1 port map( A => n13939, ZN => n11637);
   U5883 : AOI22_X1 port map( A1 => n2473, A2 => n3639, B1 => n4104, B2 => 
                           n3673, ZN => n13939);
   U5884 : INV_X1 port map( A => n14193, ZN => n11725);
   U5885 : AOI22_X1 port map( A1 => n2462, A2 => n3751, B1 => n4039, B2 => 
                           n3784, ZN => n14193);
   U5886 : INV_X1 port map( A => n14194, ZN => n11685);
   U5887 : AOI22_X1 port map( A1 => n2468, A2 => n3751, B1 => n4045, B2 => 
                           n3785, ZN => n14194);
   U5888 : INV_X1 port map( A => n14195, ZN => n11645);
   U5889 : AOI22_X1 port map( A1 => n2474, A2 => n3751, B1 => n4105, B2 => 
                           n3785, ZN => n14195);
   U5890 : INV_X1 port map( A => n13019, ZN => n12569);
   U5891 : AOI22_X1 port map( A1 => n2327, A2 => n3297, B1 => n3916, B2 => 
                           n3349, ZN => n13019);
   U5892 : INV_X1 port map( A => n13020, ZN => n12529);
   U5893 : AOI22_X1 port map( A1 => n2333, A2 => n3298, B1 => n3922, B2 => 
                           n3349, ZN => n13020);
   U5894 : INV_X1 port map( A => n13148, ZN => n12533);
   U5895 : AOI22_X1 port map( A1 => n2333, A2 => n3304, B1 => n3922, B2 => 
                           n3325, ZN => n13148);
   U5896 : INV_X1 port map( A => n13022, ZN => n12449);
   U5897 : AOI22_X1 port map( A1 => n2345, A2 => n3296, B1 => n3928, B2 => 
                           n3350, ZN => n13022);
   U5898 : INV_X1 port map( A => n13150, ZN => n12453);
   U5899 : AOI22_X1 port map( A1 => n2345, A2 => n3301, B1 => n3928, B2 => 
                           n3324, ZN => n13150);
   U5900 : INV_X1 port map( A => n13023, ZN => n12409);
   U5901 : AOI22_X1 port map( A1 => n2351, A2 => n3299, B1 => n3934, B2 => 
                           n3350, ZN => n13023);
   U5902 : INV_X1 port map( A => n13151, ZN => n12413);
   U5903 : AOI22_X1 port map( A1 => n2351, A2 => n3297, B1 => n3934, B2 => 
                           n3326, ZN => n13151);
   U5904 : INV_X1 port map( A => n13024, ZN => n12369);
   U5905 : AOI22_X1 port map( A1 => n2357, A2 => n3300, B1 => n3940, B2 => 
                           n3350, ZN => n13024);
   U5906 : INV_X1 port map( A => n13152, ZN => n12373);
   U5907 : AOI22_X1 port map( A1 => n2357, A2 => n3298, B1 => n3940, B2 => 
                           n3325, ZN => n13152);
   U5908 : INV_X1 port map( A => n13025, ZN => n12329);
   U5909 : AOI22_X1 port map( A1 => n2363, A2 => n3302, B1 => n3946, B2 => 
                           n3351, ZN => n13025);
   U5910 : INV_X1 port map( A => n13153, ZN => n12333);
   U5911 : AOI22_X1 port map( A1 => n2363, A2 => n3302, B1 => n3946, B2 => 
                           n3325, ZN => n13153);
   U5912 : INV_X1 port map( A => n13026, ZN => n12289);
   U5913 : AOI22_X1 port map( A1 => n2369, A2 => n3297, B1 => n3952, B2 => 
                           n3351, ZN => n13026);
   U5914 : INV_X1 port map( A => n13154, ZN => n12293);
   U5915 : AOI22_X1 port map( A1 => n2369, A2 => n3302, B1 => n3952, B2 => 
                           n3327, ZN => n13154);
   U5916 : INV_X1 port map( A => n13027, ZN => n12249);
   U5917 : AOI22_X1 port map( A1 => n2375, A2 => n3298, B1 => n3958, B2 => 
                           n3351, ZN => n13027);
   U5918 : INV_X1 port map( A => n13155, ZN => n12253);
   U5919 : AOI22_X1 port map( A1 => n2375, A2 => n3302, B1 => n3958, B2 => 
                           n3326, ZN => n13155);
   U5920 : INV_X1 port map( A => n13028, ZN => n12209);
   U5921 : AOI22_X1 port map( A1 => n2381, A2 => n3296, B1 => n3964, B2 => 
                           n3351, ZN => n13028);
   U5922 : INV_X1 port map( A => n13156, ZN => n12213);
   U5923 : AOI22_X1 port map( A1 => n2381, A2 => n3302, B1 => n3964, B2 => 
                           n3326, ZN => n13156);
   U5924 : INV_X1 port map( A => n13029, ZN => n12169);
   U5925 : AOI22_X1 port map( A1 => n2387, A2 => n3297, B1 => n3970, B2 => 
                           n3352, ZN => n13029);
   U5926 : INV_X1 port map( A => n13157, ZN => n12173);
   U5927 : AOI22_X1 port map( A1 => n2387, A2 => n3302, B1 => n3970, B2 => 
                           n3327, ZN => n13157);
   U5928 : INV_X1 port map( A => n13030, ZN => n12129);
   U5929 : AOI22_X1 port map( A1 => n2393, A2 => n3297, B1 => n3976, B2 => 
                           n3352, ZN => n13030);
   U5930 : INV_X1 port map( A => n13158, ZN => n12133);
   U5931 : AOI22_X1 port map( A1 => n2393, A2 => n3302, B1 => n3976, B2 => 
                           n3327, ZN => n13158);
   U5932 : INV_X1 port map( A => n13031, ZN => n12089);
   U5933 : AOI22_X1 port map( A1 => n2399, A2 => n3297, B1 => n3982, B2 => 
                           n3352, ZN => n13031);
   U5934 : INV_X1 port map( A => n13159, ZN => n12093);
   U5935 : AOI22_X1 port map( A1 => n2399, A2 => n3302, B1 => n3982, B2 => 
                           n3328, ZN => n13159);
   U5936 : INV_X1 port map( A => n13033, ZN => n12009);
   U5937 : AOI22_X1 port map( A1 => n2411, A2 => n3297, B1 => n3988, B2 => 
                           n3353, ZN => n13033);
   U5938 : INV_X1 port map( A => n13161, ZN => n12013);
   U5939 : AOI22_X1 port map( A1 => n2411, A2 => n3302, B1 => n3988, B2 => 
                           n3328, ZN => n13161);
   U5940 : INV_X1 port map( A => n13034, ZN => n11969);
   U5941 : AOI22_X1 port map( A1 => n2417, A2 => n3297, B1 => n3994, B2 => 
                           n3353, ZN => n13034);
   U5942 : INV_X1 port map( A => n13162, ZN => n11973);
   U5943 : AOI22_X1 port map( A1 => n2417, A2 => n3302, B1 => n3994, B2 => 
                           n3328, ZN => n13162);
   U5944 : INV_X1 port map( A => n13035, ZN => n11929);
   U5945 : AOI22_X1 port map( A1 => n2423, A2 => n3297, B1 => n4000, B2 => 
                           n3353, ZN => n13035);
   U5946 : INV_X1 port map( A => n13163, ZN => n11933);
   U5947 : AOI22_X1 port map( A1 => n2423, A2 => n3302, B1 => n4000, B2 => 
                           n3329, ZN => n13163);
   U5948 : INV_X1 port map( A => n13036, ZN => n11889);
   U5949 : AOI22_X1 port map( A1 => n2429, A2 => n3297, B1 => n4006, B2 => 
                           n3353, ZN => n13036);
   U5950 : INV_X1 port map( A => n13164, ZN => n11893);
   U5951 : AOI22_X1 port map( A1 => n2429, A2 => n3302, B1 => n4006, B2 => 
                           n3329, ZN => n13164);
   U5952 : INV_X1 port map( A => n13037, ZN => n11849);
   U5953 : AOI22_X1 port map( A1 => n2435, A2 => n3297, B1 => n4012, B2 => 
                           n3354, ZN => n13037);
   U5954 : INV_X1 port map( A => n13165, ZN => n11853);
   U5955 : AOI22_X1 port map( A1 => n2435, A2 => n3297, B1 => n4012, B2 => 
                           n3329, ZN => n13165);
   U5956 : INV_X1 port map( A => n13038, ZN => n11809);
   U5957 : AOI22_X1 port map( A1 => n2441, A2 => n3297, B1 => n4018, B2 => 
                           n3354, ZN => n13038);
   U5958 : INV_X1 port map( A => n13166, ZN => n11813);
   U5959 : AOI22_X1 port map( A1 => n2441, A2 => n3298, B1 => n4018, B2 => 
                           n3329, ZN => n13166);
   U5960 : INV_X1 port map( A => n13039, ZN => n11769);
   U5961 : AOI22_X1 port map( A1 => n2447, A2 => n3297, B1 => n4024, B2 => 
                           n3354, ZN => n13039);
   U5962 : INV_X1 port map( A => n13167, ZN => n11773);
   U5963 : AOI22_X1 port map( A1 => n2447, A2 => n3301, B1 => n4024, B2 => 
                           n3330, ZN => n13167);
   U5964 : INV_X1 port map( A => n13040, ZN => n11729);
   U5965 : AOI22_X1 port map( A1 => n2453, A2 => n3297, B1 => n4030, B2 => 
                           n3354, ZN => n13040);
   U5966 : INV_X1 port map( A => n13168, ZN => n11733);
   U5967 : AOI22_X1 port map( A1 => n2453, A2 => n3305, B1 => n4030, B2 => 
                           n3330, ZN => n13168);
   U5968 : INV_X1 port map( A => n13041, ZN => n11689);
   U5969 : AOI22_X1 port map( A1 => n2459, A2 => n3296, B1 => n4036, B2 => 
                           n3355, ZN => n13041);
   U5970 : INV_X1 port map( A => n13169, ZN => n11693);
   U5971 : AOI22_X1 port map( A1 => n2459, A2 => n3302, B1 => n4036, B2 => 
                           n3330, ZN => n13169);
   U5972 : INV_X1 port map( A => n13042, ZN => n11649);
   U5973 : AOI22_X1 port map( A1 => n2465, A2 => n3296, B1 => n4042, B2 => 
                           n3355, ZN => n13042);
   U5974 : INV_X1 port map( A => n13170, ZN => n11653);
   U5975 : AOI22_X1 port map( A1 => n2465, A2 => n3296, B1 => n4042, B2 => 
                           n3330, ZN => n13170);
   U5976 : INV_X1 port map( A => n13021, ZN => n12489);
   U5977 : AOI22_X1 port map( A1 => n2339, A2 => n3299, B1 => n4090, B2 => 
                           n3350, ZN => n13021);
   U5978 : INV_X1 port map( A => n13149, ZN => n12493);
   U5979 : AOI22_X1 port map( A1 => n2339, A2 => n3296, B1 => n4090, B2 => 
                           n3323, ZN => n13149);
   U5980 : INV_X1 port map( A => n13032, ZN => n12049);
   U5981 : AOI22_X1 port map( A1 => n2405, A2 => n3297, B1 => n4096, B2 => 
                           n3352, ZN => n13032);
   U5982 : INV_X1 port map( A => n13160, ZN => n12053);
   U5983 : AOI22_X1 port map( A1 => n2405, A2 => n3302, B1 => n4096, B2 => 
                           n3328, ZN => n13160);
   U5984 : INV_X1 port map( A => n13171, ZN => n11613);
   U5985 : AOI22_X1 port map( A1 => n2471, A2 => n3299, B1 => n4102, B2 => 
                           n3331, ZN => n13171);
   U5986 : INV_X1 port map( A => n13043, ZN => n11609);
   U5987 : AOI22_X1 port map( A1 => n2471, A2 => n3296, B1 => n4102, B2 => 
                           n3355, ZN => n13043);
   U5988 : INV_X1 port map( A => n13243, ZN => n12576);
   U5989 : AOI22_X1 port map( A1 => n2327, A2 => n3408, B1 => n3916, B2 => 
                           n3461, ZN => n13243);
   U5990 : INV_X1 port map( A => n13371, ZN => n12580);
   U5991 : AOI22_X1 port map( A1 => n2328, A2 => n3414, B1 => n3917, B2 => 
                           n3435, ZN => n13371);
   U5992 : INV_X1 port map( A => n13244, ZN => n12536);
   U5993 : AOI22_X1 port map( A1 => n2333, A2 => n3410, B1 => n3922, B2 => 
                           n3461, ZN => n13244);
   U5994 : INV_X1 port map( A => n13372, ZN => n12540);
   U5995 : AOI22_X1 port map( A1 => n2334, A2 => n3414, B1 => n3923, B2 => 
                           n3437, ZN => n13372);
   U5996 : INV_X1 port map( A => n13246, ZN => n12456);
   U5997 : AOI22_X1 port map( A1 => n2345, A2 => n3412, B1 => n3928, B2 => 
                           n3462, ZN => n13246);
   U5998 : INV_X1 port map( A => n13374, ZN => n12460);
   U5999 : AOI22_X1 port map( A1 => n2346, A2 => n3413, B1 => n3929, B2 => 
                           n3436, ZN => n13374);
   U6000 : INV_X1 port map( A => n13375, ZN => n12420);
   U6001 : AOI22_X1 port map( A1 => n2352, A2 => n3412, B1 => n3935, B2 => 
                           n3438, ZN => n13375);
   U6002 : INV_X1 port map( A => n13248, ZN => n12376);
   U6003 : AOI22_X1 port map( A1 => n2357, A2 => n3413, B1 => n3940, B2 => 
                           n3462, ZN => n13248);
   U6004 : INV_X1 port map( A => n13376, ZN => n12380);
   U6005 : AOI22_X1 port map( A1 => n2358, A2 => n3412, B1 => n3941, B2 => 
                           n3437, ZN => n13376);
   U6006 : INV_X1 port map( A => n13249, ZN => n12336);
   U6007 : AOI22_X1 port map( A1 => n2363, A2 => n3409, B1 => n3946, B2 => 
                           n3463, ZN => n13249);
   U6008 : INV_X1 port map( A => n13377, ZN => n12340);
   U6009 : AOI22_X1 port map( A1 => n2364, A2 => n3412, B1 => n3947, B2 => 
                           n3437, ZN => n13377);
   U6010 : INV_X1 port map( A => n13250, ZN => n12296);
   U6011 : AOI22_X1 port map( A1 => n2369, A2 => n3414, B1 => n3952, B2 => 
                           n3463, ZN => n13250);
   U6012 : INV_X1 port map( A => n13378, ZN => n12300);
   U6013 : AOI22_X1 port map( A1 => n2370, A2 => n3412, B1 => n3953, B2 => 
                           n3439, ZN => n13378);
   U6014 : INV_X1 port map( A => n13251, ZN => n12256);
   U6015 : AOI22_X1 port map( A1 => n2375, A2 => n3411, B1 => n3958, B2 => 
                           n3463, ZN => n13251);
   U6016 : INV_X1 port map( A => n13379, ZN => n12260);
   U6017 : AOI22_X1 port map( A1 => n2376, A2 => n3412, B1 => n3959, B2 => 
                           n3438, ZN => n13379);
   U6018 : INV_X1 port map( A => n13252, ZN => n12216);
   U6019 : AOI22_X1 port map( A1 => n2381, A2 => n3413, B1 => n3964, B2 => 
                           n3463, ZN => n13252);
   U6020 : INV_X1 port map( A => n13380, ZN => n12220);
   U6021 : AOI22_X1 port map( A1 => n2382, A2 => n3413, B1 => n3965, B2 => 
                           n3438, ZN => n13380);
   U6022 : INV_X1 port map( A => n13253, ZN => n12176);
   U6023 : AOI22_X1 port map( A1 => n2387, A2 => n3412, B1 => n3970, B2 => 
                           n3464, ZN => n13253);
   U6024 : INV_X1 port map( A => n13381, ZN => n12180);
   U6025 : AOI22_X1 port map( A1 => n2388, A2 => n3413, B1 => n3971, B2 => 
                           n3439, ZN => n13381);
   U6026 : INV_X1 port map( A => n13254, ZN => n12136);
   U6027 : AOI22_X1 port map( A1 => n2393, A2 => n3411, B1 => n3976, B2 => 
                           n3464, ZN => n13254);
   U6028 : INV_X1 port map( A => n13382, ZN => n12140);
   U6029 : AOI22_X1 port map( A1 => n2394, A2 => n3412, B1 => n3977, B2 => 
                           n3439, ZN => n13382);
   U6030 : INV_X1 port map( A => n13255, ZN => n12096);
   U6031 : AOI22_X1 port map( A1 => n2399, A2 => n3414, B1 => n3982, B2 => 
                           n3464, ZN => n13255);
   U6032 : INV_X1 port map( A => n13383, ZN => n12100);
   U6033 : AOI22_X1 port map( A1 => n2400, A2 => n3413, B1 => n3983, B2 => 
                           n3440, ZN => n13383);
   U6034 : INV_X1 port map( A => n13257, ZN => n12016);
   U6035 : AOI22_X1 port map( A1 => n2411, A2 => n3417, B1 => n3988, B2 => 
                           n3465, ZN => n13257);
   U6036 : INV_X1 port map( A => n13385, ZN => n12020);
   U6037 : AOI22_X1 port map( A1 => n2412, A2 => n3413, B1 => n3989, B2 => 
                           n3440, ZN => n13385);
   U6038 : INV_X1 port map( A => n13258, ZN => n11976);
   U6039 : AOI22_X1 port map( A1 => n2417, A2 => n3416, B1 => n3994, B2 => 
                           n3465, ZN => n13258);
   U6040 : INV_X1 port map( A => n13386, ZN => n11980);
   U6041 : AOI22_X1 port map( A1 => n2418, A2 => n3412, B1 => n3995, B2 => 
                           n3440, ZN => n13386);
   U6042 : INV_X1 port map( A => n13259, ZN => n11936);
   U6043 : AOI22_X1 port map( A1 => n2423, A2 => n3416, B1 => n4000, B2 => 
                           n3465, ZN => n13259);
   U6044 : INV_X1 port map( A => n13387, ZN => n11940);
   U6045 : AOI22_X1 port map( A1 => n2424, A2 => n3413, B1 => n4001, B2 => 
                           n3441, ZN => n13387);
   U6046 : INV_X1 port map( A => n13260, ZN => n11896);
   U6047 : AOI22_X1 port map( A1 => n2429, A2 => n3415, B1 => n4006, B2 => 
                           n3465, ZN => n13260);
   U6048 : INV_X1 port map( A => n13388, ZN => n11900);
   U6049 : AOI22_X1 port map( A1 => n2430, A2 => n3413, B1 => n4007, B2 => 
                           n3441, ZN => n13388);
   U6050 : INV_X1 port map( A => n13261, ZN => n11856);
   U6051 : AOI22_X1 port map( A1 => n2435, A2 => n3417, B1 => n4012, B2 => 
                           n3466, ZN => n13261);
   U6052 : INV_X1 port map( A => n13262, ZN => n11816);
   U6053 : AOI22_X1 port map( A1 => n2441, A2 => n3415, B1 => n4018, B2 => 
                           n3466, ZN => n13262);
   U6054 : INV_X1 port map( A => n13390, ZN => n11820);
   U6055 : AOI22_X1 port map( A1 => n2442, A2 => n3413, B1 => n4019, B2 => 
                           n3441, ZN => n13390);
   U6056 : INV_X1 port map( A => n13263, ZN => n11776);
   U6057 : AOI22_X1 port map( A1 => n2447, A2 => n3407, B1 => n4024, B2 => 
                           n3466, ZN => n13263);
   U6058 : INV_X1 port map( A => n13391, ZN => n11780);
   U6059 : AOI22_X1 port map( A1 => n2448, A2 => n3413, B1 => n4025, B2 => 
                           n3442, ZN => n13391);
   U6060 : INV_X1 port map( A => n13264, ZN => n11736);
   U6061 : AOI22_X1 port map( A1 => n2453, A2 => n3408, B1 => n4030, B2 => 
                           n3466, ZN => n13264);
   U6062 : INV_X1 port map( A => n13392, ZN => n11740);
   U6063 : AOI22_X1 port map( A1 => n2454, A2 => n3409, B1 => n4031, B2 => 
                           n3442, ZN => n13392);
   U6064 : INV_X1 port map( A => n13265, ZN => n11696);
   U6065 : AOI22_X1 port map( A1 => n2459, A2 => n3411, B1 => n4036, B2 => 
                           n3467, ZN => n13265);
   U6066 : INV_X1 port map( A => n13393, ZN => n11700);
   U6067 : AOI22_X1 port map( A1 => n2460, A2 => n3413, B1 => n4037, B2 => 
                           n3442, ZN => n13393);
   U6068 : INV_X1 port map( A => n13266, ZN => n11656);
   U6069 : AOI22_X1 port map( A1 => n2465, A2 => n3414, B1 => n4042, B2 => 
                           n3467, ZN => n13266);
   U6070 : INV_X1 port map( A => n13394, ZN => n11660);
   U6071 : AOI22_X1 port map( A1 => n2466, A2 => n3413, B1 => n4043, B2 => 
                           n3442, ZN => n13394);
   U6072 : INV_X1 port map( A => n13245, ZN => n12496);
   U6073 : AOI22_X1 port map( A1 => n2339, A2 => n3412, B1 => n4090, B2 => 
                           n3462, ZN => n13245);
   U6074 : INV_X1 port map( A => n13373, ZN => n12500);
   U6075 : AOI22_X1 port map( A1 => n2340, A2 => n3412, B1 => n4091, B2 => 
                           n3435, ZN => n13373);
   U6076 : INV_X1 port map( A => n13256, ZN => n12056);
   U6077 : AOI22_X1 port map( A1 => n2405, A2 => n3417, B1 => n4096, B2 => 
                           n3464, ZN => n13256);
   U6078 : INV_X1 port map( A => n13384, ZN => n12060);
   U6079 : AOI22_X1 port map( A1 => n2406, A2 => n3413, B1 => n4097, B2 => 
                           n3440, ZN => n13384);
   U6080 : INV_X1 port map( A => n13267, ZN => n11616);
   U6081 : AOI22_X1 port map( A1 => n2471, A2 => n3410, B1 => n4102, B2 => 
                           n3467, ZN => n13267);
   U6082 : INV_X1 port map( A => n13395, ZN => n11620);
   U6083 : AOI22_X1 port map( A1 => n2472, A2 => n3412, B1 => n4103, B2 => 
                           n3443, ZN => n13395);
   U6084 : INV_X1 port map( A => n13499, ZN => n12584);
   U6085 : AOI22_X1 port map( A1 => n2328, A2 => n3519, B1 => n3917, B2 => 
                           n3573, ZN => n13499);
   U6086 : INV_X1 port map( A => n13627, ZN => n12588);
   U6087 : AOI22_X1 port map( A1 => n2328, A2 => n3526, B1 => n3917, B2 => 
                           n3547, ZN => n13627);
   U6088 : INV_X1 port map( A => n13500, ZN => n12544);
   U6089 : AOI22_X1 port map( A1 => n2334, A2 => n3522, B1 => n3923, B2 => 
                           n3573, ZN => n13500);
   U6090 : INV_X1 port map( A => n13628, ZN => n12548);
   U6091 : AOI22_X1 port map( A1 => n2334, A2 => n3526, B1 => n3923, B2 => 
                           n3549, ZN => n13628);
   U6092 : INV_X1 port map( A => n13502, ZN => n12464);
   U6093 : AOI22_X1 port map( A1 => n2346, A2 => n3524, B1 => n3929, B2 => 
                           n3574, ZN => n13502);
   U6094 : INV_X1 port map( A => n13630, ZN => n12468);
   U6095 : AOI22_X1 port map( A1 => n2346, A2 => n3525, B1 => n3929, B2 => 
                           n3548, ZN => n13630);
   U6096 : INV_X1 port map( A => n13631, ZN => n12428);
   U6097 : AOI22_X1 port map( A1 => n2352, A2 => n3524, B1 => n3935, B2 => 
                           n3550, ZN => n13631);
   U6098 : INV_X1 port map( A => n13504, ZN => n12384);
   U6099 : AOI22_X1 port map( A1 => n2358, A2 => n3525, B1 => n3941, B2 => 
                           n3574, ZN => n13504);
   U6100 : INV_X1 port map( A => n13632, ZN => n12388);
   U6101 : AOI22_X1 port map( A1 => n2358, A2 => n3524, B1 => n3941, B2 => 
                           n3549, ZN => n13632);
   U6102 : INV_X1 port map( A => n13505, ZN => n12344);
   U6103 : AOI22_X1 port map( A1 => n2364, A2 => n3521, B1 => n3947, B2 => 
                           n3575, ZN => n13505);
   U6104 : INV_X1 port map( A => n13633, ZN => n12348);
   U6105 : AOI22_X1 port map( A1 => n2364, A2 => n3524, B1 => n3947, B2 => 
                           n3549, ZN => n13633);
   U6106 : INV_X1 port map( A => n13506, ZN => n12304);
   U6107 : AOI22_X1 port map( A1 => n2370, A2 => n3526, B1 => n3953, B2 => 
                           n3575, ZN => n13506);
   U6108 : INV_X1 port map( A => n13634, ZN => n12308);
   U6109 : AOI22_X1 port map( A1 => n2370, A2 => n3524, B1 => n3953, B2 => 
                           n3551, ZN => n13634);
   U6110 : INV_X1 port map( A => n13507, ZN => n12264);
   U6111 : AOI22_X1 port map( A1 => n2376, A2 => n3523, B1 => n3959, B2 => 
                           n3575, ZN => n13507);
   U6112 : INV_X1 port map( A => n13635, ZN => n12268);
   U6113 : AOI22_X1 port map( A1 => n2376, A2 => n3524, B1 => n3959, B2 => 
                           n3550, ZN => n13635);
   U6114 : INV_X1 port map( A => n13508, ZN => n12224);
   U6115 : AOI22_X1 port map( A1 => n2382, A2 => n3525, B1 => n3965, B2 => 
                           n3575, ZN => n13508);
   U6116 : INV_X1 port map( A => n13636, ZN => n12228);
   U6117 : AOI22_X1 port map( A1 => n2382, A2 => n3525, B1 => n3965, B2 => 
                           n3550, ZN => n13636);
   U6118 : INV_X1 port map( A => n13509, ZN => n12184);
   U6119 : AOI22_X1 port map( A1 => n2388, A2 => n3524, B1 => n3971, B2 => 
                           n3576, ZN => n13509);
   U6120 : INV_X1 port map( A => n13637, ZN => n12188);
   U6121 : AOI22_X1 port map( A1 => n2388, A2 => n3525, B1 => n3971, B2 => 
                           n3551, ZN => n13637);
   U6122 : INV_X1 port map( A => n13510, ZN => n12144);
   U6123 : AOI22_X1 port map( A1 => n2394, A2 => n3523, B1 => n3977, B2 => 
                           n3576, ZN => n13510);
   U6124 : INV_X1 port map( A => n13638, ZN => n12148);
   U6125 : AOI22_X1 port map( A1 => n2394, A2 => n3524, B1 => n3977, B2 => 
                           n3551, ZN => n13638);
   U6126 : INV_X1 port map( A => n13511, ZN => n12104);
   U6127 : AOI22_X1 port map( A1 => n2400, A2 => n3526, B1 => n3983, B2 => 
                           n3576, ZN => n13511);
   U6128 : INV_X1 port map( A => n13639, ZN => n12108);
   U6129 : AOI22_X1 port map( A1 => n2400, A2 => n3525, B1 => n3983, B2 => 
                           n3552, ZN => n13639);
   U6130 : INV_X1 port map( A => n13513, ZN => n12024);
   U6131 : AOI22_X1 port map( A1 => n2412, A2 => n3528, B1 => n3989, B2 => 
                           n3577, ZN => n13513);
   U6132 : INV_X1 port map( A => n13641, ZN => n12028);
   U6133 : AOI22_X1 port map( A1 => n2412, A2 => n3525, B1 => n3989, B2 => 
                           n3552, ZN => n13641);
   U6134 : INV_X1 port map( A => n13514, ZN => n11984);
   U6135 : AOI22_X1 port map( A1 => n2418, A2 => n3529, B1 => n3995, B2 => 
                           n3577, ZN => n13514);
   U6136 : INV_X1 port map( A => n13642, ZN => n11988);
   U6137 : AOI22_X1 port map( A1 => n2418, A2 => n3524, B1 => n3995, B2 => 
                           n3552, ZN => n13642);
   U6138 : INV_X1 port map( A => n13515, ZN => n11944);
   U6139 : AOI22_X1 port map( A1 => n2424, A2 => n3528, B1 => n4001, B2 => 
                           n3577, ZN => n13515);
   U6140 : INV_X1 port map( A => n13643, ZN => n11948);
   U6141 : AOI22_X1 port map( A1 => n2424, A2 => n3525, B1 => n4001, B2 => 
                           n3553, ZN => n13643);
   U6142 : INV_X1 port map( A => n13516, ZN => n11904);
   U6143 : AOI22_X1 port map( A1 => n2430, A2 => n3528, B1 => n4007, B2 => 
                           n3577, ZN => n13516);
   U6144 : INV_X1 port map( A => n13644, ZN => n11908);
   U6145 : AOI22_X1 port map( A1 => n2430, A2 => n3525, B1 => n4007, B2 => 
                           n3553, ZN => n13644);
   U6146 : INV_X1 port map( A => n13517, ZN => n11864);
   U6147 : AOI22_X1 port map( A1 => n2436, A2 => n3529, B1 => n4013, B2 => 
                           n3578, ZN => n13517);
   U6148 : INV_X1 port map( A => n13518, ZN => n11824);
   U6149 : AOI22_X1 port map( A1 => n2442, A2 => n3527, B1 => n4019, B2 => 
                           n3578, ZN => n13518);
   U6150 : INV_X1 port map( A => n13646, ZN => n11828);
   U6151 : AOI22_X1 port map( A1 => n2442, A2 => n3525, B1 => n4019, B2 => 
                           n3553, ZN => n13646);
   U6152 : INV_X1 port map( A => n13519, ZN => n11784);
   U6153 : AOI22_X1 port map( A1 => n2448, A2 => n3520, B1 => n4025, B2 => 
                           n3578, ZN => n13519);
   U6154 : INV_X1 port map( A => n13647, ZN => n11788);
   U6155 : AOI22_X1 port map( A1 => n2448, A2 => n3525, B1 => n4025, B2 => 
                           n3554, ZN => n13647);
   U6156 : INV_X1 port map( A => n13520, ZN => n11744);
   U6157 : AOI22_X1 port map( A1 => n2454, A2 => n3519, B1 => n4031, B2 => 
                           n3578, ZN => n13520);
   U6158 : INV_X1 port map( A => n13648, ZN => n11748);
   U6159 : AOI22_X1 port map( A1 => n2454, A2 => n3521, B1 => n4031, B2 => 
                           n3554, ZN => n13648);
   U6160 : INV_X1 port map( A => n13521, ZN => n11704);
   U6161 : AOI22_X1 port map( A1 => n2460, A2 => n3523, B1 => n4037, B2 => 
                           n3579, ZN => n13521);
   U6162 : INV_X1 port map( A => n13649, ZN => n11708);
   U6163 : AOI22_X1 port map( A1 => n2460, A2 => n3525, B1 => n4037, B2 => 
                           n3554, ZN => n13649);
   U6164 : INV_X1 port map( A => n13522, ZN => n11664);
   U6165 : AOI22_X1 port map( A1 => n2466, A2 => n3526, B1 => n4043, B2 => 
                           n3579, ZN => n13522);
   U6166 : INV_X1 port map( A => n13650, ZN => n11668);
   U6167 : AOI22_X1 port map( A1 => n2466, A2 => n3525, B1 => n4043, B2 => 
                           n3554, ZN => n13650);
   U6168 : INV_X1 port map( A => n13501, ZN => n12504);
   U6169 : AOI22_X1 port map( A1 => n2340, A2 => n3524, B1 => n4091, B2 => 
                           n3574, ZN => n13501);
   U6170 : INV_X1 port map( A => n13629, ZN => n12508);
   U6171 : AOI22_X1 port map( A1 => n2340, A2 => n3524, B1 => n4091, B2 => 
                           n3547, ZN => n13629);
   U6172 : INV_X1 port map( A => n13512, ZN => n12064);
   U6173 : AOI22_X1 port map( A1 => n2406, A2 => n3527, B1 => n4097, B2 => 
                           n3576, ZN => n13512);
   U6174 : INV_X1 port map( A => n13640, ZN => n12068);
   U6175 : AOI22_X1 port map( A1 => n2406, A2 => n3525, B1 => n4097, B2 => 
                           n3552, ZN => n13640);
   U6176 : INV_X1 port map( A => n13523, ZN => n11624);
   U6177 : AOI22_X1 port map( A1 => n2472, A2 => n3522, B1 => n4103, B2 => 
                           n3579, ZN => n13523);
   U6178 : INV_X1 port map( A => n13651, ZN => n11628);
   U6179 : AOI22_X1 port map( A1 => n2472, A2 => n3524, B1 => n4103, B2 => 
                           n3555, ZN => n13651);
   U6180 : INV_X1 port map( A => n13755, ZN => n12592);
   U6181 : AOI22_X1 port map( A1 => n2329, A2 => n3634, B1 => n3918, B2 => 
                           n3685, ZN => n13755);
   U6182 : INV_X1 port map( A => n13883, ZN => n12596);
   U6183 : AOI22_X1 port map( A1 => n2329, A2 => n3638, B1 => n3918, B2 => 
                           n3659, ZN => n13883);
   U6184 : INV_X1 port map( A => n13756, ZN => n12552);
   U6185 : AOI22_X1 port map( A1 => n2335, A2 => n3633, B1 => n3924, B2 => 
                           n3685, ZN => n13756);
   U6186 : INV_X1 port map( A => n13884, ZN => n12556);
   U6187 : AOI22_X1 port map( A1 => n2335, A2 => n3638, B1 => n3924, B2 => 
                           n3661, ZN => n13884);
   U6188 : INV_X1 port map( A => n13758, ZN => n12472);
   U6189 : AOI22_X1 port map( A1 => n2347, A2 => n3636, B1 => n3930, B2 => 
                           n3686, ZN => n13758);
   U6190 : INV_X1 port map( A => n13886, ZN => n12476);
   U6191 : AOI22_X1 port map( A1 => n2347, A2 => n3637, B1 => n3930, B2 => 
                           n3660, ZN => n13886);
   U6192 : INV_X1 port map( A => n13887, ZN => n12436);
   U6193 : AOI22_X1 port map( A1 => n2353, A2 => n3636, B1 => n3936, B2 => 
                           n3662, ZN => n13887);
   U6194 : INV_X1 port map( A => n13760, ZN => n12392);
   U6195 : AOI22_X1 port map( A1 => n2359, A2 => n3637, B1 => n3942, B2 => 
                           n3686, ZN => n13760);
   U6196 : INV_X1 port map( A => n13888, ZN => n12396);
   U6197 : AOI22_X1 port map( A1 => n2359, A2 => n3636, B1 => n3942, B2 => 
                           n3661, ZN => n13888);
   U6198 : INV_X1 port map( A => n13761, ZN => n12352);
   U6199 : AOI22_X1 port map( A1 => n2365, A2 => n3632, B1 => n3948, B2 => 
                           n3687, ZN => n13761);
   U6200 : INV_X1 port map( A => n13889, ZN => n12356);
   U6201 : AOI22_X1 port map( A1 => n2365, A2 => n3636, B1 => n3948, B2 => 
                           n3661, ZN => n13889);
   U6202 : INV_X1 port map( A => n13762, ZN => n12312);
   U6203 : AOI22_X1 port map( A1 => n2371, A2 => n3638, B1 => n3954, B2 => 
                           n3687, ZN => n13762);
   U6204 : INV_X1 port map( A => n13890, ZN => n12316);
   U6205 : AOI22_X1 port map( A1 => n2371, A2 => n3636, B1 => n3954, B2 => 
                           n3663, ZN => n13890);
   U6206 : INV_X1 port map( A => n13763, ZN => n12272);
   U6207 : AOI22_X1 port map( A1 => n2377, A2 => n3635, B1 => n3960, B2 => 
                           n3687, ZN => n13763);
   U6208 : INV_X1 port map( A => n13891, ZN => n12276);
   U6209 : AOI22_X1 port map( A1 => n2377, A2 => n3636, B1 => n3960, B2 => 
                           n3662, ZN => n13891);
   U6210 : INV_X1 port map( A => n13764, ZN => n12232);
   U6211 : AOI22_X1 port map( A1 => n2383, A2 => n3637, B1 => n3966, B2 => 
                           n3687, ZN => n13764);
   U6212 : INV_X1 port map( A => n13892, ZN => n12236);
   U6213 : AOI22_X1 port map( A1 => n2383, A2 => n3637, B1 => n3966, B2 => 
                           n3662, ZN => n13892);
   U6214 : INV_X1 port map( A => n13765, ZN => n12192);
   U6215 : AOI22_X1 port map( A1 => n2389, A2 => n3634, B1 => n3972, B2 => 
                           n3688, ZN => n13765);
   U6216 : INV_X1 port map( A => n13893, ZN => n12196);
   U6217 : AOI22_X1 port map( A1 => n2389, A2 => n3637, B1 => n3972, B2 => 
                           n3663, ZN => n13893);
   U6218 : INV_X1 port map( A => n13766, ZN => n12152);
   U6219 : AOI22_X1 port map( A1 => n2395, A2 => n3634, B1 => n3978, B2 => 
                           n3688, ZN => n13766);
   U6220 : INV_X1 port map( A => n13894, ZN => n12156);
   U6221 : AOI22_X1 port map( A1 => n2395, A2 => n3636, B1 => n3978, B2 => 
                           n3663, ZN => n13894);
   U6222 : INV_X1 port map( A => n13767, ZN => n12112);
   U6223 : AOI22_X1 port map( A1 => n2401, A2 => n3634, B1 => n3984, B2 => 
                           n3688, ZN => n13767);
   U6224 : INV_X1 port map( A => n13895, ZN => n12116);
   U6225 : AOI22_X1 port map( A1 => n2401, A2 => n3637, B1 => n3984, B2 => 
                           n3664, ZN => n13895);
   U6226 : INV_X1 port map( A => n13769, ZN => n12032);
   U6227 : AOI22_X1 port map( A1 => n2413, A2 => n3634, B1 => n3990, B2 => 
                           n3689, ZN => n13769);
   U6228 : INV_X1 port map( A => n13897, ZN => n12036);
   U6229 : AOI22_X1 port map( A1 => n2413, A2 => n3637, B1 => n3990, B2 => 
                           n3664, ZN => n13897);
   U6230 : INV_X1 port map( A => n13770, ZN => n11992);
   U6231 : AOI22_X1 port map( A1 => n2419, A2 => n3634, B1 => n3996, B2 => 
                           n3689, ZN => n13770);
   U6232 : INV_X1 port map( A => n13898, ZN => n11996);
   U6233 : AOI22_X1 port map( A1 => n2419, A2 => n3636, B1 => n3996, B2 => 
                           n3664, ZN => n13898);
   U6234 : INV_X1 port map( A => n13771, ZN => n11952);
   U6235 : AOI22_X1 port map( A1 => n2425, A2 => n3634, B1 => n4002, B2 => 
                           n3689, ZN => n13771);
   U6236 : INV_X1 port map( A => n13899, ZN => n11956);
   U6237 : AOI22_X1 port map( A1 => n2425, A2 => n3637, B1 => n4002, B2 => 
                           n3665, ZN => n13899);
   U6238 : INV_X1 port map( A => n13772, ZN => n11912);
   U6239 : AOI22_X1 port map( A1 => n2431, A2 => n3634, B1 => n4008, B2 => 
                           n3689, ZN => n13772);
   U6240 : INV_X1 port map( A => n13900, ZN => n11916);
   U6241 : AOI22_X1 port map( A1 => n2431, A2 => n3637, B1 => n4008, B2 => 
                           n3665, ZN => n13900);
   U6242 : INV_X1 port map( A => n13773, ZN => n11872);
   U6243 : AOI22_X1 port map( A1 => n2437, A2 => n3634, B1 => n4014, B2 => 
                           n3690, ZN => n13773);
   U6244 : INV_X1 port map( A => n13774, ZN => n11832);
   U6245 : AOI22_X1 port map( A1 => n2443, A2 => n3634, B1 => n4020, B2 => 
                           n3690, ZN => n13774);
   U6246 : INV_X1 port map( A => n13902, ZN => n11836);
   U6247 : AOI22_X1 port map( A1 => n2443, A2 => n3637, B1 => n4020, B2 => 
                           n3665, ZN => n13902);
   U6248 : INV_X1 port map( A => n13775, ZN => n11792);
   U6249 : AOI22_X1 port map( A1 => n2449, A2 => n3634, B1 => n4026, B2 => 
                           n3690, ZN => n13775);
   U6250 : INV_X1 port map( A => n13903, ZN => n11796);
   U6251 : AOI22_X1 port map( A1 => n2449, A2 => n3637, B1 => n4026, B2 => 
                           n3666, ZN => n13903);
   U6252 : INV_X1 port map( A => n13776, ZN => n11752);
   U6253 : AOI22_X1 port map( A1 => n2455, A2 => n3634, B1 => n4032, B2 => 
                           n3690, ZN => n13776);
   U6254 : INV_X1 port map( A => n13904, ZN => n11756);
   U6255 : AOI22_X1 port map( A1 => n2455, A2 => n3632, B1 => n4032, B2 => 
                           n3666, ZN => n13904);
   U6256 : INV_X1 port map( A => n13777, ZN => n11712);
   U6257 : AOI22_X1 port map( A1 => n2461, A2 => n3635, B1 => n4038, B2 => 
                           n3691, ZN => n13777);
   U6258 : INV_X1 port map( A => n13905, ZN => n11716);
   U6259 : AOI22_X1 port map( A1 => n2461, A2 => n3637, B1 => n4038, B2 => 
                           n3666, ZN => n13905);
   U6260 : INV_X1 port map( A => n13778, ZN => n11672);
   U6261 : AOI22_X1 port map( A1 => n2467, A2 => n3638, B1 => n4044, B2 => 
                           n3691, ZN => n13778);
   U6262 : INV_X1 port map( A => n13906, ZN => n11676);
   U6263 : AOI22_X1 port map( A1 => n2467, A2 => n3637, B1 => n4044, B2 => 
                           n3666, ZN => n13906);
   U6264 : INV_X1 port map( A => n13757, ZN => n12512);
   U6265 : AOI22_X1 port map( A1 => n2341, A2 => n3636, B1 => n4092, B2 => 
                           n3686, ZN => n13757);
   U6266 : INV_X1 port map( A => n13885, ZN => n12516);
   U6267 : AOI22_X1 port map( A1 => n2341, A2 => n3636, B1 => n4092, B2 => 
                           n3659, ZN => n13885);
   U6268 : INV_X1 port map( A => n13768, ZN => n12072);
   U6269 : AOI22_X1 port map( A1 => n2407, A2 => n3634, B1 => n4098, B2 => 
                           n3688, ZN => n13768);
   U6270 : INV_X1 port map( A => n13896, ZN => n12076);
   U6271 : AOI22_X1 port map( A1 => n2407, A2 => n3637, B1 => n4098, B2 => 
                           n3664, ZN => n13896);
   U6272 : INV_X1 port map( A => n13779, ZN => n11632);
   U6273 : AOI22_X1 port map( A1 => n2473, A2 => n3633, B1 => n4104, B2 => 
                           n3691, ZN => n13779);
   U6274 : INV_X1 port map( A => n13907, ZN => n11636);
   U6275 : AOI22_X1 port map( A1 => n2473, A2 => n3636, B1 => n4104, B2 => 
                           n3667, ZN => n13907);
   U6276 : INV_X1 port map( A => n14011, ZN => n12600);
   U6277 : AOI22_X1 port map( A1 => n2329, A2 => n3745, B1 => n3918, B2 => 
                           n3797, ZN => n14011);
   U6278 : INV_X1 port map( A => n14139, ZN => n12604);
   U6279 : AOI22_X1 port map( A1 => n2330, A2 => n3747, B1 => n3919, B2 => 
                           n3771, ZN => n14139);
   U6280 : INV_X1 port map( A => n14012, ZN => n12560);
   U6281 : AOI22_X1 port map( A1 => n2335, A2 => n3743, B1 => n3924, B2 => 
                           n3797, ZN => n14012);
   U6282 : INV_X1 port map( A => n14140, ZN => n12564);
   U6283 : AOI22_X1 port map( A1 => n2336, A2 => n3747, B1 => n3925, B2 => 
                           n3773, ZN => n14140);
   U6284 : INV_X1 port map( A => n14014, ZN => n12480);
   U6285 : AOI22_X1 port map( A1 => n2347, A2 => n3750, B1 => n3930, B2 => 
                           n3798, ZN => n14014);
   U6286 : INV_X1 port map( A => n14142, ZN => n12484);
   U6287 : AOI22_X1 port map( A1 => n2348, A2 => n3747, B1 => n3931, B2 => 
                           n3772, ZN => n14142);
   U6288 : INV_X1 port map( A => n14143, ZN => n12444);
   U6289 : AOI22_X1 port map( A1 => n2354, A2 => n3748, B1 => n3937, B2 => 
                           n3774, ZN => n14143);
   U6290 : INV_X1 port map( A => n14016, ZN => n12400);
   U6291 : AOI22_X1 port map( A1 => n2359, A2 => n3747, B1 => n3942, B2 => 
                           n3798, ZN => n14016);
   U6292 : INV_X1 port map( A => n14144, ZN => n12404);
   U6293 : AOI22_X1 port map( A1 => n2360, A2 => n3748, B1 => n3943, B2 => 
                           n3773, ZN => n14144);
   U6294 : INV_X1 port map( A => n14017, ZN => n12360);
   U6295 : AOI22_X1 port map( A1 => n2365, A2 => n3746, B1 => n3948, B2 => 
                           n3799, ZN => n14017);
   U6296 : INV_X1 port map( A => n14145, ZN => n12364);
   U6297 : AOI22_X1 port map( A1 => n2366, A2 => n3748, B1 => n3949, B2 => 
                           n3773, ZN => n14145);
   U6298 : INV_X1 port map( A => n14018, ZN => n12320);
   U6299 : AOI22_X1 port map( A1 => n2371, A2 => n3744, B1 => n3954, B2 => 
                           n3799, ZN => n14018);
   U6300 : INV_X1 port map( A => n14146, ZN => n12324);
   U6301 : AOI22_X1 port map( A1 => n2372, A2 => n3748, B1 => n3955, B2 => 
                           n3775, ZN => n14146);
   U6302 : INV_X1 port map( A => n14019, ZN => n12280);
   U6303 : AOI22_X1 port map( A1 => n2377, A2 => n3745, B1 => n3960, B2 => 
                           n3799, ZN => n14019);
   U6304 : INV_X1 port map( A => n14147, ZN => n12284);
   U6305 : AOI22_X1 port map( A1 => n2378, A2 => n3748, B1 => n3961, B2 => 
                           n3774, ZN => n14147);
   U6306 : INV_X1 port map( A => n14020, ZN => n12240);
   U6307 : AOI22_X1 port map( A1 => n2383, A2 => n3743, B1 => n3966, B2 => 
                           n3799, ZN => n14020);
   U6308 : INV_X1 port map( A => n14148, ZN => n12244);
   U6309 : AOI22_X1 port map( A1 => n2384, A2 => n3748, B1 => n3967, B2 => 
                           n3774, ZN => n14148);
   U6310 : INV_X1 port map( A => n14021, ZN => n12200);
   U6311 : AOI22_X1 port map( A1 => n2389, A2 => n3744, B1 => n3972, B2 => 
                           n3800, ZN => n14021);
   U6312 : INV_X1 port map( A => n14149, ZN => n12204);
   U6313 : AOI22_X1 port map( A1 => n2390, A2 => n3747, B1 => n3973, B2 => 
                           n3775, ZN => n14149);
   U6314 : INV_X1 port map( A => n14022, ZN => n12160);
   U6315 : AOI22_X1 port map( A1 => n2395, A2 => n3744, B1 => n3978, B2 => 
                           n3800, ZN => n14022);
   U6316 : INV_X1 port map( A => n14150, ZN => n12164);
   U6317 : AOI22_X1 port map( A1 => n2396, A2 => n3748, B1 => n3979, B2 => 
                           n3775, ZN => n14150);
   U6318 : INV_X1 port map( A => n14023, ZN => n12120);
   U6319 : AOI22_X1 port map( A1 => n2401, A2 => n3744, B1 => n3984, B2 => 
                           n3800, ZN => n14023);
   U6320 : INV_X1 port map( A => n14151, ZN => n12124);
   U6321 : AOI22_X1 port map( A1 => n2402, A2 => n3746, B1 => n3985, B2 => 
                           n3776, ZN => n14151);
   U6322 : INV_X1 port map( A => n14025, ZN => n12040);
   U6323 : AOI22_X1 port map( A1 => n2413, A2 => n3744, B1 => n3990, B2 => 
                           n3801, ZN => n14025);
   U6324 : INV_X1 port map( A => n14153, ZN => n12044);
   U6325 : AOI22_X1 port map( A1 => n2414, A2 => n3744, B1 => n3991, B2 => 
                           n3776, ZN => n14153);
   U6326 : INV_X1 port map( A => n14026, ZN => n12000);
   U6327 : AOI22_X1 port map( A1 => n2419, A2 => n3744, B1 => n3996, B2 => 
                           n3801, ZN => n14026);
   U6328 : INV_X1 port map( A => n14154, ZN => n12004);
   U6329 : AOI22_X1 port map( A1 => n2420, A2 => n3748, B1 => n3997, B2 => 
                           n3776, ZN => n14154);
   U6330 : INV_X1 port map( A => n14027, ZN => n11960);
   U6331 : AOI22_X1 port map( A1 => n2425, A2 => n3744, B1 => n4002, B2 => 
                           n3801, ZN => n14027);
   U6332 : INV_X1 port map( A => n14155, ZN => n11964);
   U6333 : AOI22_X1 port map( A1 => n2426, A2 => n3745, B1 => n4003, B2 => 
                           n3777, ZN => n14155);
   U6334 : INV_X1 port map( A => n14028, ZN => n11920);
   U6335 : AOI22_X1 port map( A1 => n2431, A2 => n3744, B1 => n4008, B2 => 
                           n3801, ZN => n14028);
   U6336 : INV_X1 port map( A => n14156, ZN => n11924);
   U6337 : AOI22_X1 port map( A1 => n2432, A2 => n3749, B1 => n4009, B2 => 
                           n3777, ZN => n14156);
   U6338 : INV_X1 port map( A => n14029, ZN => n11880);
   U6339 : AOI22_X1 port map( A1 => n2437, A2 => n3744, B1 => n4014, B2 => 
                           n3802, ZN => n14029);
   U6340 : INV_X1 port map( A => n14030, ZN => n11840);
   U6341 : AOI22_X1 port map( A1 => n2443, A2 => n3744, B1 => n4020, B2 => 
                           n3802, ZN => n14030);
   U6342 : INV_X1 port map( A => n14158, ZN => n11844);
   U6343 : AOI22_X1 port map( A1 => n2444, A2 => n3750, B1 => n4021, B2 => 
                           n3777, ZN => n14158);
   U6344 : INV_X1 port map( A => n14031, ZN => n11800);
   U6345 : AOI22_X1 port map( A1 => n2449, A2 => n3744, B1 => n4026, B2 => 
                           n3802, ZN => n14031);
   U6346 : INV_X1 port map( A => n14159, ZN => n11804);
   U6347 : AOI22_X1 port map( A1 => n2450, A2 => n3748, B1 => n4027, B2 => 
                           n3778, ZN => n14159);
   U6348 : INV_X1 port map( A => n14032, ZN => n11760);
   U6349 : AOI22_X1 port map( A1 => n2455, A2 => n3744, B1 => n4032, B2 => 
                           n3802, ZN => n14032);
   U6350 : INV_X1 port map( A => n14160, ZN => n11764);
   U6351 : AOI22_X1 port map( A1 => n2456, A2 => n3750, B1 => n4033, B2 => 
                           n3778, ZN => n14160);
   U6352 : INV_X1 port map( A => n14033, ZN => n11720);
   U6353 : AOI22_X1 port map( A1 => n2461, A2 => n3743, B1 => n4038, B2 => 
                           n3803, ZN => n14033);
   U6354 : INV_X1 port map( A => n14161, ZN => n11724);
   U6355 : AOI22_X1 port map( A1 => n2462, A2 => n3753, B1 => n4039, B2 => 
                           n3778, ZN => n14161);
   U6356 : INV_X1 port map( A => n14034, ZN => n11680);
   U6357 : AOI22_X1 port map( A1 => n2467, A2 => n3743, B1 => n4044, B2 => 
                           n3803, ZN => n14034);
   U6358 : INV_X1 port map( A => n14162, ZN => n11684);
   U6359 : AOI22_X1 port map( A1 => n2468, A2 => n3743, B1 => n4045, B2 => 
                           n3778, ZN => n14162);
   U6360 : INV_X1 port map( A => n14013, ZN => n12520);
   U6361 : AOI22_X1 port map( A1 => n2341, A2 => n3753, B1 => n4092, B2 => 
                           n3798, ZN => n14013);
   U6362 : INV_X1 port map( A => n14141, ZN => n12524);
   U6363 : AOI22_X1 port map( A1 => n2342, A2 => n3747, B1 => n4093, B2 => 
                           n3771, ZN => n14141);
   U6364 : INV_X1 port map( A => n14024, ZN => n12080);
   U6365 : AOI22_X1 port map( A1 => n2407, A2 => n3744, B1 => n4098, B2 => 
                           n3800, ZN => n14024);
   U6366 : INV_X1 port map( A => n14152, ZN => n12084);
   U6367 : AOI22_X1 port map( A1 => n2408, A2 => n3749, B1 => n4099, B2 => 
                           n3776, ZN => n14152);
   U6368 : INV_X1 port map( A => n14035, ZN => n11640);
   U6369 : AOI22_X1 port map( A1 => n2473, A2 => n3743, B1 => n4104, B2 => 
                           n3803, ZN => n14035);
   U6370 : INV_X1 port map( A => n14163, ZN => n11644);
   U6371 : AOI22_X1 port map( A1 => n2474, A2 => n3752, B1 => n4105, B2 => 
                           n3779, ZN => n14163);
   U6372 : INV_X1 port map( A => n13147, ZN => n12573);
   U6373 : AOI22_X1 port map( A1 => n2327, A2 => n3305, B1 => n3916, B2 => 
                           n3323, ZN => n13147);
   U6374 : INV_X1 port map( A => n12998, ZN => n12128);
   U6375 : AOI22_X1 port map( A1 => n2393, A2 => n3298, B1 => n3976, B2 => 
                           n3346, ZN => n12998);
   U6376 : INV_X1 port map( A => n12999, ZN => n12088);
   U6377 : AOI22_X1 port map( A1 => n2399, A2 => n3298, B1 => n3982, B2 => 
                           n3346, ZN => n12999);
   U6378 : INV_X1 port map( A => n13001, ZN => n12008);
   U6379 : AOI22_X1 port map( A1 => n2411, A2 => n3298, B1 => n3988, B2 => 
                           n3346, ZN => n13001);
   U6380 : INV_X1 port map( A => n13002, ZN => n11968);
   U6381 : AOI22_X1 port map( A1 => n2417, A2 => n3298, B1 => n3994, B2 => 
                           n3347, ZN => n13002);
   U6382 : INV_X1 port map( A => n13003, ZN => n11928);
   U6383 : AOI22_X1 port map( A1 => n2423, A2 => n3298, B1 => n4000, B2 => 
                           n3347, ZN => n13003);
   U6384 : INV_X1 port map( A => n13004, ZN => n11888);
   U6385 : AOI22_X1 port map( A1 => n2429, A2 => n3298, B1 => n4006, B2 => 
                           n3347, ZN => n13004);
   U6386 : INV_X1 port map( A => n13005, ZN => n11848);
   U6387 : AOI22_X1 port map( A1 => n2435, A2 => n3298, B1 => n4012, B2 => 
                           n3347, ZN => n13005);
   U6388 : INV_X1 port map( A => n13006, ZN => n11808);
   U6389 : AOI22_X1 port map( A1 => n2441, A2 => n3298, B1 => n4018, B2 => 
                           n3348, ZN => n13006);
   U6390 : INV_X1 port map( A => n13007, ZN => n11768);
   U6391 : AOI22_X1 port map( A1 => n2447, A2 => n3298, B1 => n4024, B2 => 
                           n3348, ZN => n13007);
   U6392 : INV_X1 port map( A => n13008, ZN => n11728);
   U6393 : AOI22_X1 port map( A1 => n2453, A2 => n3298, B1 => n4030, B2 => 
                           n3348, ZN => n13008);
   U6394 : INV_X1 port map( A => n13009, ZN => n11688);
   U6395 : AOI22_X1 port map( A1 => n2459, A2 => n3298, B1 => n4036, B2 => 
                           n3348, ZN => n13009);
   U6396 : INV_X1 port map( A => n13010, ZN => n11648);
   U6397 : AOI22_X1 port map( A1 => n2465, A2 => n3300, B1 => n4042, B2 => 
                           n3349, ZN => n13010);
   U6398 : INV_X1 port map( A => n13000, ZN => n12048);
   U6399 : AOI22_X1 port map( A1 => n2405, A2 => n3298, B1 => n4096, B2 => 
                           n3346, ZN => n13000);
   U6400 : INV_X1 port map( A => n13011, ZN => n11608);
   U6401 : AOI22_X1 port map( A1 => n2471, A2 => n3302, B1 => n4102, B2 => 
                           n3349, ZN => n13011);
   U6402 : INV_X1 port map( A => n13222, ZN => n12135);
   U6403 : AOI22_X1 port map( A1 => n2393, A2 => n3410, B1 => n3976, B2 => 
                           n3458, ZN => n13222);
   U6404 : INV_X1 port map( A => n13223, ZN => n12095);
   U6405 : AOI22_X1 port map( A1 => n2399, A2 => n3412, B1 => n3982, B2 => 
                           n3458, ZN => n13223);
   U6406 : INV_X1 port map( A => n13225, ZN => n12015);
   U6407 : AOI22_X1 port map( A1 => n2411, A2 => n3416, B1 => n3988, B2 => 
                           n3458, ZN => n13225);
   U6408 : INV_X1 port map( A => n13226, ZN => n11975);
   U6409 : AOI22_X1 port map( A1 => n2417, A2 => n3411, B1 => n3994, B2 => 
                           n3459, ZN => n13226);
   U6410 : INV_X1 port map( A => n13227, ZN => n11935);
   U6411 : AOI22_X1 port map( A1 => n2423, A2 => n3409, B1 => n4000, B2 => 
                           n3459, ZN => n13227);
   U6412 : INV_X1 port map( A => n13228, ZN => n11895);
   U6413 : AOI22_X1 port map( A1 => n2429, A2 => n3409, B1 => n4006, B2 => 
                           n3459, ZN => n13228);
   U6414 : INV_X1 port map( A => n13229, ZN => n11855);
   U6415 : AOI22_X1 port map( A1 => n2435, A2 => n3414, B1 => n4012, B2 => 
                           n3459, ZN => n13229);
   U6416 : INV_X1 port map( A => n13230, ZN => n11815);
   U6417 : AOI22_X1 port map( A1 => n2441, A2 => n3409, B1 => n4018, B2 => 
                           n3460, ZN => n13230);
   U6418 : INV_X1 port map( A => n13231, ZN => n11775);
   U6419 : AOI22_X1 port map( A1 => n2447, A2 => n3413, B1 => n4024, B2 => 
                           n3460, ZN => n13231);
   U6420 : INV_X1 port map( A => n13232, ZN => n11735);
   U6421 : AOI22_X1 port map( A1 => n2453, A2 => n3412, B1 => n4030, B2 => 
                           n3460, ZN => n13232);
   U6422 : INV_X1 port map( A => n13233, ZN => n11695);
   U6423 : AOI22_X1 port map( A1 => n2459, A2 => n3415, B1 => n4036, B2 => 
                           n3460, ZN => n13233);
   U6424 : INV_X1 port map( A => n13234, ZN => n11655);
   U6425 : AOI22_X1 port map( A1 => n2465, A2 => n3411, B1 => n4042, B2 => 
                           n3461, ZN => n13234);
   U6426 : INV_X1 port map( A => n13224, ZN => n12055);
   U6427 : AOI22_X1 port map( A1 => n2405, A2 => n3410, B1 => n4096, B2 => 
                           n3458, ZN => n13224);
   U6428 : INV_X1 port map( A => n13235, ZN => n11615);
   U6429 : AOI22_X1 port map( A1 => n2471, A2 => n3413, B1 => n4102, B2 => 
                           n3461, ZN => n13235);
   U6430 : INV_X1 port map( A => n13478, ZN => n12143);
   U6431 : AOI22_X1 port map( A1 => n2394, A2 => n3522, B1 => n3977, B2 => 
                           n3570, ZN => n13478);
   U6432 : INV_X1 port map( A => n13479, ZN => n12103);
   U6433 : AOI22_X1 port map( A1 => n2400, A2 => n3524, B1 => n3983, B2 => 
                           n3570, ZN => n13479);
   U6434 : INV_X1 port map( A => n13481, ZN => n12023);
   U6435 : AOI22_X1 port map( A1 => n2412, A2 => n3528, B1 => n3989, B2 => 
                           n3570, ZN => n13481);
   U6436 : INV_X1 port map( A => n13482, ZN => n11983);
   U6437 : AOI22_X1 port map( A1 => n2418, A2 => n3523, B1 => n3995, B2 => 
                           n3571, ZN => n13482);
   U6438 : INV_X1 port map( A => n13483, ZN => n11943);
   U6439 : AOI22_X1 port map( A1 => n2424, A2 => n3521, B1 => n4001, B2 => 
                           n3571, ZN => n13483);
   U6440 : INV_X1 port map( A => n13484, ZN => n11903);
   U6441 : AOI22_X1 port map( A1 => n2430, A2 => n3521, B1 => n4007, B2 => 
                           n3571, ZN => n13484);
   U6442 : INV_X1 port map( A => n13485, ZN => n11863);
   U6443 : AOI22_X1 port map( A1 => n2436, A2 => n3526, B1 => n4013, B2 => 
                           n3571, ZN => n13485);
   U6444 : INV_X1 port map( A => n13486, ZN => n11823);
   U6445 : AOI22_X1 port map( A1 => n2442, A2 => n3521, B1 => n4019, B2 => 
                           n3572, ZN => n13486);
   U6446 : INV_X1 port map( A => n13487, ZN => n11783);
   U6447 : AOI22_X1 port map( A1 => n2448, A2 => n3525, B1 => n4025, B2 => 
                           n3572, ZN => n13487);
   U6448 : INV_X1 port map( A => n13488, ZN => n11743);
   U6449 : AOI22_X1 port map( A1 => n2454, A2 => n3524, B1 => n4031, B2 => 
                           n3572, ZN => n13488);
   U6450 : INV_X1 port map( A => n13489, ZN => n11703);
   U6451 : AOI22_X1 port map( A1 => n2460, A2 => n3527, B1 => n4037, B2 => 
                           n3572, ZN => n13489);
   U6452 : INV_X1 port map( A => n13490, ZN => n11663);
   U6453 : AOI22_X1 port map( A1 => n2466, A2 => n3523, B1 => n4043, B2 => 
                           n3573, ZN => n13490);
   U6454 : INV_X1 port map( A => n13480, ZN => n12063);
   U6455 : AOI22_X1 port map( A1 => n2406, A2 => n3522, B1 => n4097, B2 => 
                           n3570, ZN => n13480);
   U6456 : INV_X1 port map( A => n13491, ZN => n11623);
   U6457 : AOI22_X1 port map( A1 => n2472, A2 => n3525, B1 => n4103, B2 => 
                           n3573, ZN => n13491);
   U6458 : INV_X1 port map( A => n13734, ZN => n12151);
   U6459 : AOI22_X1 port map( A1 => n2394, A2 => n3633, B1 => n3977, B2 => 
                           n3682, ZN => n13734);
   U6460 : INV_X1 port map( A => n13735, ZN => n12111);
   U6461 : AOI22_X1 port map( A1 => n2400, A2 => n3636, B1 => n3983, B2 => 
                           n3682, ZN => n13735);
   U6462 : INV_X1 port map( A => n13737, ZN => n12031);
   U6463 : AOI22_X1 port map( A1 => n2412, A2 => n3634, B1 => n3989, B2 => 
                           n3682, ZN => n13737);
   U6464 : INV_X1 port map( A => n13738, ZN => n11991);
   U6465 : AOI22_X1 port map( A1 => n2418, A2 => n3635, B1 => n3995, B2 => 
                           n3683, ZN => n13738);
   U6466 : INV_X1 port map( A => n13739, ZN => n11951);
   U6467 : AOI22_X1 port map( A1 => n2424, A2 => n3632, B1 => n4001, B2 => 
                           n3683, ZN => n13739);
   U6468 : INV_X1 port map( A => n13740, ZN => n11911);
   U6469 : AOI22_X1 port map( A1 => n2430, A2 => n3632, B1 => n4007, B2 => 
                           n3683, ZN => n13740);
   U6470 : INV_X1 port map( A => n13741, ZN => n11871);
   U6471 : AOI22_X1 port map( A1 => n2436, A2 => n3638, B1 => n4013, B2 => 
                           n3683, ZN => n13741);
   U6472 : INV_X1 port map( A => n13742, ZN => n11831);
   U6473 : AOI22_X1 port map( A1 => n2442, A2 => n3632, B1 => n4019, B2 => 
                           n3684, ZN => n13742);
   U6474 : INV_X1 port map( A => n13743, ZN => n11791);
   U6475 : AOI22_X1 port map( A1 => n2448, A2 => n3637, B1 => n4025, B2 => 
                           n3684, ZN => n13743);
   U6476 : INV_X1 port map( A => n13744, ZN => n11751);
   U6477 : AOI22_X1 port map( A1 => n2454, A2 => n3636, B1 => n4031, B2 => 
                           n3684, ZN => n13744);
   U6478 : INV_X1 port map( A => n13745, ZN => n11711);
   U6479 : AOI22_X1 port map( A1 => n2460, A2 => n3634, B1 => n4037, B2 => 
                           n3684, ZN => n13745);
   U6480 : INV_X1 port map( A => n13746, ZN => n11671);
   U6481 : AOI22_X1 port map( A1 => n2466, A2 => n3635, B1 => n4043, B2 => 
                           n3685, ZN => n13746);
   U6482 : INV_X1 port map( A => n13736, ZN => n12071);
   U6483 : AOI22_X1 port map( A1 => n2406, A2 => n3633, B1 => n4097, B2 => 
                           n3682, ZN => n13736);
   U6484 : INV_X1 port map( A => n13747, ZN => n11631);
   U6485 : AOI22_X1 port map( A1 => n2472, A2 => n3637, B1 => n4103, B2 => 
                           n3685, ZN => n13747);
   U6486 : INV_X1 port map( A => n13990, ZN => n12159);
   U6487 : AOI22_X1 port map( A1 => n2395, A2 => n3745, B1 => n3978, B2 => 
                           n3794, ZN => n13990);
   U6488 : INV_X1 port map( A => n13991, ZN => n12119);
   U6489 : AOI22_X1 port map( A1 => n2401, A2 => n3745, B1 => n3984, B2 => 
                           n3794, ZN => n13991);
   U6490 : INV_X1 port map( A => n13993, ZN => n12039);
   U6491 : AOI22_X1 port map( A1 => n2413, A2 => n3745, B1 => n3990, B2 => 
                           n3794, ZN => n13993);
   U6492 : INV_X1 port map( A => n13994, ZN => n11999);
   U6493 : AOI22_X1 port map( A1 => n2419, A2 => n3745, B1 => n3996, B2 => 
                           n3795, ZN => n13994);
   U6494 : INV_X1 port map( A => n13995, ZN => n11959);
   U6495 : AOI22_X1 port map( A1 => n2425, A2 => n3745, B1 => n4002, B2 => 
                           n3795, ZN => n13995);
   U6496 : INV_X1 port map( A => n13996, ZN => n11919);
   U6497 : AOI22_X1 port map( A1 => n2431, A2 => n3745, B1 => n4008, B2 => 
                           n3795, ZN => n13996);
   U6498 : INV_X1 port map( A => n13997, ZN => n11879);
   U6499 : AOI22_X1 port map( A1 => n2437, A2 => n3745, B1 => n4014, B2 => 
                           n3795, ZN => n13997);
   U6500 : INV_X1 port map( A => n13998, ZN => n11839);
   U6501 : AOI22_X1 port map( A1 => n2443, A2 => n3745, B1 => n4020, B2 => 
                           n3796, ZN => n13998);
   U6502 : INV_X1 port map( A => n13999, ZN => n11799);
   U6503 : AOI22_X1 port map( A1 => n2449, A2 => n3745, B1 => n4026, B2 => 
                           n3796, ZN => n13999);
   U6504 : INV_X1 port map( A => n14000, ZN => n11759);
   U6505 : AOI22_X1 port map( A1 => n2455, A2 => n3745, B1 => n4032, B2 => 
                           n3796, ZN => n14000);
   U6506 : INV_X1 port map( A => n14001, ZN => n11719);
   U6507 : AOI22_X1 port map( A1 => n2461, A2 => n3745, B1 => n4038, B2 => 
                           n3796, ZN => n14001);
   U6508 : INV_X1 port map( A => n14002, ZN => n11679);
   U6509 : AOI22_X1 port map( A1 => n2467, A2 => n3747, B1 => n4044, B2 => 
                           n3797, ZN => n14002);
   U6510 : INV_X1 port map( A => n13992, ZN => n12079);
   U6511 : AOI22_X1 port map( A1 => n2407, A2 => n3745, B1 => n4098, B2 => 
                           n3794, ZN => n13992);
   U6512 : INV_X1 port map( A => n14003, ZN => n11639);
   U6513 : AOI22_X1 port map( A1 => n2473, A2 => n3746, B1 => n4104, B2 => 
                           n3797, ZN => n14003);
   U6514 : INV_X1 port map( A => n12987, ZN => n12568);
   U6515 : AOI22_X1 port map( A1 => n2327, A2 => n3300, B1 => n3916, B2 => 
                           n3343, ZN => n12987);
   U6516 : INV_X1 port map( A => n13211, ZN => n12575);
   U6517 : AOI22_X1 port map( A1 => n2327, A2 => n3407, B1 => n3916, B2 => 
                           n3455, ZN => n13211);
   U6518 : INV_X1 port map( A => n13343, ZN => n12419);
   U6519 : AOI22_X1 port map( A1 => n2351, A2 => n3408, B1 => n3934, B2 => 
                           n3430, ZN => n13343);
   U6520 : INV_X1 port map( A => n13467, ZN => n12583);
   U6521 : AOI22_X1 port map( A1 => n2328, A2 => n3519, B1 => n3917, B2 => 
                           n3567, ZN => n13467);
   U6522 : INV_X1 port map( A => n13599, ZN => n12427);
   U6523 : AOI22_X1 port map( A1 => n2352, A2 => n3520, B1 => n3935, B2 => 
                           n3542, ZN => n13599);
   U6524 : INV_X1 port map( A => n13723, ZN => n12591);
   U6525 : AOI22_X1 port map( A1 => n2328, A2 => n3631, B1 => n3917, B2 => 
                           n3679, ZN => n13723);
   U6526 : INV_X1 port map( A => n13855, ZN => n12435);
   U6527 : AOI22_X1 port map( A1 => n2353, A2 => n3640, B1 => n3936, B2 => 
                           n3654, ZN => n13855);
   U6528 : INV_X1 port map( A => n13979, ZN => n12599);
   U6529 : AOI22_X1 port map( A1 => n2329, A2 => n3751, B1 => n3918, B2 => 
                           n3791, ZN => n13979);
   U6530 : INV_X1 port map( A => n14111, ZN => n12443);
   U6531 : AOI22_X1 port map( A1 => n2353, A2 => n3745, B1 => n3936, B2 => 
                           n3766, ZN => n14111);
   U6532 : INV_X1 port map( A => n13139, ZN => n11612);
   U6533 : AOI22_X1 port map( A1 => n2471, A2 => n3304, B1 => n4102, B2 => 
                           n3326, ZN => n13139);
   U6534 : NOR3_X1 port map( A1 => n12904, A2 => n12906, A3 => n12903, ZN => 
                           n12905);
   U6535 : INV_X1 port map( A => n8026, ZN => n8315);
   U6536 : INV_X1 port map( A => n3278, ZN => n3269);
   U6537 : INV_X1 port map( A => n2252, ZN => n2258);
   U6538 : NOR2_X1 port map( A1 => n14230, A2 => n4183, ZN => n14229);
   U6539 : NAND2_X1 port map( A1 => n4106, A2 => n4260, ZN => CU_I_n22);
   U6540 : INV_X1 port map( A => DataPath_LDSTR_n64, ZN => n11575);
   U6541 : NOR2_X1 port map( A1 => n2497, A2 => n4182, ZN => n14294);
   U6542 : NOR2_X1 port map( A1 => n2503, A2 => n4181, ZN => n14328);
   U6543 : BUF_X1 port map( A => n14261, Z => n2491);
   U6544 : BUF_X1 port map( A => n14261, Z => n2490);
   U6545 : BUF_X1 port map( A => n14261, Z => n2489);
   U6546 : AOI22_X1 port map( A1 => n3889, A2 => n12905, B1 => n3890, B2 => 
                           n12906, ZN => n12901);
   U6547 : BUF_X1 port map( A => n3395, Z => n3306);
   U6548 : BUF_X1 port map( A => n3291, Z => n3395);
   U6549 : BUF_X1 port map( A => n3507, Z => n3418);
   U6550 : BUF_X1 port map( A => n3403, Z => n3507);
   U6551 : BUF_X1 port map( A => n3619, Z => n3530);
   U6552 : BUF_X1 port map( A => n3515, Z => n3619);
   U6553 : BUF_X1 port map( A => n3843, Z => n3754);
   U6554 : BUF_X1 port map( A => n3739, Z => n3843);
   U6555 : BUF_X1 port map( A => n7970, Z => n2186);
   U6556 : NOR2_X1 port map( A1 => n2133, A2 => n4107, ZN => CU_I_n127);
   U6557 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_3_0_port, Z => 
                           n3629);
   U6558 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_3_0_port, Z => 
                           n3628);
   U6559 : BUF_X1 port map( A => n3290, Z => n3393);
   U6560 : BUF_X1 port map( A => n3290, Z => n3392);
   U6561 : BUF_X1 port map( A => n3290, Z => n3391);
   U6562 : BUF_X1 port map( A => n3287, Z => n3382);
   U6563 : BUF_X1 port map( A => n3289, Z => n3389);
   U6564 : BUF_X1 port map( A => n3284, Z => n3375);
   U6565 : BUF_X1 port map( A => n3285, Z => n3377);
   U6566 : BUF_X1 port map( A => n3286, Z => n3379);
   U6567 : BUF_X1 port map( A => n3286, Z => n3381);
   U6568 : BUF_X1 port map( A => n3287, Z => n3383);
   U6569 : BUF_X1 port map( A => n3288, Z => n3385);
   U6570 : BUF_X1 port map( A => n3288, Z => n3387);
   U6571 : BUF_X1 port map( A => n3287, Z => n3384);
   U6572 : BUF_X1 port map( A => n3288, Z => n3386);
   U6573 : BUF_X1 port map( A => n3289, Z => n3388);
   U6574 : BUF_X1 port map( A => n3285, Z => n3376);
   U6575 : BUF_X1 port map( A => n3285, Z => n3378);
   U6576 : BUF_X1 port map( A => n3286, Z => n3380);
   U6577 : BUF_X1 port map( A => n3289, Z => n3390);
   U6578 : BUF_X1 port map( A => n3402, Z => n3505);
   U6579 : BUF_X1 port map( A => n3402, Z => n3504);
   U6580 : BUF_X1 port map( A => n3402, Z => n3503);
   U6581 : BUF_X1 port map( A => n3399, Z => n3494);
   U6582 : BUF_X1 port map( A => n3401, Z => n3501);
   U6583 : BUF_X1 port map( A => n3396, Z => n3487);
   U6584 : BUF_X1 port map( A => n3397, Z => n3489);
   U6585 : BUF_X1 port map( A => n3398, Z => n3491);
   U6586 : BUF_X1 port map( A => n3398, Z => n3493);
   U6587 : BUF_X1 port map( A => n3399, Z => n3495);
   U6588 : BUF_X1 port map( A => n3400, Z => n3497);
   U6589 : BUF_X1 port map( A => n3400, Z => n3499);
   U6590 : BUF_X1 port map( A => n3397, Z => n3488);
   U6591 : BUF_X1 port map( A => n3398, Z => n3492);
   U6592 : BUF_X1 port map( A => n3401, Z => n3502);
   U6593 : BUF_X1 port map( A => n3397, Z => n3490);
   U6594 : BUF_X1 port map( A => n3399, Z => n3496);
   U6595 : BUF_X1 port map( A => n3400, Z => n3498);
   U6596 : BUF_X1 port map( A => n3401, Z => n3500);
   U6597 : BUF_X1 port map( A => n3514, Z => n3617);
   U6598 : BUF_X1 port map( A => n3514, Z => n3616);
   U6599 : BUF_X1 port map( A => n3514, Z => n3615);
   U6600 : BUF_X1 port map( A => n3511, Z => n3606);
   U6601 : BUF_X1 port map( A => n3513, Z => n3613);
   U6602 : BUF_X1 port map( A => n3508, Z => n3599);
   U6603 : BUF_X1 port map( A => n3509, Z => n3601);
   U6604 : BUF_X1 port map( A => n3510, Z => n3603);
   U6605 : BUF_X1 port map( A => n3510, Z => n3605);
   U6606 : BUF_X1 port map( A => n3511, Z => n3607);
   U6607 : BUF_X1 port map( A => n3512, Z => n3609);
   U6608 : BUF_X1 port map( A => n3512, Z => n3611);
   U6609 : BUF_X1 port map( A => n3509, Z => n3600);
   U6610 : BUF_X1 port map( A => n3510, Z => n3604);
   U6611 : BUF_X1 port map( A => n3513, Z => n3614);
   U6612 : BUF_X1 port map( A => n3509, Z => n3602);
   U6613 : BUF_X1 port map( A => n3511, Z => n3608);
   U6614 : BUF_X1 port map( A => n3512, Z => n3610);
   U6615 : BUF_X1 port map( A => n3513, Z => n3612);
   U6616 : BUF_X1 port map( A => n3738, Z => n3841);
   U6617 : BUF_X1 port map( A => n3738, Z => n3840);
   U6618 : BUF_X1 port map( A => n3738, Z => n3839);
   U6619 : BUF_X1 port map( A => n3735, Z => n3830);
   U6620 : BUF_X1 port map( A => n3737, Z => n3837);
   U6621 : BUF_X1 port map( A => n3732, Z => n3823);
   U6622 : BUF_X1 port map( A => n3733, Z => n3825);
   U6623 : BUF_X1 port map( A => n3734, Z => n3827);
   U6624 : BUF_X1 port map( A => n3734, Z => n3829);
   U6625 : BUF_X1 port map( A => n3735, Z => n3831);
   U6626 : BUF_X1 port map( A => n3736, Z => n3833);
   U6627 : BUF_X1 port map( A => n3736, Z => n3835);
   U6628 : BUF_X1 port map( A => n3733, Z => n3824);
   U6629 : BUF_X1 port map( A => n3734, Z => n3828);
   U6630 : BUF_X1 port map( A => n3737, Z => n3838);
   U6631 : BUF_X1 port map( A => n3733, Z => n3826);
   U6632 : BUF_X1 port map( A => n3735, Z => n3832);
   U6633 : BUF_X1 port map( A => n3736, Z => n3834);
   U6634 : BUF_X1 port map( A => n3737, Z => n3836);
   U6635 : BUF_X1 port map( A => n3291, Z => n3394);
   U6636 : BUF_X1 port map( A => n3403, Z => n3506);
   U6637 : BUF_X1 port map( A => n3515, Z => n3618);
   U6638 : BUF_X1 port map( A => n3739, Z => n3842);
   U6639 : BUF_X1 port map( A => n3254, Z => n3207);
   U6640 : BUF_X1 port map( A => n3254, Z => n3210);
   U6641 : BUF_X1 port map( A => n3251, Z => n3225);
   U6642 : BUF_X1 port map( A => n3250, Z => n3231);
   U6643 : BUF_X1 port map( A => n3250, Z => n3228);
   U6644 : BUF_X1 port map( A => n3249, Z => n3234);
   U6645 : BUF_X1 port map( A => n3253, Z => n3213);
   U6646 : BUF_X1 port map( A => n3248, Z => n3237);
   U6647 : BUF_X1 port map( A => n3248, Z => n3240);
   U6648 : BUF_X1 port map( A => n3253, Z => n3216);
   U6649 : BUF_X1 port map( A => n3254, Z => n3208);
   U6650 : BUF_X1 port map( A => n3253, Z => n3214);
   U6651 : BUF_X1 port map( A => n3254, Z => n3211);
   U6652 : BUF_X1 port map( A => n3252, Z => n3219);
   U6653 : BUF_X1 port map( A => n3252, Z => n3217);
   U6654 : BUF_X1 port map( A => n3252, Z => n3220);
   U6655 : BUF_X1 port map( A => n3251, Z => n3226);
   U6656 : BUF_X1 port map( A => n3249, Z => n3232);
   U6657 : BUF_X1 port map( A => n3250, Z => n3229);
   U6658 : BUF_X1 port map( A => n3251, Z => n3222);
   U6659 : BUF_X1 port map( A => n3249, Z => n3235);
   U6660 : BUF_X1 port map( A => n3248, Z => n3241);
   U6661 : BUF_X1 port map( A => n3251, Z => n3223);
   U6662 : BUF_X1 port map( A => n3248, Z => n3238);
   U6663 : BUF_X1 port map( A => n3253, Z => n3215);
   U6664 : BUF_X1 port map( A => n3253, Z => n3212);
   U6665 : BUF_X1 port map( A => n3254, Z => n3209);
   U6666 : BUF_X1 port map( A => n3252, Z => n3218);
   U6667 : BUF_X1 port map( A => n3249, Z => n3236);
   U6668 : BUF_X1 port map( A => n3250, Z => n3227);
   U6669 : BUF_X1 port map( A => n3252, Z => n3221);
   U6670 : BUF_X1 port map( A => n3249, Z => n3233);
   U6671 : BUF_X1 port map( A => n3251, Z => n3224);
   U6672 : BUF_X1 port map( A => n3250, Z => n3230);
   U6673 : BUF_X1 port map( A => n3248, Z => n3239);
   U6674 : BUF_X1 port map( A => n3247, Z => n3244);
   U6675 : BUF_X1 port map( A => n3247, Z => n3245);
   U6676 : BUF_X1 port map( A => n3247, Z => n3243);
   U6677 : BUF_X1 port map( A => n3247, Z => n3242);
   U6678 : BUF_X1 port map( A => n3255, Z => n3204);
   U6679 : BUF_X1 port map( A => n3255, Z => n3205);
   U6680 : BUF_X1 port map( A => n3255, Z => n3206);
   U6681 : BUF_X1 port map( A => n3091, Z => n3103);
   U6682 : BUF_X1 port map( A => n3091, Z => n3106);
   U6683 : BUF_X1 port map( A => n3092, Z => n3109);
   U6684 : BUF_X1 port map( A => n3095, Z => n3124);
   U6685 : BUF_X1 port map( A => n3096, Z => n3130);
   U6686 : BUF_X1 port map( A => n3095, Z => n3127);
   U6687 : BUF_X1 port map( A => n3097, Z => n3133);
   U6688 : BUF_X1 port map( A => n3092, Z => n3112);
   U6689 : BUF_X1 port map( A => n3097, Z => n3136);
   U6690 : BUF_X1 port map( A => n3098, Z => n3139);
   U6691 : BUF_X1 port map( A => n3093, Z => n3115);
   U6692 : BUF_X1 port map( A => n3091, Z => n3104);
   U6693 : BUF_X1 port map( A => n3091, Z => n3107);
   U6694 : BUF_X1 port map( A => n3093, Z => n3113);
   U6695 : BUF_X1 port map( A => n3092, Z => n3110);
   U6696 : BUF_X1 port map( A => n3094, Z => n3118);
   U6697 : BUF_X1 port map( A => n3093, Z => n3116);
   U6698 : BUF_X1 port map( A => n3094, Z => n3119);
   U6699 : BUF_X1 port map( A => n3095, Z => n3125);
   U6700 : BUF_X1 port map( A => n3096, Z => n3131);
   U6701 : BUF_X1 port map( A => n3096, Z => n3128);
   U6702 : BUF_X1 port map( A => n3094, Z => n3121);
   U6703 : BUF_X1 port map( A => n3097, Z => n3134);
   U6704 : BUF_X1 port map( A => n3098, Z => n3140);
   U6705 : BUF_X1 port map( A => n3094, Z => n3122);
   U6706 : BUF_X1 port map( A => n3097, Z => n3137);
   U6707 : BUF_X1 port map( A => n3093, Z => n3114);
   U6708 : BUF_X1 port map( A => n3091, Z => n3105);
   U6709 : BUF_X1 port map( A => n3098, Z => n3142);
   U6710 : BUF_X1 port map( A => n3092, Z => n3111);
   U6711 : BUF_X1 port map( A => n3092, Z => n3108);
   U6712 : BUF_X1 port map( A => n3093, Z => n3117);
   U6713 : BUF_X1 port map( A => n3097, Z => n3135);
   U6714 : BUF_X1 port map( A => n3095, Z => n3126);
   U6715 : BUF_X1 port map( A => n3094, Z => n3120);
   U6716 : BUF_X1 port map( A => n3096, Z => n3132);
   U6717 : BUF_X1 port map( A => n3095, Z => n3123);
   U6718 : BUF_X1 port map( A => n3096, Z => n3129);
   U6719 : BUF_X1 port map( A => n3098, Z => n3138);
   U6720 : BUF_X1 port map( A => n3098, Z => n3141);
   U6721 : BUF_X1 port map( A => n3099, Z => n3143);
   U6722 : BUF_X1 port map( A => n3099, Z => n3144);
   U6723 : BUF_X1 port map( A => n3199, Z => n3152);
   U6724 : BUF_X1 port map( A => n3199, Z => n3155);
   U6725 : BUF_X1 port map( A => n3196, Z => n3170);
   U6726 : BUF_X1 port map( A => n3195, Z => n3176);
   U6727 : BUF_X1 port map( A => n3195, Z => n3173);
   U6728 : BUF_X1 port map( A => n3194, Z => n3179);
   U6729 : BUF_X1 port map( A => n3198, Z => n3158);
   U6730 : BUF_X1 port map( A => n3193, Z => n3182);
   U6731 : BUF_X1 port map( A => n3193, Z => n3185);
   U6732 : BUF_X1 port map( A => n3198, Z => n3161);
   U6733 : BUF_X1 port map( A => n3199, Z => n3153);
   U6734 : BUF_X1 port map( A => n3198, Z => n3159);
   U6735 : BUF_X1 port map( A => n3199, Z => n3156);
   U6736 : BUF_X1 port map( A => n3197, Z => n3164);
   U6737 : BUF_X1 port map( A => n3197, Z => n3162);
   U6738 : BUF_X1 port map( A => n3197, Z => n3165);
   U6739 : BUF_X1 port map( A => n3196, Z => n3171);
   U6740 : BUF_X1 port map( A => n3194, Z => n3177);
   U6741 : BUF_X1 port map( A => n3195, Z => n3174);
   U6742 : BUF_X1 port map( A => n3196, Z => n3167);
   U6743 : BUF_X1 port map( A => n3194, Z => n3180);
   U6744 : BUF_X1 port map( A => n3193, Z => n3186);
   U6745 : BUF_X1 port map( A => n3196, Z => n3168);
   U6746 : BUF_X1 port map( A => n3193, Z => n3183);
   U6747 : BUF_X1 port map( A => n3198, Z => n3160);
   U6748 : BUF_X1 port map( A => n3198, Z => n3157);
   U6749 : BUF_X1 port map( A => n3199, Z => n3154);
   U6750 : BUF_X1 port map( A => n3197, Z => n3163);
   U6751 : BUF_X1 port map( A => n3194, Z => n3181);
   U6752 : BUF_X1 port map( A => n3195, Z => n3172);
   U6753 : BUF_X1 port map( A => n3197, Z => n3166);
   U6754 : BUF_X1 port map( A => n3194, Z => n3178);
   U6755 : BUF_X1 port map( A => n3196, Z => n3169);
   U6756 : BUF_X1 port map( A => n3195, Z => n3175);
   U6757 : BUF_X1 port map( A => n3193, Z => n3184);
   U6758 : BUF_X1 port map( A => n3192, Z => n3189);
   U6759 : BUF_X1 port map( A => n3192, Z => n3190);
   U6760 : BUF_X1 port map( A => n3192, Z => n3188);
   U6761 : BUF_X1 port map( A => n3192, Z => n3187);
   U6762 : BUF_X1 port map( A => n3200, Z => n3149);
   U6763 : BUF_X1 port map( A => n3200, Z => n3150);
   U6764 : BUF_X1 port map( A => n3200, Z => n3151);
   U6765 : BUF_X1 port map( A => n3036, Z => n3048);
   U6766 : BUF_X1 port map( A => n3036, Z => n3051);
   U6767 : BUF_X1 port map( A => n3037, Z => n3054);
   U6768 : BUF_X1 port map( A => n3040, Z => n3069);
   U6769 : BUF_X1 port map( A => n3041, Z => n3075);
   U6770 : BUF_X1 port map( A => n3040, Z => n3072);
   U6771 : BUF_X1 port map( A => n3042, Z => n3078);
   U6772 : BUF_X1 port map( A => n3037, Z => n3057);
   U6773 : BUF_X1 port map( A => n3042, Z => n3081);
   U6774 : BUF_X1 port map( A => n3043, Z => n3084);
   U6775 : BUF_X1 port map( A => n3038, Z => n3060);
   U6776 : BUF_X1 port map( A => n3036, Z => n3049);
   U6777 : BUF_X1 port map( A => n3036, Z => n3052);
   U6778 : BUF_X1 port map( A => n3038, Z => n3058);
   U6779 : BUF_X1 port map( A => n3037, Z => n3055);
   U6780 : BUF_X1 port map( A => n3039, Z => n3063);
   U6781 : BUF_X1 port map( A => n3038, Z => n3061);
   U6782 : BUF_X1 port map( A => n3039, Z => n3064);
   U6783 : BUF_X1 port map( A => n3040, Z => n3070);
   U6784 : BUF_X1 port map( A => n3041, Z => n3076);
   U6785 : BUF_X1 port map( A => n3041, Z => n3073);
   U6786 : BUF_X1 port map( A => n3039, Z => n3066);
   U6787 : BUF_X1 port map( A => n3042, Z => n3079);
   U6788 : BUF_X1 port map( A => n3043, Z => n3085);
   U6789 : BUF_X1 port map( A => n3039, Z => n3067);
   U6790 : BUF_X1 port map( A => n3042, Z => n3082);
   U6791 : BUF_X1 port map( A => n3038, Z => n3059);
   U6792 : BUF_X1 port map( A => n3036, Z => n3050);
   U6793 : BUF_X1 port map( A => n3043, Z => n3087);
   U6794 : BUF_X1 port map( A => n3037, Z => n3056);
   U6795 : BUF_X1 port map( A => n3037, Z => n3053);
   U6796 : BUF_X1 port map( A => n3038, Z => n3062);
   U6797 : BUF_X1 port map( A => n3042, Z => n3080);
   U6798 : BUF_X1 port map( A => n3040, Z => n3071);
   U6799 : BUF_X1 port map( A => n3039, Z => n3065);
   U6800 : BUF_X1 port map( A => n3041, Z => n3077);
   U6801 : BUF_X1 port map( A => n3040, Z => n3068);
   U6802 : BUF_X1 port map( A => n3041, Z => n3074);
   U6803 : BUF_X1 port map( A => n3043, Z => n3083);
   U6804 : BUF_X1 port map( A => n3043, Z => n3086);
   U6805 : BUF_X1 port map( A => n3044, Z => n3088);
   U6806 : BUF_X1 port map( A => n3044, Z => n3089);
   U6807 : NOR2_X1 port map( A1 => n11433, A2 => n11434, ZN => 
                           DataPath_RF_RDPORT_SPILL_n341);
   U6808 : BUF_X1 port map( A => n4223, Z => n4220);
   U6809 : NAND2_X1 port map( A1 => n4259, A2 => n4155, ZN => 
                           DataPath_WRF_CUhw_n112);
   U6810 : BUF_X1 port map( A => n4223, Z => n4219);
   U6811 : BUF_X1 port map( A => n4223, Z => n4218);
   U6812 : BUF_X1 port map( A => n4222, Z => n4221);
   U6813 : BUF_X1 port map( A => n4229, Z => n4202);
   U6814 : BUF_X1 port map( A => n4224, Z => n4216);
   U6815 : BUF_X1 port map( A => n4224, Z => n4215);
   U6816 : BUF_X1 port map( A => n4225, Z => n4214);
   U6817 : BUF_X1 port map( A => n4225, Z => n4213);
   U6818 : BUF_X1 port map( A => n4225, Z => n4212);
   U6819 : BUF_X1 port map( A => n4226, Z => n4211);
   U6820 : BUF_X1 port map( A => n4226, Z => n4210);
   U6821 : BUF_X1 port map( A => n4226, Z => n4209);
   U6822 : BUF_X1 port map( A => n4227, Z => n4208);
   U6823 : BUF_X1 port map( A => n4227, Z => n4207);
   U6824 : BUF_X1 port map( A => n4227, Z => n4206);
   U6825 : BUF_X1 port map( A => n4228, Z => n4205);
   U6826 : BUF_X1 port map( A => n4228, Z => n4204);
   U6827 : BUF_X1 port map( A => n4228, Z => n4203);
   U6828 : BUF_X1 port map( A => n4235, Z => n4182);
   U6829 : BUF_X1 port map( A => n4236, Z => n4181);
   U6830 : BUF_X1 port map( A => n4237, Z => n4180);
   U6831 : BUF_X1 port map( A => n4237, Z => n4179);
   U6832 : BUF_X1 port map( A => n4238, Z => n4178);
   U6833 : BUF_X1 port map( A => n4238, Z => n4177);
   U6834 : BUF_X1 port map( A => n4238, Z => n4176);
   U6835 : BUF_X1 port map( A => n4239, Z => n4175);
   U6836 : BUF_X1 port map( A => n4239, Z => n4174);
   U6837 : BUF_X1 port map( A => n4239, Z => n4173);
   U6838 : BUF_X1 port map( A => n4240, Z => n4171);
   U6839 : BUF_X1 port map( A => n4240, Z => n4170);
   U6840 : BUF_X1 port map( A => n4241, Z => n4169);
   U6841 : BUF_X1 port map( A => n4241, Z => n4168);
   U6842 : BUF_X1 port map( A => n4241, Z => n4167);
   U6843 : BUF_X1 port map( A => n4242, Z => n4166);
   U6844 : BUF_X1 port map( A => n4242, Z => n4165);
   U6845 : BUF_X1 port map( A => n4242, Z => n4164);
   U6846 : BUF_X1 port map( A => n4243, Z => n4163);
   U6847 : BUF_X1 port map( A => n4243, Z => n4162);
   U6848 : BUF_X1 port map( A => n4243, Z => n4161);
   U6849 : BUF_X1 port map( A => n4244, Z => n4160);
   U6850 : BUF_X1 port map( A => n4244, Z => n4159);
   U6851 : BUF_X1 port map( A => n4244, Z => n4158);
   U6852 : BUF_X1 port map( A => n4240, Z => n4172);
   U6853 : BUF_X1 port map( A => n4229, Z => n4201);
   U6854 : BUF_X1 port map( A => n4229, Z => n4200);
   U6855 : BUF_X1 port map( A => n4230, Z => n4199);
   U6856 : BUF_X1 port map( A => n4230, Z => n4198);
   U6857 : BUF_X1 port map( A => n4230, Z => n4197);
   U6858 : BUF_X1 port map( A => n4231, Z => n4196);
   U6859 : BUF_X1 port map( A => n4231, Z => n4195);
   U6860 : BUF_X1 port map( A => n4231, Z => n4194);
   U6861 : BUF_X1 port map( A => n4232, Z => n4193);
   U6862 : BUF_X1 port map( A => n4232, Z => n4192);
   U6863 : BUF_X1 port map( A => n4232, Z => n4191);
   U6864 : BUF_X1 port map( A => n4233, Z => n4190);
   U6865 : BUF_X1 port map( A => n4233, Z => n4189);
   U6866 : BUF_X1 port map( A => n4233, Z => n4188);
   U6867 : BUF_X1 port map( A => n4234, Z => n4187);
   U6868 : BUF_X1 port map( A => n4234, Z => n4186);
   U6869 : BUF_X1 port map( A => n4234, Z => n4185);
   U6870 : BUF_X1 port map( A => n4235, Z => n4184);
   U6871 : BUF_X1 port map( A => n4235, Z => n4183);
   U6872 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n338, A2 => 
                           DataPath_RF_RDPORT_SPILL_n339, ZN => 
                           DataPath_RF_RDPORT_SPILL_n10);
   U6873 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n341, A2 => 
                           DataPath_RF_RDPORT_SPILL_n339, ZN => 
                           DataPath_RF_RDPORT_SPILL_n17);
   U6874 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n346, A2 => 
                           DataPath_RF_RDPORT_SPILL_n341, ZN => 
                           DataPath_RF_RDPORT_SPILL_n23);
   U6875 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n346, A2 => 
                           DataPath_RF_RDPORT_SPILL_n338, ZN => 
                           DataPath_RF_RDPORT_SPILL_n24);
   U6876 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n346, A2 => 
                           DataPath_RF_RDPORT_SPILL_n336, ZN => 
                           DataPath_RF_RDPORT_SPILL_n26);
   U6877 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n346, A2 => 
                           DataPath_RF_RDPORT_SPILL_n340, ZN => 
                           DataPath_RF_RDPORT_SPILL_n27);
   U6878 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n340, A2 => 
                           DataPath_RF_RDPORT_SPILL_n337, ZN => 
                           DataPath_RF_RDPORT_SPILL_n12);
   U6879 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n340, A2 => 
                           DataPath_RF_RDPORT_SPILL_n339, ZN => 
                           DataPath_RF_RDPORT_SPILL_n13);
   U6880 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n336, A2 => 
                           DataPath_RF_RDPORT_SPILL_n337, ZN => 
                           DataPath_RF_RDPORT_SPILL_n11);
   U6881 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n336, A2 => 
                           DataPath_RF_RDPORT_SPILL_n339, ZN => 
                           DataPath_RF_RDPORT_SPILL_n16);
   U6882 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n347, A2 => 
                           DataPath_RF_RDPORT_SPILL_n336, ZN => 
                           DataPath_RF_RDPORT_SPILL_n22);
   U6883 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n347, A2 => 
                           DataPath_RF_RDPORT_SPILL_n338, ZN => 
                           DataPath_RF_RDPORT_SPILL_n25);
   U6884 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n347, A2 => 
                           DataPath_RF_RDPORT_SPILL_n340, ZN => 
                           DataPath_RF_RDPORT_SPILL_n28);
   U6885 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n347, A2 => 
                           DataPath_RF_RDPORT_SPILL_n341, ZN => 
                           DataPath_RF_RDPORT_SPILL_n29);
   U6886 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n337, A2 => 
                           DataPath_RF_RDPORT_SPILL_n338, ZN => 
                           DataPath_RF_RDPORT_SPILL_n14);
   U6887 : AND2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n337, A2 => 
                           DataPath_RF_RDPORT_SPILL_n341, ZN => 
                           DataPath_RF_RDPORT_SPILL_n15);
   U6888 : BUF_X1 port map( A => n4224, Z => n4217);
   U6889 : AND2_X1 port map( A1 => n6848, A2 => n6959, ZN => n1862);
   U6890 : XNOR2_X1 port map( A => n7298, B => n7367, ZN => n1863);
   U6891 : XNOR2_X1 port map( A => n5259, B => n5237, ZN => n5239);
   U6892 : XNOR2_X1 port map( A => n688, B => n5229, ZN => n4984);
   U6893 : XNOR2_X1 port map( A => n5040, B => n1864, ZN => n5374);
   U6894 : XNOR2_X1 port map( A => n5039, B => n5038, ZN => n1864);
   U6895 : XNOR2_X1 port map( A => n6791, B => n1865, ZN => n6977);
   U6896 : XNOR2_X1 port map( A => n6790, B => n6789, ZN => n1865);
   U6897 : XNOR2_X1 port map( A => n7299, B => n1329, ZN => n7366);
   U6898 : OAI211_X1 port map( C1 => n6156, C2 => n6155, A => n6154, B => n6153
                           , ZN => n6167);
   U6899 : XNOR2_X1 port map( A => n7321, B => n1866, ZN => n7325);
   U6900 : XNOR2_X1 port map( A => n7320, B => n7319, ZN => n1866);
   U6901 : XNOR2_X1 port map( A => n753, B => n1141, ZN => n5135);
   U6903 : XNOR2_X1 port map( A => n6620, B => n1692, ZN => n1869);
   U6904 : INV_X1 port map( A => n2212, ZN => n2208);
   U6905 : INV_X1 port map( A => n2202, ZN => n2199);
   U6906 : INV_X1 port map( A => n1899, ZN => n2219);
   U6907 : INV_X1 port map( A => n2211, ZN => n2209);
   U6908 : INV_X1 port map( A => n2207, ZN => n2205);
   U6909 : NAND2_X1 port map( A1 => n5298, A2 => n5299, ZN => n5300);
   U6910 : XNOR2_X1 port map( A => n6951, B => n7292, ZN => n6953);
   U6911 : CLKBUF_X1 port map( A => n2239, Z => n2138);
   U6912 : XNOR2_X1 port map( A => n5009, B => n5007, ZN => n5011);
   U6913 : XNOR2_X1 port map( A => n4753, B => n4751, ZN => n4755);
   U6914 : XNOR2_X1 port map( A => n6817, B => n6998, ZN => n6826);
   U6915 : XNOR2_X1 port map( A => n215, B => n6244, ZN => n6248);
   U6916 : XNOR2_X1 port map( A => n6744, B => n6922, ZN => n6750);
   U6917 : XNOR2_X1 port map( A => n4585, B => n4561, ZN => n1870);
   U6918 : XNOR2_X1 port map( A => n7490, B => n1871, ZN => n7491);
   U6919 : INV_X1 port map( A => n8208, ZN => n2263);
   U6920 : AND2_X1 port map( A1 => n1898, A2 => n2154, ZN => n1872);
   U6921 : XNOR2_X1 port map( A => n5016, B => n5014, ZN => n5018);
   U6922 : XNOR2_X1 port map( A => n5775, B => n6732, ZN => n5777);
   U6923 : XNOR2_X1 port map( A => n6264, B => n1194, ZN => n6270);
   U6924 : XNOR2_X1 port map( A => n7325, B => n7332, ZN => n7333);
   U6925 : XNOR2_X1 port map( A => n6873, B => n7322, ZN => n6875);
   U6926 : XNOR2_X1 port map( A => n1263, B => n6682, ZN => n1874);
   U6927 : XNOR2_X1 port map( A => n4740, B => n4746, ZN => n4747);
   U6928 : INV_X1 port map( A => n8208, ZN => n2264);
   U6929 : XNOR2_X1 port map( A => n5021, B => n5023, ZN => n5025);
   U6930 : AND2_X1 port map( A1 => n4899, A2 => n1135, ZN => n1875);
   U6931 : XNOR2_X1 port map( A => n7048, B => n667, ZN => n7049);
   U6932 : AND2_X1 port map( A1 => n6773, A2 => n6765, ZN => n1876);
   U6933 : AND2_X1 port map( A1 => n6773, A2 => n6774, ZN => n1877);
   U6934 : AND2_X1 port map( A1 => n4559, A2 => n1135, ZN => n1878);
   U6935 : XNOR2_X1 port map( A => n5764, B => n6719, ZN => n5766);
   U6936 : XNOR2_X1 port map( A => n6727, B => n6865, ZN => n6729);
   U6937 : XNOR2_X1 port map( A => n6342, B => n1303, ZN => n6368);
   U6938 : XNOR2_X1 port map( A => n6960, B => n1372, ZN => n1879);
   U6939 : XNOR2_X1 port map( A => n7411, B => n7410, ZN => n1880);
   U6940 : XNOR2_X1 port map( A => n7456, B => n7457, ZN => n1882);
   U6941 : AND2_X1 port map( A1 => n5334, A2 => n5304, ZN => n1883);
   U6942 : XNOR2_X1 port map( A => n7470, B => n7469, ZN => n1884);
   U6943 : OR2_X1 port map( A1 => n6077, A2 => n6076, ZN => n6250);
   U6944 : XNOR2_X1 port map( A => n6450, B => n6452, ZN => n6453);
   U6945 : NAND2_X1 port map( A1 => n7510, A2 => n7509, ZN => n7511);
   U6946 : NAND2_X1 port map( A1 => n7506, A2 => n7505, ZN => n7512);
   U6947 : AND2_X1 port map( A1 => n600, A2 => n5824, ZN => n1885);
   U6948 : XNOR2_X1 port map( A => n2161, B => n624, ZN => n6331);
   U6949 : XNOR2_X1 port map( A => n6320, B => n6318, ZN => n6321);
   U6950 : AND2_X1 port map( A1 => n867, A2 => n5887, ZN => n1886);
   U6951 : AND2_X1 port map( A1 => n5797, A2 => n5796, ZN => n1887);
   U6952 : XNOR2_X1 port map( A => n17154, B => n6302, ZN => n1889);
   U6953 : OR2_X1 port map( A1 => n6159, A2 => n6163, ZN => n6154);
   U6954 : INV_X1 port map( A => n1374, ZN => n2197);
   U6955 : AND2_X1 port map( A1 => n5962, A2 => n2154, ZN => n1892);
   U6956 : CLKBUF_X1 port map( A => n799, Z => n2249);
   U6957 : AND2_X1 port map( A1 => n5716, A2 => n2154, ZN => n1893);
   U6958 : INV_X1 port map( A => n4134, ZN => n4129);
   U6959 : NOR3_X1 port map( A1 => n4155, A2 => n11607, A3 => 
                           DataPath_i_DONE_SPILL_EX, ZN => 
                           DataPath_WRF_CUhw_N217);
   U6960 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n2, A2 => 
                           DataPath_ALUhw_MUXOUT_n3, ZN => 
                           DataPath_i_ALU_OUT_9_port);
   U6961 : AOI22_X1 port map( A1 => n11508, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_105_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n2);
   U6962 : INV_X1 port map( A => n12897, ZN => n11508);
   U6963 : BUF_X1 port map( A => n3910, Z => n3902);
   U6964 : AND2_X1 port map( A1 => n6332, A2 => n2154, ZN => n1894);
   U6965 : BUF_X1 port map( A => n3910, Z => n3901);
   U6966 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n54, A2 => 
                           DataPath_ALUhw_MUXOUT_n55, ZN => 
                           DataPath_i_ALU_OUT_16_port);
   U6967 : AOI22_X1 port map( A1 => n11501, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_112_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n54);
   U6968 : AOI22_X1 port map( A1 => DataPath_ALUhw_i_Q_EXTENDED_80_port, A2 => 
                           n8322, B1 => n11584, B2 => n2258, ZN => 
                           DataPath_ALUhw_MUXOUT_n55);
   U6969 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n58, A2 => 
                           DataPath_ALUhw_MUXOUT_n59, ZN => 
                           DataPath_i_ALU_OUT_14_port);
   U6970 : AOI22_X1 port map( A1 => n11504, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_110_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n58);
   U6971 : AOI22_X1 port map( A1 => DataPath_ALUhw_i_Q_EXTENDED_78_port, A2 => 
                           n8322, B1 => n11586, B2 => n2258, ZN => 
                           DataPath_ALUhw_MUXOUT_n59);
   U6972 : INV_X1 port map( A => n12899, ZN => n11504);
   U6973 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n60, A2 => 
                           DataPath_ALUhw_MUXOUT_n61, ZN => 
                           DataPath_i_ALU_OUT_13_port);
   U6974 : AOI22_X1 port map( A1 => n11503, A2 => n2272, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_109_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n60);
   U6975 : INV_X1 port map( A => n12900, ZN => n11503);
   U6976 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n56, A2 => 
                           DataPath_ALUhw_MUXOUT_n57, ZN => 
                           DataPath_i_ALU_OUT_15_port);
   U6977 : AOI22_X1 port map( A1 => n11505, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_111_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n56);
   U6978 : AOI22_X1 port map( A1 => DataPath_ALUhw_i_Q_EXTENDED_79_port, A2 => 
                           n8322, B1 => n11585, B2 => n2258, ZN => 
                           DataPath_ALUhw_MUXOUT_n57);
   U6979 : INV_X1 port map( A => n12898, ZN => n11505);
   U6980 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n62, A2 => 
                           DataPath_ALUhw_MUXOUT_n63, ZN => 
                           DataPath_i_ALU_OUT_12_port);
   U6981 : AOI22_X1 port map( A1 => n11502, A2 => n2272, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_108_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n62);
   U6982 : AOI22_X1 port map( A1 => DataPath_ALUhw_i_Q_EXTENDED_76_port, A2 => 
                           n8322, B1 => n11587, B2 => n2258, ZN => 
                           DataPath_ALUhw_MUXOUT_n63);
   U6983 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n64, A2 => 
                           DataPath_ALUhw_MUXOUT_n65, ZN => 
                           DataPath_i_ALU_OUT_11_port);
   U6984 : AOI22_X1 port map( A1 => n11510, A2 => n2272, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_107_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n64);
   U6985 : INV_X1 port map( A => n12895, ZN => n11510);
   U6986 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n66, A2 => 
                           DataPath_ALUhw_MUXOUT_n67, ZN => 
                           DataPath_i_ALU_OUT_10_port);
   U6987 : AOI22_X1 port map( A1 => n11509, A2 => n2272, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_106_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n66);
   U6988 : INV_X1 port map( A => n12896, ZN => n11509);
   U6989 : NAND3_X1 port map( A1 => n7747, A2 => n17175, A3 => n2260, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n191);
   U6990 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n600, ZN => n8073);
   U6991 : INV_X1 port map( A => n4134, ZN => n4130);
   U6992 : INV_X1 port map( A => n4134, ZN => n4131);
   U6993 : AOI21_X1 port map( B1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_8_port, B2 
                           => n11516, A => n11534, ZN => n12927);
   U6994 : AND2_X1 port map( A1 => n374, A2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_6_port, ZN 
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_8_port);
   U6995 : OAI22_X1 port map( A1 => n8318, A2 => DataPath_ALUhw_SHIFTER_HW_n191
                           , B1 => n8308, B2 => DataPath_ALUhw_SHIFTER_HW_n192,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n282);
   U6996 : OAI22_X1 port map( A1 => n8316, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8317, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n275);
   U6997 : INV_X1 port map( A => n11539, ZN => n7207);
   U6998 : OAI221_X1 port map( B1 => n11363, B2 => n11577, C1 => n11578, C2 => 
                           DataPath_LDSTR_n39, A => DataPath_LDSTR_n38, ZN => 
                           DRAM_DATA_OUT_8_port);
   U6999 : OAI221_X1 port map( B1 => n11361, B2 => n11577, C1 => 
                           DataPath_LDSTR_n37, C2 => n11578, A => 
                           DataPath_LDSTR_n38, ZN => DRAM_DATA_OUT_9_port);
   U7000 : OAI221_X1 port map( B1 => n11359, B2 => n11577, C1 => n11578, C2 => 
                           DataPath_LDSTR_n54, A => DataPath_LDSTR_n38, ZN => 
                           DRAM_DATA_OUT_10_port);
   U7001 : OAI221_X1 port map( B1 => n11357, B2 => n11577, C1 => n11578, C2 => 
                           DataPath_LDSTR_n52, A => DataPath_LDSTR_n38, ZN => 
                           DRAM_DATA_OUT_11_port);
   U7002 : OAI221_X1 port map( B1 => n11355, B2 => n11577, C1 => n11578, C2 => 
                           DataPath_LDSTR_n50, A => DataPath_LDSTR_n38, ZN => 
                           DRAM_DATA_OUT_12_port);
   U7003 : OAI221_X1 port map( B1 => n11353, B2 => n11577, C1 => n11578, C2 => 
                           DataPath_LDSTR_n48, A => DataPath_LDSTR_n38, ZN => 
                           DRAM_DATA_OUT_13_port);
   U7004 : OAI221_X1 port map( B1 => n11351, B2 => n11577, C1 => n11578, C2 => 
                           DataPath_LDSTR_n43, A => DataPath_LDSTR_n38, ZN => 
                           DRAM_DATA_OUT_14_port);
   U7005 : AND2_X1 port map( A1 => DataPath_LDSTR_n78, A2 => n11580, ZN => 
                           DataPath_LDSTR_n58);
   U7006 : OR2_X1 port map( A1 => DataPath_LDSTR_n62, A2 => n4128, ZN => 
                           DataPath_LDSTR_n38);
   U7007 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n8, A2 => 
                           DataPath_ALUhw_MUXOUT_n9, ZN => 
                           DataPath_i_ALU_OUT_8_port);
   U7008 : AOI22_X1 port map( A1 => n11507, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_104_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n8);
   U7009 : INV_X1 port map( A => n12959, ZN => n11399);
   U7010 : OAI211_X1 port map( C1 => DataPath_ALUhw_SHIFTER_HW_n529, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n600, A => 
                           DataPath_ALUhw_SHIFTER_HW_n621, B => 
                           DataPath_ALUhw_SHIFTER_HW_n622, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n269);
   U7011 : OAI211_X1 port map( C1 => DataPath_ALUhw_SHIFTER_HW_n540, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n600, A => 
                           DataPath_ALUhw_SHIFTER_HW_n625, B => 
                           DataPath_ALUhw_SHIFTER_HW_n626, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n419);
   U7012 : OAI211_X1 port map( C1 => DataPath_ALUhw_SHIFTER_HW_n411, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n600, A => 
                           DataPath_ALUhw_SHIFTER_HW_n635, B => 
                           DataPath_ALUhw_SHIFTER_HW_n636, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n588);
   U7013 : NAND2_X1 port map( A1 => n1896, A2 => n4134, ZN => n8031);
   U7014 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n548, ZN => n7989);
   U7015 : BUF_X1 port map( A => n14397, Z => n2515);
   U7016 : BUF_X1 port map( A => n14907, Z => n2605);
   U7017 : BUF_X1 port map( A => n14941, Z => n2611);
   U7018 : BUF_X1 port map( A => n14975, Z => n2617);
   U7019 : BUF_X1 port map( A => n15009, Z => n2623);
   U7020 : BUF_X1 port map( A => n15043, Z => n2629);
   U7021 : BUF_X1 port map( A => n15077, Z => n2635);
   U7022 : BUF_X1 port map( A => n15111, Z => n2641);
   U7023 : BUF_X1 port map( A => n15145, Z => n2647);
   U7024 : BUF_X1 port map( A => n15451, Z => n2701);
   U7025 : BUF_X1 port map( A => n15485, Z => n2707);
   U7026 : BUF_X1 port map( A => n15519, Z => n2713);
   U7027 : BUF_X1 port map( A => n15553, Z => n2719);
   U7028 : BUF_X1 port map( A => n15587, Z => n2725);
   U7029 : BUF_X1 port map( A => n15621, Z => n2731);
   U7030 : BUF_X1 port map( A => n15655, Z => n2737);
   U7031 : BUF_X1 port map( A => n15689, Z => n2743);
   U7032 : BUF_X1 port map( A => n15995, Z => n2797);
   U7033 : BUF_X1 port map( A => n16029, Z => n2803);
   U7034 : BUF_X1 port map( A => n16063, Z => n2809);
   U7035 : BUF_X1 port map( A => n16097, Z => n2815);
   U7036 : BUF_X1 port map( A => n16131, Z => n2821);
   U7037 : BUF_X1 port map( A => n16165, Z => n2827);
   U7038 : BUF_X1 port map( A => n16199, Z => n2833);
   U7039 : BUF_X1 port map( A => n16233, Z => n2839);
   U7040 : BUF_X1 port map( A => n16539, Z => n2893);
   U7041 : BUF_X1 port map( A => n16573, Z => n2899);
   U7042 : BUF_X1 port map( A => n14363, Z => n2509);
   U7043 : BUF_X1 port map( A => n14431, Z => n2521);
   U7044 : BUF_X1 port map( A => n14465, Z => n2527);
   U7045 : BUF_X1 port map( A => n14499, Z => n2533);
   U7046 : BUF_X1 port map( A => n14533, Z => n2539);
   U7047 : BUF_X1 port map( A => n14567, Z => n2545);
   U7048 : BUF_X1 port map( A => n14601, Z => n2551);
   U7049 : BUF_X1 port map( A => n16607, Z => n2905);
   U7050 : BUF_X1 port map( A => n16641, Z => n2911);
   U7051 : BUF_X1 port map( A => n16675, Z => n2917);
   U7052 : BUF_X1 port map( A => n16709, Z => n2923);
   U7053 : BUF_X1 port map( A => n16743, Z => n2929);
   U7054 : BUF_X1 port map( A => n16777, Z => n2935);
   U7055 : BUF_X1 port map( A => n14635, Z => n2557);
   U7056 : BUF_X1 port map( A => n14669, Z => n2563);
   U7057 : BUF_X1 port map( A => n14703, Z => n2569);
   U7058 : BUF_X1 port map( A => n14737, Z => n2575);
   U7059 : BUF_X1 port map( A => n14771, Z => n2581);
   U7060 : BUF_X1 port map( A => n14805, Z => n2587);
   U7061 : BUF_X1 port map( A => n14839, Z => n2593);
   U7062 : BUF_X1 port map( A => n14873, Z => n2599);
   U7063 : BUF_X1 port map( A => n15179, Z => n2653);
   U7064 : BUF_X1 port map( A => n15213, Z => n2659);
   U7065 : BUF_X1 port map( A => n15247, Z => n2665);
   U7066 : BUF_X1 port map( A => n15281, Z => n2671);
   U7067 : BUF_X1 port map( A => n15315, Z => n2677);
   U7068 : BUF_X1 port map( A => n15349, Z => n2683);
   U7069 : BUF_X1 port map( A => n15383, Z => n2689);
   U7070 : BUF_X1 port map( A => n15417, Z => n2695);
   U7071 : BUF_X1 port map( A => n15723, Z => n2749);
   U7072 : BUF_X1 port map( A => n15757, Z => n2755);
   U7073 : BUF_X1 port map( A => n15791, Z => n2761);
   U7074 : BUF_X1 port map( A => n15825, Z => n2767);
   U7075 : BUF_X1 port map( A => n15859, Z => n2773);
   U7076 : BUF_X1 port map( A => n15893, Z => n2779);
   U7077 : BUF_X1 port map( A => n15927, Z => n2785);
   U7078 : BUF_X1 port map( A => n15961, Z => n2791);
   U7079 : BUF_X1 port map( A => n16267, Z => n2845);
   U7080 : BUF_X1 port map( A => n16301, Z => n2851);
   U7081 : BUF_X1 port map( A => n16335, Z => n2857);
   U7082 : BUF_X1 port map( A => n16369, Z => n2863);
   U7083 : BUF_X1 port map( A => n16403, Z => n2869);
   U7084 : BUF_X1 port map( A => n16437, Z => n2875);
   U7085 : BUF_X1 port map( A => n16471, Z => n2881);
   U7086 : BUF_X1 port map( A => n16505, Z => n2887);
   U7087 : BUF_X1 port map( A => n16811, Z => n2941);
   U7088 : BUF_X1 port map( A => n16845, Z => n2947);
   U7089 : BUF_X1 port map( A => n16879, Z => n2953);
   U7090 : BUF_X1 port map( A => n16913, Z => n2959);
   U7091 : BUF_X1 port map( A => n16947, Z => n2965);
   U7092 : BUF_X1 port map( A => n16981, Z => n2971);
   U7093 : BUF_X1 port map( A => n17015, Z => n2977);
   U7094 : BUF_X1 port map( A => n17049, Z => n2983);
   U7095 : BUF_X1 port map( A => n14397, Z => n2514);
   U7096 : BUF_X1 port map( A => n14397, Z => n2513);
   U7097 : BUF_X1 port map( A => n14907, Z => n2604);
   U7098 : BUF_X1 port map( A => n14907, Z => n2603);
   U7099 : BUF_X1 port map( A => n14941, Z => n2610);
   U7100 : BUF_X1 port map( A => n14941, Z => n2609);
   U7101 : BUF_X1 port map( A => n14975, Z => n2616);
   U7102 : BUF_X1 port map( A => n14975, Z => n2615);
   U7103 : BUF_X1 port map( A => n15009, Z => n2622);
   U7104 : BUF_X1 port map( A => n15009, Z => n2621);
   U7105 : BUF_X1 port map( A => n15043, Z => n2628);
   U7106 : BUF_X1 port map( A => n15043, Z => n2627);
   U7107 : BUF_X1 port map( A => n15077, Z => n2634);
   U7108 : BUF_X1 port map( A => n15077, Z => n2633);
   U7109 : BUF_X1 port map( A => n15111, Z => n2640);
   U7110 : BUF_X1 port map( A => n15111, Z => n2639);
   U7111 : BUF_X1 port map( A => n15145, Z => n2646);
   U7112 : BUF_X1 port map( A => n15145, Z => n2645);
   U7113 : BUF_X1 port map( A => n15451, Z => n2700);
   U7114 : BUF_X1 port map( A => n15451, Z => n2699);
   U7115 : BUF_X1 port map( A => n15485, Z => n2706);
   U7116 : BUF_X1 port map( A => n15485, Z => n2705);
   U7117 : BUF_X1 port map( A => n15519, Z => n2712);
   U7118 : BUF_X1 port map( A => n15519, Z => n2711);
   U7119 : BUF_X1 port map( A => n15553, Z => n2718);
   U7120 : BUF_X1 port map( A => n15553, Z => n2717);
   U7121 : BUF_X1 port map( A => n15587, Z => n2724);
   U7122 : BUF_X1 port map( A => n15587, Z => n2723);
   U7123 : BUF_X1 port map( A => n15621, Z => n2730);
   U7124 : BUF_X1 port map( A => n15621, Z => n2729);
   U7125 : BUF_X1 port map( A => n15655, Z => n2736);
   U7126 : BUF_X1 port map( A => n15655, Z => n2735);
   U7127 : BUF_X1 port map( A => n15689, Z => n2742);
   U7128 : BUF_X1 port map( A => n15689, Z => n2741);
   U7129 : BUF_X1 port map( A => n15995, Z => n2796);
   U7130 : BUF_X1 port map( A => n15995, Z => n2795);
   U7131 : BUF_X1 port map( A => n16029, Z => n2802);
   U7132 : BUF_X1 port map( A => n16029, Z => n2801);
   U7133 : BUF_X1 port map( A => n16063, Z => n2808);
   U7134 : BUF_X1 port map( A => n16063, Z => n2807);
   U7135 : BUF_X1 port map( A => n16097, Z => n2814);
   U7136 : BUF_X1 port map( A => n16097, Z => n2813);
   U7137 : BUF_X1 port map( A => n16131, Z => n2820);
   U7138 : BUF_X1 port map( A => n16131, Z => n2819);
   U7139 : BUF_X1 port map( A => n16165, Z => n2826);
   U7140 : BUF_X1 port map( A => n16165, Z => n2825);
   U7141 : BUF_X1 port map( A => n16199, Z => n2832);
   U7142 : BUF_X1 port map( A => n16199, Z => n2831);
   U7143 : BUF_X1 port map( A => n16233, Z => n2838);
   U7144 : BUF_X1 port map( A => n16233, Z => n2837);
   U7145 : BUF_X1 port map( A => n16539, Z => n2892);
   U7146 : BUF_X1 port map( A => n16539, Z => n2891);
   U7147 : BUF_X1 port map( A => n16573, Z => n2898);
   U7148 : BUF_X1 port map( A => n16573, Z => n2897);
   U7149 : BUF_X1 port map( A => n14363, Z => n2508);
   U7150 : BUF_X1 port map( A => n14363, Z => n2507);
   U7151 : BUF_X1 port map( A => n14431, Z => n2520);
   U7152 : BUF_X1 port map( A => n14431, Z => n2519);
   U7153 : BUF_X1 port map( A => n14465, Z => n2526);
   U7154 : BUF_X1 port map( A => n14465, Z => n2525);
   U7155 : BUF_X1 port map( A => n14499, Z => n2532);
   U7156 : BUF_X1 port map( A => n14499, Z => n2531);
   U7157 : BUF_X1 port map( A => n14533, Z => n2538);
   U7158 : BUF_X1 port map( A => n14533, Z => n2537);
   U7159 : BUF_X1 port map( A => n14567, Z => n2544);
   U7160 : BUF_X1 port map( A => n14567, Z => n2543);
   U7161 : BUF_X1 port map( A => n14601, Z => n2550);
   U7162 : BUF_X1 port map( A => n14601, Z => n2549);
   U7163 : BUF_X1 port map( A => n16607, Z => n2904);
   U7164 : BUF_X1 port map( A => n16607, Z => n2903);
   U7165 : BUF_X1 port map( A => n16641, Z => n2910);
   U7166 : BUF_X1 port map( A => n16641, Z => n2909);
   U7167 : BUF_X1 port map( A => n16675, Z => n2916);
   U7168 : BUF_X1 port map( A => n16675, Z => n2915);
   U7169 : BUF_X1 port map( A => n16709, Z => n2922);
   U7170 : BUF_X1 port map( A => n16709, Z => n2921);
   U7171 : BUF_X1 port map( A => n16743, Z => n2928);
   U7172 : BUF_X1 port map( A => n16743, Z => n2927);
   U7173 : BUF_X1 port map( A => n16777, Z => n2934);
   U7174 : BUF_X1 port map( A => n16777, Z => n2933);
   U7175 : OAI22_X1 port map( A1 => n11492, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n181, B1 => n8316, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n182, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n250);
   U7176 : BUF_X1 port map( A => n2325, Z => n2327);
   U7177 : BUF_X1 port map( A => n2331, Z => n2333);
   U7178 : BUF_X1 port map( A => n2343, Z => n2345);
   U7179 : BUF_X1 port map( A => n2349, Z => n2351);
   U7180 : BUF_X1 port map( A => n2355, Z => n2357);
   U7181 : BUF_X1 port map( A => n2361, Z => n2363);
   U7182 : BUF_X1 port map( A => n2367, Z => n2369);
   U7183 : BUF_X1 port map( A => n2373, Z => n2375);
   U7184 : BUF_X1 port map( A => n2379, Z => n2381);
   U7185 : BUF_X1 port map( A => n2385, Z => n2387);
   U7186 : BUF_X1 port map( A => n2391, Z => n2393);
   U7187 : BUF_X1 port map( A => n2397, Z => n2399);
   U7188 : BUF_X1 port map( A => n2409, Z => n2411);
   U7189 : BUF_X1 port map( A => n2415, Z => n2417);
   U7190 : BUF_X1 port map( A => n2421, Z => n2423);
   U7191 : BUF_X1 port map( A => n2427, Z => n2429);
   U7192 : BUF_X1 port map( A => n2433, Z => n2435);
   U7193 : BUF_X1 port map( A => n2439, Z => n2441);
   U7194 : BUF_X1 port map( A => n2445, Z => n2447);
   U7195 : BUF_X1 port map( A => n2451, Z => n2453);
   U7196 : BUF_X1 port map( A => n2457, Z => n2459);
   U7197 : BUF_X1 port map( A => n2463, Z => n2465);
   U7198 : BUF_X1 port map( A => n2337, Z => n2339);
   U7199 : BUF_X1 port map( A => n2403, Z => n2405);
   U7200 : BUF_X1 port map( A => n2469, Z => n2471);
   U7201 : BUF_X1 port map( A => n2325, Z => n2328);
   U7202 : BUF_X1 port map( A => n2331, Z => n2334);
   U7203 : BUF_X1 port map( A => n2343, Z => n2346);
   U7204 : BUF_X1 port map( A => n2349, Z => n2352);
   U7205 : BUF_X1 port map( A => n2355, Z => n2358);
   U7206 : BUF_X1 port map( A => n2361, Z => n2364);
   U7207 : BUF_X1 port map( A => n2367, Z => n2370);
   U7208 : BUF_X1 port map( A => n2373, Z => n2376);
   U7209 : BUF_X1 port map( A => n2379, Z => n2382);
   U7210 : BUF_X1 port map( A => n2385, Z => n2388);
   U7211 : BUF_X1 port map( A => n2391, Z => n2394);
   U7212 : BUF_X1 port map( A => n2397, Z => n2400);
   U7213 : BUF_X1 port map( A => n2409, Z => n2412);
   U7214 : BUF_X1 port map( A => n2415, Z => n2418);
   U7215 : BUF_X1 port map( A => n2421, Z => n2424);
   U7216 : BUF_X1 port map( A => n2427, Z => n2430);
   U7217 : BUF_X1 port map( A => n2433, Z => n2436);
   U7218 : BUF_X1 port map( A => n2439, Z => n2442);
   U7219 : BUF_X1 port map( A => n2445, Z => n2448);
   U7220 : BUF_X1 port map( A => n2451, Z => n2454);
   U7221 : BUF_X1 port map( A => n2457, Z => n2460);
   U7222 : BUF_X1 port map( A => n2463, Z => n2466);
   U7223 : BUF_X1 port map( A => n2337, Z => n2340);
   U7224 : BUF_X1 port map( A => n2403, Z => n2406);
   U7225 : BUF_X1 port map( A => n2469, Z => n2472);
   U7226 : BUF_X1 port map( A => n2326, Z => n2329);
   U7227 : BUF_X1 port map( A => n2332, Z => n2335);
   U7228 : BUF_X1 port map( A => n2344, Z => n2347);
   U7229 : BUF_X1 port map( A => n2350, Z => n2353);
   U7230 : BUF_X1 port map( A => n2356, Z => n2359);
   U7231 : BUF_X1 port map( A => n2362, Z => n2365);
   U7232 : BUF_X1 port map( A => n2368, Z => n2371);
   U7233 : BUF_X1 port map( A => n2374, Z => n2377);
   U7234 : BUF_X1 port map( A => n2380, Z => n2383);
   U7235 : BUF_X1 port map( A => n2386, Z => n2389);
   U7236 : BUF_X1 port map( A => n2392, Z => n2395);
   U7237 : BUF_X1 port map( A => n2398, Z => n2401);
   U7238 : BUF_X1 port map( A => n2410, Z => n2413);
   U7239 : BUF_X1 port map( A => n2416, Z => n2419);
   U7240 : BUF_X1 port map( A => n2422, Z => n2425);
   U7241 : BUF_X1 port map( A => n2428, Z => n2431);
   U7242 : BUF_X1 port map( A => n2434, Z => n2437);
   U7243 : BUF_X1 port map( A => n2440, Z => n2443);
   U7244 : BUF_X1 port map( A => n2446, Z => n2449);
   U7245 : BUF_X1 port map( A => n2452, Z => n2455);
   U7246 : BUF_X1 port map( A => n2458, Z => n2461);
   U7247 : BUF_X1 port map( A => n2464, Z => n2467);
   U7248 : BUF_X1 port map( A => n2338, Z => n2341);
   U7249 : BUF_X1 port map( A => n2404, Z => n2407);
   U7250 : BUF_X1 port map( A => n2470, Z => n2473);
   U7251 : OAI221_X2 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n600, B2 => 
                           n8011, C1 => n8010, C2 => n8037, A => n8009, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n151);
   U7252 : OAI221_X2 port map( B1 => n8002, B2 => n8037, C1 => 
                           DataPath_ALUhw_SHIFTER_HW_n411, C2 => n2134, A => 
                           n8001, ZN => DataPath_ALUhw_SHIFTER_HW_n171);
   U7253 : BUF_X1 port map( A => n2284, Z => n2288);
   U7254 : BUF_X1 port map( A => n2290, Z => n2294);
   U7255 : BUF_X1 port map( A => n2296, Z => n2300);
   U7256 : BUF_X1 port map( A => n2302, Z => n2306);
   U7257 : BUF_X1 port map( A => n2308, Z => n2312);
   U7258 : BUF_X1 port map( A => n2314, Z => n2318);
   U7259 : BUF_X1 port map( A => n2320, Z => n2324);
   U7260 : BUF_X1 port map( A => n2284, Z => n2287);
   U7261 : BUF_X1 port map( A => n2290, Z => n2293);
   U7262 : BUF_X1 port map( A => n2296, Z => n2299);
   U7263 : BUF_X1 port map( A => n2302, Z => n2305);
   U7264 : BUF_X1 port map( A => n2308, Z => n2311);
   U7265 : BUF_X1 port map( A => n2314, Z => n2317);
   U7266 : BUF_X1 port map( A => n2320, Z => n2323);
   U7267 : BUF_X1 port map( A => n2283, Z => n2286);
   U7268 : BUF_X1 port map( A => n2289, Z => n2292);
   U7269 : BUF_X1 port map( A => n2295, Z => n2298);
   U7270 : BUF_X1 port map( A => n2301, Z => n2304);
   U7271 : BUF_X1 port map( A => n2307, Z => n2310);
   U7272 : BUF_X1 port map( A => n2313, Z => n2316);
   U7273 : BUF_X1 port map( A => n2319, Z => n2322);
   U7274 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_1_port
                           , A2 => n11506, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_1_port
                           , B2 => n12928, ZN => n12900);
   U7275 : BUF_X1 port map( A => n2326, Z => n2330);
   U7276 : BUF_X1 port map( A => n2283, Z => n2285);
   U7277 : BUF_X1 port map( A => n2289, Z => n2291);
   U7278 : BUF_X1 port map( A => n2295, Z => n2297);
   U7279 : BUF_X1 port map( A => n2301, Z => n2303);
   U7280 : BUF_X1 port map( A => n2307, Z => n2309);
   U7281 : BUF_X1 port map( A => n2313, Z => n2315);
   U7282 : BUF_X1 port map( A => n2319, Z => n2321);
   U7283 : AOI21_X1 port map( B1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_20_port, B2
                           => n8326, A => n11525, ZN => n12930);
   U7284 : AND2_X1 port map( A1 => n7979, A2 => n4265, ZN => n1895);
   U7285 : NAND4_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n582, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n583, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n584, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n585, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_96_port);
   U7286 : AOI222_X1 port map( A1 => n8306, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n588, B1 => n8307, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, C1 => n8312, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n419, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n582);
   U7287 : AOI221_X1 port map( B1 => n8300, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, C1 => n8299, C2 => 
                           n523, A => DataPath_ALUhw_SHIFTER_HW_n586, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n585);
   U7288 : AOI221_X1 port map( B1 => n8314, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n201, C1 => n8309, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n211, A => 
                           DataPath_ALUhw_SHIFTER_HW_n603, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n584);
   U7289 : AOI21_X1 port map( B1 => n11537, B2 => n373, A => n11519, ZN => 
                           n12918);
   U7290 : AOI21_X1 port map( B1 => n11535, B2 => n374, A => n11536, ZN => 
                           n12917);
   U7291 : BUF_X1 port map( A => CU_I_n104, Z => n4127);
   U7292 : BUF_X1 port map( A => n3903, Z => n3904);
   U7293 : BUF_X1 port map( A => n3910, Z => n3903);
   U7294 : BUF_X1 port map( A => n409, Z => n4117);
   U7295 : AND3_X1 port map( A1 => n2261, A2 => n17179, A3 => n2130, ZN => 
                           n1896);
   U7296 : BUF_X1 port map( A => n3907, Z => n3905);
   U7297 : BUF_X1 port map( A => n3909, Z => n3906);
   U7298 : BUF_X1 port map( A => n3903, Z => n3908);
   U7299 : BUF_X1 port map( A => n3903, Z => n3907);
   U7300 : BUF_X1 port map( A => n3903, Z => n3909);
   U7301 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n10, A2 => 
                           DataPath_ALUhw_MUXOUT_n11, ZN => 
                           DataPath_i_ALU_OUT_7_port);
   U7302 : AOI22_X1 port map( A1 => n11515, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_103_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n10);
   U7303 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n16, A2 => 
                           DataPath_ALUhw_MUXOUT_n17, ZN => 
                           DataPath_i_ALU_OUT_4_port);
   U7304 : AOI22_X1 port map( A1 => n11512, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_100_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n16);
   U7305 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n18, A2 => 
                           DataPath_ALUhw_MUXOUT_n19, ZN => 
                           DataPath_i_ALU_OUT_3_port);
   U7306 : AOI22_X1 port map( A1 => n11485, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_99_port, B2 => n8321, ZN
                           => DataPath_ALUhw_MUXOUT_n18);
   U7307 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n24, A2 => 
                           DataPath_ALUhw_MUXOUT_n25, ZN => 
                           DataPath_i_ALU_OUT_2_port);
   U7308 : AOI22_X1 port map( A1 => n11486, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_98_port, B2 => n8321, ZN
                           => DataPath_ALUhw_MUXOUT_n24);
   U7309 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n46, A2 => 
                           DataPath_ALUhw_MUXOUT_n47, ZN => 
                           DataPath_i_ALU_OUT_1_port);
   U7310 : AOI22_X1 port map( A1 => n11487, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_97_port, B2 => n8321, ZN
                           => DataPath_ALUhw_MUXOUT_n46);
   U7311 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n68, A2 => 
                           DataPath_ALUhw_MUXOUT_n69, ZN => 
                           DataPath_i_ALU_OUT_0_port);
   U7312 : AOI22_X1 port map( A1 => n11488, A2 => n2272, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_96_port, B2 => n8321, ZN
                           => DataPath_ALUhw_MUXOUT_n68);
   U7313 : INV_X1 port map( A => DataPath_LDSTR_n70, ZN => n11349);
   U7314 : BUF_X1 port map( A => n7991, Z => n2281);
   U7315 : AND2_X1 port map( A1 => n3890, A2 => n11607, ZN => 
                           DataPath_RF_c_swin_masked_1bit_3_0_port);
   U7316 : AND2_X1 port map( A1 => n372, A2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_14_port, ZN
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_16_port)
                           ;
   U7317 : INV_X1 port map( A => n12924, ZN => n11524);
   U7318 : AOI21_X1 port map( B1 => n11525, B2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_2_24_port, A 
                           => n11528, ZN => n12924);
   U7319 : INV_X1 port map( A => n12921, ZN => n11528);
   U7320 : AOI21_X1 port map( B1 => n11529, B2 => n375, A => n11530, ZN => 
                           n12921);
   U7321 : BUF_X1 port map( A => n7991, Z => n2280);
   U7322 : INV_X1 port map( A => n12889, ZN => n11485);
   U7323 : AOI22_X1 port map( A1 => n4129, A2 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_3_port
                           , B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_3_port
                           , B2 => n4133, ZN => n12889);
   U7324 : BUF_X1 port map( A => n3294, Z => n3284);
   U7325 : BUF_X1 port map( A => n3406, Z => n3396);
   U7326 : BUF_X1 port map( A => n3518, Z => n3508);
   U7327 : BUF_X1 port map( A => n3742, Z => n3732);
   U7328 : INV_X1 port map( A => n12890, ZN => n11486);
   U7329 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_2_port
                           , A2 => n4129, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_2_port
                           , B2 => n4133, ZN => n12890);
   U7330 : INV_X1 port map( A => n12891, ZN => n11487);
   U7331 : AOI22_X1 port map( A1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_1_port
                           , A2 => n4129, B1 => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_1_port
                           , B2 => n4133, ZN => n12891);
   U7332 : INV_X1 port map( A => n12919, ZN => n11520);
   U7333 : AOI21_X1 port map( B1 => n11521, B2 => n372, A => n11522, ZN => 
                           n12919);
   U7334 : INV_X1 port map( A => n12922, ZN => n11531);
   U7335 : AOI21_X1 port map( B1 => n11532, B2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_28_port, A 
                           => n11533, ZN => n12922);
   U7336 : INV_X1 port map( A => n12916, ZN => n11533);
   U7337 : INV_X1 port map( A => n12915, ZN => n11532);
   U7338 : NOR3_X1 port map( A1 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7, A3 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n6);
   U7339 : NOR2_X1 port map( A1 => n11400, A2 => DataPath_i_DONE_FILL_EX, ZN =>
                           n12904);
   U7340 : NOR2_X1 port map( A1 => i_EN2, A2 => n4183, ZN => n14230);
   U7341 : INV_X1 port map( A => n303, ZN => n3265);
   U7342 : INV_X1 port map( A => n303, ZN => n3266);
   U7343 : INV_X1 port map( A => n1932, ZN => n4107);
   U7344 : NOR2_X1 port map( A1 => n14237, A2 => n4183, ZN => n14236);
   U7345 : INV_X1 port map( A => DataPath_LDSTR_n40, ZN => n11576);
   U7346 : INV_X1 port map( A => DataPath_LDSTR_n47, ZN => n11577);
   U7347 : INV_X1 port map( A => DataPath_RF_PUSH_ADDRGEN_n34, ZN => n11446);
   U7348 : BUF_X1 port map( A => n410, Z => n2272);
   U7349 : AND2_X1 port map( A1 => DataPath_i_DONE_FILL_EX, A2 => n11400, ZN =>
                           n12903);
   U7350 : AND2_X1 port map( A1 => DataPath_i_DONE_SPILL_EX, A2 => 
                           DataPath_i_DONE_FILL_EX, ZN => n12906);
   U7351 : BUF_X1 port map( A => n14295, Z => n2497);
   U7352 : BUF_X1 port map( A => n14329, Z => n2503);
   U7353 : BUF_X1 port map( A => n410, Z => n2271);
   U7354 : BUF_X1 port map( A => n4046, Z => n4048);
   U7355 : BUF_X1 port map( A => n4046, Z => n4049);
   U7356 : BUF_X1 port map( A => n4047, Z => n4050);
   U7357 : BUF_X1 port map( A => n14295, Z => n2496);
   U7358 : BUF_X1 port map( A => n14295, Z => n2495);
   U7359 : BUF_X1 port map( A => n14329, Z => n2502);
   U7360 : BUF_X1 port map( A => n14329, Z => n2501);
   U7361 : BUF_X1 port map( A => n14635, Z => n2556);
   U7362 : BUF_X1 port map( A => n14635, Z => n2555);
   U7363 : BUF_X1 port map( A => n14669, Z => n2562);
   U7364 : BUF_X1 port map( A => n14669, Z => n2561);
   U7365 : BUF_X1 port map( A => n14703, Z => n2568);
   U7366 : BUF_X1 port map( A => n14703, Z => n2567);
   U7367 : BUF_X1 port map( A => n14737, Z => n2574);
   U7368 : BUF_X1 port map( A => n14737, Z => n2573);
   U7369 : BUF_X1 port map( A => n14771, Z => n2580);
   U7370 : BUF_X1 port map( A => n14771, Z => n2579);
   U7371 : BUF_X1 port map( A => n14805, Z => n2586);
   U7372 : BUF_X1 port map( A => n14805, Z => n2585);
   U7373 : BUF_X1 port map( A => n14839, Z => n2592);
   U7374 : BUF_X1 port map( A => n14839, Z => n2591);
   U7375 : BUF_X1 port map( A => n14873, Z => n2598);
   U7376 : BUF_X1 port map( A => n14873, Z => n2597);
   U7377 : BUF_X1 port map( A => n15179, Z => n2652);
   U7378 : BUF_X1 port map( A => n15179, Z => n2651);
   U7379 : BUF_X1 port map( A => n15213, Z => n2658);
   U7380 : BUF_X1 port map( A => n15213, Z => n2657);
   U7381 : BUF_X1 port map( A => n15247, Z => n2664);
   U7382 : BUF_X1 port map( A => n15247, Z => n2663);
   U7383 : BUF_X1 port map( A => n15281, Z => n2670);
   U7384 : BUF_X1 port map( A => n15281, Z => n2669);
   U7385 : BUF_X1 port map( A => n15315, Z => n2676);
   U7386 : BUF_X1 port map( A => n15315, Z => n2675);
   U7387 : BUF_X1 port map( A => n15349, Z => n2682);
   U7388 : BUF_X1 port map( A => n15349, Z => n2681);
   U7389 : BUF_X1 port map( A => n15383, Z => n2688);
   U7390 : BUF_X1 port map( A => n15383, Z => n2687);
   U7391 : BUF_X1 port map( A => n15417, Z => n2694);
   U7392 : BUF_X1 port map( A => n15417, Z => n2693);
   U7393 : BUF_X1 port map( A => n15723, Z => n2748);
   U7394 : BUF_X1 port map( A => n15723, Z => n2747);
   U7395 : BUF_X1 port map( A => n15757, Z => n2754);
   U7396 : BUF_X1 port map( A => n15757, Z => n2753);
   U7397 : BUF_X1 port map( A => n15791, Z => n2760);
   U7398 : BUF_X1 port map( A => n15791, Z => n2759);
   U7399 : BUF_X1 port map( A => n15825, Z => n2766);
   U7400 : BUF_X1 port map( A => n15825, Z => n2765);
   U7401 : BUF_X1 port map( A => n15859, Z => n2772);
   U7402 : BUF_X1 port map( A => n15859, Z => n2771);
   U7403 : BUF_X1 port map( A => n15893, Z => n2778);
   U7404 : BUF_X1 port map( A => n15893, Z => n2777);
   U7405 : BUF_X1 port map( A => n15927, Z => n2784);
   U7406 : BUF_X1 port map( A => n15927, Z => n2783);
   U7407 : BUF_X1 port map( A => n15961, Z => n2790);
   U7408 : BUF_X1 port map( A => n15961, Z => n2789);
   U7409 : BUF_X1 port map( A => n16267, Z => n2844);
   U7410 : BUF_X1 port map( A => n16267, Z => n2843);
   U7411 : BUF_X1 port map( A => n16301, Z => n2850);
   U7412 : BUF_X1 port map( A => n16301, Z => n2849);
   U7413 : BUF_X1 port map( A => n16335, Z => n2856);
   U7414 : BUF_X1 port map( A => n16335, Z => n2855);
   U7415 : BUF_X1 port map( A => n16369, Z => n2862);
   U7416 : BUF_X1 port map( A => n16369, Z => n2861);
   U7417 : BUF_X1 port map( A => n16403, Z => n2868);
   U7418 : BUF_X1 port map( A => n16403, Z => n2867);
   U7419 : BUF_X1 port map( A => n16437, Z => n2874);
   U7420 : BUF_X1 port map( A => n16437, Z => n2873);
   U7421 : BUF_X1 port map( A => n16471, Z => n2880);
   U7422 : BUF_X1 port map( A => n16471, Z => n2879);
   U7423 : BUF_X1 port map( A => n16505, Z => n2886);
   U7424 : BUF_X1 port map( A => n16505, Z => n2885);
   U7425 : BUF_X1 port map( A => n16811, Z => n2940);
   U7426 : BUF_X1 port map( A => n16811, Z => n2939);
   U7427 : BUF_X1 port map( A => n16845, Z => n2946);
   U7428 : BUF_X1 port map( A => n16845, Z => n2945);
   U7429 : BUF_X1 port map( A => n16879, Z => n2952);
   U7430 : BUF_X1 port map( A => n16879, Z => n2951);
   U7431 : BUF_X1 port map( A => n16913, Z => n2958);
   U7432 : BUF_X1 port map( A => n16913, Z => n2957);
   U7433 : BUF_X1 port map( A => n16947, Z => n2964);
   U7434 : BUF_X1 port map( A => n16947, Z => n2963);
   U7435 : BUF_X1 port map( A => n16981, Z => n2970);
   U7436 : BUF_X1 port map( A => n16981, Z => n2969);
   U7437 : BUF_X1 port map( A => n17015, Z => n2976);
   U7438 : BUF_X1 port map( A => n17015, Z => n2975);
   U7439 : BUF_X1 port map( A => n17049, Z => n2982);
   U7440 : BUF_X1 port map( A => n17049, Z => n2981);
   U7441 : BUF_X1 port map( A => n3891, Z => n3889);
   U7442 : NOR2_X1 port map( A1 => i_EN2, A2 => n4182, ZN => n14261);
   U7443 : BUF_X1 port map( A => n11590, Z => n2477);
   U7444 : INV_X1 port map( A => n1932, ZN => n4106);
   U7445 : BUF_X1 port map( A => n11590, Z => n2475);
   U7446 : BUF_X1 port map( A => n11590, Z => n2476);
   U7447 : BUF_X1 port map( A => n4052, Z => n4054);
   U7448 : BUF_X1 port map( A => n4058, Z => n4060);
   U7449 : BUF_X1 port map( A => n4064, Z => n4066);
   U7450 : BUF_X1 port map( A => n4070, Z => n4072);
   U7451 : BUF_X1 port map( A => n4076, Z => n4078);
   U7452 : BUF_X1 port map( A => n4082, Z => n4084);
   U7453 : BUF_X1 port map( A => n4052, Z => n4055);
   U7454 : BUF_X1 port map( A => n4058, Z => n4061);
   U7455 : BUF_X1 port map( A => n4064, Z => n4067);
   U7456 : BUF_X1 port map( A => n4070, Z => n4073);
   U7457 : BUF_X1 port map( A => n4076, Z => n4079);
   U7458 : BUF_X1 port map( A => n4082, Z => n4085);
   U7459 : BUF_X1 port map( A => n4053, Z => n4056);
   U7460 : BUF_X1 port map( A => n4059, Z => n4062);
   U7461 : BUF_X1 port map( A => n4065, Z => n4068);
   U7462 : BUF_X1 port map( A => n4071, Z => n4074);
   U7463 : BUF_X1 port map( A => n4077, Z => n4080);
   U7464 : BUF_X1 port map( A => n4083, Z => n4086);
   U7465 : BUF_X1 port map( A => n3914, Z => n3916);
   U7466 : BUF_X1 port map( A => n3920, Z => n3922);
   U7467 : BUF_X1 port map( A => n3926, Z => n3928);
   U7468 : BUF_X1 port map( A => n3932, Z => n3934);
   U7469 : BUF_X1 port map( A => n3938, Z => n3940);
   U7470 : BUF_X1 port map( A => n3944, Z => n3946);
   U7471 : BUF_X1 port map( A => n3950, Z => n3952);
   U7472 : BUF_X1 port map( A => n3956, Z => n3958);
   U7473 : BUF_X1 port map( A => n3962, Z => n3964);
   U7474 : BUF_X1 port map( A => n3968, Z => n3970);
   U7475 : BUF_X1 port map( A => n3974, Z => n3976);
   U7476 : BUF_X1 port map( A => n3980, Z => n3982);
   U7477 : BUF_X1 port map( A => n3986, Z => n3988);
   U7478 : BUF_X1 port map( A => n3992, Z => n3994);
   U7479 : BUF_X1 port map( A => n3998, Z => n4000);
   U7480 : BUF_X1 port map( A => n4004, Z => n4006);
   U7481 : BUF_X1 port map( A => n4010, Z => n4012);
   U7482 : BUF_X1 port map( A => n4016, Z => n4018);
   U7483 : BUF_X1 port map( A => n4022, Z => n4024);
   U7484 : BUF_X1 port map( A => n4028, Z => n4030);
   U7485 : BUF_X1 port map( A => n4034, Z => n4036);
   U7486 : BUF_X1 port map( A => n4040, Z => n4042);
   U7487 : BUF_X1 port map( A => n4088, Z => n4090);
   U7488 : BUF_X1 port map( A => n4094, Z => n4096);
   U7489 : BUF_X1 port map( A => n4100, Z => n4102);
   U7490 : BUF_X1 port map( A => n3914, Z => n3917);
   U7491 : BUF_X1 port map( A => n3920, Z => n3923);
   U7492 : BUF_X1 port map( A => n3926, Z => n3929);
   U7493 : BUF_X1 port map( A => n3932, Z => n3935);
   U7494 : BUF_X1 port map( A => n3938, Z => n3941);
   U7495 : BUF_X1 port map( A => n3944, Z => n3947);
   U7496 : BUF_X1 port map( A => n3950, Z => n3953);
   U7497 : BUF_X1 port map( A => n3956, Z => n3959);
   U7498 : BUF_X1 port map( A => n3962, Z => n3965);
   U7499 : BUF_X1 port map( A => n3968, Z => n3971);
   U7500 : BUF_X1 port map( A => n3974, Z => n3977);
   U7501 : BUF_X1 port map( A => n3980, Z => n3983);
   U7502 : BUF_X1 port map( A => n3986, Z => n3989);
   U7503 : BUF_X1 port map( A => n3992, Z => n3995);
   U7504 : BUF_X1 port map( A => n3998, Z => n4001);
   U7505 : BUF_X1 port map( A => n4004, Z => n4007);
   U7506 : BUF_X1 port map( A => n4010, Z => n4013);
   U7507 : BUF_X1 port map( A => n4016, Z => n4019);
   U7508 : BUF_X1 port map( A => n4022, Z => n4025);
   U7509 : BUF_X1 port map( A => n4028, Z => n4031);
   U7510 : BUF_X1 port map( A => n4034, Z => n4037);
   U7511 : BUF_X1 port map( A => n4040, Z => n4043);
   U7512 : BUF_X1 port map( A => n4088, Z => n4091);
   U7513 : BUF_X1 port map( A => n4094, Z => n4097);
   U7514 : BUF_X1 port map( A => n4100, Z => n4103);
   U7515 : BUF_X1 port map( A => n3915, Z => n3918);
   U7516 : BUF_X1 port map( A => n3921, Z => n3924);
   U7517 : BUF_X1 port map( A => n3927, Z => n3930);
   U7518 : BUF_X1 port map( A => n3933, Z => n3936);
   U7519 : BUF_X1 port map( A => n3939, Z => n3942);
   U7520 : BUF_X1 port map( A => n3945, Z => n3948);
   U7521 : BUF_X1 port map( A => n3951, Z => n3954);
   U7522 : BUF_X1 port map( A => n3957, Z => n3960);
   U7523 : BUF_X1 port map( A => n3963, Z => n3966);
   U7524 : BUF_X1 port map( A => n3969, Z => n3972);
   U7525 : BUF_X1 port map( A => n3975, Z => n3978);
   U7526 : BUF_X1 port map( A => n3981, Z => n3984);
   U7527 : BUF_X1 port map( A => n3987, Z => n3990);
   U7528 : BUF_X1 port map( A => n3993, Z => n3996);
   U7529 : BUF_X1 port map( A => n3999, Z => n4002);
   U7530 : BUF_X1 port map( A => n4005, Z => n4008);
   U7531 : BUF_X1 port map( A => n4011, Z => n4014);
   U7532 : BUF_X1 port map( A => n4017, Z => n4020);
   U7533 : BUF_X1 port map( A => n4023, Z => n4026);
   U7534 : BUF_X1 port map( A => n4029, Z => n4032);
   U7535 : BUF_X1 port map( A => n4035, Z => n4038);
   U7536 : BUF_X1 port map( A => n4041, Z => n4044);
   U7537 : BUF_X1 port map( A => n4089, Z => n4092);
   U7538 : BUF_X1 port map( A => n4095, Z => n4098);
   U7539 : BUF_X1 port map( A => n4101, Z => n4104);
   U7540 : AOI22_X1 port map( A1 => n3269, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n6, B1 => n3270, 
                           B2 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n2);
   U7541 : NOR2_X1 port map( A1 => DataPath_LDSTR_n71, A2 => n4118, ZN => 
                           DataPath_LDSTR_n64);
   U7542 : BUF_X1 port map( A => n2332, Z => n2336);
   U7543 : BUF_X1 port map( A => n2344, Z => n2348);
   U7544 : BUF_X1 port map( A => n2350, Z => n2354);
   U7545 : BUF_X1 port map( A => n2356, Z => n2360);
   U7546 : BUF_X1 port map( A => n2362, Z => n2366);
   U7547 : BUF_X1 port map( A => n2368, Z => n2372);
   U7548 : BUF_X1 port map( A => n2374, Z => n2378);
   U7549 : BUF_X1 port map( A => n2380, Z => n2384);
   U7550 : BUF_X1 port map( A => n2386, Z => n2390);
   U7551 : BUF_X1 port map( A => n2392, Z => n2396);
   U7552 : BUF_X1 port map( A => n2398, Z => n2402);
   U7553 : BUF_X1 port map( A => n2410, Z => n2414);
   U7554 : BUF_X1 port map( A => n2416, Z => n2420);
   U7555 : BUF_X1 port map( A => n2422, Z => n2426);
   U7556 : BUF_X1 port map( A => n2428, Z => n2432);
   U7557 : BUF_X1 port map( A => n2434, Z => n2438);
   U7558 : BUF_X1 port map( A => n2440, Z => n2444);
   U7559 : BUF_X1 port map( A => n2446, Z => n2450);
   U7560 : BUF_X1 port map( A => n2452, Z => n2456);
   U7561 : BUF_X1 port map( A => n2458, Z => n2462);
   U7562 : BUF_X1 port map( A => n2464, Z => n2468);
   U7563 : BUF_X1 port map( A => n2338, Z => n2342);
   U7564 : BUF_X1 port map( A => n2404, Z => n2408);
   U7565 : BUF_X1 port map( A => n2470, Z => n2474);
   U7566 : INV_X1 port map( A => DataPath_i_DONE_SPILL_EX, ZN => n11400);
   U7567 : BUF_X1 port map( A => n3279, Z => n3278);
   U7568 : BUF_X1 port map( A => n3280, Z => n3277);
   U7569 : NAND2_X1 port map( A1 => n12955, A2 => n4260, ZN => n12952);
   U7570 : NAND2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n30, A2 => n4260, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_n27);
   U7571 : INV_X1 port map( A => DataPath_i_DONE_FILL_EX, ZN => n11382);
   U7572 : BUF_X1 port map( A => n2257, Z => n2252);
   U7573 : BUF_X1 port map( A => n4047, Z => n4051);
   U7574 : BUF_X1 port map( A => n4128, Z => n4119);
   U7575 : BUF_X1 port map( A => n4128, Z => n4125);
   U7576 : BUF_X1 port map( A => n4128, Z => n4120);
   U7577 : BUF_X1 port map( A => n4124, Z => n4122);
   U7578 : BUF_X1 port map( A => n4128, Z => n4126);
   U7579 : BUF_X1 port map( A => n4126, Z => n4121);
   U7580 : BUF_X1 port map( A => n4128, Z => n4124);
   U7581 : BUF_X1 port map( A => n4128, Z => n4123);
   U7582 : BUF_X1 port map( A => n409, Z => n4112);
   U7583 : BUF_X1 port map( A => n409, Z => n4113);
   U7584 : BUF_X1 port map( A => n4109, Z => n4115);
   U7585 : BUF_X1 port map( A => n409, Z => n4109);
   U7586 : BUF_X1 port map( A => n409, Z => n4110);
   U7587 : BUF_X1 port map( A => n409, Z => n4111);
   U7588 : BUF_X1 port map( A => n409, Z => n4114);
   U7589 : BUF_X1 port map( A => n4110, Z => n4116);
   U7590 : BUF_X1 port map( A => n3283, Z => n3271);
   U7591 : BUF_X1 port map( A => n3283, Z => n3272);
   U7592 : BUF_X1 port map( A => n3282, Z => n3273);
   U7593 : BUF_X1 port map( A => n3282, Z => n3274);
   U7594 : BUF_X1 port map( A => n2257, Z => n2253);
   U7595 : BUF_X1 port map( A => n2256, Z => n2254);
   U7596 : BUF_X1 port map( A => n4053, Z => n4057);
   U7597 : BUF_X1 port map( A => n4059, Z => n4063);
   U7598 : BUF_X1 port map( A => n4065, Z => n4069);
   U7599 : BUF_X1 port map( A => n4071, Z => n4075);
   U7600 : BUF_X1 port map( A => n4077, Z => n4081);
   U7601 : BUF_X1 port map( A => n4083, Z => n4087);
   U7602 : BUF_X1 port map( A => n3281, Z => n3275);
   U7603 : BUF_X1 port map( A => n3281, Z => n3276);
   U7604 : BUF_X1 port map( A => n3915, Z => n3919);
   U7605 : BUF_X1 port map( A => n3921, Z => n3925);
   U7606 : BUF_X1 port map( A => n3927, Z => n3931);
   U7607 : BUF_X1 port map( A => n3933, Z => n3937);
   U7608 : BUF_X1 port map( A => n3939, Z => n3943);
   U7609 : BUF_X1 port map( A => n3945, Z => n3949);
   U7610 : BUF_X1 port map( A => n3951, Z => n3955);
   U7611 : BUF_X1 port map( A => n3957, Z => n3961);
   U7612 : BUF_X1 port map( A => n3963, Z => n3967);
   U7613 : BUF_X1 port map( A => n3969, Z => n3973);
   U7614 : BUF_X1 port map( A => n3975, Z => n3979);
   U7615 : BUF_X1 port map( A => n3981, Z => n3985);
   U7616 : BUF_X1 port map( A => n3987, Z => n3991);
   U7617 : BUF_X1 port map( A => n3993, Z => n3997);
   U7618 : BUF_X1 port map( A => n3999, Z => n4003);
   U7619 : BUF_X1 port map( A => n4005, Z => n4009);
   U7620 : BUF_X1 port map( A => n4011, Z => n4015);
   U7621 : BUF_X1 port map( A => n4017, Z => n4021);
   U7622 : BUF_X1 port map( A => n4023, Z => n4027);
   U7623 : BUF_X1 port map( A => n4029, Z => n4033);
   U7624 : BUF_X1 port map( A => n4035, Z => n4039);
   U7625 : BUF_X1 port map( A => n4041, Z => n4045);
   U7626 : BUF_X1 port map( A => n4089, Z => n4093);
   U7627 : BUF_X1 port map( A => n4095, Z => n4099);
   U7628 : BUF_X1 port map( A => n4101, Z => n4105);
   U7629 : BUF_X1 port map( A => CU_I_n104, Z => n4128);
   U7630 : BUF_X1 port map( A => n2256, Z => n2255);
   U7631 : BUF_X1 port map( A => n3292, Z => n3290);
   U7632 : BUF_X1 port map( A => n3293, Z => n3287);
   U7633 : BUF_X1 port map( A => n3293, Z => n3288);
   U7634 : BUF_X1 port map( A => n3293, Z => n3286);
   U7635 : BUF_X1 port map( A => n3292, Z => n3289);
   U7636 : BUF_X1 port map( A => n3404, Z => n3402);
   U7637 : BUF_X1 port map( A => n3405, Z => n3398);
   U7638 : BUF_X1 port map( A => n3405, Z => n3399);
   U7639 : BUF_X1 port map( A => n3405, Z => n3400);
   U7640 : BUF_X1 port map( A => n3404, Z => n3401);
   U7641 : BUF_X1 port map( A => n3516, Z => n3514);
   U7642 : BUF_X1 port map( A => n3517, Z => n3510);
   U7643 : BUF_X1 port map( A => n3517, Z => n3511);
   U7644 : BUF_X1 port map( A => n3517, Z => n3512);
   U7645 : BUF_X1 port map( A => n3516, Z => n3513);
   U7646 : BUF_X1 port map( A => n3740, Z => n3738);
   U7647 : BUF_X1 port map( A => n3741, Z => n3734);
   U7648 : BUF_X1 port map( A => n3741, Z => n3735);
   U7649 : BUF_X1 port map( A => n3741, Z => n3736);
   U7650 : BUF_X1 port map( A => n3740, Z => n3737);
   U7651 : BUF_X1 port map( A => n3294, Z => n3285);
   U7652 : BUF_X1 port map( A => n3406, Z => n3397);
   U7653 : BUF_X1 port map( A => n3518, Z => n3509);
   U7654 : BUF_X1 port map( A => n3742, Z => n3733);
   U7655 : BUF_X1 port map( A => n3292, Z => n3291);
   U7656 : BUF_X1 port map( A => n3404, Z => n3403);
   U7657 : BUF_X1 port map( A => n3516, Z => n3515);
   U7658 : BUF_X1 port map( A => n3740, Z => n3739);
   U7659 : INV_X1 port map( A => n4144, ZN => n4155);
   U7660 : INV_X1 port map( A => n4145, ZN => n4156);
   U7661 : BUF_X1 port map( A => n3896, Z => n3857);
   U7662 : BUF_X1 port map( A => n3893, Z => n3876);
   U7663 : BUF_X1 port map( A => n3892, Z => n3884);
   U7664 : BUF_X1 port map( A => n3892, Z => n3881);
   U7665 : BUF_X1 port map( A => n3894, Z => n3869);
   U7666 : BUF_X1 port map( A => n3894, Z => n3872);
   U7667 : BUF_X1 port map( A => n3896, Z => n3858);
   U7668 : BUF_X1 port map( A => n3895, Z => n3864);
   U7669 : BUF_X1 port map( A => n3895, Z => n3861);
   U7670 : BUF_X1 port map( A => n3894, Z => n3867);
   U7671 : BUF_X1 port map( A => n3892, Z => n3879);
   U7672 : BUF_X1 port map( A => n3894, Z => n3868);
   U7673 : BUF_X1 port map( A => n3893, Z => n3877);
   U7674 : BUF_X1 port map( A => n3892, Z => n3882);
   U7675 : BUF_X1 port map( A => n3897, Z => n3849);
   U7676 : BUF_X1 port map( A => n3894, Z => n3870);
   U7677 : BUF_X1 port map( A => n3897, Z => n3851);
   U7678 : BUF_X1 port map( A => n3897, Z => n3852);
   U7679 : BUF_X1 port map( A => n3896, Z => n3859);
   U7680 : BUF_X1 port map( A => n3895, Z => n3865);
   U7681 : BUF_X1 port map( A => n3897, Z => n3854);
   U7682 : BUF_X1 port map( A => n3895, Z => n3862);
   U7683 : BUF_X1 port map( A => n3896, Z => n3855);
   U7684 : BUF_X1 port map( A => n3896, Z => n3860);
   U7685 : BUF_X1 port map( A => n3893, Z => n3875);
   U7686 : BUF_X1 port map( A => n3895, Z => n3866);
   U7687 : BUF_X1 port map( A => n3893, Z => n3878);
   U7688 : BUF_X1 port map( A => n3895, Z => n3863);
   U7689 : BUF_X1 port map( A => n3897, Z => n3850);
   U7690 : BUF_X1 port map( A => n3893, Z => n3873);
   U7691 : BUF_X1 port map( A => n3892, Z => n3880);
   U7692 : BUF_X1 port map( A => n3897, Z => n3853);
   U7693 : BUF_X1 port map( A => n3896, Z => n3856);
   U7694 : BUF_X1 port map( A => n3892, Z => n3883);
   U7695 : BUF_X1 port map( A => n3894, Z => n3871);
   U7696 : BUF_X1 port map( A => n3893, Z => n3874);
   U7697 : BUF_X1 port map( A => n3891, Z => n3885);
   U7698 : BUF_X1 port map( A => n3891, Z => n3888);
   U7699 : BUF_X1 port map( A => n3891, Z => n3887);
   U7700 : BUF_X1 port map( A => n3891, Z => n3886);
   U7701 : BUF_X1 port map( A => n3898, Z => n3848);
   U7702 : BUF_X1 port map( A => n3898, Z => n3847);
   U7703 : NOR2_X1 port map( A1 => n11434, A2 => 
                           DataPath_RF_spill_address_1_port, ZN => 
                           DataPath_RF_RDPORT_SPILL_n338);
   U7704 : NOR2_X1 port map( A1 => DataPath_RF_spill_address_1_port, A2 => 
                           DataPath_RF_spill_address_0_port, ZN => 
                           DataPath_RF_RDPORT_SPILL_n340);
   U7705 : NOR2_X1 port map( A1 => DataPath_RF_spill_address_3_port, A2 => 
                           DataPath_RF_spill_address_2_port, ZN => 
                           DataPath_RF_RDPORT_SPILL_n346);
   U7706 : NOR2_X1 port map( A1 => n11433, A2 => 
                           DataPath_RF_spill_address_0_port, ZN => 
                           DataPath_RF_RDPORT_SPILL_n336);
   U7707 : NOR2_X1 port map( A1 => n11432, A2 => 
                           DataPath_RF_spill_address_3_port, ZN => 
                           DataPath_RF_RDPORT_SPILL_n347);
   U7708 : BUF_X1 port map( A => n3203, Z => n3253);
   U7709 : BUF_X1 port map( A => n3203, Z => n3254);
   U7710 : BUF_X1 port map( A => n3202, Z => n3252);
   U7711 : BUF_X1 port map( A => n3201, Z => n3249);
   U7712 : BUF_X1 port map( A => n3202, Z => n3251);
   U7713 : BUF_X1 port map( A => n3202, Z => n3250);
   U7714 : BUF_X1 port map( A => n3201, Z => n3248);
   U7715 : BUF_X1 port map( A => n3102, Z => n3091);
   U7716 : BUF_X1 port map( A => n3047, Z => n3036);
   U7717 : BUF_X1 port map( A => n3148, Z => n3198);
   U7718 : BUF_X1 port map( A => n3102, Z => n3092);
   U7719 : BUF_X1 port map( A => n3148, Z => n3199);
   U7720 : BUF_X1 port map( A => n3047, Z => n3037);
   U7721 : BUF_X1 port map( A => n3102, Z => n3093);
   U7722 : BUF_X1 port map( A => n3047, Z => n3038);
   U7723 : BUF_X1 port map( A => n3100, Z => n3097);
   U7724 : BUF_X1 port map( A => n3045, Z => n3042);
   U7725 : BUF_X1 port map( A => n3101, Z => n3094);
   U7726 : BUF_X1 port map( A => n3147, Z => n3197);
   U7727 : BUF_X1 port map( A => n3046, Z => n3039);
   U7728 : BUF_X1 port map( A => n3146, Z => n3194);
   U7729 : BUF_X1 port map( A => n3101, Z => n3095);
   U7730 : BUF_X1 port map( A => n3147, Z => n3196);
   U7731 : BUF_X1 port map( A => n3046, Z => n3040);
   U7732 : BUF_X1 port map( A => n3101, Z => n3096);
   U7733 : BUF_X1 port map( A => n3147, Z => n3195);
   U7734 : BUF_X1 port map( A => n3046, Z => n3041);
   U7735 : BUF_X1 port map( A => n3146, Z => n3193);
   U7736 : BUF_X1 port map( A => n3100, Z => n3098);
   U7737 : BUF_X1 port map( A => n3045, Z => n3043);
   U7738 : BUF_X1 port map( A => n3201, Z => n3247);
   U7739 : BUF_X1 port map( A => n3146, Z => n3192);
   U7740 : BUF_X1 port map( A => n3203, Z => n3255);
   U7741 : BUF_X1 port map( A => n3148, Z => n3200);
   U7742 : BUF_X1 port map( A => n4245, Z => n4157);
   U7743 : BUF_X1 port map( A => n4246, Z => n4245);
   U7744 : AND2_X1 port map( A1 => DataPath_RF_spill_address_3_port, A2 => 
                           DataPath_RF_spill_address_2_port, ZN => 
                           DataPath_RF_RDPORT_SPILL_n339);
   U7745 : AND2_X1 port map( A1 => DataPath_RF_spill_address_3_port, A2 => 
                           n11432, ZN => DataPath_RF_RDPORT_SPILL_n337);
   U7746 : INV_X1 port map( A => DataPath_RF_spill_address_1_port, ZN => n11433
                           );
   U7747 : BUF_X1 port map( A => n3100, Z => n3099);
   U7748 : BUF_X1 port map( A => n3045, Z => n3044);
   U7749 : INV_X1 port map( A => DataPath_RF_spill_address_0_port, ZN => n11434
                           );
   U7750 : INV_X1 port map( A => DataPath_RF_spill_address_2_port, ZN => n11432
                           );
   U7751 : BUF_X1 port map( A => n4249, Z => n4236);
   U7752 : BUF_X1 port map( A => n4248, Z => n4237);
   U7753 : BUF_X1 port map( A => n4248, Z => n4238);
   U7754 : BUF_X1 port map( A => n4248, Z => n4239);
   U7755 : BUF_X1 port map( A => n4247, Z => n4241);
   U7756 : BUF_X1 port map( A => n4247, Z => n4242);
   U7757 : BUF_X1 port map( A => n4246, Z => n4243);
   U7758 : BUF_X1 port map( A => n4246, Z => n4244);
   U7759 : BUF_X1 port map( A => n4247, Z => n4240);
   U7760 : BUF_X1 port map( A => n4251, Z => n4229);
   U7761 : BUF_X1 port map( A => n4251, Z => n4230);
   U7762 : BUF_X1 port map( A => n4250, Z => n4231);
   U7763 : BUF_X1 port map( A => n4250, Z => n4232);
   U7764 : BUF_X1 port map( A => n4250, Z => n4233);
   U7765 : BUF_X1 port map( A => n4249, Z => n4234);
   U7766 : BUF_X1 port map( A => n4249, Z => n4235);
   U7767 : BUF_X1 port map( A => n4253, Z => n4223);
   U7768 : BUF_X1 port map( A => n4253, Z => n4224);
   U7769 : BUF_X1 port map( A => n4252, Z => n4225);
   U7770 : BUF_X1 port map( A => n4252, Z => n4226);
   U7771 : BUF_X1 port map( A => n4252, Z => n4227);
   U7772 : BUF_X1 port map( A => n4253, Z => n4222);
   U7773 : BUF_X1 port map( A => n4251, Z => n4228);
   U7774 : OR2_X1 port map( A1 => DRAMRF_READNOTWRITE_port, A2 => i_RF_MEM_WM, 
                           ZN => DRAMRF_ISSUE);
   U7775 : NOR2_X1 port map( A1 => DataPath_i_DONE_SPILL_EX, A2 => n3900, ZN =>
                           i_RF_MEM_WM);
   U7776 : XNOR2_X1 port map( A => n5804, B => n1897, ZN => n6773);
   U7777 : XNOR2_X1 port map( A => n6754, B => n6755, ZN => n1897);
   U7778 : XNOR2_X1 port map( A => n8143, B => n2245, ZN => n1898);
   U7779 : OAI21_X1 port map( B1 => n5578, B2 => n2244, A => n5577, ZN => n5856
                           );
   U7780 : XNOR2_X1 port map( A => n6890, B => n8166, ZN => n1899);
   U7781 : BUF_X2 port map( A => n7286, Z => n2179);
   U7782 : BUF_X2 port map( A => n7275, Z => n2175);
   U7783 : CLKBUF_X1 port map( A => n7275, Z => n2176);
   U7784 : BUF_X2 port map( A => n7273, Z => n2177);
   U7785 : CLKBUF_X1 port map( A => n7273, Z => n2178);
   U7786 : XNOR2_X1 port map( A => n7375, B => n7374, ZN => n1901);
   U7787 : XNOR2_X1 port map( A => n7363, B => n7362, ZN => n1902);
   U7788 : XNOR2_X1 port map( A => n7348, B => n7347, ZN => n1903);
   U7789 : XNOR2_X1 port map( A => n7336, B => n7335, ZN => n1904);
   U7790 : OAI21_X1 port map( B1 => n7501, B2 => n7507, A => n7502, ZN => n7506
                           );
   U7791 : AND2_X1 port map( A1 => n4444, A2 => n4443, ZN => n1906);
   U7792 : XNOR2_X1 port map( A => n6563, B => n6562, ZN => n6564);
   U7793 : OR2_X1 port map( A1 => n6160, A2 => n6967, ZN => n6155);
   U7794 : NOR3_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n32, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_n35, A3 => n4155, ZN => 
                           DataPath_i_DONE_SPILL_EX);
   U7795 : INV_X1 port map( A => n12957, ZN => n11607);
   U7796 : BUF_X1 port map( A => n4140, Z => n4134);
   U7797 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n597, ZN => n11539);
   U7798 : INV_X1 port map( A => DataPath_RF_PUSH_ADDRGEN_n32, ZN => n11597);
   U7799 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n639, A2 => n4132
                           , ZN => DataPath_ALUhw_SHIFTER_HW_n548);
   U7800 : NOR2_X1 port map( A1 => n4214, A2 => DataPath_WRF_CUhw_n114, ZN => 
                           DataPath_WRF_CUhw_N177_port);
   U7801 : NOR2_X1 port map( A1 => n4214, A2 => DataPath_WRF_CUhw_n115, ZN => 
                           DataPath_WRF_CUhw_N176_port);
   U7802 : NOR2_X1 port map( A1 => n4212, A2 => DataPath_WRF_CUhw_n120, ZN => 
                           DataPath_WRF_CUhw_N171_port);
   U7803 : NOR2_X1 port map( A1 => n4213, A2 => DataPath_WRF_CUhw_n119, ZN => 
                           DataPath_WRF_CUhw_N172_port);
   U7804 : NOR2_X1 port map( A1 => n4213, A2 => DataPath_WRF_CUhw_n116, ZN => 
                           DataPath_WRF_CUhw_N175_port);
   U7805 : NOR2_X1 port map( A1 => n4213, A2 => DataPath_WRF_CUhw_n117, ZN => 
                           DataPath_WRF_CUhw_N174_port);
   U7806 : NOR2_X1 port map( A1 => n4213, A2 => DataPath_WRF_CUhw_n118, ZN => 
                           DataPath_WRF_CUhw_N173_port);
   U7807 : NOR2_X1 port map( A1 => n4210, A2 => DataPath_WRF_CUhw_n129, ZN => 
                           DataPath_WRF_CUhw_N162_port);
   U7808 : NOR2_X1 port map( A1 => n4210, A2 => DataPath_WRF_CUhw_n128, ZN => 
                           DataPath_WRF_CUhw_N163_port);
   U7809 : NOR2_X1 port map( A1 => n4211, A2 => DataPath_WRF_CUhw_n127, ZN => 
                           DataPath_WRF_CUhw_N164_port);
   U7810 : NOR2_X1 port map( A1 => n4211, A2 => DataPath_WRF_CUhw_n126, ZN => 
                           DataPath_WRF_CUhw_N165_port);
   U7811 : NOR2_X1 port map( A1 => n4211, A2 => DataPath_WRF_CUhw_n125, ZN => 
                           DataPath_WRF_CUhw_N166_port);
   U7812 : NOR2_X1 port map( A1 => n4211, A2 => DataPath_WRF_CUhw_n124, ZN => 
                           DataPath_WRF_CUhw_N167_port);
   U7813 : NOR2_X1 port map( A1 => n4210, A2 => DataPath_WRF_CUhw_n123, ZN => 
                           DataPath_WRF_CUhw_N168_port);
   U7814 : NOR2_X1 port map( A1 => n4212, A2 => DataPath_WRF_CUhw_n122, ZN => 
                           DataPath_WRF_CUhw_N169_port);
   U7815 : NOR2_X1 port map( A1 => n4212, A2 => DataPath_WRF_CUhw_n121, ZN => 
                           DataPath_WRF_CUhw_N170_port);
   U7816 : INV_X1 port map( A => n3899, ZN => n3910);
   U7817 : OAI21_X2 port map( B1 => n12960, B2 => n12957, A => n12951, ZN => 
                           n12977);
   U7818 : OAI21_X1 port map( B1 => DataPath_LDSTR_n84, B2 => 
                           DataPath_LDSTR_n78, A => n11580, ZN => 
                           DataPath_LDSTR_n66);
   U7819 : INV_X1 port map( A => DataPath_LDSTR_n80, ZN => n11578);
   U7820 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_8_port, A2 => n4179, ZN 
                           => n14363);
   U7821 : OAI222_X1 port map( A1 => n3273, A2 => n1925, B1 => n3295, B2 => 
                           n11398, C1 => n2478, C2 => n1909, ZN => 
                           DataPath_RF_en_regi_8_port);
   U7822 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_11_port, A2 => n4178, ZN
                           => n14465);
   U7823 : OAI222_X1 port map( A1 => n2478, A2 => n1928, B1 => n3303, B2 => 
                           n11395, C1 => n3273, C2 => n1921, ZN => 
                           DataPath_RF_en_regi_11_port);
   U7824 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_12_port, A2 => n4177, ZN
                           => n14499);
   U7825 : OAI222_X1 port map( A1 => n2478, A2 => n1929, B1 => n3304, B2 => 
                           n11394, C1 => n3271, C2 => n1922, ZN => 
                           DataPath_RF_en_regi_12_port);
   U7826 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_13_port, A2 => n4177, ZN
                           => n14533);
   U7827 : OAI222_X1 port map( A1 => n2479, A2 => n1930, B1 => n3295, B2 => 
                           n11393, C1 => n3272, C2 => n1923, ZN => 
                           DataPath_RF_en_regi_13_port);
   U7828 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_14_port, A2 => n4176, ZN
                           => n14567);
   U7829 : OAI222_X1 port map( A1 => n2478, A2 => n1931, B1 => n3305, B2 => 
                           n11392, C1 => n3272, C2 => n1924, ZN => 
                           DataPath_RF_en_regi_14_port);
   U7830 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_15_port, A2 => n4176, ZN
                           => n14601);
   U7831 : OAI222_X1 port map( A1 => n2478, A2 => n1926, B1 => n3303, B2 => 
                           n11391, C1 => n3271, C2 => n1910, ZN => 
                           DataPath_RF_en_regi_15_port);
   U7832 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_24_port, A2 => n4171, ZN
                           => n14907);
   U7833 : OAI222_X1 port map( A1 => n2479, A2 => n1925, B1 => n11398, B2 => 
                           n3415, C1 => n1909, C2 => n2480, ZN => 
                           DataPath_RF_en_regi_24_port);
   U7834 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_25_port, A2 => n4171, ZN
                           => n14941);
   U7835 : OAI222_X1 port map( A1 => n1919, A2 => n2479, B1 => n11397, B2 => 
                           n3417, C1 => n1908, C2 => n2480, ZN => 
                           DataPath_RF_en_regi_25_port);
   U7836 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_27_port, A2 => n4170, ZN
                           => n15009);
   U7837 : OAI222_X1 port map( A1 => n1928, A2 => n2481, B1 => n11395, B2 => 
                           n3408, C1 => n2478, C2 => n1921, ZN => 
                           DataPath_RF_en_regi_27_port);
   U7838 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_28_port, A2 => n4169, ZN
                           => n15043);
   U7839 : OAI222_X1 port map( A1 => n1929, A2 => n2481, B1 => n11394, B2 => 
                           n3407, C1 => n2478, C2 => n1922, ZN => 
                           DataPath_RF_en_regi_28_port);
   U7840 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_29_port, A2 => n4169, ZN
                           => n15077);
   U7841 : OAI222_X1 port map( A1 => n1930, A2 => n2481, B1 => n11393, B2 => 
                           n3417, C1 => n2478, C2 => n1923, ZN => 
                           DataPath_RF_en_regi_29_port);
   U7842 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_30_port, A2 => n4168, ZN
                           => n15111);
   U7843 : OAI222_X1 port map( A1 => n1931, A2 => n2481, B1 => n11392, B2 => 
                           n3415, C1 => n2478, C2 => n1924, ZN => 
                           DataPath_RF_en_regi_30_port);
   U7844 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_31_port, A2 => n4168, ZN
                           => n15145);
   U7845 : OAI222_X1 port map( A1 => n1926, A2 => n2481, B1 => n11391, B2 => 
                           n3416, C1 => n2478, C2 => n1910, ZN => 
                           DataPath_RF_en_regi_31_port);
   U7846 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_40_port, A2 => n4163, ZN
                           => n15451);
   U7847 : OAI222_X1 port map( A1 => n1925, A2 => n2481, B1 => n11398, B2 => 
                           n3529, C1 => n1909, C2 => n2482, ZN => 
                           DataPath_RF_en_regi_40_port);
   U7848 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_41_port, A2 => n4163, ZN
                           => n15485);
   U7849 : OAI222_X1 port map( A1 => n1919, A2 => n2481, B1 => n11397, B2 => 
                           n3527, C1 => n1908, C2 => n2482, ZN => 
                           DataPath_RF_en_regi_41_port);
   U7850 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_42_port, A2 => n4162, ZN
                           => n15519);
   U7851 : OAI222_X1 port map( A1 => n1927, A2 => n2483, B1 => n11396, B2 => 
                           n3520, C1 => n1920, C2 => n2481, ZN => 
                           DataPath_RF_en_regi_42_port);
   U7852 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_44_port, A2 => n4161, ZN
                           => n15587);
   U7853 : OAI222_X1 port map( A1 => n1929, A2 => n2483, B1 => n11394, B2 => 
                           n3519, C1 => n1922, C2 => n2480, ZN => 
                           DataPath_RF_en_regi_44_port);
   U7854 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_45_port, A2 => n4161, ZN
                           => n15621);
   U7855 : OAI222_X1 port map( A1 => n1930, A2 => n2483, B1 => n11393, B2 => 
                           n3529, C1 => n1923, C2 => n2481, ZN => 
                           DataPath_RF_en_regi_45_port);
   U7856 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_46_port, A2 => n4160, ZN
                           => n15655);
   U7857 : OAI222_X1 port map( A1 => n1931, A2 => n2483, B1 => n11392, B2 => 
                           n3527, C1 => n1924, C2 => n2481, ZN => 
                           DataPath_RF_en_regi_46_port);
   U7858 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_10_port, A2 => n4178, ZN
                           => n14431);
   U7859 : OAI222_X1 port map( A1 => n2478, A2 => n1927, B1 => n3295, B2 => 
                           n11396, C1 => n3271, C2 => n1920, ZN => 
                           DataPath_RF_en_regi_10_port);
   U7860 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_26_port, A2 => n4170, ZN
                           => n14975);
   U7861 : OAI222_X1 port map( A1 => n1927, A2 => n2481, B1 => n11396, B2 => 
                           n3415, C1 => n2478, C2 => n1920, ZN => 
                           DataPath_RF_en_regi_26_port);
   U7862 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_43_port, A2 => n4162, ZN
                           => n15553);
   U7863 : OAI222_X1 port map( A1 => n1928, A2 => n2483, B1 => n11395, B2 => 
                           n3528, C1 => n1921, C2 => n2481, ZN => 
                           DataPath_RF_en_regi_43_port);
   U7864 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_47_port, A2 => n4160, ZN
                           => n15689);
   U7865 : OAI222_X1 port map( A1 => n1926, A2 => n2483, B1 => n11391, B2 => 
                           n3527, C1 => n1910, C2 => n2480, ZN => 
                           DataPath_RF_en_regi_47_port);
   U7866 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_56_port, A2 => n4200, ZN
                           => n15995);
   U7867 : OAI222_X1 port map( A1 => n1925, A2 => n2483, B1 => n11398, B2 => 
                           n3631, C1 => n1909, C2 => n2485, ZN => 
                           DataPath_RF_en_regi_56_port);
   U7868 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_57_port, A2 => n4199, ZN
                           => n16029);
   U7869 : OAI222_X1 port map( A1 => n1919, A2 => n2483, B1 => n11397, B2 => 
                           n3640, C1 => n1908, C2 => n2485, ZN => 
                           DataPath_RF_en_regi_57_port);
   U7870 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_58_port, A2 => n4199, ZN
                           => n16063);
   U7871 : OAI222_X1 port map( A1 => n2485, A2 => n1927, B1 => n11396, B2 => 
                           n3641, C1 => n1920, C2 => n2483, ZN => 
                           DataPath_RF_en_regi_58_port);
   U7872 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_59_port, A2 => n4198, ZN
                           => n16097);
   U7873 : OAI222_X1 port map( A1 => n2485, A2 => n1928, B1 => n11395, B2 => 
                           n3640, C1 => n1921, C2 => n2483, ZN => 
                           DataPath_RF_en_regi_59_port);
   U7874 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_60_port, A2 => n4198, ZN
                           => n16131);
   U7875 : OAI222_X1 port map( A1 => n2485, A2 => n1929, B1 => n11394, B2 => 
                           n3641, C1 => n1922, C2 => n2483, ZN => 
                           DataPath_RF_en_regi_60_port);
   U7876 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_61_port, A2 => n4197, ZN
                           => n16165);
   U7877 : OAI222_X1 port map( A1 => n2485, A2 => n1930, B1 => n11393, B2 => 
                           n3640, C1 => n1923, C2 => n2483, ZN => 
                           DataPath_RF_en_regi_61_port);
   U7878 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_62_port, A2 => n4197, ZN
                           => n16199);
   U7879 : OAI222_X1 port map( A1 => n2485, A2 => n1931, B1 => n11392, B2 => 
                           n3639, C1 => n1924, C2 => n2483, ZN => 
                           DataPath_RF_en_regi_62_port);
   U7880 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_63_port, A2 => n4196, ZN
                           => n16233);
   U7881 : OAI222_X1 port map( A1 => n1926, A2 => n2485, B1 => n11391, B2 => 
                           n3641, C1 => n1910, C2 => n2482, ZN => 
                           DataPath_RF_en_regi_63_port);
   U7882 : NAND2_X1 port map( A1 => n7077, A2 => n4257, ZN => n7979);
   U7883 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n549, ZN => n7991);
   U7884 : NAND2_X1 port map( A1 => n11580, A2 => DataPath_LDSTR_n79, ZN => 
                           DataPath_LDSTR_n57);
   U7885 : OAI221_X1 port map( B1 => n11348, B2 => n11577, C1 => n11578, C2 => 
                           DataPath_LDSTR_n70, A => DataPath_LDSTR_n62, ZN => 
                           DRAM_DATA_OUT_15_port);
   U7886 : INV_X1 port map( A => DRAM_DATA_OUT_7_port, ZN => n11348);
   U7887 : OAI221_X1 port map( B1 => n11363, B2 => n11575, C1 => n17106, C2 => 
                           DataPath_LDSTR_n40, A => DataPath_LDSTR_n45, ZN => 
                           DRAM_DATA_OUT_16_port);
   U7888 : OAI221_X1 port map( B1 => n11361, B2 => n11575, C1 => n17105, C2 => 
                           DataPath_LDSTR_n40, A => DataPath_LDSTR_n45, ZN => 
                           DRAM_DATA_OUT_17_port);
   U7889 : OAI221_X1 port map( B1 => n11359, B2 => n11575, C1 => 
                           DataPath_LDSTR_n40, C2 => n17104, A => 
                           DataPath_LDSTR_n45, ZN => DRAM_DATA_OUT_18_port);
   U7890 : OAI221_X1 port map( B1 => n11357, B2 => n11575, C1 => n17103, C2 => 
                           DataPath_LDSTR_n40, A => DataPath_LDSTR_n45, ZN => 
                           DRAM_DATA_OUT_19_port);
   U7891 : OAI221_X1 port map( B1 => n11355, B2 => n11575, C1 => n17101, C2 => 
                           DataPath_LDSTR_n40, A => DataPath_LDSTR_n45, ZN => 
                           DRAM_DATA_OUT_20_port);
   U7892 : OAI221_X1 port map( B1 => n11353, B2 => n11575, C1 => n17100, C2 => 
                           DataPath_LDSTR_n40, A => DataPath_LDSTR_n45, ZN => 
                           DRAM_DATA_OUT_21_port);
   U7893 : OAI221_X1 port map( B1 => n11351, B2 => n11575, C1 => n17099, C2 => 
                           DataPath_LDSTR_n40, A => DataPath_LDSTR_n45, ZN => 
                           DRAM_DATA_OUT_22_port);
   U7894 : AND2_X1 port map( A1 => n4136, A2 => n7196, ZN => n1907);
   U7895 : AOI22_X1 port map( A1 => n11349, A2 => DataPath_LDSTR_n60, B1 => 
                           DRAM_DATA_OUT_7_port, B2 => n11578, ZN => 
                           DataPath_LDSTR_n41);
   U7896 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11366, B1 => 
                           n11350, B2 => DataPath_LDSTR_n58, ZN => 
                           DataPath_LDSTR_n70);
   U7897 : INV_X1 port map( A => n17107, ZN => n11366);
   U7898 : INV_X1 port map( A => n4436, ZN => n7712);
   U7899 : OAI22_X1 port map( A1 => n17089, A2 => DataPath_LDSTR_n40, B1 => 
                           DataPath_LDSTR_n41, B2 => DataPath_LDSTR_n42, ZN => 
                           DRAM_DATA_OUT_31_port);
   U7900 : NOR2_X1 port map( A1 => n4127, A2 => n11480, ZN => 
                           DataPath_LDSTR_n42);
   U7901 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_23_port, A2 => n4172, ZN
                           => n14873);
   U7902 : OAI22_X1 port map( A1 => n2479, A2 => n1918, B1 => n3305, B2 => 
                           n11383, ZN => DataPath_RF_en_regi_23_port);
   U7903 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_80_port, A2 => n4188, ZN
                           => n16811);
   U7904 : OAI22_X1 port map( A1 => n3276, A2 => n1911, B1 => n3743, B2 => 
                           n11390, ZN => DataPath_RF_en_regi_80_port);
   U7905 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_81_port, A2 => n4187, ZN
                           => n16845);
   U7906 : OAI22_X1 port map( A1 => n3275, A2 => n1912, B1 => n3743, B2 => 
                           n11389, ZN => DataPath_RF_en_regi_81_port);
   U7907 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_82_port, A2 => n4187, ZN
                           => n16879);
   U7908 : OAI22_X1 port map( A1 => n3275, A2 => n1913, B1 => n3752, B2 => 
                           n11388, ZN => DataPath_RF_en_regi_82_port);
   U7909 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_83_port, A2 => n4186, ZN
                           => n16913);
   U7910 : OAI22_X1 port map( A1 => n3276, A2 => n1914, B1 => n3753, B2 => 
                           n11387, ZN => DataPath_RF_en_regi_83_port);
   U7911 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_84_port, A2 => n4186, ZN
                           => n16947);
   U7912 : OAI22_X1 port map( A1 => n3275, A2 => n1915, B1 => n3751, B2 => 
                           n11386, ZN => DataPath_RF_en_regi_84_port);
   U7913 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_86_port, A2 => n4185, ZN
                           => n17015);
   U7914 : OAI22_X1 port map( A1 => n3275, A2 => n1917, B1 => n3752, B2 => 
                           n11384, ZN => DataPath_RF_en_regi_86_port);
   U7915 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_16_port, A2 => n4175, ZN
                           => n14635);
   U7916 : OAI22_X1 port map( A1 => n2479, A2 => n1911, B1 => n3295, B2 => 
                           n11390, ZN => DataPath_RF_en_regi_16_port);
   U7917 : OAI22_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n587, A2 => n2984
                           , B1 => n11496, B2 => DataPath_ALUhw_SHIFTER_HW_n150
                           , ZN => DataPath_ALUhw_SHIFTER_HW_n586);
   U7918 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_39_port, A2 => n4164, ZN
                           => n15417);
   U7919 : OAI22_X1 port map( A1 => n1918, A2 => n2480, B1 => n11383, B2 => 
                           n3416, ZN => DataPath_RF_en_regi_39_port);
   U7920 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_55_port, A2 => n4200, ZN
                           => n15961);
   U7921 : OAI22_X1 port map( A1 => n1918, A2 => n2482, B1 => n11383, B2 => 
                           n3528, ZN => DataPath_RF_en_regi_55_port);
   U7922 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_64_port, A2 => n4196, ZN
                           => n16267);
   U7923 : OAI22_X1 port map( A1 => n1911, A2 => n2484, B1 => n11390, B2 => 
                           n3641, ZN => DataPath_RF_en_regi_64_port);
   U7924 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_65_port, A2 => n4195, ZN
                           => n16301);
   U7925 : OAI22_X1 port map( A1 => n1912, A2 => n2484, B1 => n11389, B2 => 
                           n3639, ZN => DataPath_RF_en_regi_65_port);
   U7926 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_66_port, A2 => n4195, ZN
                           => n16335);
   U7927 : OAI22_X1 port map( A1 => n1913, A2 => n2484, B1 => n11388, B2 => 
                           n3639, ZN => DataPath_RF_en_regi_66_port);
   U7928 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_67_port, A2 => n4194, ZN
                           => n16369);
   U7929 : OAI22_X1 port map( A1 => n1914, A2 => n2484, B1 => n11387, B2 => 
                           n3639, ZN => DataPath_RF_en_regi_67_port);
   U7930 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_68_port, A2 => n4194, ZN
                           => n16403);
   U7931 : OAI22_X1 port map( A1 => n1915, A2 => n2484, B1 => n11386, B2 => 
                           n3631, ZN => DataPath_RF_en_regi_68_port);
   U7932 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_69_port, A2 => n4193, ZN
                           => n16437);
   U7933 : OAI22_X1 port map( A1 => n1916, A2 => n2484, B1 => n11385, B2 => 
                           n3640, ZN => DataPath_RF_en_regi_69_port);
   U7934 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_70_port, A2 => n4193, ZN
                           => n16471);
   U7935 : OAI22_X1 port map( A1 => n1917, A2 => n2484, B1 => n11384, B2 => 
                           n3641, ZN => DataPath_RF_en_regi_70_port);
   U7936 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_71_port, A2 => n4192, ZN
                           => n16505);
   U7937 : OAI22_X1 port map( A1 => n1918, A2 => n2484, B1 => n11383, B2 => 
                           n3641, ZN => DataPath_RF_en_regi_71_port);
   U7938 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_87_port, A2 => n4184, ZN
                           => n17049);
   U7939 : OAI22_X1 port map( A1 => n3276, A2 => n1918, B1 => n11383, B2 => 
                           n3753, ZN => DataPath_RF_en_regi_87_port);
   U7940 : OAI22_X1 port map( A1 => n8313, A2 => DataPath_ALUhw_SHIFTER_HW_n181
                           , B1 => n8319, B2 => DataPath_ALUhw_SHIFTER_HW_n182,
                           ZN => DataPath_ALUhw_SHIFTER_HW_n331);
   U7941 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_9_port, A2 => n4179, ZN 
                           => n14397);
   U7942 : OAI222_X1 port map( A1 => n1919, A2 => n3277, B1 => n11397, B2 => 
                           n3304, C1 => n1908, C2 => n2479, ZN => 
                           DataPath_RF_en_regi_9_port);
   U7943 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_72_port, A2 => n4192, ZN
                           => n16539);
   U7944 : OAI222_X1 port map( A1 => n1925, A2 => n2485, B1 => n11398, B2 => 
                           n3753, C1 => n3272, C2 => n1909, ZN => 
                           DataPath_RF_en_regi_72_port);
   U7945 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_73_port, A2 => n4191, ZN
                           => n16573);
   U7946 : OAI222_X1 port map( A1 => n1919, A2 => n2485, B1 => n11397, B2 => 
                           n3752, C1 => n3272, C2 => n1908, ZN => 
                           DataPath_RF_en_regi_73_port);
   U7947 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_74_port, A2 => n4191, ZN
                           => n16607);
   U7948 : OAI222_X1 port map( A1 => n3273, A2 => n1927, B1 => n3752, B2 => 
                           n11396, C1 => n2484, C2 => n1920, ZN => 
                           DataPath_RF_en_regi_74_port);
   U7949 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_75_port, A2 => n4190, ZN
                           => n16641);
   U7950 : OAI222_X1 port map( A1 => n3274, A2 => n1928, B1 => n3753, B2 => 
                           n11395, C1 => n2485, C2 => n1921, ZN => 
                           DataPath_RF_en_regi_75_port);
   U7951 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_76_port, A2 => n4190, ZN
                           => n16675);
   U7952 : OAI222_X1 port map( A1 => n3274, A2 => n1929, B1 => n3751, B2 => 
                           n11394, C1 => n2484, C2 => n1922, ZN => 
                           DataPath_RF_en_regi_76_port);
   U7953 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_77_port, A2 => n4189, ZN
                           => n16709);
   U7954 : OAI222_X1 port map( A1 => n3273, A2 => n1930, B1 => n3751, B2 => 
                           n11393, C1 => n2484, C2 => n1923, ZN => 
                           DataPath_RF_en_regi_77_port);
   U7955 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_78_port, A2 => n4189, ZN
                           => n16743);
   U7956 : OAI222_X1 port map( A1 => n3274, A2 => n1931, B1 => n3753, B2 => 
                           n11392, C1 => n2484, C2 => n1924, ZN => 
                           DataPath_RF_en_regi_78_port);
   U7957 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_79_port, A2 => n4188, ZN
                           => n16777);
   U7958 : OAI222_X1 port map( A1 => n3274, A2 => n1926, B1 => n3751, B2 => 
                           n11391, C1 => n1910, C2 => n2485, ZN => 
                           DataPath_RF_en_regi_79_port);
   U7959 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_17_port, A2 => n4175, ZN
                           => n14669);
   U7960 : OAI22_X1 port map( A1 => n2479, A2 => n1912, B1 => n3304, B2 => 
                           n11389, ZN => DataPath_RF_en_regi_17_port);
   U7961 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_18_port, A2 => n4174, ZN
                           => n14703);
   U7962 : OAI22_X1 port map( A1 => n2479, A2 => n1913, B1 => n3303, B2 => 
                           n11388, ZN => DataPath_RF_en_regi_18_port);
   U7963 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_19_port, A2 => n4174, ZN
                           => n14737);
   U7964 : OAI22_X1 port map( A1 => n2479, A2 => n1914, B1 => n3305, B2 => 
                           n11387, ZN => DataPath_RF_en_regi_19_port);
   U7965 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_20_port, A2 => n4173, ZN
                           => n14771);
   U7966 : OAI22_X1 port map( A1 => n2479, A2 => n1915, B1 => n3303, B2 => 
                           n11386, ZN => DataPath_RF_en_regi_20_port);
   U7967 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_21_port, A2 => n4173, ZN
                           => n14805);
   U7968 : OAI22_X1 port map( A1 => n2479, A2 => n1916, B1 => n3304, B2 => 
                           n11385, ZN => DataPath_RF_en_regi_21_port);
   U7969 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_22_port, A2 => n4172, ZN
                           => n14839);
   U7970 : OAI22_X1 port map( A1 => n2479, A2 => n1917, B1 => n3303, B2 => 
                           n11384, ZN => DataPath_RF_en_regi_22_port);
   U7971 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_32_port, A2 => n4167, ZN
                           => n15179);
   U7972 : OAI22_X1 port map( A1 => n1911, A2 => n2480, B1 => n11390, B2 => 
                           n3417, ZN => DataPath_RF_en_regi_32_port);
   U7973 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_33_port, A2 => n4167, ZN
                           => n15213);
   U7974 : OAI22_X1 port map( A1 => n1912, A2 => n2480, B1 => n11389, B2 => 
                           n3407, ZN => DataPath_RF_en_regi_33_port);
   U7975 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_34_port, A2 => n4166, ZN
                           => n15247);
   U7976 : OAI22_X1 port map( A1 => n1913, A2 => n2480, B1 => n11388, B2 => 
                           n3415, ZN => DataPath_RF_en_regi_34_port);
   U7977 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_35_port, A2 => n4166, ZN
                           => n15281);
   U7978 : OAI22_X1 port map( A1 => n1914, A2 => n2480, B1 => n11387, B2 => 
                           n3417, ZN => DataPath_RF_en_regi_35_port);
   U7979 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_36_port, A2 => n4165, ZN
                           => n15315);
   U7980 : OAI22_X1 port map( A1 => n1915, A2 => n2480, B1 => n11386, B2 => 
                           n3416, ZN => DataPath_RF_en_regi_36_port);
   U7981 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_37_port, A2 => n4165, ZN
                           => n15349);
   U7982 : OAI22_X1 port map( A1 => n1916, A2 => n2480, B1 => n11385, B2 => 
                           n3415, ZN => DataPath_RF_en_regi_37_port);
   U7983 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_38_port, A2 => n4164, ZN
                           => n15383);
   U7984 : OAI22_X1 port map( A1 => n1917, A2 => n2480, B1 => n11384, B2 => 
                           n3408, ZN => DataPath_RF_en_regi_38_port);
   U7985 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_48_port, A2 => n4159, ZN
                           => n15723);
   U7986 : OAI22_X1 port map( A1 => n1911, A2 => n2482, B1 => n11390, B2 => 
                           n3529, ZN => DataPath_RF_en_regi_48_port);
   U7987 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_49_port, A2 => n4159, ZN
                           => n15757);
   U7988 : OAI22_X1 port map( A1 => n1912, A2 => n2482, B1 => n11389, B2 => 
                           n3520, ZN => DataPath_RF_en_regi_49_port);
   U7989 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_50_port, A2 => n4158, ZN
                           => n15791);
   U7990 : OAI22_X1 port map( A1 => n1913, A2 => n2482, B1 => n11388, B2 => 
                           n3527, ZN => DataPath_RF_en_regi_50_port);
   U7991 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_51_port, A2 => n4158, ZN
                           => n15825);
   U7992 : OAI22_X1 port map( A1 => n1914, A2 => n2482, B1 => n11387, B2 => 
                           n3529, ZN => DataPath_RF_en_regi_51_port);
   U7993 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_52_port, A2 => n4172, ZN
                           => n15859);
   U7994 : OAI22_X1 port map( A1 => n1915, A2 => n2482, B1 => n11386, B2 => 
                           n3528, ZN => DataPath_RF_en_regi_52_port);
   U7995 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_53_port, A2 => n4201, ZN
                           => n15893);
   U7996 : OAI22_X1 port map( A1 => n1916, A2 => n2482, B1 => n11385, B2 => 
                           n3527, ZN => DataPath_RF_en_regi_53_port);
   U7997 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_54_port, A2 => n4201, ZN
                           => n15927);
   U7998 : OAI22_X1 port map( A1 => n1917, A2 => n2482, B1 => n11384, B2 => 
                           n3519, ZN => DataPath_RF_en_regi_54_port);
   U7999 : NOR2_X1 port map( A1 => DataPath_RF_en_regi_85_port, A2 => n4185, ZN
                           => n16981);
   U8000 : OAI22_X1 port map( A1 => n3276, A2 => n1916, B1 => n3743, B2 => 
                           n11385, ZN => DataPath_RF_en_regi_85_port);
   U8001 : NAND2_X1 port map( A1 => n11498, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n641, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n598);
   U8002 : NOR2_X1 port map( A1 => n408, A2 => DataPath_LDSTR_n80, ZN => 
                           DataPath_LDSTR_n83);
   U8003 : OAI211_X1 port map( C1 => DataPath_LDSTR_n39, C2 => 
                           DataPath_LDSTR_n44, A => DataPath_LDSTR_n45, B => 
                           DataPath_LDSTR_n59, ZN => DRAM_DATA_OUT_24_port);
   U8004 : AOI22_X1 port map( A1 => n11576, A2 => n11364, B1 => 
                           DataPath_LDSTR_n47, B2 => DRAM_DATA_OUT_0_port, ZN 
                           => DataPath_LDSTR_n59);
   U8005 : OAI211_X1 port map( C1 => DataPath_LDSTR_n37, C2 => 
                           DataPath_LDSTR_n44, A => DataPath_LDSTR_n45, B => 
                           DataPath_LDSTR_n56, ZN => DRAM_DATA_OUT_25_port);
   U8006 : AOI22_X1 port map( A1 => n11576, A2 => n11362, B1 => 
                           DataPath_LDSTR_n47, B2 => DRAM_DATA_OUT_1_port, ZN 
                           => DataPath_LDSTR_n56);
   U8007 : OAI211_X1 port map( C1 => DataPath_LDSTR_n54, C2 => 
                           DataPath_LDSTR_n44, A => DataPath_LDSTR_n45, B => 
                           DataPath_LDSTR_n55, ZN => DRAM_DATA_OUT_26_port);
   U8008 : AOI22_X1 port map( A1 => n11360, A2 => n11576, B1 => 
                           DataPath_LDSTR_n47, B2 => DRAM_DATA_OUT_2_port, ZN 
                           => DataPath_LDSTR_n55);
   U8009 : OAI211_X1 port map( C1 => DataPath_LDSTR_n52, C2 => 
                           DataPath_LDSTR_n44, A => DataPath_LDSTR_n45, B => 
                           DataPath_LDSTR_n53, ZN => DRAM_DATA_OUT_27_port);
   U8010 : AOI22_X1 port map( A1 => n11576, A2 => n11358, B1 => 
                           DataPath_LDSTR_n47, B2 => DRAM_DATA_OUT_3_port, ZN 
                           => DataPath_LDSTR_n53);
   U8011 : OAI211_X1 port map( C1 => DataPath_LDSTR_n50, C2 => 
                           DataPath_LDSTR_n44, A => DataPath_LDSTR_n45, B => 
                           DataPath_LDSTR_n51, ZN => DRAM_DATA_OUT_28_port);
   U8012 : AOI22_X1 port map( A1 => n11576, A2 => n11356, B1 => 
                           DataPath_LDSTR_n47, B2 => DRAM_DATA_OUT_4_port, ZN 
                           => DataPath_LDSTR_n51);
   U8013 : OAI211_X1 port map( C1 => DataPath_LDSTR_n48, C2 => 
                           DataPath_LDSTR_n44, A => DataPath_LDSTR_n45, B => 
                           DataPath_LDSTR_n49, ZN => DRAM_DATA_OUT_29_port);
   U8014 : AOI22_X1 port map( A1 => n11576, A2 => n11354, B1 => 
                           DataPath_LDSTR_n47, B2 => DRAM_DATA_OUT_5_port, ZN 
                           => DataPath_LDSTR_n49);
   U8015 : OAI211_X1 port map( C1 => DataPath_LDSTR_n43, C2 => 
                           DataPath_LDSTR_n44, A => DataPath_LDSTR_n45, B => 
                           DataPath_LDSTR_n46, ZN => DRAM_DATA_OUT_30_port);
   U8016 : AOI22_X1 port map( A1 => n11576, A2 => n11352, B1 => 
                           DataPath_LDSTR_n47, B2 => DRAM_DATA_OUT_6_port, ZN 
                           => DataPath_LDSTR_n46);
   U8017 : AOI21_X1 port map( B1 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_27_port, B2
                           => n364, A => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_28_port, ZN
                           => n12916);
   U8018 : BUF_X1 port map( A => DataPath_ALUhw_BWISE_n70, Z => n2985);
   U8019 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n349, ZN => n11497);
   U8020 : NAND4_X1 port map( A1 => DataPath_LDSTR_n60, A2 => n4118, A3 => 
                           n11349, A4 => n11480, ZN => DataPath_LDSTR_n61);
   U8021 : AOI22_X1 port map( A1 => DataPath_LDSTR_n64, A2 => 
                           DRAM_DATA_OUT_7_port, B1 => n11576, B2 => n11365, ZN
                           => DataPath_LDSTR_n63);
   U8022 : INV_X1 port map( A => n17098, ZN => n11365);
   U8023 : BUF_X1 port map( A => n3844, Z => n3891);
   U8024 : AOI21_X1 port map( B1 => n11526, B2 => n376, A => n11527, ZN => 
                           n12920);
   U8025 : NAND2_X1 port map( A1 => n12960, A2 => n11607, ZN => n12959);
   U8026 : INV_X1 port map( A => DataPath_LDSTR_n72, ZN => n11580);
   U8027 : BUF_X1 port map( A => n4140, Z => n4135);
   U8028 : BUF_X1 port map( A => n4135, Z => n4132);
   U8029 : BUF_X1 port map( A => n4138, Z => n4136);
   U8030 : INV_X1 port map( A => DRAM_DATA_OUT_0_port, ZN => n11363);
   U8031 : INV_X1 port map( A => DRAM_DATA_OUT_1_port, ZN => n11361);
   U8032 : INV_X1 port map( A => DRAM_DATA_OUT_2_port, ZN => n11359);
   U8033 : INV_X1 port map( A => DRAM_DATA_OUT_3_port, ZN => n11357);
   U8034 : INV_X1 port map( A => DRAM_DATA_OUT_4_port, ZN => n11355);
   U8035 : INV_X1 port map( A => DRAM_DATA_OUT_5_port, ZN => n11353);
   U8036 : INV_X1 port map( A => DRAM_DATA_OUT_6_port, ZN => n11351);
   U8037 : BUF_X1 port map( A => n4135, Z => n4138);
   U8038 : BUF_X1 port map( A => n4138, Z => n4137);
   U8039 : BUF_X1 port map( A => n4136, Z => n4139);
   U8040 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n576, ZN => n11498);
   U8041 : NOR2_X1 port map( A1 => n4207, A2 => DataPath_WRF_CUhw_n141, ZN => 
                           DataPath_WRF_CUhw_N150_port);
   U8042 : NOR2_X1 port map( A1 => n4207, A2 => DataPath_WRF_CUhw_n140, ZN => 
                           DataPath_WRF_CUhw_N151);
   U8043 : NOR2_X1 port map( A1 => n4207, A2 => DataPath_WRF_CUhw_n139, ZN => 
                           DataPath_WRF_CUhw_N152_port);
   U8044 : NOR2_X1 port map( A1 => n4208, A2 => DataPath_WRF_CUhw_n138, ZN => 
                           DataPath_WRF_CUhw_N153_port);
   U8045 : NOR2_X1 port map( A1 => n4208, A2 => DataPath_WRF_CUhw_n137, ZN => 
                           DataPath_WRF_CUhw_N154_port);
   U8046 : NOR2_X1 port map( A1 => n4208, A2 => DataPath_WRF_CUhw_n136, ZN => 
                           DataPath_WRF_CUhw_N155_port);
   U8047 : NOR2_X1 port map( A1 => n4208, A2 => DataPath_WRF_CUhw_n135, ZN => 
                           DataPath_WRF_CUhw_N156_port);
   U8048 : NOR2_X1 port map( A1 => n4209, A2 => DataPath_WRF_CUhw_n134, ZN => 
                           DataPath_WRF_CUhw_N157_port);
   U8049 : NOR2_X1 port map( A1 => n4209, A2 => DataPath_WRF_CUhw_n133, ZN => 
                           DataPath_WRF_CUhw_N158_port);
   U8050 : NOR2_X1 port map( A1 => n4209, A2 => DataPath_WRF_CUhw_n132, ZN => 
                           DataPath_WRF_CUhw_N159_port);
   U8051 : NOR2_X1 port map( A1 => n4209, A2 => DataPath_WRF_CUhw_n131, ZN => 
                           DataPath_WRF_CUhw_N160_port);
   U8052 : NOR2_X1 port map( A1 => n4210, A2 => DataPath_WRF_CUhw_n130, ZN => 
                           DataPath_WRF_CUhw_N161_port);
   U8053 : NAND2_X1 port map( A1 => DataPath_LDSTR_n83, A2 => n11574, ZN => 
                           DataPath_LDSTR_n65);
   U8054 : INV_X1 port map( A => DataPath_LDSTR_n69, ZN => n11574);
   U8055 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n12, A2 => 
                           DataPath_ALUhw_MUXOUT_n13, ZN => 
                           DataPath_i_ALU_OUT_6_port);
   U8056 : AOI22_X1 port map( A1 => n11514, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_102_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n12);
   U8057 : NAND2_X1 port map( A1 => DataPath_ALUhw_MUXOUT_n14, A2 => 
                           DataPath_ALUhw_MUXOUT_n15, ZN => 
                           DataPath_i_ALU_OUT_5_port);
   U8058 : AOI22_X1 port map( A1 => n11513, A2 => n2271, B1 => 
                           DataPath_ALUhw_i_Q_EXTENDED_101_port, B2 => n8321, 
                           ZN => DataPath_ALUhw_MUXOUT_n14);
   U8059 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n478, ZN => n11499);
   U8060 : BUF_X1 port map( A => n11542, Z => n2284);
   U8061 : BUF_X1 port map( A => n11542, Z => n2283);
   U8062 : BUF_X1 port map( A => n11549, Z => n2325);
   U8063 : BUF_X1 port map( A => n11543, Z => n2290);
   U8064 : BUF_X1 port map( A => n11544, Z => n2296);
   U8065 : BUF_X1 port map( A => n11545, Z => n2302);
   U8066 : BUF_X1 port map( A => n11546, Z => n2308);
   U8067 : BUF_X1 port map( A => n11547, Z => n2314);
   U8068 : BUF_X1 port map( A => n11548, Z => n2320);
   U8069 : BUF_X1 port map( A => n11549, Z => n2326);
   U8070 : BUF_X1 port map( A => n11543, Z => n2289);
   U8071 : BUF_X1 port map( A => n11544, Z => n2295);
   U8072 : BUF_X1 port map( A => n11545, Z => n2301);
   U8073 : BUF_X1 port map( A => n11546, Z => n2307);
   U8074 : BUF_X1 port map( A => n11547, Z => n2313);
   U8075 : BUF_X1 port map( A => n11548, Z => n2319);
   U8076 : BUF_X1 port map( A => n11550, Z => n2331);
   U8077 : BUF_X1 port map( A => n11552, Z => n2343);
   U8078 : BUF_X1 port map( A => n11553, Z => n2349);
   U8079 : BUF_X1 port map( A => n11554, Z => n2355);
   U8080 : BUF_X1 port map( A => n11555, Z => n2361);
   U8081 : BUF_X1 port map( A => n11556, Z => n2367);
   U8082 : BUF_X1 port map( A => n11557, Z => n2373);
   U8083 : BUF_X1 port map( A => n11558, Z => n2379);
   U8084 : BUF_X1 port map( A => n11559, Z => n2385);
   U8085 : BUF_X1 port map( A => n11560, Z => n2391);
   U8086 : BUF_X1 port map( A => n11561, Z => n2397);
   U8087 : BUF_X1 port map( A => n11563, Z => n2409);
   U8088 : BUF_X1 port map( A => n11564, Z => n2415);
   U8089 : BUF_X1 port map( A => n11565, Z => n2421);
   U8090 : BUF_X1 port map( A => n11566, Z => n2427);
   U8091 : BUF_X1 port map( A => n11567, Z => n2433);
   U8092 : BUF_X1 port map( A => n11568, Z => n2439);
   U8093 : BUF_X1 port map( A => n11569, Z => n2445);
   U8094 : BUF_X1 port map( A => n11570, Z => n2451);
   U8095 : BUF_X1 port map( A => n11571, Z => n2457);
   U8096 : BUF_X1 port map( A => n11572, Z => n2463);
   U8097 : BUF_X1 port map( A => n11551, Z => n2337);
   U8098 : BUF_X1 port map( A => n11562, Z => n2403);
   U8099 : BUF_X1 port map( A => n11573, Z => n2469);
   U8100 : BUF_X1 port map( A => n11550, Z => n2332);
   U8101 : BUF_X1 port map( A => n11552, Z => n2344);
   U8102 : BUF_X1 port map( A => n11553, Z => n2350);
   U8103 : BUF_X1 port map( A => n11554, Z => n2356);
   U8104 : BUF_X1 port map( A => n11555, Z => n2362);
   U8105 : BUF_X1 port map( A => n11556, Z => n2368);
   U8106 : BUF_X1 port map( A => n11557, Z => n2374);
   U8107 : BUF_X1 port map( A => n11558, Z => n2380);
   U8108 : BUF_X1 port map( A => n11559, Z => n2386);
   U8109 : BUF_X1 port map( A => n11560, Z => n2392);
   U8110 : BUF_X1 port map( A => n11561, Z => n2398);
   U8111 : BUF_X1 port map( A => n11563, Z => n2410);
   U8112 : BUF_X1 port map( A => n11564, Z => n2416);
   U8113 : BUF_X1 port map( A => n11565, Z => n2422);
   U8114 : BUF_X1 port map( A => n11566, Z => n2428);
   U8115 : BUF_X1 port map( A => n11567, Z => n2434);
   U8116 : BUF_X1 port map( A => n11568, Z => n2440);
   U8117 : BUF_X1 port map( A => n11569, Z => n2446);
   U8118 : BUF_X1 port map( A => n11570, Z => n2452);
   U8119 : BUF_X1 port map( A => n11571, Z => n2458);
   U8120 : BUF_X1 port map( A => n11572, Z => n2464);
   U8121 : BUF_X1 port map( A => n11551, Z => n2338);
   U8122 : BUF_X1 port map( A => n11562, Z => n2404);
   U8123 : BUF_X1 port map( A => n11573, Z => n2470);
   U8124 : INV_X1 port map( A => DataPath_ALUhw_BWISE_n137, ZN => n11500);
   U8125 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n639, ZN => n11538);
   U8126 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_1_0_port, Z => 
                           n3406);
   U8127 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_0_0_port, Z => 
                           n3294);
   U8128 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_4_0_port, Z => 
                           n3742);
   U8129 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_2_0_port, Z => 
                           n3518);
   U8130 : OAI21_X2 port map( B1 => DataPath_RF_PUSH_ADDRGEN_n35, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_n32, A => 
                           DataPath_RF_PUSH_ADDRGEN_n26, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n52);
   U8131 : NOR2_X1 port map( A1 => DataPath_RF_n9, A2 => 
                           DataPath_i_DONE_FILL_EX, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5);
   U8132 : NOR2_X1 port map( A1 => i_EN3, A2 => n4182, ZN => n14237);
   U8133 : NAND2_X1 port map( A1 => DataPath_LDSTR_n71, A2 => 
                           DataPath_LDSTR_n72, ZN => DataPath_LDSTR_n40);
   U8134 : NAND2_X1 port map( A1 => DataPath_LDSTR_n60, A2 => n4119, ZN => 
                           DataPath_LDSTR_n44);
   U8135 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11373, B1 => 
                           DataPath_LDSTR_n58, B2 => n11364, ZN => 
                           DataPath_LDSTR_n39);
   U8136 : INV_X1 port map( A => n17083, ZN => n11373);
   U8137 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11371, B1 => 
                           DataPath_LDSTR_n58, B2 => n11360, ZN => 
                           DataPath_LDSTR_n54);
   U8138 : INV_X1 port map( A => n17112, ZN => n11371);
   U8139 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11370, B1 => 
                           DataPath_LDSTR_n58, B2 => n11358, ZN => 
                           DataPath_LDSTR_n52);
   U8140 : INV_X1 port map( A => n17111, ZN => n11370);
   U8141 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11369, B1 => 
                           DataPath_LDSTR_n58, B2 => n11356, ZN => 
                           DataPath_LDSTR_n50);
   U8142 : INV_X1 port map( A => n17110, ZN => n11369);
   U8143 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11368, B1 => 
                           DataPath_LDSTR_n58, B2 => n11354, ZN => 
                           DataPath_LDSTR_n48);
   U8144 : INV_X1 port map( A => n17109, ZN => n11368);
   U8145 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11367, B1 => 
                           DataPath_LDSTR_n58, B2 => n11352, ZN => 
                           DataPath_LDSTR_n43);
   U8146 : INV_X1 port map( A => n17108, ZN => n11367);
   U8147 : INV_X1 port map( A => n7083, ZN => n8322);
   U8148 : AOI22_X1 port map( A1 => DataPath_LDSTR_n57, A2 => n11372, B1 => 
                           n11362, B2 => DataPath_LDSTR_n58, ZN => 
                           DataPath_LDSTR_n37);
   U8149 : INV_X1 port map( A => n17082, ZN => n11372);
   U8150 : AND2_X1 port map( A1 => DataPath_i_DONE_FILL_EX, A2 => 
                           DataPath_RF_n9, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4);
   U8151 : AND2_X1 port map( A1 => n11431, A2 => DataPath_i_DONE_FILL_EX, ZN =>
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7);
   U8152 : INV_X1 port map( A => DataPath_RF_n9, ZN => n11431);
   U8153 : BUF_X1 port map( A => n11595, Z => n2485);
   U8154 : BUF_X1 port map( A => n11541, Z => n2282);
   U8155 : BUF_X1 port map( A => DataPath_WRF_CUhw_n148, Z => n3263);
   U8156 : BUF_X1 port map( A => DataPath_WRF_CUhw_n148, Z => n3262);
   U8157 : NOR2_X1 port map( A1 => i_EN3, A2 => n4181, ZN => n14295);
   U8158 : NOR2_X1 port map( A1 => i_EN3, A2 => n4181, ZN => n14329);
   U8159 : BUF_X1 port map( A => n11595, Z => n2484);
   U8160 : BUF_X1 port map( A => n11594, Z => n2483);
   U8161 : BUF_X1 port map( A => n11594, Z => n2482);
   U8162 : BUF_X1 port map( A => n11592, Z => n2478);
   U8163 : BUF_X1 port map( A => n11593, Z => n2480);
   U8164 : BUF_X1 port map( A => n11593, Z => n2481);
   U8165 : BUF_X1 port map( A => n11592, Z => n2479);
   U8166 : BUF_X1 port map( A => DataPath_WRF_CUhw_n148, Z => n3264);
   U8167 : NOR2_X1 port map( A1 => n11578, A2 => DataPath_LDSTR_n60, ZN => 
                           DataPath_LDSTR_n71);
   U8168 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_9_port, A2 => n3911,
                           ZN => n1908);
   U8169 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_8_port, A2 => n3911,
                           ZN => n1909);
   U8170 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_31_port, A2 => n3911
                           , ZN => n1910);
   U8171 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_16_port, A2 => n3913
                           , ZN => n1911);
   U8172 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_17_port, A2 => n3912
                           , ZN => n1912);
   U8173 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_18_port, A2 => n3912
                           , ZN => n1913);
   U8174 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_19_port, A2 => n3912
                           , ZN => n1914);
   U8175 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_20_port, A2 => n3912
                           , ZN => n1915);
   U8176 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_21_port, A2 => n3912
                           , ZN => n1916);
   U8177 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_22_port, A2 => n3912
                           , ZN => n1917);
   U8178 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_23_port, A2 => n3912
                           , ZN => n1918);
   U8179 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_25_port, A2 => n3912
                           , ZN => n1919);
   U8180 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_26_port, A2 => n3912
                           , ZN => n1920);
   U8181 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_27_port, A2 => n3912
                           , ZN => n1921);
   U8182 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_28_port, A2 => n3911
                           , ZN => n1922);
   U8183 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_29_port, A2 => n3911
                           , ZN => n1923);
   U8184 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_30_port, A2 => n3911
                           , ZN => n1924);
   U8185 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_24_port, A2 => n3912
                           , ZN => n1925);
   U8186 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_15_port, A2 => n3913
                           , ZN => n1926);
   U8187 : NAND2_X1 port map( A1 => n4261, A2 => n12958, ZN => n12955);
   U8188 : OAI21_X1 port map( B1 => n11607, B2 => n12951, A => n12959, ZN => 
                           n12958);
   U8189 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_10_port, A2 => n3913
                           , ZN => n1927);
   U8190 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_11_port, A2 => n3913
                           , ZN => n1928);
   U8191 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_12_port, A2 => n3913
                           , ZN => n1929);
   U8192 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_13_port, A2 => n3913
                           , ZN => n1930);
   U8193 : NAND2_X1 port map( A1 => DataPath_RF_dec_output_14_port, A2 => n3913
                           , ZN => n1931);
   U8194 : BUF_X1 port map( A => DataPath_ALUhw_BWISE_n70, Z => n2986);
   U8195 : MUX2_X1 port map( A => n7517, B => n7518, S => n7516, Z => n7519);
   U8196 : BUF_X1 port map( A => DataPath_i_WF, Z => n3911);
   U8197 : BUF_X1 port map( A => DataPath_i_WF, Z => n3912);
   U8198 : NOR2_X1 port map( A1 => n12970, A2 => n4157, ZN => 
                           DataPath_RF_POP_ADDRGEN_N61);
   U8199 : NOR2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n45, A2 => n4184, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N61);
   U8200 : AND2_X1 port map( A1 => CU_I_n71, A2 => n4260, ZN => n1932);
   U8201 : OAI21_X1 port map( B1 => DataPath_WRF_CUhw_N26_port, B2 => n303, A 
                           => DataPath_WRF_CUhw_n150, ZN => 
                           DataPath_WRF_CUhw_n154);
   U8202 : NAND2_X1 port map( A1 => n4262, A2 => DataPath_RF_PUSH_ADDRGEN_n33, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_n30);
   U8203 : OAI21_X1 port map( B1 => n3909, B2 => DataPath_RF_PUSH_ADDRGEN_n26, 
                           A => DataPath_RF_PUSH_ADDRGEN_n34, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n33);
   U8204 : NAND2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n35, A2 => n11597,
                           ZN => DataPath_RF_PUSH_ADDRGEN_n34);
   U8205 : BUF_X1 port map( A => DataPath_i_WF, Z => n3913);
   U8206 : AOI21_X1 port map( B1 => DataPath_WRF_CUhw_n146, B2 => 
                           DataPath_WRF_CUhw_n147, A => n4218, ZN => 
                           DataPath_WRF_CUhw_N145_port);
   U8207 : AOI221_X1 port map( B1 => n3264, B2 => n11382, C1 => n2477, C2 => 
                           n11400, A => DataPath_WRF_CUhw_n149, ZN => 
                           DataPath_WRF_CUhw_n147);
   U8208 : AOI22_X1 port map( A1 => n3264, A2 => n3901, B1 => 
                           DataPath_WRF_CUhw_N26_port, B2 => n3265, ZN => 
                           DataPath_WRF_CUhw_n146);
   U8209 : AOI21_X1 port map( B1 => n303, B2 => DataPath_WRF_CUhw_n150, A => 
                           n12957, ZN => DataPath_WRF_CUhw_n149);
   U8210 : BUF_X1 port map( A => n4139, Z => n4133);
   U8211 : INV_X1 port map( A => DataPath_WRF_CUhw_n150, ZN => n11590);
   U8212 : NOR2_X1 port map( A1 => n4107, A2 => n11481, ZN => CU_I_n151);
   U8213 : NOR2_X1 port map( A1 => n4207, A2 => DataPath_WRF_CUhw_n142, ZN => 
                           DataPath_WRF_CUhw_N149_port);
   U8214 : NOR2_X1 port map( A1 => n4202, A2 => DataPath_WRF_CUhw_n145, ZN => 
                           DataPath_WRF_CUhw_N146_port);
   U8215 : NOR2_X1 port map( A1 => n4206, A2 => DataPath_WRF_CUhw_n144, ZN => 
                           DataPath_WRF_CUhw_N147_port);
   U8216 : NOR2_X1 port map( A1 => n4206, A2 => DataPath_WRF_CUhw_n143, ZN => 
                           DataPath_WRF_CUhw_N148_port);
   U8217 : NOR2_X1 port map( A1 => n4206, A2 => n12969, ZN => 
                           DataPath_RF_POP_ADDRGEN_N47);
   U8218 : NOR2_X1 port map( A1 => n4206, A2 => n12968, ZN => 
                           DataPath_RF_POP_ADDRGEN_N48);
   U8219 : NOR2_X1 port map( A1 => n4205, A2 => n12967, ZN => 
                           DataPath_RF_POP_ADDRGEN_N49);
   U8220 : NOR2_X1 port map( A1 => n4205, A2 => n12966, ZN => 
                           DataPath_RF_POP_ADDRGEN_N50);
   U8221 : NOR2_X1 port map( A1 => n4205, A2 => n12965, ZN => 
                           DataPath_RF_POP_ADDRGEN_N51);
   U8222 : NOR2_X1 port map( A1 => n4205, A2 => n12964, ZN => 
                           DataPath_RF_POP_ADDRGEN_N52);
   U8223 : NOR2_X1 port map( A1 => n4204, A2 => n12963, ZN => 
                           DataPath_RF_POP_ADDRGEN_N53);
   U8224 : NOR2_X1 port map( A1 => n4204, A2 => n12962, ZN => 
                           DataPath_RF_POP_ADDRGEN_N54);
   U8225 : NOR2_X1 port map( A1 => n4204, A2 => n12961, ZN => 
                           DataPath_RF_POP_ADDRGEN_N55);
   U8226 : NOR2_X1 port map( A1 => n4204, A2 => n12975, ZN => 
                           DataPath_RF_POP_ADDRGEN_N56);
   U8227 : NOR2_X1 port map( A1 => n4203, A2 => n12974, ZN => 
                           DataPath_RF_POP_ADDRGEN_N57);
   U8228 : NOR2_X1 port map( A1 => n4203, A2 => n12973, ZN => 
                           DataPath_RF_POP_ADDRGEN_N58);
   U8229 : NOR2_X1 port map( A1 => n4203, A2 => n12972, ZN => 
                           DataPath_RF_POP_ADDRGEN_N59);
   U8230 : NOR2_X1 port map( A1 => n4203, A2 => n12971, ZN => 
                           DataPath_RF_POP_ADDRGEN_N60);
   U8231 : NOR2_X1 port map( A1 => n4214, A2 => DataPath_RF_PUSH_ADDRGEN_n44, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N47_port);
   U8232 : NOR2_X1 port map( A1 => n4214, A2 => DataPath_RF_PUSH_ADDRGEN_n43, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N48_port);
   U8233 : NOR2_X1 port map( A1 => n4215, A2 => DataPath_RF_PUSH_ADDRGEN_n42, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N49_port);
   U8234 : NOR2_X1 port map( A1 => n4215, A2 => DataPath_RF_PUSH_ADDRGEN_n41, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N50_port);
   U8235 : NOR2_X1 port map( A1 => n4215, A2 => DataPath_RF_PUSH_ADDRGEN_n40, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N51_port);
   U8236 : NOR2_X1 port map( A1 => n4215, A2 => DataPath_RF_PUSH_ADDRGEN_n39, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N52_port);
   U8237 : NOR2_X1 port map( A1 => n4216, A2 => DataPath_RF_PUSH_ADDRGEN_n38, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N53_port);
   U8238 : NOR2_X1 port map( A1 => n4216, A2 => DataPath_RF_PUSH_ADDRGEN_n37, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N54_port);
   U8239 : NOR2_X1 port map( A1 => n4216, A2 => DataPath_RF_PUSH_ADDRGEN_n36, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N55);
   U8240 : NOR2_X1 port map( A1 => n4216, A2 => DataPath_RF_PUSH_ADDRGEN_n50, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N56);
   U8241 : NOR2_X1 port map( A1 => n4217, A2 => DataPath_RF_PUSH_ADDRGEN_n49, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N57);
   U8242 : NOR2_X1 port map( A1 => n4217, A2 => DataPath_RF_PUSH_ADDRGEN_n48, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N58);
   U8243 : NOR2_X1 port map( A1 => n4212, A2 => DataPath_RF_PUSH_ADDRGEN_n47, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N59);
   U8244 : NOR2_X1 port map( A1 => n4202, A2 => DataPath_RF_PUSH_ADDRGEN_n46, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N60);
   U8245 : NOR2_X1 port map( A1 => n1438, A2 => n4107, ZN => CU_I_n128);
   U8246 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_31_port, Z => 
                           n3914);
   U8247 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_30_port, Z => 
                           n3920);
   U8248 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_29_port, Z => 
                           n3926);
   U8249 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_28_port, Z => 
                           n3932);
   U8250 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_27_port, Z => 
                           n3938);
   U8251 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_26_port, Z => 
                           n3944);
   U8252 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_25_port, Z => 
                           n3950);
   U8253 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_24_port, Z => 
                           n3956);
   U8254 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_23_port, Z => 
                           n3962);
   U8255 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_22_port, Z => 
                           n3968);
   U8256 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_21_port, Z => 
                           n3974);
   U8257 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_20_port, Z => 
                           n3980);
   U8258 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_19_port, Z => 
                           n3986);
   U8259 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_18_port, Z => 
                           n3992);
   U8260 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_17_port, Z => 
                           n3998);
   U8261 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_16_port, Z => 
                           n4004);
   U8262 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_15_port, Z => 
                           n4010);
   U8263 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_14_port, Z => 
                           n4016);
   U8264 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_13_port, Z => 
                           n4022);
   U8265 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_12_port, Z => 
                           n4028);
   U8266 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_10_port, Z => 
                           n4040);
   U8267 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_9_port, Z => 
                           n4046);
   U8268 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_8_port, Z => 
                           n4052);
   U8269 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_7_port, Z => 
                           n4058);
   U8270 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_6_port, Z => 
                           n4064);
   U8271 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_5_port, Z => 
                           n4070);
   U8272 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_4_port, Z => 
                           n4076);
   U8273 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_3_port, Z => 
                           n4082);
   U8274 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_2_port, Z => 
                           n4088);
   U8275 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_1_port, Z => 
                           n4094);
   U8276 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_0_port, Z => 
                           n4100);
   U8277 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_11_port, Z => 
                           n4034);
   U8278 : AND2_X1 port map( A1 => DataPath_LDSTR_n60, A2 => n408, ZN => 
                           DataPath_LDSTR_n78);
   U8279 : INV_X1 port map( A => n17089, ZN => n11350);
   U8280 : INV_X1 port map( A => n12956, ZN => n8647);
   U8281 : OAI21_X1 port map( B1 => n12957, B2 => n12952, A => n12955, ZN => 
                           n12956);
   U8282 : INV_X1 port map( A => DataPath_RF_PUSH_ADDRGEN_n31, ZN => n8648);
   U8283 : OAI21_X1 port map( B1 => DataPath_RF_PUSH_ADDRGEN_n32, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_n27, A => 
                           DataPath_RF_PUSH_ADDRGEN_n30, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n31);
   U8284 : NAND2_X1 port map( A1 => n12976, A2 => n4266, ZN => 
                           DataPath_RF_POP_ADDRGEN_N46);
   U8285 : NAND2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n51, A2 => n4260, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_N46_port);
   U8286 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_10_port, Z => 
                           n4041);
   U8287 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_9_port, Z => 
                           n4047);
   U8288 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_8_port, Z => 
                           n4053);
   U8289 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_7_port, Z => 
                           n4059);
   U8290 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_6_port, Z => 
                           n4065);
   U8291 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_5_port, Z => 
                           n4071);
   U8292 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_4_port, Z => 
                           n4077);
   U8293 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_31_port, Z => 
                           n3915);
   U8294 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_30_port, Z => 
                           n3921);
   U8295 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_29_port, Z => 
                           n3927);
   U8296 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_28_port, Z => 
                           n3933);
   U8297 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_27_port, Z => 
                           n3939);
   U8298 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_26_port, Z => 
                           n3945);
   U8299 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_25_port, Z => 
                           n3951);
   U8300 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_24_port, Z => 
                           n3957);
   U8301 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_23_port, Z => 
                           n3963);
   U8302 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_22_port, Z => 
                           n3969);
   U8303 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_21_port, Z => 
                           n3975);
   U8304 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_20_port, Z => 
                           n3981);
   U8305 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_19_port, Z => 
                           n3987);
   U8306 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_18_port, Z => 
                           n3993);
   U8307 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_17_port, Z => 
                           n3999);
   U8308 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_16_port, Z => 
                           n4005);
   U8309 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_15_port, Z => 
                           n4011);
   U8310 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_14_port, Z => 
                           n4017);
   U8311 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_13_port, Z => 
                           n4023);
   U8312 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_12_port, Z => 
                           n4029);
   U8313 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_3_port, Z => 
                           n4083);
   U8314 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_2_port, Z => 
                           n4089);
   U8315 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_1_port, Z => 
                           n4095);
   U8316 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_0_port, Z => 
                           n4101);
   U8317 : BUF_X1 port map( A => DataPath_i_RF_BUS_FROM_RF_CU_11_port, Z => 
                           n4035);
   U8318 : BUF_X1 port map( A => DataPath_ALUhw_BWISE_n70, Z => n2987);
   U8319 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_1_0_port, Z => 
                           n3405);
   U8320 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_1_0_port, Z => 
                           n3404);
   U8321 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_0_0_port, Z => 
                           n3293);
   U8322 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_0_0_port, Z => 
                           n3292);
   U8323 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_4_0_port, Z => 
                           n3741);
   U8324 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_4_0_port, Z => 
                           n3740);
   U8325 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_2_0_port, Z => 
                           n3517);
   U8326 : BUF_X1 port map( A => DataPath_RF_c_swin_masked_1bit_2_0_port, Z => 
                           n3516);
   U8327 : INV_X1 port map( A => n3268, ZN => n3280);
   U8328 : INV_X1 port map( A => n3267, ZN => n3279);
   U8329 : INV_X1 port map( A => n3268, ZN => n3283);
   U8330 : INV_X1 port map( A => n3268, ZN => n3282);
   U8331 : INV_X1 port map( A => n3268, ZN => n3281);
   U8332 : BUF_X1 port map( A => n8205, Z => n2256);
   U8333 : BUF_X1 port map( A => n8205, Z => n2257);
   U8334 : OR3_X1 port map( A1 => DataPath_RF_spill_address_ext_6_port, A2 => 
                           DataPath_RF_spill_address_ext_7_port, A3 => 
                           DataPath_RF_spill_address_ext_5_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n12);
   U8335 : NOR3_X1 port map( A1 => DataPath_RF_SPILLADDR_ENC_n15, A2 => 
                           DataPath_RF_spill_address_ext_10_port, A3 => n11443,
                           ZN => DataPath_RF_SPILLADDR_ENC_n14);
   U8336 : INV_X1 port map( A => DataPath_RF_SPILLADDR_ENC_n16, ZN => n11443);
   U8337 : NOR3_X1 port map( A1 => DataPath_RF_SPILLADDR_ENC_n22, A2 => 
                           DataPath_RF_spill_address_ext_1_port, A3 => 
                           DataPath_RF_spill_address_ext_0_port, ZN => 
                           DataPath_RF_spill_address_1_port);
   U8338 : AOI211_X1 port map( C1 => DataPath_RF_SPILLADDR_ENC_n23, C2 => 
                           DataPath_RF_SPILLADDR_ENC_n24, A => 
                           DataPath_RF_spill_address_ext_3_port, B => 
                           DataPath_RF_spill_address_ext_2_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n22);
   U8339 : NOR2_X1 port map( A1 => DataPath_RF_spill_address_ext_5_port, A2 => 
                           DataPath_RF_spill_address_ext_4_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n23);
   U8340 : NOR3_X1 port map( A1 => DataPath_RF_spill_address_ext_12_port, A2 =>
                           DataPath_RF_spill_address_ext_13_port, A3 => n11445,
                           ZN => DataPath_RF_SPILLADDR_ENC_n16);
   U8341 : INV_X1 port map( A => DataPath_RF_SPILLADDR_ENC_n21, ZN => n11445);
   U8342 : AOI21_X1 port map( B1 => DataPath_RF_SPILLADDR_ENC_n17, B2 => 
                           DataPath_RF_SPILLADDR_ENC_n18, A => 
                           DataPath_RF_SPILLADDR_ENC_n13, ZN => 
                           DataPath_RF_spill_address_2_port);
   U8343 : AOI21_X1 port map( B1 => DataPath_RF_SPILLADDR_ENC_n19, B2 => 
                           DataPath_RF_SPILLADDR_ENC_n20, A => 
                           DataPath_RF_spill_address_ext_4_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n17);
   U8344 : NOR3_X1 port map( A1 => DataPath_RF_spill_address_ext_5_port, A2 => 
                           DataPath_RF_spill_address_ext_7_port, A3 => 
                           DataPath_RF_spill_address_ext_6_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n18);
   U8345 : NOR2_X1 port map( A1 => DataPath_RF_spill_address_ext_10_port, A2 =>
                           DataPath_RF_SPILLADDR_ENC_n16, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n19);
   U8346 : NOR2_X1 port map( A1 => DataPath_RF_spill_address_ext_0_port, A2 => 
                           DataPath_RF_SPILLADDR_ENC_n28, ZN => 
                           DataPath_RF_spill_address_0_port);
   U8347 : AOI21_X1 port map( B1 => DataPath_RF_SPILLADDR_ENC_n29, B2 => n11435
                           , A => DataPath_RF_spill_address_ext_1_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n28);
   U8348 : INV_X1 port map( A => DataPath_RF_spill_address_ext_2_port, ZN => 
                           n11435);
   U8349 : OAI21_X1 port map( B1 => DataPath_RF_spill_address_ext_4_port, B2 =>
                           DataPath_RF_SPILLADDR_ENC_n30, A => n11436, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n29);
   U8350 : NOR3_X1 port map( A1 => DataPath_RF_spill_address_ext_11_port, A2 =>
                           DataPath_RF_spill_address_ext_9_port, A3 => 
                           DataPath_RF_spill_address_ext_8_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n20);
   U8351 : NOR2_X1 port map( A1 => DataPath_RF_spill_address_ext_15_port, A2 =>
                           DataPath_RF_spill_address_ext_14_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n21);
   U8352 : AOI21_X1 port map( B1 => DataPath_RF_SPILLADDR_ENC_n31, B2 => n11437
                           , A => DataPath_RF_spill_address_ext_5_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n30);
   U8353 : OAI21_X1 port map( B1 => DataPath_RF_spill_address_ext_8_port, B2 =>
                           DataPath_RF_SPILLADDR_ENC_n32, A => n11438, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n31);
   U8354 : AOI21_X1 port map( B1 => DataPath_RF_SPILLADDR_ENC_n33, B2 => n11441
                           , A => DataPath_RF_spill_address_ext_9_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n32);
   U8355 : OAI21_X1 port map( B1 => DataPath_RF_spill_address_ext_12_port, B2 
                           => DataPath_RF_SPILLADDR_ENC_n34, A => n11442, ZN =>
                           DataPath_RF_SPILLADDR_ENC_n33);
   U8356 : AOI21_X1 port map( B1 => DataPath_RF_spill_address_ext_15_port, B2 
                           => n11444, A => 
                           DataPath_RF_spill_address_ext_13_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n34);
   U8357 : INV_X1 port map( A => DataPath_RF_spill_address_ext_14_port, ZN => 
                           n11444);
   U8358 : BUF_X1 port map( A => n3845, Z => n3895);
   U8359 : BUF_X1 port map( A => n3845, Z => n3896);
   U8360 : BUF_X1 port map( A => n3844, Z => n3892);
   U8361 : BUF_X1 port map( A => n3845, Z => n3894);
   U8362 : BUF_X1 port map( A => n3844, Z => n3893);
   U8363 : BUF_X1 port map( A => n3846, Z => n3897);
   U8364 : NOR2_X1 port map( A1 => DataPath_i_DONE_FILL_EX, A2 => n12957, ZN =>
                           DRAMRF_READNOTWRITE_port);
   U8365 : OR4_X1 port map( A1 => DataPath_RF_spill_address_ext_0_port, A2 => 
                           DataPath_RF_spill_address_ext_1_port, A3 => 
                           DataPath_RF_spill_address_ext_2_port, A4 => 
                           DataPath_RF_spill_address_ext_3_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n13);
   U8366 : OAI211_X1 port map( C1 => DataPath_RF_SPILLADDR_ENC_n26, C2 => 
                           DataPath_RF_SPILLADDR_ENC_n27, A => n11439, B => 
                           n11440, ZN => DataPath_RF_SPILLADDR_ENC_n25);
   U8367 : NAND2_X1 port map( A1 => n11441, A2 => n11442, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n27);
   U8368 : NOR3_X1 port map( A1 => DataPath_RF_SPILLADDR_ENC_n21, A2 => 
                           DataPath_RF_spill_address_ext_13_port, A3 => 
                           DataPath_RF_spill_address_ext_12_port, ZN => 
                           DataPath_RF_SPILLADDR_ENC_n26);
   U8369 : BUF_X1 port map( A => n4154, Z => n4144);
   U8370 : BUF_X1 port map( A => n4153, Z => n4146);
   U8371 : BUF_X1 port map( A => n4154, Z => n4145);
   U8372 : BUF_X1 port map( A => n4153, Z => n4147);
   U8373 : BUF_X1 port map( A => n4154, Z => n4143);
   U8374 : BUF_X1 port map( A => n4152, Z => n4149);
   U8375 : BUF_X1 port map( A => n4152, Z => n4150);
   U8376 : BUF_X1 port map( A => n4153, Z => n4148);
   U8377 : INV_X1 port map( A => DataPath_RF_spill_address_ext_10_port, ZN => 
                           n11441);
   U8378 : INV_X1 port map( A => DataPath_RF_spill_address_ext_11_port, ZN => 
                           n11442);
   U8379 : INV_X1 port map( A => DataPath_RF_spill_address_ext_6_port, ZN => 
                           n11437);
   U8380 : INV_X1 port map( A => DataPath_RF_spill_address_ext_7_port, ZN => 
                           n11438);
   U8381 : INV_X1 port map( A => DataPath_RF_spill_address_ext_8_port, ZN => 
                           n11439);
   U8382 : INV_X1 port map( A => DataPath_RF_spill_address_ext_9_port, ZN => 
                           n11440);
   U8383 : INV_X1 port map( A => DataPath_WRF_CUhw_n142, ZN => 
                           DRAMRF_ADDRESS(3));
   U8384 : INV_X1 port map( A => DataPath_WRF_CUhw_n141, ZN => 
                           DRAMRF_ADDRESS(4));
   U8385 : INV_X1 port map( A => DataPath_WRF_CUhw_n140, ZN => 
                           DRAMRF_ADDRESS(5));
   U8386 : INV_X1 port map( A => DataPath_WRF_CUhw_n139, ZN => 
                           DRAMRF_ADDRESS(6));
   U8387 : INV_X1 port map( A => DataPath_WRF_CUhw_n138, ZN => 
                           DRAMRF_ADDRESS(7));
   U8388 : INV_X1 port map( A => DataPath_WRF_CUhw_n137, ZN => 
                           DRAMRF_ADDRESS(8));
   U8389 : INV_X1 port map( A => DataPath_WRF_CUhw_n136, ZN => 
                           DRAMRF_ADDRESS(9));
   U8390 : INV_X1 port map( A => DataPath_WRF_CUhw_n114, ZN => 
                           DRAMRF_ADDRESS(31));
   U8391 : INV_X1 port map( A => DataPath_WRF_CUhw_n145, ZN => 
                           DRAMRF_ADDRESS(0));
   U8392 : INV_X1 port map( A => DataPath_WRF_CUhw_n144, ZN => 
                           DRAMRF_ADDRESS(1));
   U8393 : INV_X1 port map( A => DataPath_WRF_CUhw_n143, ZN => 
                           DRAMRF_ADDRESS(2));
   U8394 : INV_X1 port map( A => DataPath_WRF_CUhw_n135, ZN => 
                           DRAMRF_ADDRESS(10));
   U8395 : INV_X1 port map( A => DataPath_WRF_CUhw_n134, ZN => 
                           DRAMRF_ADDRESS(11));
   U8396 : INV_X1 port map( A => DataPath_WRF_CUhw_n133, ZN => 
                           DRAMRF_ADDRESS(12));
   U8397 : INV_X1 port map( A => DataPath_WRF_CUhw_n132, ZN => 
                           DRAMRF_ADDRESS(13));
   U8398 : INV_X1 port map( A => DataPath_WRF_CUhw_n131, ZN => 
                           DRAMRF_ADDRESS(14));
   U8399 : INV_X1 port map( A => DataPath_WRF_CUhw_n130, ZN => 
                           DRAMRF_ADDRESS(15));
   U8400 : INV_X1 port map( A => DataPath_WRF_CUhw_n129, ZN => 
                           DRAMRF_ADDRESS(16));
   U8401 : INV_X1 port map( A => DataPath_WRF_CUhw_n128, ZN => 
                           DRAMRF_ADDRESS(17));
   U8402 : INV_X1 port map( A => DataPath_WRF_CUhw_n127, ZN => 
                           DRAMRF_ADDRESS(18));
   U8403 : INV_X1 port map( A => DataPath_WRF_CUhw_n126, ZN => 
                           DRAMRF_ADDRESS(19));
   U8404 : INV_X1 port map( A => DataPath_WRF_CUhw_n125, ZN => 
                           DRAMRF_ADDRESS(20));
   U8405 : INV_X1 port map( A => DataPath_WRF_CUhw_n124, ZN => 
                           DRAMRF_ADDRESS(21));
   U8406 : INV_X1 port map( A => DataPath_WRF_CUhw_n123, ZN => 
                           DRAMRF_ADDRESS(22));
   U8407 : INV_X1 port map( A => DataPath_WRF_CUhw_n122, ZN => 
                           DRAMRF_ADDRESS(23));
   U8408 : INV_X1 port map( A => DataPath_WRF_CUhw_n121, ZN => 
                           DRAMRF_ADDRESS(24));
   U8409 : INV_X1 port map( A => DataPath_WRF_CUhw_n120, ZN => 
                           DRAMRF_ADDRESS(25));
   U8410 : INV_X1 port map( A => DataPath_WRF_CUhw_n119, ZN => 
                           DRAMRF_ADDRESS(26));
   U8411 : INV_X1 port map( A => DataPath_WRF_CUhw_n118, ZN => 
                           DRAMRF_ADDRESS(27));
   U8412 : INV_X1 port map( A => DataPath_WRF_CUhw_n117, ZN => 
                           DRAMRF_ADDRESS(28));
   U8413 : INV_X1 port map( A => DataPath_WRF_CUhw_n116, ZN => 
                           DRAMRF_ADDRESS(29));
   U8414 : INV_X1 port map( A => DataPath_WRF_CUhw_n115, ZN => 
                           DRAMRF_ADDRESS(30));
   U8415 : INV_X1 port map( A => DataPath_RF_spill_address_ext_3_port, ZN => 
                           n11436);
   U8416 : BUF_X1 port map( A => n3846, Z => n3898);
   U8417 : BUF_X1 port map( A => n4152, Z => n4151);
   U8418 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n9, Z => n3203);
   U8419 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n9, Z => n3202);
   U8420 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n9, Z => n3201);
   U8421 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n8, Z => n3148);
   U8422 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n8, Z => n3147);
   U8423 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n8, Z => n3146);
   U8424 : BUF_X1 port map( A => n4255, Z => n4248);
   U8425 : BUF_X1 port map( A => n4254, Z => n4251);
   U8426 : BUF_X1 port map( A => n4255, Z => n4250);
   U8427 : BUF_X1 port map( A => n4255, Z => n4249);
   U8428 : BUF_X1 port map( A => n4254, Z => n4253);
   U8429 : BUF_X1 port map( A => n4254, Z => n4252);
   U8430 : BUF_X1 port map( A => n4256, Z => n4246);
   U8431 : BUF_X1 port map( A => n4256, Z => n4247);
   U8432 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n6, Z => n3047);
   U8433 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n6, Z => n3046);
   U8434 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n6, Z => n3045);
   U8435 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n7, Z => n3102);
   U8436 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n7, Z => n3101);
   U8437 : BUF_X1 port map( A => DataPath_RF_SELBLOCK_INLOC_n7, Z => n3100);
   U8438 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n330, A2 => 
                           DataPath_RF_RDPORT_SPILL_n331, ZN => 
                           DRAMRF_DATA_OUT(0));
   U8439 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n332, A2 => 
                           DataPath_RF_RDPORT_SPILL_n333, A3 => 
                           DataPath_RF_RDPORT_SPILL_n334, A4 => 
                           DataPath_RF_RDPORT_SPILL_n335, ZN => 
                           DataPath_RF_RDPORT_SPILL_n331);
   U8440 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n342, A2 => 
                           DataPath_RF_RDPORT_SPILL_n343, A3 => 
                           DataPath_RF_RDPORT_SPILL_n344, A4 => 
                           DataPath_RF_RDPORT_SPILL_n345, ZN => 
                           DataPath_RF_RDPORT_SPILL_n330);
   U8441 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_448_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_480_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n332);
   U8442 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n220, A2 => 
                           DataPath_RF_RDPORT_SPILL_n221, ZN => 
                           DRAMRF_DATA_OUT(1));
   U8443 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n222, A2 => 
                           DataPath_RF_RDPORT_SPILL_n223, A3 => 
                           DataPath_RF_RDPORT_SPILL_n224, A4 => 
                           DataPath_RF_RDPORT_SPILL_n225, ZN => 
                           DataPath_RF_RDPORT_SPILL_n221);
   U8444 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n226, A2 => 
                           DataPath_RF_RDPORT_SPILL_n227, A3 => 
                           DataPath_RF_RDPORT_SPILL_n228, A4 => 
                           DataPath_RF_RDPORT_SPILL_n229, ZN => 
                           DataPath_RF_RDPORT_SPILL_n220);
   U8445 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_449_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_481_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n222);
   U8446 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n110, A2 => 
                           DataPath_RF_RDPORT_SPILL_n111, ZN => 
                           DRAMRF_DATA_OUT(2));
   U8447 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n112, A2 => 
                           DataPath_RF_RDPORT_SPILL_n113, A3 => 
                           DataPath_RF_RDPORT_SPILL_n114, A4 => 
                           DataPath_RF_RDPORT_SPILL_n115, ZN => 
                           DataPath_RF_RDPORT_SPILL_n111);
   U8448 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n116, A2 => 
                           DataPath_RF_RDPORT_SPILL_n117, A3 => 
                           DataPath_RF_RDPORT_SPILL_n118, A4 => 
                           DataPath_RF_RDPORT_SPILL_n119, ZN => 
                           DataPath_RF_RDPORT_SPILL_n110);
   U8449 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_450_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_482_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n112);
   U8450 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n80, A2 => 
                           DataPath_RF_RDPORT_SPILL_n81, ZN => 
                           DRAMRF_DATA_OUT(3));
   U8451 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n82, A2 => 
                           DataPath_RF_RDPORT_SPILL_n83, A3 => 
                           DataPath_RF_RDPORT_SPILL_n84, A4 => 
                           DataPath_RF_RDPORT_SPILL_n85, ZN => 
                           DataPath_RF_RDPORT_SPILL_n81);
   U8452 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n86, A2 => 
                           DataPath_RF_RDPORT_SPILL_n87, A3 => 
                           DataPath_RF_RDPORT_SPILL_n88, A4 => 
                           DataPath_RF_RDPORT_SPILL_n89, ZN => 
                           DataPath_RF_RDPORT_SPILL_n80);
   U8453 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_451_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_483_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n82);
   U8454 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n70, A2 => 
                           DataPath_RF_RDPORT_SPILL_n71, ZN => 
                           DRAMRF_DATA_OUT(4));
   U8455 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n72, A2 => 
                           DataPath_RF_RDPORT_SPILL_n73, A3 => 
                           DataPath_RF_RDPORT_SPILL_n74, A4 => 
                           DataPath_RF_RDPORT_SPILL_n75, ZN => 
                           DataPath_RF_RDPORT_SPILL_n71);
   U8456 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n76, A2 => 
                           DataPath_RF_RDPORT_SPILL_n77, A3 => 
                           DataPath_RF_RDPORT_SPILL_n78, A4 => 
                           DataPath_RF_RDPORT_SPILL_n79, ZN => 
                           DataPath_RF_RDPORT_SPILL_n70);
   U8457 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_452_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_484_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n72);
   U8458 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n60, A2 => 
                           DataPath_RF_RDPORT_SPILL_n61, ZN => 
                           DRAMRF_DATA_OUT(5));
   U8459 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n62, A2 => 
                           DataPath_RF_RDPORT_SPILL_n63, A3 => 
                           DataPath_RF_RDPORT_SPILL_n64, A4 => 
                           DataPath_RF_RDPORT_SPILL_n65, ZN => 
                           DataPath_RF_RDPORT_SPILL_n61);
   U8460 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n66, A2 => 
                           DataPath_RF_RDPORT_SPILL_n67, A3 => 
                           DataPath_RF_RDPORT_SPILL_n68, A4 => 
                           DataPath_RF_RDPORT_SPILL_n69, ZN => 
                           DataPath_RF_RDPORT_SPILL_n60);
   U8461 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_453_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_485_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n62);
   U8462 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n50, A2 => 
                           DataPath_RF_RDPORT_SPILL_n51, ZN => 
                           DRAMRF_DATA_OUT(6));
   U8463 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n52, A2 => 
                           DataPath_RF_RDPORT_SPILL_n53, A3 => 
                           DataPath_RF_RDPORT_SPILL_n54, A4 => 
                           DataPath_RF_RDPORT_SPILL_n55, ZN => 
                           DataPath_RF_RDPORT_SPILL_n51);
   U8464 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n56, A2 => 
                           DataPath_RF_RDPORT_SPILL_n57, A3 => 
                           DataPath_RF_RDPORT_SPILL_n58, A4 => 
                           DataPath_RF_RDPORT_SPILL_n59, ZN => 
                           DataPath_RF_RDPORT_SPILL_n50);
   U8465 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_454_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_486_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n52);
   U8466 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n40, A2 => 
                           DataPath_RF_RDPORT_SPILL_n41, ZN => 
                           DRAMRF_DATA_OUT(7));
   U8467 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n42, A2 => 
                           DataPath_RF_RDPORT_SPILL_n43, A3 => 
                           DataPath_RF_RDPORT_SPILL_n44, A4 => 
                           DataPath_RF_RDPORT_SPILL_n45, ZN => 
                           DataPath_RF_RDPORT_SPILL_n41);
   U8468 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n46, A2 => 
                           DataPath_RF_RDPORT_SPILL_n47, A3 => 
                           DataPath_RF_RDPORT_SPILL_n48, A4 => 
                           DataPath_RF_RDPORT_SPILL_n49, ZN => 
                           DataPath_RF_RDPORT_SPILL_n40);
   U8469 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_455_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_487_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n42);
   U8470 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n30, A2 => 
                           DataPath_RF_RDPORT_SPILL_n31, ZN => 
                           DRAMRF_DATA_OUT(8));
   U8471 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n32, A2 => 
                           DataPath_RF_RDPORT_SPILL_n33, A3 => 
                           DataPath_RF_RDPORT_SPILL_n34, A4 => 
                           DataPath_RF_RDPORT_SPILL_n35, ZN => 
                           DataPath_RF_RDPORT_SPILL_n31);
   U8472 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n36, A2 => 
                           DataPath_RF_RDPORT_SPILL_n37, A3 => 
                           DataPath_RF_RDPORT_SPILL_n38, A4 => 
                           DataPath_RF_RDPORT_SPILL_n39, ZN => 
                           DataPath_RF_RDPORT_SPILL_n30);
   U8473 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_456_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_488_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n32);
   U8474 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n4, A2 => 
                           DataPath_RF_RDPORT_SPILL_n5, ZN => 
                           DRAMRF_DATA_OUT(9));
   U8475 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n6, A2 => 
                           DataPath_RF_RDPORT_SPILL_n7, A3 => 
                           DataPath_RF_RDPORT_SPILL_n8, A4 => 
                           DataPath_RF_RDPORT_SPILL_n9, ZN => 
                           DataPath_RF_RDPORT_SPILL_n5);
   U8476 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n18, A2 => 
                           DataPath_RF_RDPORT_SPILL_n19, A3 => 
                           DataPath_RF_RDPORT_SPILL_n20, A4 => 
                           DataPath_RF_RDPORT_SPILL_n21, ZN => 
                           DataPath_RF_RDPORT_SPILL_n4);
   U8477 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_457_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_489_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n6);
   U8478 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n320, A2 => 
                           DataPath_RF_RDPORT_SPILL_n321, ZN => 
                           DRAMRF_DATA_OUT(10));
   U8479 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n322, A2 => 
                           DataPath_RF_RDPORT_SPILL_n323, A3 => 
                           DataPath_RF_RDPORT_SPILL_n324, A4 => 
                           DataPath_RF_RDPORT_SPILL_n325, ZN => 
                           DataPath_RF_RDPORT_SPILL_n321);
   U8480 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n326, A2 => 
                           DataPath_RF_RDPORT_SPILL_n327, A3 => 
                           DataPath_RF_RDPORT_SPILL_n328, A4 => 
                           DataPath_RF_RDPORT_SPILL_n329, ZN => 
                           DataPath_RF_RDPORT_SPILL_n320);
   U8481 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_458_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_490_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n322);
   U8482 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n310, A2 => 
                           DataPath_RF_RDPORT_SPILL_n311, ZN => 
                           DRAMRF_DATA_OUT(11));
   U8483 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n312, A2 => 
                           DataPath_RF_RDPORT_SPILL_n313, A3 => 
                           DataPath_RF_RDPORT_SPILL_n314, A4 => 
                           DataPath_RF_RDPORT_SPILL_n315, ZN => 
                           DataPath_RF_RDPORT_SPILL_n311);
   U8484 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n316, A2 => 
                           DataPath_RF_RDPORT_SPILL_n317, A3 => 
                           DataPath_RF_RDPORT_SPILL_n318, A4 => 
                           DataPath_RF_RDPORT_SPILL_n319, ZN => 
                           DataPath_RF_RDPORT_SPILL_n310);
   U8485 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_459_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_491_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n312);
   U8486 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n300, A2 => 
                           DataPath_RF_RDPORT_SPILL_n301, ZN => 
                           DRAMRF_DATA_OUT(12));
   U8487 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n302, A2 => 
                           DataPath_RF_RDPORT_SPILL_n303, A3 => 
                           DataPath_RF_RDPORT_SPILL_n304, A4 => 
                           DataPath_RF_RDPORT_SPILL_n305, ZN => 
                           DataPath_RF_RDPORT_SPILL_n301);
   U8488 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n306, A2 => 
                           DataPath_RF_RDPORT_SPILL_n307, A3 => 
                           DataPath_RF_RDPORT_SPILL_n308, A4 => 
                           DataPath_RF_RDPORT_SPILL_n309, ZN => 
                           DataPath_RF_RDPORT_SPILL_n300);
   U8489 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_460_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_492_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n302);
   U8490 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n290, A2 => 
                           DataPath_RF_RDPORT_SPILL_n291, ZN => 
                           DRAMRF_DATA_OUT(13));
   U8491 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n292, A2 => 
                           DataPath_RF_RDPORT_SPILL_n293, A3 => 
                           DataPath_RF_RDPORT_SPILL_n294, A4 => 
                           DataPath_RF_RDPORT_SPILL_n295, ZN => 
                           DataPath_RF_RDPORT_SPILL_n291);
   U8492 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n296, A2 => 
                           DataPath_RF_RDPORT_SPILL_n297, A3 => 
                           DataPath_RF_RDPORT_SPILL_n298, A4 => 
                           DataPath_RF_RDPORT_SPILL_n299, ZN => 
                           DataPath_RF_RDPORT_SPILL_n290);
   U8493 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_461_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_493_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n292);
   U8494 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n280, A2 => 
                           DataPath_RF_RDPORT_SPILL_n281, ZN => 
                           DRAMRF_DATA_OUT(14));
   U8495 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n282, A2 => 
                           DataPath_RF_RDPORT_SPILL_n283, A3 => 
                           DataPath_RF_RDPORT_SPILL_n284, A4 => 
                           DataPath_RF_RDPORT_SPILL_n285, ZN => 
                           DataPath_RF_RDPORT_SPILL_n281);
   U8496 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n286, A2 => 
                           DataPath_RF_RDPORT_SPILL_n287, A3 => 
                           DataPath_RF_RDPORT_SPILL_n288, A4 => 
                           DataPath_RF_RDPORT_SPILL_n289, ZN => 
                           DataPath_RF_RDPORT_SPILL_n280);
   U8497 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_462_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_494_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n282);
   U8498 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n270, A2 => 
                           DataPath_RF_RDPORT_SPILL_n271, ZN => 
                           DRAMRF_DATA_OUT(15));
   U8499 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n272, A2 => 
                           DataPath_RF_RDPORT_SPILL_n273, A3 => 
                           DataPath_RF_RDPORT_SPILL_n274, A4 => 
                           DataPath_RF_RDPORT_SPILL_n275, ZN => 
                           DataPath_RF_RDPORT_SPILL_n271);
   U8500 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n276, A2 => 
                           DataPath_RF_RDPORT_SPILL_n277, A3 => 
                           DataPath_RF_RDPORT_SPILL_n278, A4 => 
                           DataPath_RF_RDPORT_SPILL_n279, ZN => 
                           DataPath_RF_RDPORT_SPILL_n270);
   U8501 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_463_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_495_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n272);
   U8502 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n260, A2 => 
                           DataPath_RF_RDPORT_SPILL_n261, ZN => 
                           DRAMRF_DATA_OUT(16));
   U8503 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n262, A2 => 
                           DataPath_RF_RDPORT_SPILL_n263, A3 => 
                           DataPath_RF_RDPORT_SPILL_n264, A4 => 
                           DataPath_RF_RDPORT_SPILL_n265, ZN => 
                           DataPath_RF_RDPORT_SPILL_n261);
   U8504 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n266, A2 => 
                           DataPath_RF_RDPORT_SPILL_n267, A3 => 
                           DataPath_RF_RDPORT_SPILL_n268, A4 => 
                           DataPath_RF_RDPORT_SPILL_n269, ZN => 
                           DataPath_RF_RDPORT_SPILL_n260);
   U8505 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_464_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_496_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n262);
   U8506 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n250, A2 => 
                           DataPath_RF_RDPORT_SPILL_n251, ZN => 
                           DRAMRF_DATA_OUT(17));
   U8507 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n252, A2 => 
                           DataPath_RF_RDPORT_SPILL_n253, A3 => 
                           DataPath_RF_RDPORT_SPILL_n254, A4 => 
                           DataPath_RF_RDPORT_SPILL_n255, ZN => 
                           DataPath_RF_RDPORT_SPILL_n251);
   U8508 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n256, A2 => 
                           DataPath_RF_RDPORT_SPILL_n257, A3 => 
                           DataPath_RF_RDPORT_SPILL_n258, A4 => 
                           DataPath_RF_RDPORT_SPILL_n259, ZN => 
                           DataPath_RF_RDPORT_SPILL_n250);
   U8509 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_465_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_497_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n252);
   U8510 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n240, A2 => 
                           DataPath_RF_RDPORT_SPILL_n241, ZN => 
                           DRAMRF_DATA_OUT(18));
   U8511 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n242, A2 => 
                           DataPath_RF_RDPORT_SPILL_n243, A3 => 
                           DataPath_RF_RDPORT_SPILL_n244, A4 => 
                           DataPath_RF_RDPORT_SPILL_n245, ZN => 
                           DataPath_RF_RDPORT_SPILL_n241);
   U8512 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n246, A2 => 
                           DataPath_RF_RDPORT_SPILL_n247, A3 => 
                           DataPath_RF_RDPORT_SPILL_n248, A4 => 
                           DataPath_RF_RDPORT_SPILL_n249, ZN => 
                           DataPath_RF_RDPORT_SPILL_n240);
   U8513 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_466_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_498_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n242);
   U8514 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n230, A2 => 
                           DataPath_RF_RDPORT_SPILL_n231, ZN => 
                           DRAMRF_DATA_OUT(19));
   U8515 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n232, A2 => 
                           DataPath_RF_RDPORT_SPILL_n233, A3 => 
                           DataPath_RF_RDPORT_SPILL_n234, A4 => 
                           DataPath_RF_RDPORT_SPILL_n235, ZN => 
                           DataPath_RF_RDPORT_SPILL_n231);
   U8516 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n236, A2 => 
                           DataPath_RF_RDPORT_SPILL_n237, A3 => 
                           DataPath_RF_RDPORT_SPILL_n238, A4 => 
                           DataPath_RF_RDPORT_SPILL_n239, ZN => 
                           DataPath_RF_RDPORT_SPILL_n230);
   U8517 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_467_port,
                           A2 => n3006, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_499_port, B2 => 
                           n3009, ZN => DataPath_RF_RDPORT_SPILL_n232);
   U8518 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n210, A2 => 
                           DataPath_RF_RDPORT_SPILL_n211, ZN => 
                           DRAMRF_DATA_OUT(20));
   U8519 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n212, A2 => 
                           DataPath_RF_RDPORT_SPILL_n213, A3 => 
                           DataPath_RF_RDPORT_SPILL_n214, A4 => 
                           DataPath_RF_RDPORT_SPILL_n215, ZN => 
                           DataPath_RF_RDPORT_SPILL_n211);
   U8520 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n216, A2 => 
                           DataPath_RF_RDPORT_SPILL_n217, A3 => 
                           DataPath_RF_RDPORT_SPILL_n218, A4 => 
                           DataPath_RF_RDPORT_SPILL_n219, ZN => 
                           DataPath_RF_RDPORT_SPILL_n210);
   U8521 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_468_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_500_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n212);
   U8522 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n200, A2 => 
                           DataPath_RF_RDPORT_SPILL_n201, ZN => 
                           DRAMRF_DATA_OUT(21));
   U8523 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n202, A2 => 
                           DataPath_RF_RDPORT_SPILL_n203, A3 => 
                           DataPath_RF_RDPORT_SPILL_n204, A4 => 
                           DataPath_RF_RDPORT_SPILL_n205, ZN => 
                           DataPath_RF_RDPORT_SPILL_n201);
   U8524 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n206, A2 => 
                           DataPath_RF_RDPORT_SPILL_n207, A3 => 
                           DataPath_RF_RDPORT_SPILL_n208, A4 => 
                           DataPath_RF_RDPORT_SPILL_n209, ZN => 
                           DataPath_RF_RDPORT_SPILL_n200);
   U8525 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_469_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_501_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n202);
   U8526 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n190, A2 => 
                           DataPath_RF_RDPORT_SPILL_n191, ZN => 
                           DRAMRF_DATA_OUT(22));
   U8527 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n192, A2 => 
                           DataPath_RF_RDPORT_SPILL_n193, A3 => 
                           DataPath_RF_RDPORT_SPILL_n194, A4 => 
                           DataPath_RF_RDPORT_SPILL_n195, ZN => 
                           DataPath_RF_RDPORT_SPILL_n191);
   U8528 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n196, A2 => 
                           DataPath_RF_RDPORT_SPILL_n197, A3 => 
                           DataPath_RF_RDPORT_SPILL_n198, A4 => 
                           DataPath_RF_RDPORT_SPILL_n199, ZN => 
                           DataPath_RF_RDPORT_SPILL_n190);
   U8529 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_470_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_502_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n192);
   U8530 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n180, A2 => 
                           DataPath_RF_RDPORT_SPILL_n181, ZN => 
                           DRAMRF_DATA_OUT(23));
   U8531 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n182, A2 => 
                           DataPath_RF_RDPORT_SPILL_n183, A3 => 
                           DataPath_RF_RDPORT_SPILL_n184, A4 => 
                           DataPath_RF_RDPORT_SPILL_n185, ZN => 
                           DataPath_RF_RDPORT_SPILL_n181);
   U8532 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n186, A2 => 
                           DataPath_RF_RDPORT_SPILL_n187, A3 => 
                           DataPath_RF_RDPORT_SPILL_n188, A4 => 
                           DataPath_RF_RDPORT_SPILL_n189, ZN => 
                           DataPath_RF_RDPORT_SPILL_n180);
   U8533 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_471_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_503_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n182);
   U8534 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n170, A2 => 
                           DataPath_RF_RDPORT_SPILL_n171, ZN => 
                           DRAMRF_DATA_OUT(24));
   U8535 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n172, A2 => 
                           DataPath_RF_RDPORT_SPILL_n173, A3 => 
                           DataPath_RF_RDPORT_SPILL_n174, A4 => 
                           DataPath_RF_RDPORT_SPILL_n175, ZN => 
                           DataPath_RF_RDPORT_SPILL_n171);
   U8536 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n176, A2 => 
                           DataPath_RF_RDPORT_SPILL_n177, A3 => 
                           DataPath_RF_RDPORT_SPILL_n178, A4 => 
                           DataPath_RF_RDPORT_SPILL_n179, ZN => 
                           DataPath_RF_RDPORT_SPILL_n170);
   U8537 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_472_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_504_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n172);
   U8538 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n160, A2 => 
                           DataPath_RF_RDPORT_SPILL_n161, ZN => 
                           DRAMRF_DATA_OUT(25));
   U8539 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n162, A2 => 
                           DataPath_RF_RDPORT_SPILL_n163, A3 => 
                           DataPath_RF_RDPORT_SPILL_n164, A4 => 
                           DataPath_RF_RDPORT_SPILL_n165, ZN => 
                           DataPath_RF_RDPORT_SPILL_n161);
   U8540 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n166, A2 => 
                           DataPath_RF_RDPORT_SPILL_n167, A3 => 
                           DataPath_RF_RDPORT_SPILL_n168, A4 => 
                           DataPath_RF_RDPORT_SPILL_n169, ZN => 
                           DataPath_RF_RDPORT_SPILL_n160);
   U8541 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_473_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_505_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n162);
   U8542 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n150, A2 => 
                           DataPath_RF_RDPORT_SPILL_n151, ZN => 
                           DRAMRF_DATA_OUT(26));
   U8543 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n152, A2 => 
                           DataPath_RF_RDPORT_SPILL_n153, A3 => 
                           DataPath_RF_RDPORT_SPILL_n154, A4 => 
                           DataPath_RF_RDPORT_SPILL_n155, ZN => 
                           DataPath_RF_RDPORT_SPILL_n151);
   U8544 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n156, A2 => 
                           DataPath_RF_RDPORT_SPILL_n157, A3 => 
                           DataPath_RF_RDPORT_SPILL_n158, A4 => 
                           DataPath_RF_RDPORT_SPILL_n159, ZN => 
                           DataPath_RF_RDPORT_SPILL_n150);
   U8545 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_474_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_506_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n152);
   U8546 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n140, A2 => 
                           DataPath_RF_RDPORT_SPILL_n141, ZN => 
                           DRAMRF_DATA_OUT(27));
   U8547 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n142, A2 => 
                           DataPath_RF_RDPORT_SPILL_n143, A3 => 
                           DataPath_RF_RDPORT_SPILL_n144, A4 => 
                           DataPath_RF_RDPORT_SPILL_n145, ZN => 
                           DataPath_RF_RDPORT_SPILL_n141);
   U8548 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n146, A2 => 
                           DataPath_RF_RDPORT_SPILL_n147, A3 => 
                           DataPath_RF_RDPORT_SPILL_n148, A4 => 
                           DataPath_RF_RDPORT_SPILL_n149, ZN => 
                           DataPath_RF_RDPORT_SPILL_n140);
   U8549 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_475_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_507_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n142);
   U8550 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n130, A2 => 
                           DataPath_RF_RDPORT_SPILL_n131, ZN => 
                           DRAMRF_DATA_OUT(28));
   U8551 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n132, A2 => 
                           DataPath_RF_RDPORT_SPILL_n133, A3 => 
                           DataPath_RF_RDPORT_SPILL_n134, A4 => 
                           DataPath_RF_RDPORT_SPILL_n135, ZN => 
                           DataPath_RF_RDPORT_SPILL_n131);
   U8552 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n136, A2 => 
                           DataPath_RF_RDPORT_SPILL_n137, A3 => 
                           DataPath_RF_RDPORT_SPILL_n138, A4 => 
                           DataPath_RF_RDPORT_SPILL_n139, ZN => 
                           DataPath_RF_RDPORT_SPILL_n130);
   U8553 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_476_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_508_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n132);
   U8554 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n120, A2 => 
                           DataPath_RF_RDPORT_SPILL_n121, ZN => 
                           DRAMRF_DATA_OUT(29));
   U8555 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n122, A2 => 
                           DataPath_RF_RDPORT_SPILL_n123, A3 => 
                           DataPath_RF_RDPORT_SPILL_n124, A4 => 
                           DataPath_RF_RDPORT_SPILL_n125, ZN => 
                           DataPath_RF_RDPORT_SPILL_n121);
   U8556 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n126, A2 => 
                           DataPath_RF_RDPORT_SPILL_n127, A3 => 
                           DataPath_RF_RDPORT_SPILL_n128, A4 => 
                           DataPath_RF_RDPORT_SPILL_n129, ZN => 
                           DataPath_RF_RDPORT_SPILL_n120);
   U8557 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_477_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_509_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n122);
   U8558 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n100, A2 => 
                           DataPath_RF_RDPORT_SPILL_n101, ZN => 
                           DRAMRF_DATA_OUT(30));
   U8559 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n102, A2 => 
                           DataPath_RF_RDPORT_SPILL_n103, A3 => 
                           DataPath_RF_RDPORT_SPILL_n104, A4 => 
                           DataPath_RF_RDPORT_SPILL_n105, ZN => 
                           DataPath_RF_RDPORT_SPILL_n101);
   U8560 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n106, A2 => 
                           DataPath_RF_RDPORT_SPILL_n107, A3 => 
                           DataPath_RF_RDPORT_SPILL_n108, A4 => 
                           DataPath_RF_RDPORT_SPILL_n109, ZN => 
                           DataPath_RF_RDPORT_SPILL_n100);
   U8561 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_478_port,
                           A2 => n3007, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_510_port, B2 => 
                           n3010, ZN => DataPath_RF_RDPORT_SPILL_n102);
   U8562 : OR2_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n90, A2 => 
                           DataPath_RF_RDPORT_SPILL_n91, ZN => 
                           DRAMRF_DATA_OUT(31));
   U8563 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n92, A2 => 
                           DataPath_RF_RDPORT_SPILL_n93, A3 => 
                           DataPath_RF_RDPORT_SPILL_n94, A4 => 
                           DataPath_RF_RDPORT_SPILL_n95, ZN => 
                           DataPath_RF_RDPORT_SPILL_n91);
   U8564 : NAND4_X1 port map( A1 => DataPath_RF_RDPORT_SPILL_n96, A2 => 
                           DataPath_RF_RDPORT_SPILL_n97, A3 => 
                           DataPath_RF_RDPORT_SPILL_n98, A4 => 
                           DataPath_RF_RDPORT_SPILL_n99, ZN => 
                           DataPath_RF_RDPORT_SPILL_n90);
   U8565 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_479_port,
                           A2 => n3008, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_511_port, B2 => 
                           n3011, ZN => DataPath_RF_RDPORT_SPILL_n92);
   U8567 : MUX2_X1 port map( A => DataPath_i_PIPLIN_A_12_port, B => 
                           DataPath_i_PIPLIN_IN1_12_port, S => n2150, Z => 
                           n1934);
   U8568 : MUX2_X1 port map( A => DataPath_i_PIPLIN_A_13_port, B => 
                           DataPath_i_PIPLIN_IN1_13_port, S => n2151, Z => 
                           n1935);
   U8569 : NOR2_X1 port map( A1 => n318, A2 => CU_I_n108, ZN => n4451);
   U8570 : AOI222_X1 port map( A1 => n270, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N140_port, B2 => n3262, C1 => n407
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n114);
   U8571 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_31_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_31_port, ZN => 
                           DataPath_WRF_CUhw_N140_port);
   U8572 : AOI222_X1 port map( A1 => n267, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N139_port, B2 => n3262, C1 => n387
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n115);
   U8573 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_30_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_30_port, ZN => 
                           DataPath_WRF_CUhw_N139_port);
   U8574 : AOI222_X1 port map( A1 => n283, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N134_port, B2 => n3263, C1 => n388
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n120);
   U8575 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_25_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_25_port, ZN => 
                           DataPath_WRF_CUhw_N134_port);
   U8576 : AOI222_X1 port map( A1 => n284, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N135_port, B2 => n3263, C1 => n389
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n119);
   U8577 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_26_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_26_port, ZN => 
                           DataPath_WRF_CUhw_N135_port);
   U8578 : AOI222_X1 port map( A1 => n268, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N138_port, B2 => n3262, C1 => n390
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n116);
   U8579 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_29_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_29_port, ZN => 
                           DataPath_WRF_CUhw_N138_port);
   U8580 : AOI222_X1 port map( A1 => n269, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N137_port, B2 => n3262, C1 => n391
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n117);
   U8581 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_28_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_28_port, ZN => 
                           DataPath_WRF_CUhw_N137_port);
   U8582 : AOI222_X1 port map( A1 => n285, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N136_port, B2 => n3263, C1 => n392
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n118);
   U8583 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_27_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_27_port, ZN => 
                           DataPath_WRF_CUhw_N136_port);
   U8584 : AOI222_X1 port map( A1 => n286, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N126_port, B2 => n3264, C1 => n393
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n128);
   U8585 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_17_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_17_port, ZN => 
                           DataPath_WRF_CUhw_N126_port);
   U8586 : AOI222_X1 port map( A1 => n287, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N127_port, B2 => n3263, C1 => n394
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n127);
   U8587 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_18_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_18_port, ZN => 
                           DataPath_WRF_CUhw_N127_port);
   U8588 : AOI222_X1 port map( A1 => n288, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N128_port, B2 => n3263, C1 => n395
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n126);
   U8589 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_19_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_19_port, ZN => 
                           DataPath_WRF_CUhw_N128_port);
   U8590 : AOI222_X1 port map( A1 => n289, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N129_port, B2 => n3263, C1 => n396
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n125);
   U8591 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_20_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_20_port, ZN => 
                           DataPath_WRF_CUhw_N129_port);
   U8592 : AOI222_X1 port map( A1 => n290, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N130_port, B2 => n3263, C1 => n397
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n124);
   U8593 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_21_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_21_port, ZN => 
                           DataPath_WRF_CUhw_N130_port);
   U8594 : AOI222_X1 port map( A1 => n291, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N131_port, B2 => n3263, C1 => n398
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n123);
   U8595 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_22_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_22_port, ZN => 
                           DataPath_WRF_CUhw_N131_port);
   U8596 : AOI222_X1 port map( A1 => n292, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N132_port, B2 => n3263, C1 => n399
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n122);
   U8597 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_23_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_23_port, ZN => 
                           DataPath_WRF_CUhw_N132_port);
   U8598 : AOI222_X1 port map( A1 => n293, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N133_port, B2 => n3263, C1 => n400
                           , C2 => n2476, ZN => DataPath_WRF_CUhw_n121);
   U8599 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_24_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_24_port, ZN => 
                           DataPath_WRF_CUhw_N133_port);
   U8600 : NAND2_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_state_1_port, 
                           A2 => n12950, ZN => n12957);
   U8601 : NAND2_X1 port map( A1 => n4129, A2 => i_ALU_OP_4_port, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n597);
   U8602 : NOR2_X1 port map( A1 => n4155, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n35);
   U8603 : AOI21_X1 port map( B1 => i_ALU_OP_3_port, B2 => i_ALU_OP_4_port, A 
                           => n11539, ZN => DataPath_ALUhw_SHIFTER_HW_n639);
   U8604 : NAND2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_state_1_port,
                           A2 => DataPath_RF_PUSH_ADDRGEN_n22, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n32);
   U8605 : NAND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_30_port, A2 => 
                           n1987, ZN => n2127);
   U8606 : NAND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_30_port, A2 => 
                           n1989, ZN => n2128);
   U8607 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_18_port, A2 => 
                           n1958, ZN => n1936);
   U8608 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_19_port, A2 => 
                           n1936, ZN => n1937);
   U8609 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_20_port, A2 => 
                           n1937, ZN => n1938);
   U8610 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_21_port, A2 => 
                           n1938, ZN => n1939);
   U8611 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_22_port, A2 => 
                           n1939, ZN => n1940);
   U8612 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_20_port, A2 => 
                           n1976, ZN => n1941);
   U8613 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_21_port, A2 => 
                           n1941, ZN => n1942);
   U8614 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_22_port, A2 => 
                           n1942, ZN => n1943);
   U8615 : OR2_X1 port map( A1 => n1855, A2 => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_3_port);
   U8616 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_3_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_3_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_4_port);
   U8617 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_4_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_4_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_5_port);
   U8618 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_5_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_5_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_6_port);
   U8619 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_6_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_6_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_7_port);
   U8620 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_7_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_7_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_8_port);
   U8621 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_8_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_8_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_9_port);
   U8622 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_9_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_9_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_10_port);
   U8623 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_10_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_10_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_11_port);
   U8624 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_11_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_11_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_12_port);
   U8625 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_12_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_12_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_13_port);
   U8626 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_13_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_13_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_14_port);
   U8627 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_14_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_14_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_15_port);
   U8628 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_15_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_15_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_16_port);
   U8629 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_16_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_16_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_17_port);
   U8630 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_17_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_17_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_18_port);
   U8631 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_18_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_18_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_19_port);
   U8632 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_19_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_19_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_20_port);
   U8633 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_20_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_20_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_21_port);
   U8634 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_21_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_21_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_22_port);
   U8635 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_22_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_22_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_23_port);
   U8636 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_23_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_23_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_24_port);
   U8637 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_24_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_24_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_25_port);
   U8638 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_25_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_25_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_26_port);
   U8639 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_26_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_26_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_27_port);
   U8640 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_27_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_27_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_28_port);
   U8641 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_28_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_28_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_29_port);
   U8642 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_29_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_29_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_30_port);
   U8643 : BUF_X1 port map( A => DataPath_RF_n10, Z => n3899);
   U8644 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_4_port, A2 => 
                           n1955, ZN => n1944);
   U8645 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_5_port, A2 => 
                           n1944, ZN => n1945);
   U8646 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_6_port, A2 => 
                           n1945, ZN => n1946);
   U8647 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_7_port, A2 => 
                           n1946, ZN => n1947);
   U8648 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_8_port, A2 => 
                           n1947, ZN => n1948);
   U8649 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_9_port, A2 => 
                           n1948, ZN => n1949);
   U8650 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_10_port, A2 => 
                           n1949, ZN => n1950);
   U8651 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_11_port, A2 => 
                           n1950, ZN => n1951);
   U8652 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_12_port, A2 => 
                           n1951, ZN => n1952);
   U8653 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_13_port, A2 => 
                           n1952, ZN => n1953);
   U8654 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_14_port, A2 => 
                           n1953, ZN => n1954);
   U8655 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_3_port, A2 => 
                           n1991, ZN => n1955);
   U8656 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_15_port, A2 => 
                           n1954, ZN => n1956);
   U8657 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_16_port, A2 => 
                           n1956, ZN => n1957);
   U8658 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_17_port, A2 => 
                           n1957, ZN => n1958);
   U8659 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_4_port, A2 => 
                           n1978, ZN => n1959);
   U8660 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_5_port, A2 => 
                           n1959, ZN => n1960);
   U8661 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_6_port, A2 => 
                           n1960, ZN => n1961);
   U8662 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_7_port, A2 => 
                           n1961, ZN => n1962);
   U8663 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_8_port, A2 => 
                           n1962, ZN => n1963);
   U8664 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_9_port, A2 => 
                           n1963, ZN => n1964);
   U8665 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_10_port, A2 => 
                           n1964, ZN => n1965);
   U8666 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_11_port, A2 => 
                           n1965, ZN => n1966);
   U8667 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_12_port, A2 => 
                           n1966, ZN => n1967);
   U8668 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_13_port, A2 => 
                           n1967, ZN => n1968);
   U8669 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_14_port, A2 => 
                           n1968, ZN => n1969);
   U8670 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_15_port, A2 => 
                           n1969, ZN => n1970);
   U8671 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_23_port, A2 => 
                           n1940, ZN => n1971);
   U8672 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_16_port, A2 => 
                           n1970, ZN => n1972);
   U8673 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_17_port, A2 => 
                           n1972, ZN => n1973);
   U8674 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_24_port, A2 => 
                           n1971, ZN => n1974);
   U8675 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_18_port, A2 => 
                           n1973, ZN => n1975);
   U8676 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_19_port, A2 => 
                           n1975, ZN => n1976);
   U8677 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_25_port, A2 => 
                           n1974, ZN => n1977);
   U8678 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_3_port, A2 => 
                           n1990, ZN => n1978);
   U8679 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_26_port, A2 => 
                           n1977, ZN => n1979);
   U8680 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_23_port, A2 => 
                           n1943, ZN => n1980);
   U8681 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_27_port, A2 => 
                           n1979, ZN => n1981);
   U8682 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_24_port, A2 => 
                           n1980, ZN => n1982);
   U8683 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_25_port, A2 => 
                           n1982, ZN => n1983);
   U8684 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_28_port, A2 => 
                           n1981, ZN => n1984);
   U8685 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_26_port, A2 => 
                           n1983, ZN => n1985);
   U8686 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_27_port, A2 => 
                           n1985, ZN => n1986);
   U8687 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_29_port, A2 => 
                           n1984, ZN => n1987);
   U8688 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_28_port, A2 => 
                           n1986, ZN => n1988);
   U8689 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_29_port, A2 => 
                           n1988, ZN => n1989);
   U8690 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_N217, A2 => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => n1990);
   U8691 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_N26_port, A2 => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => n1991);
   U8692 : OR2_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_30_port, A2 => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_30_port, ZN => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_31_port);
   U8693 : INV_X1 port map( A => n14258, ZN => n8675);
   U8694 : AOI22_X1 port map( A1 => n343, A2 => n1895, B1 => 
                           DRAM_ADDRESS_16_port, B2 => n8323, ZN => n14258);
   U8695 : INV_X1 port map( A => n14256, ZN => n8677);
   U8696 : AOI22_X1 port map( A1 => n1770, A2 => n1895, B1 => 
                           DRAM_ADDRESS_14_port, B2 => n8323, ZN => n14256);
   U8697 : INV_X1 port map( A => n14255, ZN => n8678);
   U8698 : AOI22_X1 port map( A1 => n1771, A2 => n1895, B1 => 
                           DRAM_ADDRESS_13_port, B2 => n8323, ZN => n14255);
   U8699 : INV_X1 port map( A => n14257, ZN => n8676);
   U8700 : AOI22_X1 port map( A1 => n344, A2 => n1895, B1 => 
                           DRAM_ADDRESS_15_port, B2 => n8323, ZN => n14257);
   U8701 : INV_X1 port map( A => n14254, ZN => n8679);
   U8702 : AOI22_X1 port map( A1 => n345, A2 => n1895, B1 => 
                           DRAM_ADDRESS_12_port, B2 => n8323, ZN => n14254);
   U8703 : INV_X1 port map( A => n14253, ZN => n8680);
   U8704 : AOI22_X1 port map( A1 => n346, A2 => n1895, B1 => 
                           DRAM_ADDRESS_11_port, B2 => n8323, ZN => n14253);
   U8705 : INV_X1 port map( A => n14252, ZN => n8681);
   U8706 : AOI22_X1 port map( A1 => n377, A2 => n1895, B1 => 
                           DRAM_ADDRESS_10_port, B2 => n8323, ZN => n14252);
   U8707 : INV_X1 port map( A => n14251, ZN => n8682);
   U8708 : AOI22_X1 port map( A1 => n378, A2 => n1895, B1 => 
                           DRAM_ADDRESS_9_port, B2 => n8323, ZN => n14251);
   U8709 : AOI222_X1 port map( A1 => n294, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N125_port, B2 => n3264, C1 => n401
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n129);
   U8710 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_16_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_16_port, ZN => 
                           DataPath_WRF_CUhw_N125_port);
   U8711 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17107, C1 => 
                           DataPath_LDSTR_n66, C2 => n17098, A => 
                           DataPath_LDSTR_n77, ZN => DRAM_DATA_OUT_7_port);
   U8712 : AOI22_X1 port map( A1 => n11350, A2 => DataPath_LDSTR_n68, B1 => 
                           n11374, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n77);
   U8713 : INV_X1 port map( A => n17084, ZN => n11374);
   U8714 : AOI22_X1 port map( A1 => DRAM_DATA_IN(7), A2 => n4118, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_7_port, B2 => n4119, 
                           ZN => n17084);
   U8715 : NOR2_X1 port map( A1 => DRAM_READY, A2 => n11582, ZN => CU_I_n71);
   U8716 : INV_X1 port map( A => DRAM_ISSUE_port, ZN => n11582);
   U8717 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17083, C1 => 
                           DataPath_LDSTR_n66, C2 => n17106, A => 
                           DataPath_LDSTR_n82, ZN => DRAM_DATA_OUT_0_port);
   U8718 : AOI22_X1 port map( A1 => n11364, A2 => DataPath_LDSTR_n68, B1 => 
                           n11381, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n82);
   U8719 : INV_X1 port map( A => n17113, ZN => n11381);
   U8720 : AOI22_X1 port map( A1 => DRAM_DATA_IN(0), A2 => i_DATAMEM_RM, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_0_port, B2 => n4127, 
                           ZN => n17113);
   U8721 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17112, C1 => 
                           DataPath_LDSTR_n66, C2 => n17104, A => 
                           DataPath_LDSTR_n81, ZN => DRAM_DATA_OUT_2_port);
   U8722 : AOI22_X1 port map( A1 => n11360, A2 => DataPath_LDSTR_n68, B1 => 
                           n11379, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n81);
   U8723 : INV_X1 port map( A => n17091, ZN => n11379);
   U8724 : AOI22_X1 port map( A1 => DRAM_DATA_IN(2), A2 => i_DATAMEM_RM, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_2_port, B2 => n4121, 
                           ZN => n17091);
   U8725 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17111, C1 => 
                           DataPath_LDSTR_n66, C2 => n17103, A => 
                           DataPath_LDSTR_n76, ZN => DRAM_DATA_OUT_3_port);
   U8726 : AOI22_X1 port map( A1 => n11358, A2 => DataPath_LDSTR_n68, B1 => 
                           n11378, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n76);
   U8727 : INV_X1 port map( A => n17088, ZN => n11378);
   U8728 : AOI22_X1 port map( A1 => DRAM_DATA_IN(3), A2 => n4118, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_3_port, B2 => n4120, 
                           ZN => n17088);
   U8729 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17110, C1 => 
                           DataPath_LDSTR_n66, C2 => n17101, A => 
                           DataPath_LDSTR_n75, ZN => DRAM_DATA_OUT_4_port);
   U8730 : AOI22_X1 port map( A1 => n11356, A2 => DataPath_LDSTR_n68, B1 => 
                           n11377, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n75);
   U8731 : INV_X1 port map( A => n17087, ZN => n11377);
   U8732 : AOI22_X1 port map( A1 => DRAM_DATA_IN(4), A2 => n4118, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_4_port, B2 => n4120, 
                           ZN => n17087);
   U8733 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17109, C1 => 
                           DataPath_LDSTR_n66, C2 => n17100, A => 
                           DataPath_LDSTR_n74, ZN => DRAM_DATA_OUT_5_port);
   U8734 : AOI22_X1 port map( A1 => n11354, A2 => DataPath_LDSTR_n68, B1 => 
                           n11376, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n74);
   U8735 : INV_X1 port map( A => n17086, ZN => n11376);
   U8736 : AOI22_X1 port map( A1 => DRAM_DATA_IN(5), A2 => n4118, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_5_port, B2 => n4120, 
                           ZN => n17086);
   U8737 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17108, C1 => 
                           DataPath_LDSTR_n66, C2 => n17099, A => 
                           DataPath_LDSTR_n73, ZN => DRAM_DATA_OUT_6_port);
   U8738 : AOI22_X1 port map( A1 => n11352, A2 => DataPath_LDSTR_n68, B1 => 
                           n11375, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n73);
   U8739 : INV_X1 port map( A => n17085, ZN => n11375);
   U8740 : AOI22_X1 port map( A1 => DRAM_DATA_IN(6), A2 => n4118, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_6_port, B2 => n4119, 
                           ZN => n17085);
   U8741 : OAI221_X1 port map( B1 => DataPath_LDSTR_n65, B2 => n17082, C1 => 
                           DataPath_LDSTR_n66, C2 => n17105, A => 
                           DataPath_LDSTR_n67, ZN => DRAM_DATA_OUT_1_port);
   U8742 : AOI22_X1 port map( A1 => n11362, A2 => DataPath_LDSTR_n68, B1 => 
                           n11380, B2 => DataPath_LDSTR_n69, ZN => 
                           DataPath_LDSTR_n67);
   U8743 : INV_X1 port map( A => n17102, ZN => n11380);
   U8744 : AOI22_X1 port map( A1 => DRAM_DATA_IN(1), A2 => i_DATAMEM_RM, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_1_port, B2 => n4124, 
                           ZN => n17102);
   U8745 : NOR2_X1 port map( A1 => n11579, A2 => DATA_SIZE_1_port, ZN => 
                           DataPath_LDSTR_n60);
   U8746 : NAND2_X1 port map( A1 => n11580, A2 => DataPath_LDSTR_n85, ZN => 
                           DataPath_LDSTR_n69);
   U8747 : AND2_X1 port map( A1 => DataPath_LDSTR_n79, A2 => DataPath_LDSTR_n86
                           , ZN => DataPath_LDSTR_n85);
   U8748 : NOR2_X1 port map( A1 => n4155, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, ZN => 
                           n12960);
   U8749 : OAI21_X1 port map( B1 => i_ALU_OP_3_port, B2 => n4129, A => n11499, 
                           ZN => DataPath_ALUhw_SHIFTER_HW_n549);
   U8750 : OR3_X1 port map( A1 => DataPath_LDSTR_n41, A2 => i_UNSIG_SIGN_N, A3 
                           => n4127, ZN => DataPath_LDSTR_n45);
   U8751 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_14_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_13_port, ZN => 
                           n12971);
   U8752 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_13_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_12_port, ZN => 
                           n12972);
   U8753 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_12_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_11_port, ZN => 
                           n12973);
   U8754 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_11_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_10_port, ZN => 
                           n12974);
   U8755 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_10_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_9_port, ZN => 
                           n12975);
   U8756 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_9_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_8_port, ZN => 
                           n12961);
   U8757 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_8_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_7_port, ZN => 
                           n12962);
   U8758 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_7_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_6_port, ZN => 
                           n12963);
   U8759 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_6_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_5_port, ZN => 
                           n12964);
   U8760 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_5_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_4_port, ZN => 
                           n12965);
   U8761 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_4_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_3_port, ZN => 
                           n12966);
   U8762 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_3_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_2_port, ZN => 
                           n12967);
   U8763 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_2_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_1_port, ZN => 
                           n12968);
   U8764 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_1_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_0_port, ZN => 
                           n12969);
   U8765 : AOI22_X1 port map( A1 => n12977, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, B1 => 
                           n11399, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_14_port, ZN => 
                           n12970);
   U8766 : NAND2_X1 port map( A1 => i_ALU_OP_4_port, A2 => n4132, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n576);
   U8767 : AOI21_X1 port map( B1 => n12977, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_0_port, A => 
                           n11606, ZN => n12976);
   U8768 : INV_X1 port map( A => n12953, ZN => n11606);
   U8769 : OAI21_X1 port map( B1 => DATA_SIZE_1_port, B2 => DATA_SIZE_0_port, A
                           => n4118, ZN => DataPath_LDSTR_n72);
   U8770 : OAI21_X1 port map( B1 => i_ALU_OP_4_port, B2 => 
                           DataPath_ALUhw_BWISE_n135, A => 
                           DataPath_ALUhw_BWISE_n136, ZN => 
                           DataPath_ALUhw_BWISE_n70);
   U8771 : AOI21_X1 port map( B1 => i_ALU_OP_3_port, B2 => n4132, A => 
                           DataPath_ALUhw_BWISE_n137, ZN => 
                           DataPath_ALUhw_BWISE_n135);
   U8772 : OR3_X1 port map( A1 => n4129, A2 => i_ALU_OP_3_port, A3 => n11540, 
                           ZN => DataPath_ALUhw_BWISE_n136);
   U8773 : NOR2_X1 port map( A1 => n4134, A2 => i_ALU_OP_3_port, ZN => 
                           DataPath_ALUhw_BWISE_n137);
   U8774 : INV_X1 port map( A => DataPath_RF_fill_address_ext_14_port, ZN => 
                           n11397);
   U8775 : OAI22_X1 port map( A1 => n3907, A2 => n12934, B1 => n12971, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_14_port);
   U8776 : INV_X1 port map( A => DataPath_RF_fill_address_ext_15_port, ZN => 
                           n11398);
   U8777 : OAI22_X1 port map( A1 => n3906, A2 => n12933, B1 => n12970, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_15_port);
   U8778 : INV_X1 port map( A => DataPath_RF_fill_address_ext_7_port, ZN => 
                           n11390);
   U8779 : OAI22_X1 port map( A1 => n3909, A2 => n12941, B1 => n12963, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_7_port);
   U8780 : INV_X1 port map( A => DataPath_RF_fill_address_ext_6_port, ZN => 
                           n11389);
   U8781 : OAI22_X1 port map( A1 => n3908, A2 => n12942, B1 => n12964, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_6_port);
   U8782 : INV_X1 port map( A => DataPath_RF_fill_address_ext_5_port, ZN => 
                           n11388);
   U8783 : OAI22_X1 port map( A1 => n3908, A2 => n12943, B1 => n12965, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_5_port);
   U8784 : INV_X1 port map( A => DataPath_RF_fill_address_ext_4_port, ZN => 
                           n11387);
   U8785 : OAI22_X1 port map( A1 => n3908, A2 => n12944, B1 => n12966, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_4_port);
   U8786 : INV_X1 port map( A => DataPath_RF_fill_address_ext_3_port, ZN => 
                           n11386);
   U8787 : OAI22_X1 port map( A1 => n3907, A2 => n12945, B1 => n12967, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_3_port);
   U8788 : INV_X1 port map( A => DataPath_RF_fill_address_ext_2_port, ZN => 
                           n11385);
   U8789 : OAI22_X1 port map( A1 => n3908, A2 => n12946, B1 => n12968, B2 => 
                           n3899, ZN => DataPath_RF_fill_address_ext_2_port);
   U8790 : INV_X1 port map( A => DataPath_RF_fill_address_ext_1_port, ZN => 
                           n11384);
   U8791 : OAI22_X1 port map( A1 => n3907, A2 => n12947, B1 => n12969, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_1_port);
   U8792 : INV_X1 port map( A => DataPath_RF_fill_address_ext_0_port, ZN => 
                           n11383);
   U8793 : OAI22_X1 port map( A1 => n3905, A2 => n12948, B1 => n12976, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_0_port);
   U8794 : INV_X1 port map( A => DataPath_RF_fill_address_ext_13_port, ZN => 
                           n11396);
   U8795 : OAI22_X1 port map( A1 => n3907, A2 => n12935, B1 => n12972, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_13_port);
   U8796 : INV_X1 port map( A => DataPath_RF_fill_address_ext_12_port, ZN => 
                           n11395);
   U8797 : OAI22_X1 port map( A1 => n3906, A2 => n12936, B1 => n12973, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_12_port);
   U8798 : INV_X1 port map( A => DataPath_RF_fill_address_ext_11_port, ZN => 
                           n11394);
   U8799 : OAI22_X1 port map( A1 => n3906, A2 => n12937, B1 => n12974, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_11_port);
   U8800 : INV_X1 port map( A => DataPath_RF_fill_address_ext_10_port, ZN => 
                           n11393);
   U8801 : OAI22_X1 port map( A1 => n3906, A2 => n12938, B1 => n12975, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_10_port);
   U8802 : INV_X1 port map( A => DataPath_RF_fill_address_ext_9_port, ZN => 
                           n11392);
   U8803 : OAI22_X1 port map( A1 => n3909, A2 => n12939, B1 => n12961, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_9_port);
   U8804 : INV_X1 port map( A => DataPath_RF_fill_address_ext_8_port, ZN => 
                           n11391);
   U8805 : OAI22_X1 port map( A1 => n3909, A2 => n12940, B1 => n12962, B2 => 
                           n3900, ZN => DataPath_RF_fill_address_ext_8_port);
   U8806 : AOI21_X1 port map( B1 => DRAM_READNOTWRITE_port, B2 => CU_I_n104, A 
                           => CU_I_n98, ZN => DRAM_ISSUE_port);
   U8807 : NOR2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n576, A2 => 
                           i_ALU_OP_3_port, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n349);
   U8808 : NAND2_X1 port map( A1 => DATA_SIZE_1_port, A2 => n11579, ZN => 
                           DataPath_LDSTR_n80);
   U8809 : NAND2_X1 port map( A1 => i_ALU_OP_3_port, A2 => n4132, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n641);
   U8810 : NOR2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n641, A2 => 
                           i_ALU_OP_4_port, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n478);
   U8811 : NAND2_X1 port map( A1 => DataPath_LDSTR_n60, A2 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_1_port, ZN =>
                           DataPath_LDSTR_n79);
   U8812 : AND3_X1 port map( A1 => n11578, A2 => n408, A3 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_0_port, ZN =>
                           DataPath_LDSTR_n84);
   U8813 : AND2_X1 port map( A1 => DataPath_RF_c_swin_2_port, A2 => n11607, ZN 
                           => DataPath_RF_c_swin_masked_1bit_1_0_port);
   U8814 : AND2_X1 port map( A1 => DataPath_RF_c_swin_1_port, A2 => n11607, ZN 
                           => DataPath_RF_c_swin_masked_1bit_0_0_port);
   U8815 : AND2_X1 port map( A1 => DataPath_RF_c_swin_0_port, A2 => n11607, ZN 
                           => DataPath_RF_c_swin_masked_1bit_4_0_port);
   U8816 : AND2_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n11607, ZN 
                           => DataPath_RF_c_swin_masked_1bit_2_0_port);
   U8817 : INV_X1 port map( A => n17114, ZN => n11542);
   U8818 : AOI22_X1 port map( A1 => n256, A2 => DataPath_i_REG_LDSTR_OUT_9_port
                           , B1 => DataPath_i_REG_MEM_ALUOUT_9_port, B2 => 
                           n4109, ZN => n17114);
   U8819 : INV_X1 port map( A => n14250, ZN => n8683);
   U8820 : AOI22_X1 port map( A1 => n379, A2 => n1895, B1 => 
                           DRAM_ADDRESS_8_port, B2 => n8323, ZN => n14250);
   U8821 : INV_X1 port map( A => n14249, ZN => n8684);
   U8822 : AOI22_X1 port map( A1 => n380, A2 => n1895, B1 => 
                           DRAM_ADDRESS_7_port, B2 => n8323, ZN => n14249);
   U8823 : INV_X1 port map( A => n14248, ZN => n8685);
   U8824 : AOI22_X1 port map( A1 => n381, A2 => n1895, B1 => 
                           DRAM_ADDRESS_6_port, B2 => n8323, ZN => n14248);
   U8825 : INV_X1 port map( A => n14247, ZN => n8686);
   U8826 : AOI22_X1 port map( A1 => n382, A2 => n1895, B1 => 
                           DRAM_ADDRESS_5_port, B2 => n8323, ZN => n14247);
   U8827 : INV_X1 port map( A => n14246, ZN => n8687);
   U8828 : AOI22_X1 port map( A1 => n383, A2 => n1895, B1 => 
                           DRAM_ADDRESS_4_port, B2 => n8323, ZN => n14246);
   U8829 : INV_X1 port map( A => n14245, ZN => n8688);
   U8830 : AOI22_X1 port map( A1 => n384, A2 => n1895, B1 => 
                           DRAM_ADDRESS_3_port, B2 => n8323, ZN => n14245);
   U8831 : INV_X1 port map( A => n14244, ZN => n8689);
   U8832 : AOI22_X1 port map( A1 => n385, A2 => n1895, B1 => 
                           DRAM_ADDRESS_2_port, B2 => n8323, ZN => n14244);
   U8833 : INV_X1 port map( A => n14243, ZN => n8690);
   U8834 : AOI22_X1 port map( A1 => n386, A2 => n1895, B1 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_1_port, B2 =>
                           n8323, ZN => n14243);
   U8835 : INV_X1 port map( A => n14242, ZN => n8691);
   U8836 : AOI22_X1 port map( A1 => n11482, A2 => n1895, B1 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_0_port, B2 =>
                           n8323, ZN => n14242);
   U8837 : INV_X1 port map( A => n17081, ZN => n11482);
   U8838 : AOI22_X1 port map( A1 => DataPath_i_SETCMP_OUT_0_port, A2 => 
                           i_SEL_ALU_SETCMP, B1 => DataPath_i_ALU_OUT_0_port, 
                           B2 => n8325, ZN => n17081);
   U8839 : INV_X1 port map( A => n17121, ZN => n11549);
   U8840 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_31_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_31_port, B2 =>
                           n4110, ZN => n17121);
   U8841 : INV_X1 port map( A => n17115, ZN => n11543);
   U8842 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_8_port, A2 => n256
                           , B1 => DataPath_i_REG_MEM_ALUOUT_8_port, B2 => 
                           n4109, ZN => n17115);
   U8843 : INV_X1 port map( A => n17116, ZN => n11544);
   U8844 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_7_port, A2 => n256
                           , B1 => DataPath_i_REG_MEM_ALUOUT_7_port, B2 => 
                           n4109, ZN => n17116);
   U8845 : INV_X1 port map( A => n17117, ZN => n11545);
   U8846 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_6_port, A2 => n256
                           , B1 => DataPath_i_REG_MEM_ALUOUT_6_port, B2 => 
                           n4109, ZN => n17117);
   U8847 : INV_X1 port map( A => n17118, ZN => n11546);
   U8848 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_5_port, A2 => n256
                           , B1 => DataPath_i_REG_MEM_ALUOUT_5_port, B2 => 
                           n4110, ZN => n17118);
   U8849 : INV_X1 port map( A => n17119, ZN => n11547);
   U8850 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_4_port, A2 => n256
                           , B1 => DataPath_i_REG_MEM_ALUOUT_4_port, B2 => 
                           n4110, ZN => n17119);
   U8851 : INV_X1 port map( A => n17120, ZN => n11548);
   U8852 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_3_port, A2 => n256
                           , B1 => DataPath_i_REG_MEM_ALUOUT_3_port, B2 => 
                           n4110, ZN => n17120);
   U8853 : AOI222_X1 port map( A1 => n305, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N113_port, B2 => n3263, C1 => n413
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n141);
   U8854 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_4_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_4_port, ZN => 
                           DataPath_WRF_CUhw_N113_port);
   U8855 : AOI222_X1 port map( A1 => n306, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N114_port, B2 => n3262, C1 => n414
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n140);
   U8856 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_5_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_5_port, ZN => 
                           DataPath_WRF_CUhw_N114_port);
   U8857 : AOI222_X1 port map( A1 => n307, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N115_port, B2 => n3262, C1 => n415
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n139);
   U8858 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_6_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_6_port, ZN => 
                           DataPath_WRF_CUhw_N115_port);
   U8859 : AOI222_X1 port map( A1 => n308, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N116_port, B2 => n3262, C1 => n416
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n138);
   U8860 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_7_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_7_port, ZN => 
                           DataPath_WRF_CUhw_N116_port);
   U8861 : AOI222_X1 port map( A1 => n295, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N117_port, B2 => n3262, C1 => n417
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n137);
   U8862 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_8_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_8_port, ZN => 
                           DataPath_WRF_CUhw_N117_port);
   U8863 : AOI222_X1 port map( A1 => n296, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N118_port, B2 => n3262, C1 => n418
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n136);
   U8864 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_9_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_9_port, ZN => 
                           DataPath_WRF_CUhw_N118_port);
   U8865 : AOI222_X1 port map( A1 => n297, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N119_port, B2 => n3264, C1 => n419
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n135);
   U8866 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_10_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_10_port, ZN => 
                           DataPath_WRF_CUhw_N119_port);
   U8867 : AOI222_X1 port map( A1 => n298, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N120_port, B2 => n3264, C1 => n402
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n134);
   U8868 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_11_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_11_port, ZN => 
                           DataPath_WRF_CUhw_N120_port);
   U8869 : AOI222_X1 port map( A1 => n299, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N121_port, B2 => n3264, C1 => n403
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n133);
   U8870 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_12_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_12_port, ZN => 
                           DataPath_WRF_CUhw_N121_port);
   U8871 : AOI222_X1 port map( A1 => n300, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N122_port, B2 => n3264, C1 => n404
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n132);
   U8872 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_13_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_13_port, ZN => 
                           DataPath_WRF_CUhw_N122_port);
   U8873 : AOI222_X1 port map( A1 => n301, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N123_port, B2 => n3264, C1 => n405
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n131);
   U8874 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_14_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_14_port, ZN => 
                           DataPath_WRF_CUhw_N123_port);
   U8875 : AOI222_X1 port map( A1 => n302, A2 => n3266, B1 => 
                           DataPath_WRF_CUhw_N124_port, B2 => n3264, C1 => n406
                           , C2 => n2475, ZN => DataPath_WRF_CUhw_n130);
   U8876 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_15_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_15_port, ZN => 
                           DataPath_WRF_CUhw_N124_port);
   U8877 : BUF_X1 port map( A => DataPath_RF_c_swin_4_port, Z => n3844);
   U8878 : INV_X1 port map( A => n14394, ZN => n8788);
   U8879 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_31_port, B2 => n2509, ZN
                           => n14394);
   U8880 : INV_X1 port map( A => n14393, ZN => n8789);
   U8881 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_30_port, B2 => n2509, ZN
                           => n14393);
   U8882 : INV_X1 port map( A => n14392, ZN => n8790);
   U8883 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_29_port, B2 => n2509, ZN
                           => n14392);
   U8884 : INV_X1 port map( A => n14391, ZN => n8791);
   U8885 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_28_port, B2 => n2509, ZN
                           => n14391);
   U8886 : INV_X1 port map( A => n14390, ZN => n8792);
   U8887 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_27_port, B2 => n2509, ZN
                           => n14390);
   U8888 : INV_X1 port map( A => n14389, ZN => n8793);
   U8889 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_26_port, B2 => n2509, ZN
                           => n14389);
   U8890 : INV_X1 port map( A => n14388, ZN => n8794);
   U8891 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_25_port, B2 => n2509, ZN
                           => n14388);
   U8892 : INV_X1 port map( A => n14387, ZN => n8795);
   U8893 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_24_port, B2 => n2509, ZN
                           => n14387);
   U8894 : INV_X1 port map( A => n14386, ZN => n8796);
   U8895 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_23_port, B2 => n2508, ZN
                           => n14386);
   U8896 : INV_X1 port map( A => n14385, ZN => n8797);
   U8897 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_22_port, B2 => n2508, ZN
                           => n14385);
   U8898 : INV_X1 port map( A => n14384, ZN => n8798);
   U8899 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_21_port, B2 => n2508, ZN
                           => n14384);
   U8900 : INV_X1 port map( A => n14383, ZN => n8799);
   U8901 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2504, B1 => 
                           DataPath_RF_bus_reg_dataout_20_port, B2 => n2508, ZN
                           => n14383);
   U8902 : INV_X1 port map( A => n14382, ZN => n8800);
   U8903 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_19_port, B2 => n2508, ZN
                           => n14382);
   U8904 : INV_X1 port map( A => n14381, ZN => n8801);
   U8905 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_18_port, B2 => n2508, ZN
                           => n14381);
   U8906 : INV_X1 port map( A => n14380, ZN => n8802);
   U8907 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_17_port, B2 => n2508, ZN
                           => n14380);
   U8908 : INV_X1 port map( A => n14379, ZN => n8803);
   U8909 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_16_port, B2 => n2508, ZN
                           => n14379);
   U8910 : INV_X1 port map( A => n14378, ZN => n8804);
   U8911 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_15_port, B2 => n2508, ZN
                           => n14378);
   U8912 : INV_X1 port map( A => n14377, ZN => n8805);
   U8913 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_14_port, B2 => n2508, ZN
                           => n14377);
   U8914 : INV_X1 port map( A => n14376, ZN => n8806);
   U8915 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_13_port, B2 => n2508, ZN
                           => n14376);
   U8916 : INV_X1 port map( A => n14375, ZN => n8807);
   U8917 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_12_port, B2 => n2508, ZN
                           => n14375);
   U8918 : INV_X1 port map( A => n14374, ZN => n8808);
   U8919 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_11_port, B2 => n2507, ZN
                           => n14374);
   U8920 : INV_X1 port map( A => n14373, ZN => n8809);
   U8921 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_10_port, B2 => n2507, ZN
                           => n14373);
   U8922 : INV_X1 port map( A => n14372, ZN => n8810);
   U8923 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_9_port, B2 => n2507, ZN 
                           => n14372);
   U8924 : INV_X1 port map( A => n14371, ZN => n8811);
   U8925 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2505, B1 => 
                           DataPath_RF_bus_reg_dataout_8_port, B2 => n2507, ZN 
                           => n14371);
   U8926 : INV_X1 port map( A => n14370, ZN => n8812);
   U8927 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_7_port, B2 => n2507, ZN 
                           => n14370);
   U8928 : INV_X1 port map( A => n14369, ZN => n8813);
   U8929 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_6_port, B2 => n2507, ZN 
                           => n14369);
   U8930 : INV_X1 port map( A => n14368, ZN => n8814);
   U8931 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_5_port, B2 => n2507, ZN 
                           => n14368);
   U8932 : INV_X1 port map( A => n14367, ZN => n8815);
   U8933 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_4_port, B2 => n2507, ZN 
                           => n14367);
   U8934 : INV_X1 port map( A => n14366, ZN => n8816);
   U8935 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_3_port, B2 => n2507, ZN 
                           => n14366);
   U8936 : INV_X1 port map( A => n14365, ZN => n8817);
   U8937 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_2_port, B2 => n2507, ZN 
                           => n14365);
   U8938 : INV_X1 port map( A => n14364, ZN => n8818);
   U8939 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_1_port, B2 => n2507, ZN 
                           => n14364);
   U8940 : INV_X1 port map( A => n14361, ZN => n8819);
   U8941 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2506, B1 => 
                           DataPath_RF_bus_reg_dataout_0_port, B2 => n2507, ZN 
                           => n14361);
   U8942 : INV_X1 port map( A => n14428, ZN => n8820);
   U8943 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_63_port, B2 => n2515, ZN
                           => n14428);
   U8944 : INV_X1 port map( A => n14427, ZN => n8821);
   U8945 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_62_port, B2 => n2515, ZN
                           => n14427);
   U8946 : INV_X1 port map( A => n14426, ZN => n8822);
   U8947 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_61_port, B2 => n2515, ZN
                           => n14426);
   U8948 : INV_X1 port map( A => n14425, ZN => n8823);
   U8949 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_60_port, B2 => n2515, ZN
                           => n14425);
   U8950 : INV_X1 port map( A => n14424, ZN => n8824);
   U8951 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_59_port, B2 => n2515, ZN
                           => n14424);
   U8952 : INV_X1 port map( A => n14423, ZN => n8825);
   U8953 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_58_port, B2 => n2515, ZN
                           => n14423);
   U8954 : INV_X1 port map( A => n14422, ZN => n8826);
   U8955 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_57_port, B2 => n2515, ZN
                           => n14422);
   U8956 : INV_X1 port map( A => n14421, ZN => n8827);
   U8957 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_56_port, B2 => n2515, ZN
                           => n14421);
   U8958 : INV_X1 port map( A => n14420, ZN => n8828);
   U8959 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_55_port, B2 => n2514, ZN
                           => n14420);
   U8960 : INV_X1 port map( A => n14419, ZN => n8829);
   U8961 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_54_port, B2 => n2514, ZN
                           => n14419);
   U8962 : INV_X1 port map( A => n14418, ZN => n8830);
   U8963 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_53_port, B2 => n2514, ZN
                           => n14418);
   U8964 : INV_X1 port map( A => n14417, ZN => n8831);
   U8965 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2510, B1 => 
                           DataPath_RF_bus_reg_dataout_52_port, B2 => n2514, ZN
                           => n14417);
   U8966 : INV_X1 port map( A => n14416, ZN => n8832);
   U8967 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_51_port, B2 => n2514, ZN
                           => n14416);
   U8968 : INV_X1 port map( A => n14415, ZN => n8833);
   U8969 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_50_port, B2 => n2514, ZN
                           => n14415);
   U8970 : INV_X1 port map( A => n14414, ZN => n8834);
   U8971 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_49_port, B2 => n2514, ZN
                           => n14414);
   U8972 : INV_X1 port map( A => n14413, ZN => n8835);
   U8973 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_48_port, B2 => n2514, ZN
                           => n14413);
   U8974 : INV_X1 port map( A => n14412, ZN => n8836);
   U8975 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_47_port, B2 => n2514, ZN
                           => n14412);
   U8976 : INV_X1 port map( A => n14411, ZN => n8837);
   U8977 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_46_port, B2 => n2514, ZN
                           => n14411);
   U8978 : INV_X1 port map( A => n14410, ZN => n8838);
   U8979 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_45_port, B2 => n2514, ZN
                           => n14410);
   U8980 : INV_X1 port map( A => n14409, ZN => n8839);
   U8981 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_44_port, B2 => n2514, ZN
                           => n14409);
   U8982 : INV_X1 port map( A => n14408, ZN => n8840);
   U8983 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_43_port, B2 => n2513, ZN
                           => n14408);
   U8984 : INV_X1 port map( A => n14407, ZN => n8841);
   U8985 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_42_port, B2 => n2513, ZN
                           => n14407);
   U8986 : INV_X1 port map( A => n14406, ZN => n8842);
   U8987 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_41_port, B2 => n2513, ZN
                           => n14406);
   U8988 : INV_X1 port map( A => n14405, ZN => n8843);
   U8989 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2511, B1 => 
                           DataPath_RF_bus_reg_dataout_40_port, B2 => n2513, ZN
                           => n14405);
   U8990 : INV_X1 port map( A => n14404, ZN => n8844);
   U8991 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_39_port, B2 => n2513, ZN
                           => n14404);
   U8992 : INV_X1 port map( A => n14403, ZN => n8845);
   U8993 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_38_port, B2 => n2513, ZN
                           => n14403);
   U8994 : INV_X1 port map( A => n14402, ZN => n8846);
   U8995 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_37_port, B2 => n2513, ZN
                           => n14402);
   U8996 : INV_X1 port map( A => n14401, ZN => n8847);
   U8997 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_36_port, B2 => n2513, ZN
                           => n14401);
   U8998 : INV_X1 port map( A => n14400, ZN => n8848);
   U8999 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_35_port, B2 => n2513, ZN
                           => n14400);
   U9000 : INV_X1 port map( A => n14399, ZN => n8849);
   U9001 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_34_port, B2 => n2513, ZN
                           => n14399);
   U9002 : INV_X1 port map( A => n14398, ZN => n8850);
   U9003 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_33_port, B2 => n2513, ZN
                           => n14398);
   U9004 : INV_X1 port map( A => n14395, ZN => n8851);
   U9005 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2512, B1 => 
                           DataPath_RF_bus_reg_dataout_32_port, B2 => n2513, ZN
                           => n14395);
   U9006 : INV_X1 port map( A => n14462, ZN => n8852);
   U9007 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_95_port, B2 => n2521, ZN
                           => n14462);
   U9008 : INV_X1 port map( A => n14461, ZN => n8853);
   U9009 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_94_port, B2 => n2521, ZN
                           => n14461);
   U9010 : INV_X1 port map( A => n14460, ZN => n8854);
   U9011 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_93_port, B2 => n2521, ZN
                           => n14460);
   U9012 : INV_X1 port map( A => n14459, ZN => n8855);
   U9013 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_92_port, B2 => n2521, ZN
                           => n14459);
   U9014 : INV_X1 port map( A => n14458, ZN => n8856);
   U9015 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_91_port, B2 => n2521, ZN
                           => n14458);
   U9016 : INV_X1 port map( A => n14457, ZN => n8857);
   U9017 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_90_port, B2 => n2521, ZN
                           => n14457);
   U9018 : INV_X1 port map( A => n14456, ZN => n8858);
   U9019 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_89_port, B2 => n2521, ZN
                           => n14456);
   U9020 : INV_X1 port map( A => n14455, ZN => n8859);
   U9021 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_88_port, B2 => n2521, ZN
                           => n14455);
   U9022 : INV_X1 port map( A => n14454, ZN => n8860);
   U9023 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_87_port, B2 => n2520, ZN
                           => n14454);
   U9024 : INV_X1 port map( A => n14453, ZN => n8861);
   U9025 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_86_port, B2 => n2520, ZN
                           => n14453);
   U9026 : INV_X1 port map( A => n14452, ZN => n8862);
   U9027 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_85_port, B2 => n2520, ZN
                           => n14452);
   U9028 : INV_X1 port map( A => n14451, ZN => n8863);
   U9029 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2516, B1 => 
                           DataPath_RF_bus_reg_dataout_84_port, B2 => n2520, ZN
                           => n14451);
   U9030 : INV_X1 port map( A => n14450, ZN => n8864);
   U9031 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_83_port, B2 => n2520, ZN
                           => n14450);
   U9032 : INV_X1 port map( A => n14449, ZN => n8865);
   U9033 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_82_port, B2 => n2520, ZN
                           => n14449);
   U9034 : INV_X1 port map( A => n14448, ZN => n8866);
   U9035 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_81_port, B2 => n2520, ZN
                           => n14448);
   U9036 : INV_X1 port map( A => n14447, ZN => n8867);
   U9037 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_80_port, B2 => n2520, ZN
                           => n14447);
   U9038 : INV_X1 port map( A => n14446, ZN => n8868);
   U9039 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_79_port, B2 => n2520, ZN
                           => n14446);
   U9040 : INV_X1 port map( A => n14445, ZN => n8869);
   U9041 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_78_port, B2 => n2520, ZN
                           => n14445);
   U9042 : INV_X1 port map( A => n14444, ZN => n8870);
   U9043 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_77_port, B2 => n2520, ZN
                           => n14444);
   U9044 : INV_X1 port map( A => n14443, ZN => n8871);
   U9045 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_76_port, B2 => n2520, ZN
                           => n14443);
   U9046 : INV_X1 port map( A => n14442, ZN => n8872);
   U9047 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_75_port, B2 => n2519, ZN
                           => n14442);
   U9048 : INV_X1 port map( A => n14441, ZN => n8873);
   U9049 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_74_port, B2 => n2519, ZN
                           => n14441);
   U9050 : INV_X1 port map( A => n14440, ZN => n8874);
   U9051 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_73_port, B2 => n2519, ZN
                           => n14440);
   U9052 : INV_X1 port map( A => n14439, ZN => n8875);
   U9053 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2517, B1 => 
                           DataPath_RF_bus_reg_dataout_72_port, B2 => n2519, ZN
                           => n14439);
   U9054 : INV_X1 port map( A => n14438, ZN => n8876);
   U9055 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_71_port, B2 => n2519, ZN
                           => n14438);
   U9056 : INV_X1 port map( A => n14437, ZN => n8877);
   U9057 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_70_port, B2 => n2519, ZN
                           => n14437);
   U9058 : INV_X1 port map( A => n14436, ZN => n8878);
   U9059 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_69_port, B2 => n2519, ZN
                           => n14436);
   U9060 : INV_X1 port map( A => n14435, ZN => n8879);
   U9061 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_68_port, B2 => n2519, ZN
                           => n14435);
   U9062 : INV_X1 port map( A => n14434, ZN => n8880);
   U9063 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_67_port, B2 => n2519, ZN
                           => n14434);
   U9064 : INV_X1 port map( A => n14433, ZN => n8881);
   U9065 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_66_port, B2 => n2519, ZN
                           => n14433);
   U9066 : INV_X1 port map( A => n14432, ZN => n8882);
   U9067 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_65_port, B2 => n2519, ZN
                           => n14432);
   U9068 : INV_X1 port map( A => n14429, ZN => n8883);
   U9069 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2518, B1 => 
                           DataPath_RF_bus_reg_dataout_64_port, B2 => n2519, ZN
                           => n14429);
   U9070 : INV_X1 port map( A => n14496, ZN => n8884);
   U9071 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_127_port, B2 => n2527, 
                           ZN => n14496);
   U9072 : INV_X1 port map( A => n14495, ZN => n8885);
   U9073 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_126_port, B2 => n2527, 
                           ZN => n14495);
   U9074 : INV_X1 port map( A => n14494, ZN => n8886);
   U9075 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_125_port, B2 => n2527, 
                           ZN => n14494);
   U9076 : INV_X1 port map( A => n14493, ZN => n8887);
   U9077 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_124_port, B2 => n2527, 
                           ZN => n14493);
   U9078 : INV_X1 port map( A => n14492, ZN => n8888);
   U9079 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_123_port, B2 => n2527, 
                           ZN => n14492);
   U9080 : INV_X1 port map( A => n14491, ZN => n8889);
   U9081 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_122_port, B2 => n2527, 
                           ZN => n14491);
   U9082 : INV_X1 port map( A => n14490, ZN => n8890);
   U9083 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_121_port, B2 => n2527, 
                           ZN => n14490);
   U9084 : INV_X1 port map( A => n14489, ZN => n8891);
   U9085 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_120_port, B2 => n2527, 
                           ZN => n14489);
   U9086 : INV_X1 port map( A => n14488, ZN => n8892);
   U9087 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_119_port, B2 => n2526, 
                           ZN => n14488);
   U9088 : INV_X1 port map( A => n14487, ZN => n8893);
   U9089 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_118_port, B2 => n2526, 
                           ZN => n14487);
   U9090 : INV_X1 port map( A => n14486, ZN => n8894);
   U9091 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_117_port, B2 => n2526, 
                           ZN => n14486);
   U9092 : INV_X1 port map( A => n14485, ZN => n8895);
   U9093 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2522, B1 => 
                           DataPath_RF_bus_reg_dataout_116_port, B2 => n2526, 
                           ZN => n14485);
   U9094 : INV_X1 port map( A => n14484, ZN => n8896);
   U9095 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_115_port, B2 => n2526, 
                           ZN => n14484);
   U9096 : INV_X1 port map( A => n14483, ZN => n8897);
   U9097 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_114_port, B2 => n2526, 
                           ZN => n14483);
   U9098 : INV_X1 port map( A => n14482, ZN => n8898);
   U9099 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_113_port, B2 => n2526, 
                           ZN => n14482);
   U9100 : INV_X1 port map( A => n14481, ZN => n8899);
   U9101 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_112_port, B2 => n2526, 
                           ZN => n14481);
   U9102 : INV_X1 port map( A => n14480, ZN => n8900);
   U9103 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_111_port, B2 => n2526, 
                           ZN => n14480);
   U9104 : INV_X1 port map( A => n14479, ZN => n8901);
   U9105 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_110_port, B2 => n2526, 
                           ZN => n14479);
   U9106 : INV_X1 port map( A => n14478, ZN => n8902);
   U9107 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_109_port, B2 => n2526, 
                           ZN => n14478);
   U9108 : INV_X1 port map( A => n14477, ZN => n8903);
   U9109 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_108_port, B2 => n2526, 
                           ZN => n14477);
   U9110 : INV_X1 port map( A => n14476, ZN => n8904);
   U9111 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_107_port, B2 => n2525, 
                           ZN => n14476);
   U9112 : INV_X1 port map( A => n14475, ZN => n8905);
   U9113 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_106_port, B2 => n2525, 
                           ZN => n14475);
   U9114 : INV_X1 port map( A => n14474, ZN => n8906);
   U9115 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_105_port, B2 => n2525, 
                           ZN => n14474);
   U9116 : INV_X1 port map( A => n14473, ZN => n8907);
   U9117 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2523, B1 => 
                           DataPath_RF_bus_reg_dataout_104_port, B2 => n2525, 
                           ZN => n14473);
   U9118 : INV_X1 port map( A => n14472, ZN => n8908);
   U9119 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_103_port, B2 => n2525, 
                           ZN => n14472);
   U9120 : INV_X1 port map( A => n14471, ZN => n8909);
   U9121 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_102_port, B2 => n2525, 
                           ZN => n14471);
   U9122 : INV_X1 port map( A => n14470, ZN => n8910);
   U9123 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_101_port, B2 => n2525, 
                           ZN => n14470);
   U9124 : INV_X1 port map( A => n14469, ZN => n8911);
   U9125 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_100_port, B2 => n2525, 
                           ZN => n14469);
   U9126 : INV_X1 port map( A => n14468, ZN => n8912);
   U9127 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_99_port, B2 => n2525, ZN
                           => n14468);
   U9128 : INV_X1 port map( A => n14467, ZN => n8913);
   U9129 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_98_port, B2 => n2525, ZN
                           => n14467);
   U9130 : INV_X1 port map( A => n14466, ZN => n8914);
   U9131 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_97_port, B2 => n2525, ZN
                           => n14466);
   U9132 : INV_X1 port map( A => n14463, ZN => n8915);
   U9133 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2524, B1 => 
                           DataPath_RF_bus_reg_dataout_96_port, B2 => n2525, ZN
                           => n14463);
   U9134 : INV_X1 port map( A => n14530, ZN => n8916);
   U9135 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_159_port, B2 => n2533, 
                           ZN => n14530);
   U9136 : INV_X1 port map( A => n14529, ZN => n8917);
   U9137 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_158_port, B2 => n2533, 
                           ZN => n14529);
   U9138 : INV_X1 port map( A => n14528, ZN => n8918);
   U9139 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_157_port, B2 => n2533, 
                           ZN => n14528);
   U9140 : INV_X1 port map( A => n14527, ZN => n8919);
   U9141 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_156_port, B2 => n2533, 
                           ZN => n14527);
   U9142 : INV_X1 port map( A => n14526, ZN => n8920);
   U9143 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_155_port, B2 => n2533, 
                           ZN => n14526);
   U9144 : INV_X1 port map( A => n14525, ZN => n8921);
   U9145 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_154_port, B2 => n2533, 
                           ZN => n14525);
   U9146 : INV_X1 port map( A => n14524, ZN => n8922);
   U9147 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_153_port, B2 => n2533, 
                           ZN => n14524);
   U9148 : INV_X1 port map( A => n14523, ZN => n8923);
   U9149 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_152_port, B2 => n2533, 
                           ZN => n14523);
   U9150 : INV_X1 port map( A => n14522, ZN => n8924);
   U9151 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_151_port, B2 => n2532, 
                           ZN => n14522);
   U9152 : INV_X1 port map( A => n14521, ZN => n8925);
   U9153 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_150_port, B2 => n2532, 
                           ZN => n14521);
   U9154 : INV_X1 port map( A => n14520, ZN => n8926);
   U9155 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_149_port, B2 => n2532, 
                           ZN => n14520);
   U9156 : INV_X1 port map( A => n14519, ZN => n8927);
   U9157 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2528, B1 => 
                           DataPath_RF_bus_reg_dataout_148_port, B2 => n2532, 
                           ZN => n14519);
   U9158 : INV_X1 port map( A => n14518, ZN => n8928);
   U9159 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_147_port, B2 => n2532, 
                           ZN => n14518);
   U9160 : INV_X1 port map( A => n14517, ZN => n8929);
   U9161 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_146_port, B2 => n2532, 
                           ZN => n14517);
   U9162 : INV_X1 port map( A => n14516, ZN => n8930);
   U9163 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_145_port, B2 => n2532, 
                           ZN => n14516);
   U9164 : INV_X1 port map( A => n14515, ZN => n8931);
   U9165 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_144_port, B2 => n2532, 
                           ZN => n14515);
   U9166 : INV_X1 port map( A => n14514, ZN => n8932);
   U9167 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_143_port, B2 => n2532, 
                           ZN => n14514);
   U9168 : INV_X1 port map( A => n14513, ZN => n8933);
   U9169 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_142_port, B2 => n2532, 
                           ZN => n14513);
   U9170 : INV_X1 port map( A => n14512, ZN => n8934);
   U9171 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_141_port, B2 => n2532, 
                           ZN => n14512);
   U9172 : INV_X1 port map( A => n14511, ZN => n8935);
   U9173 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_140_port, B2 => n2532, 
                           ZN => n14511);
   U9174 : INV_X1 port map( A => n14510, ZN => n8936);
   U9175 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_139_port, B2 => n2531, 
                           ZN => n14510);
   U9176 : INV_X1 port map( A => n14509, ZN => n8937);
   U9177 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_138_port, B2 => n2531, 
                           ZN => n14509);
   U9178 : INV_X1 port map( A => n14508, ZN => n8938);
   U9179 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_137_port, B2 => n2531, 
                           ZN => n14508);
   U9180 : INV_X1 port map( A => n14507, ZN => n8939);
   U9181 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2529, B1 => 
                           DataPath_RF_bus_reg_dataout_136_port, B2 => n2531, 
                           ZN => n14507);
   U9182 : INV_X1 port map( A => n14506, ZN => n8940);
   U9183 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_135_port, B2 => n2531, 
                           ZN => n14506);
   U9184 : INV_X1 port map( A => n14505, ZN => n8941);
   U9185 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_134_port, B2 => n2531, 
                           ZN => n14505);
   U9186 : INV_X1 port map( A => n14504, ZN => n8942);
   U9187 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_133_port, B2 => n2531, 
                           ZN => n14504);
   U9188 : INV_X1 port map( A => n14503, ZN => n8943);
   U9189 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_132_port, B2 => n2531, 
                           ZN => n14503);
   U9190 : INV_X1 port map( A => n14502, ZN => n8944);
   U9191 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_131_port, B2 => n2531, 
                           ZN => n14502);
   U9192 : INV_X1 port map( A => n14501, ZN => n8945);
   U9193 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_130_port, B2 => n2531, 
                           ZN => n14501);
   U9194 : INV_X1 port map( A => n14500, ZN => n8946);
   U9195 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_129_port, B2 => n2531, 
                           ZN => n14500);
   U9196 : INV_X1 port map( A => n14497, ZN => n8947);
   U9197 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2530, B1 => 
                           DataPath_RF_bus_reg_dataout_128_port, B2 => n2531, 
                           ZN => n14497);
   U9198 : INV_X1 port map( A => n14564, ZN => n8948);
   U9199 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_191_port, B2 => n2539, 
                           ZN => n14564);
   U9200 : INV_X1 port map( A => n14563, ZN => n8949);
   U9201 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_190_port, B2 => n2539, 
                           ZN => n14563);
   U9202 : INV_X1 port map( A => n14562, ZN => n8950);
   U9203 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_189_port, B2 => n2539, 
                           ZN => n14562);
   U9204 : INV_X1 port map( A => n14561, ZN => n8951);
   U9205 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_188_port, B2 => n2539, 
                           ZN => n14561);
   U9206 : INV_X1 port map( A => n14560, ZN => n8952);
   U9207 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_187_port, B2 => n2539, 
                           ZN => n14560);
   U9208 : INV_X1 port map( A => n14559, ZN => n8953);
   U9209 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_186_port, B2 => n2539, 
                           ZN => n14559);
   U9210 : INV_X1 port map( A => n14558, ZN => n8954);
   U9211 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_185_port, B2 => n2539, 
                           ZN => n14558);
   U9212 : INV_X1 port map( A => n14557, ZN => n8955);
   U9213 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_184_port, B2 => n2539, 
                           ZN => n14557);
   U9214 : INV_X1 port map( A => n14556, ZN => n8956);
   U9215 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_183_port, B2 => n2538, 
                           ZN => n14556);
   U9216 : INV_X1 port map( A => n14555, ZN => n8957);
   U9217 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_182_port, B2 => n2538, 
                           ZN => n14555);
   U9218 : INV_X1 port map( A => n14554, ZN => n8958);
   U9219 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_181_port, B2 => n2538, 
                           ZN => n14554);
   U9220 : INV_X1 port map( A => n14553, ZN => n8959);
   U9221 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2534, B1 => 
                           DataPath_RF_bus_reg_dataout_180_port, B2 => n2538, 
                           ZN => n14553);
   U9222 : INV_X1 port map( A => n14552, ZN => n8960);
   U9223 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_179_port, B2 => n2538, 
                           ZN => n14552);
   U9224 : INV_X1 port map( A => n14551, ZN => n8961);
   U9225 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_178_port, B2 => n2538, 
                           ZN => n14551);
   U9226 : INV_X1 port map( A => n14550, ZN => n8962);
   U9227 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_177_port, B2 => n2538, 
                           ZN => n14550);
   U9228 : INV_X1 port map( A => n14549, ZN => n8963);
   U9229 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_176_port, B2 => n2538, 
                           ZN => n14549);
   U9230 : INV_X1 port map( A => n14548, ZN => n8964);
   U9231 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_175_port, B2 => n2538, 
                           ZN => n14548);
   U9232 : INV_X1 port map( A => n14547, ZN => n8965);
   U9233 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_174_port, B2 => n2538, 
                           ZN => n14547);
   U9234 : INV_X1 port map( A => n14546, ZN => n8966);
   U9235 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_173_port, B2 => n2538, 
                           ZN => n14546);
   U9236 : INV_X1 port map( A => n14545, ZN => n8967);
   U9237 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_172_port, B2 => n2538, 
                           ZN => n14545);
   U9238 : INV_X1 port map( A => n14544, ZN => n8968);
   U9239 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_171_port, B2 => n2537, 
                           ZN => n14544);
   U9240 : INV_X1 port map( A => n14543, ZN => n8969);
   U9241 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_170_port, B2 => n2537, 
                           ZN => n14543);
   U9242 : INV_X1 port map( A => n14542, ZN => n8970);
   U9243 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_169_port, B2 => n2537, 
                           ZN => n14542);
   U9244 : INV_X1 port map( A => n14541, ZN => n8971);
   U9245 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2535, B1 => 
                           DataPath_RF_bus_reg_dataout_168_port, B2 => n2537, 
                           ZN => n14541);
   U9246 : INV_X1 port map( A => n14540, ZN => n8972);
   U9247 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_167_port, B2 => n2537, 
                           ZN => n14540);
   U9248 : INV_X1 port map( A => n14539, ZN => n8973);
   U9249 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_166_port, B2 => n2537, 
                           ZN => n14539);
   U9250 : INV_X1 port map( A => n14538, ZN => n8974);
   U9251 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_165_port, B2 => n2537, 
                           ZN => n14538);
   U9252 : INV_X1 port map( A => n14537, ZN => n8975);
   U9253 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_164_port, B2 => n2537, 
                           ZN => n14537);
   U9254 : INV_X1 port map( A => n14536, ZN => n8976);
   U9255 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_163_port, B2 => n2537, 
                           ZN => n14536);
   U9256 : INV_X1 port map( A => n14535, ZN => n8977);
   U9257 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_162_port, B2 => n2537, 
                           ZN => n14535);
   U9258 : INV_X1 port map( A => n14534, ZN => n8978);
   U9259 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_161_port, B2 => n2537, 
                           ZN => n14534);
   U9260 : INV_X1 port map( A => n14531, ZN => n8979);
   U9261 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2536, B1 => 
                           DataPath_RF_bus_reg_dataout_160_port, B2 => n2537, 
                           ZN => n14531);
   U9262 : INV_X1 port map( A => n14598, ZN => n8980);
   U9263 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_223_port, B2 => n2545, 
                           ZN => n14598);
   U9264 : INV_X1 port map( A => n14597, ZN => n8981);
   U9265 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_222_port, B2 => n2545, 
                           ZN => n14597);
   U9266 : INV_X1 port map( A => n14596, ZN => n8982);
   U9267 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_221_port, B2 => n2545, 
                           ZN => n14596);
   U9268 : INV_X1 port map( A => n14595, ZN => n8983);
   U9269 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_220_port, B2 => n2545, 
                           ZN => n14595);
   U9270 : INV_X1 port map( A => n14594, ZN => n8984);
   U9271 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_219_port, B2 => n2545, 
                           ZN => n14594);
   U9272 : INV_X1 port map( A => n14593, ZN => n8985);
   U9273 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_218_port, B2 => n2545, 
                           ZN => n14593);
   U9274 : INV_X1 port map( A => n14592, ZN => n8986);
   U9275 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_217_port, B2 => n2545, 
                           ZN => n14592);
   U9276 : INV_X1 port map( A => n14591, ZN => n8987);
   U9277 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_216_port, B2 => n2545, 
                           ZN => n14591);
   U9278 : INV_X1 port map( A => n14590, ZN => n8988);
   U9279 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_215_port, B2 => n2544, 
                           ZN => n14590);
   U9280 : INV_X1 port map( A => n14589, ZN => n8989);
   U9281 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_214_port, B2 => n2544, 
                           ZN => n14589);
   U9282 : INV_X1 port map( A => n14588, ZN => n8990);
   U9283 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_213_port, B2 => n2544, 
                           ZN => n14588);
   U9284 : INV_X1 port map( A => n14587, ZN => n8991);
   U9285 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2540, B1 => 
                           DataPath_RF_bus_reg_dataout_212_port, B2 => n2544, 
                           ZN => n14587);
   U9286 : INV_X1 port map( A => n14586, ZN => n8992);
   U9287 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_211_port, B2 => n2544, 
                           ZN => n14586);
   U9288 : INV_X1 port map( A => n14585, ZN => n8993);
   U9289 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_210_port, B2 => n2544, 
                           ZN => n14585);
   U9290 : INV_X1 port map( A => n14584, ZN => n8994);
   U9291 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_209_port, B2 => n2544, 
                           ZN => n14584);
   U9292 : INV_X1 port map( A => n14583, ZN => n8995);
   U9293 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_208_port, B2 => n2544, 
                           ZN => n14583);
   U9294 : INV_X1 port map( A => n14582, ZN => n8996);
   U9295 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_207_port, B2 => n2544, 
                           ZN => n14582);
   U9296 : INV_X1 port map( A => n14581, ZN => n8997);
   U9297 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_206_port, B2 => n2544, 
                           ZN => n14581);
   U9298 : INV_X1 port map( A => n14580, ZN => n8998);
   U9299 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_205_port, B2 => n2544, 
                           ZN => n14580);
   U9300 : INV_X1 port map( A => n14579, ZN => n8999);
   U9301 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_204_port, B2 => n2544, 
                           ZN => n14579);
   U9302 : INV_X1 port map( A => n14578, ZN => n9000);
   U9303 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_203_port, B2 => n2543, 
                           ZN => n14578);
   U9304 : INV_X1 port map( A => n14577, ZN => n9001);
   U9305 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_202_port, B2 => n2543, 
                           ZN => n14577);
   U9306 : INV_X1 port map( A => n14576, ZN => n9002);
   U9307 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_201_port, B2 => n2543, 
                           ZN => n14576);
   U9308 : INV_X1 port map( A => n14575, ZN => n9003);
   U9309 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2541, B1 => 
                           DataPath_RF_bus_reg_dataout_200_port, B2 => n2543, 
                           ZN => n14575);
   U9310 : INV_X1 port map( A => n14574, ZN => n9004);
   U9311 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_199_port, B2 => n2543, 
                           ZN => n14574);
   U9312 : INV_X1 port map( A => n14573, ZN => n9005);
   U9313 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_198_port, B2 => n2543, 
                           ZN => n14573);
   U9314 : INV_X1 port map( A => n14572, ZN => n9006);
   U9315 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_197_port, B2 => n2543, 
                           ZN => n14572);
   U9316 : INV_X1 port map( A => n14571, ZN => n9007);
   U9317 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_196_port, B2 => n2543, 
                           ZN => n14571);
   U9318 : INV_X1 port map( A => n14570, ZN => n9008);
   U9319 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_195_port, B2 => n2543, 
                           ZN => n14570);
   U9320 : INV_X1 port map( A => n14569, ZN => n9009);
   U9321 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_194_port, B2 => n2543, 
                           ZN => n14569);
   U9322 : INV_X1 port map( A => n14568, ZN => n9010);
   U9323 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_193_port, B2 => n2543, 
                           ZN => n14568);
   U9324 : INV_X1 port map( A => n14565, ZN => n9011);
   U9325 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2542, B1 => 
                           DataPath_RF_bus_reg_dataout_192_port, B2 => n2543, 
                           ZN => n14565);
   U9326 : INV_X1 port map( A => n14632, ZN => n9012);
   U9327 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_255_port, B2 => n2551, 
                           ZN => n14632);
   U9328 : INV_X1 port map( A => n14631, ZN => n9013);
   U9329 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_254_port, B2 => n2551, 
                           ZN => n14631);
   U9330 : INV_X1 port map( A => n14630, ZN => n9014);
   U9331 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_253_port, B2 => n2551, 
                           ZN => n14630);
   U9332 : INV_X1 port map( A => n14629, ZN => n9015);
   U9333 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_252_port, B2 => n2551, 
                           ZN => n14629);
   U9334 : INV_X1 port map( A => n14628, ZN => n9016);
   U9335 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_251_port, B2 => n2551, 
                           ZN => n14628);
   U9336 : INV_X1 port map( A => n14627, ZN => n9017);
   U9337 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_250_port, B2 => n2551, 
                           ZN => n14627);
   U9338 : INV_X1 port map( A => n14626, ZN => n9018);
   U9339 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_249_port, B2 => n2551, 
                           ZN => n14626);
   U9340 : INV_X1 port map( A => n14625, ZN => n9019);
   U9341 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_248_port, B2 => n2551, 
                           ZN => n14625);
   U9342 : INV_X1 port map( A => n14624, ZN => n9020);
   U9343 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_247_port, B2 => n2550, 
                           ZN => n14624);
   U9344 : INV_X1 port map( A => n14623, ZN => n9021);
   U9345 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_246_port, B2 => n2550, 
                           ZN => n14623);
   U9346 : INV_X1 port map( A => n14622, ZN => n9022);
   U9347 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_245_port, B2 => n2550, 
                           ZN => n14622);
   U9348 : INV_X1 port map( A => n14621, ZN => n9023);
   U9349 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2546, B1 => 
                           DataPath_RF_bus_reg_dataout_244_port, B2 => n2550, 
                           ZN => n14621);
   U9350 : INV_X1 port map( A => n14620, ZN => n9024);
   U9351 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_243_port, B2 => n2550, 
                           ZN => n14620);
   U9352 : INV_X1 port map( A => n14619, ZN => n9025);
   U9353 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_242_port, B2 => n2550, 
                           ZN => n14619);
   U9354 : INV_X1 port map( A => n14618, ZN => n9026);
   U9355 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_241_port, B2 => n2550, 
                           ZN => n14618);
   U9356 : INV_X1 port map( A => n14617, ZN => n9027);
   U9357 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_240_port, B2 => n2550, 
                           ZN => n14617);
   U9358 : INV_X1 port map( A => n14616, ZN => n9028);
   U9359 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_239_port, B2 => n2550, 
                           ZN => n14616);
   U9360 : INV_X1 port map( A => n14615, ZN => n9029);
   U9361 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_238_port, B2 => n2550, 
                           ZN => n14615);
   U9362 : INV_X1 port map( A => n14614, ZN => n9030);
   U9363 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_237_port, B2 => n2550, 
                           ZN => n14614);
   U9364 : INV_X1 port map( A => n14613, ZN => n9031);
   U9365 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_236_port, B2 => n2550, 
                           ZN => n14613);
   U9366 : INV_X1 port map( A => n14612, ZN => n9032);
   U9367 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_235_port, B2 => n2549, 
                           ZN => n14612);
   U9368 : INV_X1 port map( A => n14611, ZN => n9033);
   U9369 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_234_port, B2 => n2549, 
                           ZN => n14611);
   U9370 : INV_X1 port map( A => n14610, ZN => n9034);
   U9371 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_233_port, B2 => n2549, 
                           ZN => n14610);
   U9372 : INV_X1 port map( A => n14609, ZN => n9035);
   U9373 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2547, B1 => 
                           DataPath_RF_bus_reg_dataout_232_port, B2 => n2549, 
                           ZN => n14609);
   U9374 : INV_X1 port map( A => n14608, ZN => n9036);
   U9375 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_231_port, B2 => n2549, 
                           ZN => n14608);
   U9376 : INV_X1 port map( A => n14607, ZN => n9037);
   U9377 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_230_port, B2 => n2549, 
                           ZN => n14607);
   U9378 : INV_X1 port map( A => n14606, ZN => n9038);
   U9379 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_229_port, B2 => n2549, 
                           ZN => n14606);
   U9380 : INV_X1 port map( A => n14605, ZN => n9039);
   U9381 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_228_port, B2 => n2549, 
                           ZN => n14605);
   U9382 : INV_X1 port map( A => n14604, ZN => n9040);
   U9383 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_227_port, B2 => n2549, 
                           ZN => n14604);
   U9384 : INV_X1 port map( A => n14603, ZN => n9041);
   U9385 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_226_port, B2 => n2549, 
                           ZN => n14603);
   U9386 : INV_X1 port map( A => n14602, ZN => n9042);
   U9387 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_225_port, B2 => n2549, 
                           ZN => n14602);
   U9388 : INV_X1 port map( A => n14599, ZN => n9043);
   U9389 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2548, B1 => 
                           DataPath_RF_bus_reg_dataout_224_port, B2 => n2549, 
                           ZN => n14599);
   U9390 : INV_X1 port map( A => n14666, ZN => n9044);
   U9391 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_287_port, B2 => n2557, 
                           ZN => n14666);
   U9392 : INV_X1 port map( A => n14665, ZN => n9045);
   U9393 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_286_port, B2 => n2557, 
                           ZN => n14665);
   U9394 : INV_X1 port map( A => n14664, ZN => n9046);
   U9395 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_285_port, B2 => n2557, 
                           ZN => n14664);
   U9396 : INV_X1 port map( A => n14663, ZN => n9047);
   U9397 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_284_port, B2 => n2557, 
                           ZN => n14663);
   U9398 : INV_X1 port map( A => n14662, ZN => n9048);
   U9399 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_283_port, B2 => n2557, 
                           ZN => n14662);
   U9400 : INV_X1 port map( A => n14661, ZN => n9049);
   U9401 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_282_port, B2 => n2557, 
                           ZN => n14661);
   U9402 : INV_X1 port map( A => n14660, ZN => n9050);
   U9403 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_281_port, B2 => n2557, 
                           ZN => n14660);
   U9404 : INV_X1 port map( A => n14659, ZN => n9051);
   U9405 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_280_port, B2 => n2557, 
                           ZN => n14659);
   U9406 : INV_X1 port map( A => n14658, ZN => n9052);
   U9407 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_279_port, B2 => n2556, 
                           ZN => n14658);
   U9408 : INV_X1 port map( A => n14657, ZN => n9053);
   U9409 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_278_port, B2 => n2556, 
                           ZN => n14657);
   U9410 : INV_X1 port map( A => n14656, ZN => n9054);
   U9411 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_277_port, B2 => n2556, 
                           ZN => n14656);
   U9412 : INV_X1 port map( A => n14655, ZN => n9055);
   U9413 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2552, B1 => 
                           DataPath_RF_bus_reg_dataout_276_port, B2 => n2556, 
                           ZN => n14655);
   U9414 : INV_X1 port map( A => n14654, ZN => n9056);
   U9415 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_275_port, B2 => n2556, 
                           ZN => n14654);
   U9416 : INV_X1 port map( A => n14653, ZN => n9057);
   U9417 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_274_port, B2 => n2556, 
                           ZN => n14653);
   U9418 : INV_X1 port map( A => n14652, ZN => n9058);
   U9419 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_273_port, B2 => n2556, 
                           ZN => n14652);
   U9420 : INV_X1 port map( A => n14651, ZN => n9059);
   U9421 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_272_port, B2 => n2556, 
                           ZN => n14651);
   U9422 : INV_X1 port map( A => n14650, ZN => n9060);
   U9423 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_271_port, B2 => n2556, 
                           ZN => n14650);
   U9424 : INV_X1 port map( A => n14649, ZN => n9061);
   U9425 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_270_port, B2 => n2556, 
                           ZN => n14649);
   U9426 : INV_X1 port map( A => n14648, ZN => n9062);
   U9427 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_269_port, B2 => n2556, 
                           ZN => n14648);
   U9428 : INV_X1 port map( A => n14647, ZN => n9063);
   U9429 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_268_port, B2 => n2556, 
                           ZN => n14647);
   U9430 : INV_X1 port map( A => n14646, ZN => n9064);
   U9431 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_267_port, B2 => n2555, 
                           ZN => n14646);
   U9432 : INV_X1 port map( A => n14645, ZN => n9065);
   U9433 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_266_port, B2 => n2555, 
                           ZN => n14645);
   U9434 : INV_X1 port map( A => n14644, ZN => n9066);
   U9435 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_265_port, B2 => n2555, 
                           ZN => n14644);
   U9436 : INV_X1 port map( A => n14643, ZN => n9067);
   U9437 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2553, B1 => 
                           DataPath_RF_bus_reg_dataout_264_port, B2 => n2555, 
                           ZN => n14643);
   U9438 : INV_X1 port map( A => n14642, ZN => n9068);
   U9439 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_263_port, B2 => n2555, 
                           ZN => n14642);
   U9440 : INV_X1 port map( A => n14641, ZN => n9069);
   U9441 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_262_port, B2 => n2555, 
                           ZN => n14641);
   U9442 : INV_X1 port map( A => n14640, ZN => n9070);
   U9443 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_261_port, B2 => n2555, 
                           ZN => n14640);
   U9444 : INV_X1 port map( A => n14639, ZN => n9071);
   U9445 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_260_port, B2 => n2555, 
                           ZN => n14639);
   U9446 : INV_X1 port map( A => n14638, ZN => n9072);
   U9447 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_259_port, B2 => n2555, 
                           ZN => n14638);
   U9448 : INV_X1 port map( A => n14637, ZN => n9073);
   U9449 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_258_port, B2 => n2555, 
                           ZN => n14637);
   U9450 : INV_X1 port map( A => n14636, ZN => n9074);
   U9451 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_257_port, B2 => n2555, 
                           ZN => n14636);
   U9452 : INV_X1 port map( A => n14633, ZN => n9075);
   U9453 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2554, B1 => 
                           DataPath_RF_bus_reg_dataout_256_port, B2 => n2555, 
                           ZN => n14633);
   U9454 : INV_X1 port map( A => n14700, ZN => n9076);
   U9455 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_319_port, B2 => n2563, 
                           ZN => n14700);
   U9456 : INV_X1 port map( A => n14699, ZN => n9077);
   U9457 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_318_port, B2 => n2563, 
                           ZN => n14699);
   U9458 : INV_X1 port map( A => n14698, ZN => n9078);
   U9459 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_317_port, B2 => n2563, 
                           ZN => n14698);
   U9460 : INV_X1 port map( A => n14697, ZN => n9079);
   U9461 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_316_port, B2 => n2563, 
                           ZN => n14697);
   U9462 : INV_X1 port map( A => n14696, ZN => n9080);
   U9463 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_315_port, B2 => n2563, 
                           ZN => n14696);
   U9464 : INV_X1 port map( A => n14695, ZN => n9081);
   U9465 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_314_port, B2 => n2563, 
                           ZN => n14695);
   U9466 : INV_X1 port map( A => n14694, ZN => n9082);
   U9467 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_313_port, B2 => n2563, 
                           ZN => n14694);
   U9468 : INV_X1 port map( A => n14693, ZN => n9083);
   U9469 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_312_port, B2 => n2563, 
                           ZN => n14693);
   U9470 : INV_X1 port map( A => n14692, ZN => n9084);
   U9471 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_311_port, B2 => n2562, 
                           ZN => n14692);
   U9472 : INV_X1 port map( A => n14691, ZN => n9085);
   U9473 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_310_port, B2 => n2562, 
                           ZN => n14691);
   U9474 : INV_X1 port map( A => n14690, ZN => n9086);
   U9475 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_309_port, B2 => n2562, 
                           ZN => n14690);
   U9476 : INV_X1 port map( A => n14689, ZN => n9087);
   U9477 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2558, B1 => 
                           DataPath_RF_bus_reg_dataout_308_port, B2 => n2562, 
                           ZN => n14689);
   U9478 : INV_X1 port map( A => n14688, ZN => n9088);
   U9479 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_307_port, B2 => n2562, 
                           ZN => n14688);
   U9480 : INV_X1 port map( A => n14687, ZN => n9089);
   U9481 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_306_port, B2 => n2562, 
                           ZN => n14687);
   U9482 : INV_X1 port map( A => n14686, ZN => n9090);
   U9483 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_305_port, B2 => n2562, 
                           ZN => n14686);
   U9484 : INV_X1 port map( A => n14685, ZN => n9091);
   U9485 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_304_port, B2 => n2562, 
                           ZN => n14685);
   U9486 : INV_X1 port map( A => n14684, ZN => n9092);
   U9487 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_303_port, B2 => n2562, 
                           ZN => n14684);
   U9488 : INV_X1 port map( A => n14683, ZN => n9093);
   U9489 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_302_port, B2 => n2562, 
                           ZN => n14683);
   U9490 : INV_X1 port map( A => n14682, ZN => n9094);
   U9491 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_301_port, B2 => n2562, 
                           ZN => n14682);
   U9492 : INV_X1 port map( A => n14681, ZN => n9095);
   U9493 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_300_port, B2 => n2562, 
                           ZN => n14681);
   U9494 : INV_X1 port map( A => n14680, ZN => n9096);
   U9495 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_299_port, B2 => n2561, 
                           ZN => n14680);
   U9496 : INV_X1 port map( A => n14679, ZN => n9097);
   U9497 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_298_port, B2 => n2561, 
                           ZN => n14679);
   U9498 : INV_X1 port map( A => n14678, ZN => n9098);
   U9499 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_297_port, B2 => n2561, 
                           ZN => n14678);
   U9500 : INV_X1 port map( A => n14677, ZN => n9099);
   U9501 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2559, B1 => 
                           DataPath_RF_bus_reg_dataout_296_port, B2 => n2561, 
                           ZN => n14677);
   U9502 : INV_X1 port map( A => n14676, ZN => n9100);
   U9503 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_295_port, B2 => n2561, 
                           ZN => n14676);
   U9504 : INV_X1 port map( A => n14675, ZN => n9101);
   U9505 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_294_port, B2 => n2561, 
                           ZN => n14675);
   U9506 : INV_X1 port map( A => n14674, ZN => n9102);
   U9507 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_293_port, B2 => n2561, 
                           ZN => n14674);
   U9508 : INV_X1 port map( A => n14673, ZN => n9103);
   U9509 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_292_port, B2 => n2561, 
                           ZN => n14673);
   U9510 : INV_X1 port map( A => n14672, ZN => n9104);
   U9511 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_291_port, B2 => n2561, 
                           ZN => n14672);
   U9512 : INV_X1 port map( A => n14671, ZN => n9105);
   U9513 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_290_port, B2 => n2561, 
                           ZN => n14671);
   U9514 : INV_X1 port map( A => n14670, ZN => n9106);
   U9515 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_289_port, B2 => n2561, 
                           ZN => n14670);
   U9516 : INV_X1 port map( A => n14667, ZN => n9107);
   U9517 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2560, B1 => 
                           DataPath_RF_bus_reg_dataout_288_port, B2 => n2561, 
                           ZN => n14667);
   U9518 : INV_X1 port map( A => n14734, ZN => n9108);
   U9519 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_351_port, B2 => n2569, 
                           ZN => n14734);
   U9520 : INV_X1 port map( A => n14733, ZN => n9109);
   U9521 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_350_port, B2 => n2569, 
                           ZN => n14733);
   U9522 : INV_X1 port map( A => n14732, ZN => n9110);
   U9523 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_349_port, B2 => n2569, 
                           ZN => n14732);
   U9524 : INV_X1 port map( A => n14731, ZN => n9111);
   U9525 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_348_port, B2 => n2569, 
                           ZN => n14731);
   U9526 : INV_X1 port map( A => n14730, ZN => n9112);
   U9527 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_347_port, B2 => n2569, 
                           ZN => n14730);
   U9528 : INV_X1 port map( A => n14729, ZN => n9113);
   U9529 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_346_port, B2 => n2569, 
                           ZN => n14729);
   U9530 : INV_X1 port map( A => n14728, ZN => n9114);
   U9531 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_345_port, B2 => n2569, 
                           ZN => n14728);
   U9532 : INV_X1 port map( A => n14727, ZN => n9115);
   U9533 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_344_port, B2 => n2569, 
                           ZN => n14727);
   U9534 : INV_X1 port map( A => n14726, ZN => n9116);
   U9535 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_343_port, B2 => n2568, 
                           ZN => n14726);
   U9536 : INV_X1 port map( A => n14725, ZN => n9117);
   U9537 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_342_port, B2 => n2568, 
                           ZN => n14725);
   U9538 : INV_X1 port map( A => n14724, ZN => n9118);
   U9539 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_341_port, B2 => n2568, 
                           ZN => n14724);
   U9540 : INV_X1 port map( A => n14723, ZN => n9119);
   U9541 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2564, B1 => 
                           DataPath_RF_bus_reg_dataout_340_port, B2 => n2568, 
                           ZN => n14723);
   U9542 : INV_X1 port map( A => n14722, ZN => n9120);
   U9543 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_339_port, B2 => n2568, 
                           ZN => n14722);
   U9544 : INV_X1 port map( A => n14721, ZN => n9121);
   U9545 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_338_port, B2 => n2568, 
                           ZN => n14721);
   U9546 : INV_X1 port map( A => n14720, ZN => n9122);
   U9547 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_337_port, B2 => n2568, 
                           ZN => n14720);
   U9548 : INV_X1 port map( A => n14719, ZN => n9123);
   U9549 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_336_port, B2 => n2568, 
                           ZN => n14719);
   U9550 : INV_X1 port map( A => n14718, ZN => n9124);
   U9551 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_335_port, B2 => n2568, 
                           ZN => n14718);
   U9552 : INV_X1 port map( A => n14717, ZN => n9125);
   U9553 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_334_port, B2 => n2568, 
                           ZN => n14717);
   U9554 : INV_X1 port map( A => n14716, ZN => n9126);
   U9555 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_333_port, B2 => n2568, 
                           ZN => n14716);
   U9556 : INV_X1 port map( A => n14715, ZN => n9127);
   U9557 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_332_port, B2 => n2568, 
                           ZN => n14715);
   U9558 : INV_X1 port map( A => n14714, ZN => n9128);
   U9559 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_331_port, B2 => n2567, 
                           ZN => n14714);
   U9560 : INV_X1 port map( A => n14713, ZN => n9129);
   U9561 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_330_port, B2 => n2567, 
                           ZN => n14713);
   U9562 : INV_X1 port map( A => n14712, ZN => n9130);
   U9563 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_329_port, B2 => n2567, 
                           ZN => n14712);
   U9564 : INV_X1 port map( A => n14711, ZN => n9131);
   U9565 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2565, B1 => 
                           DataPath_RF_bus_reg_dataout_328_port, B2 => n2567, 
                           ZN => n14711);
   U9566 : INV_X1 port map( A => n14710, ZN => n9132);
   U9567 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_327_port, B2 => n2567, 
                           ZN => n14710);
   U9568 : INV_X1 port map( A => n14709, ZN => n9133);
   U9569 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_326_port, B2 => n2567, 
                           ZN => n14709);
   U9570 : INV_X1 port map( A => n14708, ZN => n9134);
   U9571 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_325_port, B2 => n2567, 
                           ZN => n14708);
   U9572 : INV_X1 port map( A => n14707, ZN => n9135);
   U9573 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_324_port, B2 => n2567, 
                           ZN => n14707);
   U9574 : INV_X1 port map( A => n14706, ZN => n9136);
   U9575 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_323_port, B2 => n2567, 
                           ZN => n14706);
   U9576 : INV_X1 port map( A => n14705, ZN => n9137);
   U9577 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_322_port, B2 => n2567, 
                           ZN => n14705);
   U9578 : INV_X1 port map( A => n14704, ZN => n9138);
   U9579 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_321_port, B2 => n2567, 
                           ZN => n14704);
   U9580 : INV_X1 port map( A => n14701, ZN => n9139);
   U9581 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2566, B1 => 
                           DataPath_RF_bus_reg_dataout_320_port, B2 => n2567, 
                           ZN => n14701);
   U9582 : INV_X1 port map( A => n14768, ZN => n9140);
   U9583 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_383_port, B2 => n2575, 
                           ZN => n14768);
   U9584 : INV_X1 port map( A => n14767, ZN => n9141);
   U9585 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_382_port, B2 => n2575, 
                           ZN => n14767);
   U9586 : INV_X1 port map( A => n14766, ZN => n9142);
   U9587 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_381_port, B2 => n2575, 
                           ZN => n14766);
   U9588 : INV_X1 port map( A => n14765, ZN => n9143);
   U9589 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_380_port, B2 => n2575, 
                           ZN => n14765);
   U9590 : INV_X1 port map( A => n14764, ZN => n9144);
   U9591 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_379_port, B2 => n2575, 
                           ZN => n14764);
   U9592 : INV_X1 port map( A => n14763, ZN => n9145);
   U9593 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_378_port, B2 => n2575, 
                           ZN => n14763);
   U9594 : INV_X1 port map( A => n14762, ZN => n9146);
   U9595 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_377_port, B2 => n2575, 
                           ZN => n14762);
   U9596 : INV_X1 port map( A => n14761, ZN => n9147);
   U9597 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_376_port, B2 => n2575, 
                           ZN => n14761);
   U9598 : INV_X1 port map( A => n14760, ZN => n9148);
   U9599 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_375_port, B2 => n2574, 
                           ZN => n14760);
   U9600 : INV_X1 port map( A => n14759, ZN => n9149);
   U9601 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_374_port, B2 => n2574, 
                           ZN => n14759);
   U9602 : INV_X1 port map( A => n14758, ZN => n9150);
   U9603 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_373_port, B2 => n2574, 
                           ZN => n14758);
   U9604 : INV_X1 port map( A => n14757, ZN => n9151);
   U9605 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2570, B1 => 
                           DataPath_RF_bus_reg_dataout_372_port, B2 => n2574, 
                           ZN => n14757);
   U9606 : INV_X1 port map( A => n14756, ZN => n9152);
   U9607 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_371_port, B2 => n2574, 
                           ZN => n14756);
   U9608 : INV_X1 port map( A => n14755, ZN => n9153);
   U9609 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_370_port, B2 => n2574, 
                           ZN => n14755);
   U9610 : INV_X1 port map( A => n14754, ZN => n9154);
   U9611 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_369_port, B2 => n2574, 
                           ZN => n14754);
   U9612 : INV_X1 port map( A => n14753, ZN => n9155);
   U9613 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_368_port, B2 => n2574, 
                           ZN => n14753);
   U9614 : INV_X1 port map( A => n14752, ZN => n9156);
   U9615 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_367_port, B2 => n2574, 
                           ZN => n14752);
   U9616 : INV_X1 port map( A => n14751, ZN => n9157);
   U9617 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_366_port, B2 => n2574, 
                           ZN => n14751);
   U9618 : INV_X1 port map( A => n14750, ZN => n9158);
   U9619 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_365_port, B2 => n2574, 
                           ZN => n14750);
   U9620 : INV_X1 port map( A => n14749, ZN => n9159);
   U9621 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_364_port, B2 => n2574, 
                           ZN => n14749);
   U9622 : INV_X1 port map( A => n14748, ZN => n9160);
   U9623 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_363_port, B2 => n2573, 
                           ZN => n14748);
   U9624 : INV_X1 port map( A => n14747, ZN => n9161);
   U9625 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_362_port, B2 => n2573, 
                           ZN => n14747);
   U9626 : INV_X1 port map( A => n14746, ZN => n9162);
   U9627 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_361_port, B2 => n2573, 
                           ZN => n14746);
   U9628 : INV_X1 port map( A => n14745, ZN => n9163);
   U9629 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2571, B1 => 
                           DataPath_RF_bus_reg_dataout_360_port, B2 => n2573, 
                           ZN => n14745);
   U9630 : INV_X1 port map( A => n14744, ZN => n9164);
   U9631 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_359_port, B2 => n2573, 
                           ZN => n14744);
   U9632 : INV_X1 port map( A => n14743, ZN => n9165);
   U9633 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_358_port, B2 => n2573, 
                           ZN => n14743);
   U9634 : INV_X1 port map( A => n14742, ZN => n9166);
   U9635 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_357_port, B2 => n2573, 
                           ZN => n14742);
   U9636 : INV_X1 port map( A => n14741, ZN => n9167);
   U9637 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_356_port, B2 => n2573, 
                           ZN => n14741);
   U9638 : INV_X1 port map( A => n14740, ZN => n9168);
   U9639 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_355_port, B2 => n2573, 
                           ZN => n14740);
   U9640 : INV_X1 port map( A => n14739, ZN => n9169);
   U9641 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_354_port, B2 => n2573, 
                           ZN => n14739);
   U9642 : INV_X1 port map( A => n14738, ZN => n9170);
   U9643 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_353_port, B2 => n2573, 
                           ZN => n14738);
   U9644 : INV_X1 port map( A => n14735, ZN => n9171);
   U9645 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2572, B1 => 
                           DataPath_RF_bus_reg_dataout_352_port, B2 => n2573, 
                           ZN => n14735);
   U9646 : INV_X1 port map( A => n14802, ZN => n9172);
   U9647 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_415_port, B2 => n2581, 
                           ZN => n14802);
   U9648 : INV_X1 port map( A => n14801, ZN => n9173);
   U9649 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_414_port, B2 => n2581, 
                           ZN => n14801);
   U9650 : INV_X1 port map( A => n14800, ZN => n9174);
   U9651 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_413_port, B2 => n2581, 
                           ZN => n14800);
   U9652 : INV_X1 port map( A => n14799, ZN => n9175);
   U9653 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_412_port, B2 => n2581, 
                           ZN => n14799);
   U9654 : INV_X1 port map( A => n14798, ZN => n9176);
   U9655 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_411_port, B2 => n2581, 
                           ZN => n14798);
   U9656 : INV_X1 port map( A => n14797, ZN => n9177);
   U9657 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_410_port, B2 => n2581, 
                           ZN => n14797);
   U9658 : INV_X1 port map( A => n14796, ZN => n9178);
   U9659 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_409_port, B2 => n2581, 
                           ZN => n14796);
   U9660 : INV_X1 port map( A => n14795, ZN => n9179);
   U9661 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_408_port, B2 => n2581, 
                           ZN => n14795);
   U9662 : INV_X1 port map( A => n14794, ZN => n9180);
   U9663 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_407_port, B2 => n2580, 
                           ZN => n14794);
   U9664 : INV_X1 port map( A => n14793, ZN => n9181);
   U9665 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_406_port, B2 => n2580, 
                           ZN => n14793);
   U9666 : INV_X1 port map( A => n14792, ZN => n9182);
   U9667 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_405_port, B2 => n2580, 
                           ZN => n14792);
   U9668 : INV_X1 port map( A => n14791, ZN => n9183);
   U9669 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2576, B1 => 
                           DataPath_RF_bus_reg_dataout_404_port, B2 => n2580, 
                           ZN => n14791);
   U9670 : INV_X1 port map( A => n14790, ZN => n9184);
   U9671 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_403_port, B2 => n2580, 
                           ZN => n14790);
   U9672 : INV_X1 port map( A => n14789, ZN => n9185);
   U9673 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_402_port, B2 => n2580, 
                           ZN => n14789);
   U9674 : INV_X1 port map( A => n14788, ZN => n9186);
   U9675 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_401_port, B2 => n2580, 
                           ZN => n14788);
   U9676 : INV_X1 port map( A => n14787, ZN => n9187);
   U9677 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_400_port, B2 => n2580, 
                           ZN => n14787);
   U9678 : INV_X1 port map( A => n14786, ZN => n9188);
   U9679 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_399_port, B2 => n2580, 
                           ZN => n14786);
   U9680 : INV_X1 port map( A => n14785, ZN => n9189);
   U9681 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_398_port, B2 => n2580, 
                           ZN => n14785);
   U9682 : INV_X1 port map( A => n14784, ZN => n9190);
   U9683 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_397_port, B2 => n2580, 
                           ZN => n14784);
   U9684 : INV_X1 port map( A => n14783, ZN => n9191);
   U9685 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_396_port, B2 => n2580, 
                           ZN => n14783);
   U9686 : INV_X1 port map( A => n14782, ZN => n9192);
   U9687 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_395_port, B2 => n2579, 
                           ZN => n14782);
   U9688 : INV_X1 port map( A => n14781, ZN => n9193);
   U9689 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_394_port, B2 => n2579, 
                           ZN => n14781);
   U9690 : INV_X1 port map( A => n14780, ZN => n9194);
   U9691 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_393_port, B2 => n2579, 
                           ZN => n14780);
   U9692 : INV_X1 port map( A => n14779, ZN => n9195);
   U9693 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2577, B1 => 
                           DataPath_RF_bus_reg_dataout_392_port, B2 => n2579, 
                           ZN => n14779);
   U9694 : INV_X1 port map( A => n14778, ZN => n9196);
   U9695 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_391_port, B2 => n2579, 
                           ZN => n14778);
   U9696 : INV_X1 port map( A => n14777, ZN => n9197);
   U9697 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_390_port, B2 => n2579, 
                           ZN => n14777);
   U9698 : INV_X1 port map( A => n14776, ZN => n9198);
   U9699 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_389_port, B2 => n2579, 
                           ZN => n14776);
   U9700 : INV_X1 port map( A => n14775, ZN => n9199);
   U9701 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_388_port, B2 => n2579, 
                           ZN => n14775);
   U9702 : INV_X1 port map( A => n14774, ZN => n9200);
   U9703 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_387_port, B2 => n2579, 
                           ZN => n14774);
   U9704 : INV_X1 port map( A => n14773, ZN => n9201);
   U9705 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_386_port, B2 => n2579, 
                           ZN => n14773);
   U9706 : INV_X1 port map( A => n14772, ZN => n9202);
   U9707 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_385_port, B2 => n2579, 
                           ZN => n14772);
   U9708 : INV_X1 port map( A => n14769, ZN => n9203);
   U9709 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2578, B1 => 
                           DataPath_RF_bus_reg_dataout_384_port, B2 => n2579, 
                           ZN => n14769);
   U9710 : INV_X1 port map( A => n14836, ZN => n9204);
   U9711 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_447_port, B2 => n2587, 
                           ZN => n14836);
   U9712 : INV_X1 port map( A => n14835, ZN => n9205);
   U9713 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_446_port, B2 => n2587, 
                           ZN => n14835);
   U9714 : INV_X1 port map( A => n14834, ZN => n9206);
   U9715 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_445_port, B2 => n2587, 
                           ZN => n14834);
   U9716 : INV_X1 port map( A => n14833, ZN => n9207);
   U9717 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_444_port, B2 => n2587, 
                           ZN => n14833);
   U9718 : INV_X1 port map( A => n14832, ZN => n9208);
   U9719 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_443_port, B2 => n2587, 
                           ZN => n14832);
   U9720 : INV_X1 port map( A => n14831, ZN => n9209);
   U9721 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_442_port, B2 => n2587, 
                           ZN => n14831);
   U9722 : INV_X1 port map( A => n14830, ZN => n9210);
   U9723 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_441_port, B2 => n2587, 
                           ZN => n14830);
   U9724 : INV_X1 port map( A => n14829, ZN => n9211);
   U9725 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_440_port, B2 => n2587, 
                           ZN => n14829);
   U9726 : INV_X1 port map( A => n14828, ZN => n9212);
   U9727 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_439_port, B2 => n2586, 
                           ZN => n14828);
   U9728 : INV_X1 port map( A => n14827, ZN => n9213);
   U9729 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_438_port, B2 => n2586, 
                           ZN => n14827);
   U9730 : INV_X1 port map( A => n14826, ZN => n9214);
   U9731 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_437_port, B2 => n2586, 
                           ZN => n14826);
   U9732 : INV_X1 port map( A => n14825, ZN => n9215);
   U9733 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2582, B1 => 
                           DataPath_RF_bus_reg_dataout_436_port, B2 => n2586, 
                           ZN => n14825);
   U9734 : INV_X1 port map( A => n14824, ZN => n9216);
   U9735 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_435_port, B2 => n2586, 
                           ZN => n14824);
   U9736 : INV_X1 port map( A => n14823, ZN => n9217);
   U9737 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_434_port, B2 => n2586, 
                           ZN => n14823);
   U9738 : INV_X1 port map( A => n14822, ZN => n9218);
   U9739 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_433_port, B2 => n2586, 
                           ZN => n14822);
   U9740 : INV_X1 port map( A => n14821, ZN => n9219);
   U9741 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_432_port, B2 => n2586, 
                           ZN => n14821);
   U9742 : INV_X1 port map( A => n14820, ZN => n9220);
   U9743 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_431_port, B2 => n2586, 
                           ZN => n14820);
   U9744 : INV_X1 port map( A => n14819, ZN => n9221);
   U9745 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_430_port, B2 => n2586, 
                           ZN => n14819);
   U9746 : INV_X1 port map( A => n14818, ZN => n9222);
   U9747 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_429_port, B2 => n2586, 
                           ZN => n14818);
   U9748 : INV_X1 port map( A => n14817, ZN => n9223);
   U9749 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_428_port, B2 => n2586, 
                           ZN => n14817);
   U9750 : INV_X1 port map( A => n14816, ZN => n9224);
   U9751 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_427_port, B2 => n2585, 
                           ZN => n14816);
   U9752 : INV_X1 port map( A => n14815, ZN => n9225);
   U9753 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_426_port, B2 => n2585, 
                           ZN => n14815);
   U9754 : INV_X1 port map( A => n14814, ZN => n9226);
   U9755 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_425_port, B2 => n2585, 
                           ZN => n14814);
   U9756 : INV_X1 port map( A => n14813, ZN => n9227);
   U9757 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2583, B1 => 
                           DataPath_RF_bus_reg_dataout_424_port, B2 => n2585, 
                           ZN => n14813);
   U9758 : INV_X1 port map( A => n14812, ZN => n9228);
   U9759 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_423_port, B2 => n2585, 
                           ZN => n14812);
   U9760 : INV_X1 port map( A => n14811, ZN => n9229);
   U9761 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_422_port, B2 => n2585, 
                           ZN => n14811);
   U9762 : INV_X1 port map( A => n14810, ZN => n9230);
   U9763 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_421_port, B2 => n2585, 
                           ZN => n14810);
   U9764 : INV_X1 port map( A => n14809, ZN => n9231);
   U9765 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_420_port, B2 => n2585, 
                           ZN => n14809);
   U9766 : INV_X1 port map( A => n14808, ZN => n9232);
   U9767 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_419_port, B2 => n2585, 
                           ZN => n14808);
   U9768 : INV_X1 port map( A => n14807, ZN => n9233);
   U9769 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_418_port, B2 => n2585, 
                           ZN => n14807);
   U9770 : INV_X1 port map( A => n14806, ZN => n9234);
   U9771 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_417_port, B2 => n2585, 
                           ZN => n14806);
   U9772 : INV_X1 port map( A => n14803, ZN => n9235);
   U9773 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2584, B1 => 
                           DataPath_RF_bus_reg_dataout_416_port, B2 => n2585, 
                           ZN => n14803);
   U9774 : INV_X1 port map( A => n14870, ZN => n9236);
   U9775 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_479_port, B2 => n2593, 
                           ZN => n14870);
   U9776 : INV_X1 port map( A => n14869, ZN => n9237);
   U9777 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_478_port, B2 => n2593, 
                           ZN => n14869);
   U9778 : INV_X1 port map( A => n14868, ZN => n9238);
   U9779 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_477_port, B2 => n2593, 
                           ZN => n14868);
   U9780 : INV_X1 port map( A => n14867, ZN => n9239);
   U9781 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_476_port, B2 => n2593, 
                           ZN => n14867);
   U9782 : INV_X1 port map( A => n14866, ZN => n9240);
   U9783 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_475_port, B2 => n2593, 
                           ZN => n14866);
   U9784 : INV_X1 port map( A => n14865, ZN => n9241);
   U9785 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_474_port, B2 => n2593, 
                           ZN => n14865);
   U9786 : INV_X1 port map( A => n14864, ZN => n9242);
   U9787 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_473_port, B2 => n2593, 
                           ZN => n14864);
   U9788 : INV_X1 port map( A => n14863, ZN => n9243);
   U9789 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_472_port, B2 => n2593, 
                           ZN => n14863);
   U9790 : INV_X1 port map( A => n14862, ZN => n9244);
   U9791 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_471_port, B2 => n2592, 
                           ZN => n14862);
   U9792 : INV_X1 port map( A => n14861, ZN => n9245);
   U9793 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_470_port, B2 => n2592, 
                           ZN => n14861);
   U9794 : INV_X1 port map( A => n14860, ZN => n9246);
   U9795 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_469_port, B2 => n2592, 
                           ZN => n14860);
   U9796 : INV_X1 port map( A => n14859, ZN => n9247);
   U9797 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2588, B1 => 
                           DataPath_RF_bus_reg_dataout_468_port, B2 => n2592, 
                           ZN => n14859);
   U9798 : INV_X1 port map( A => n14858, ZN => n9248);
   U9799 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_467_port, B2 => n2592, 
                           ZN => n14858);
   U9800 : INV_X1 port map( A => n14857, ZN => n9249);
   U9801 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_466_port, B2 => n2592, 
                           ZN => n14857);
   U9802 : INV_X1 port map( A => n14856, ZN => n9250);
   U9803 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_465_port, B2 => n2592, 
                           ZN => n14856);
   U9804 : INV_X1 port map( A => n14855, ZN => n9251);
   U9805 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_464_port, B2 => n2592, 
                           ZN => n14855);
   U9806 : INV_X1 port map( A => n14854, ZN => n9252);
   U9807 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_463_port, B2 => n2592, 
                           ZN => n14854);
   U9808 : INV_X1 port map( A => n14853, ZN => n9253);
   U9809 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_462_port, B2 => n2592, 
                           ZN => n14853);
   U9810 : INV_X1 port map( A => n14852, ZN => n9254);
   U9811 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_461_port, B2 => n2592, 
                           ZN => n14852);
   U9812 : INV_X1 port map( A => n14851, ZN => n9255);
   U9813 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_460_port, B2 => n2592, 
                           ZN => n14851);
   U9814 : INV_X1 port map( A => n14850, ZN => n9256);
   U9815 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_459_port, B2 => n2591, 
                           ZN => n14850);
   U9816 : INV_X1 port map( A => n14849, ZN => n9257);
   U9817 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_458_port, B2 => n2591, 
                           ZN => n14849);
   U9818 : INV_X1 port map( A => n14848, ZN => n9258);
   U9819 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_457_port, B2 => n2591, 
                           ZN => n14848);
   U9820 : INV_X1 port map( A => n14847, ZN => n9259);
   U9821 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2589, B1 => 
                           DataPath_RF_bus_reg_dataout_456_port, B2 => n2591, 
                           ZN => n14847);
   U9822 : INV_X1 port map( A => n14846, ZN => n9260);
   U9823 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_455_port, B2 => n2591, 
                           ZN => n14846);
   U9824 : INV_X1 port map( A => n14845, ZN => n9261);
   U9825 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_454_port, B2 => n2591, 
                           ZN => n14845);
   U9826 : INV_X1 port map( A => n14844, ZN => n9262);
   U9827 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_453_port, B2 => n2591, 
                           ZN => n14844);
   U9828 : INV_X1 port map( A => n14843, ZN => n9263);
   U9829 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_452_port, B2 => n2591, 
                           ZN => n14843);
   U9830 : INV_X1 port map( A => n14842, ZN => n9264);
   U9831 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_451_port, B2 => n2591, 
                           ZN => n14842);
   U9832 : INV_X1 port map( A => n14841, ZN => n9265);
   U9833 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_450_port, B2 => n2591, 
                           ZN => n14841);
   U9834 : INV_X1 port map( A => n14840, ZN => n9266);
   U9835 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_449_port, B2 => n2591, 
                           ZN => n14840);
   U9836 : INV_X1 port map( A => n14837, ZN => n9267);
   U9837 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2590, B1 => 
                           DataPath_RF_bus_reg_dataout_448_port, B2 => n2591, 
                           ZN => n14837);
   U9838 : INV_X1 port map( A => n14904, ZN => n9268);
   U9839 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_31_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_511_port, B2 => n2599, 
                           ZN => n14904);
   U9840 : INV_X1 port map( A => n14903, ZN => n9269);
   U9841 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_30_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_510_port, B2 => n2599, 
                           ZN => n14903);
   U9842 : INV_X1 port map( A => n14902, ZN => n9270);
   U9843 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_29_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_509_port, B2 => n2599, 
                           ZN => n14902);
   U9844 : INV_X1 port map( A => n14901, ZN => n9271);
   U9845 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_28_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_508_port, B2 => n2599, 
                           ZN => n14901);
   U9846 : INV_X1 port map( A => n14900, ZN => n9272);
   U9847 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_27_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_507_port, B2 => n2599, 
                           ZN => n14900);
   U9848 : INV_X1 port map( A => n14899, ZN => n9273);
   U9849 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_26_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_506_port, B2 => n2599, 
                           ZN => n14899);
   U9850 : INV_X1 port map( A => n14898, ZN => n9274);
   U9851 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_25_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_505_port, B2 => n2599, 
                           ZN => n14898);
   U9852 : INV_X1 port map( A => n14897, ZN => n9275);
   U9853 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_24_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_504_port, B2 => n2599, 
                           ZN => n14897);
   U9854 : INV_X1 port map( A => n14896, ZN => n9276);
   U9855 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_23_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_503_port, B2 => n2598, 
                           ZN => n14896);
   U9856 : INV_X1 port map( A => n14895, ZN => n9277);
   U9857 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_22_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_502_port, B2 => n2598, 
                           ZN => n14895);
   U9858 : INV_X1 port map( A => n14894, ZN => n9278);
   U9859 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_21_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_501_port, B2 => n2598, 
                           ZN => n14894);
   U9860 : INV_X1 port map( A => n14893, ZN => n9279);
   U9861 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_20_port, 
                           A2 => n2594, B1 => 
                           DataPath_RF_bus_reg_dataout_500_port, B2 => n2598, 
                           ZN => n14893);
   U9862 : INV_X1 port map( A => n14892, ZN => n9280);
   U9863 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_19_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_499_port, B2 => n2598, 
                           ZN => n14892);
   U9864 : INV_X1 port map( A => n14891, ZN => n9281);
   U9865 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_18_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_498_port, B2 => n2598, 
                           ZN => n14891);
   U9866 : INV_X1 port map( A => n14890, ZN => n9282);
   U9867 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_17_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_497_port, B2 => n2598, 
                           ZN => n14890);
   U9868 : INV_X1 port map( A => n14889, ZN => n9283);
   U9869 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_16_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_496_port, B2 => n2598, 
                           ZN => n14889);
   U9870 : INV_X1 port map( A => n14888, ZN => n9284);
   U9871 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_15_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_495_port, B2 => n2598, 
                           ZN => n14888);
   U9872 : INV_X1 port map( A => n14887, ZN => n9285);
   U9873 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_14_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_494_port, B2 => n2598, 
                           ZN => n14887);
   U9874 : INV_X1 port map( A => n14886, ZN => n9286);
   U9875 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_13_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_493_port, B2 => n2598, 
                           ZN => n14886);
   U9876 : INV_X1 port map( A => n14885, ZN => n9287);
   U9877 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_12_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_492_port, B2 => n2598, 
                           ZN => n14885);
   U9878 : INV_X1 port map( A => n14884, ZN => n9288);
   U9879 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_11_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_491_port, B2 => n2597, 
                           ZN => n14884);
   U9880 : INV_X1 port map( A => n14883, ZN => n9289);
   U9881 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_10_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_490_port, B2 => n2597, 
                           ZN => n14883);
   U9882 : INV_X1 port map( A => n14882, ZN => n9290);
   U9883 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_9_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_489_port, B2 => n2597, 
                           ZN => n14882);
   U9884 : INV_X1 port map( A => n14881, ZN => n9291);
   U9885 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_8_port, 
                           A2 => n2595, B1 => 
                           DataPath_RF_bus_reg_dataout_488_port, B2 => n2597, 
                           ZN => n14881);
   U9886 : INV_X1 port map( A => n14880, ZN => n9292);
   U9887 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_7_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_487_port, B2 => n2597, 
                           ZN => n14880);
   U9888 : INV_X1 port map( A => n14879, ZN => n9293);
   U9889 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_6_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_486_port, B2 => n2597, 
                           ZN => n14879);
   U9890 : INV_X1 port map( A => n14878, ZN => n9294);
   U9891 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_5_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_485_port, B2 => n2597, 
                           ZN => n14878);
   U9892 : INV_X1 port map( A => n14877, ZN => n9295);
   U9893 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_4_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_484_port, B2 => n2597, 
                           ZN => n14877);
   U9894 : INV_X1 port map( A => n14876, ZN => n9296);
   U9895 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_3_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_483_port, B2 => n2597, 
                           ZN => n14876);
   U9896 : INV_X1 port map( A => n14875, ZN => n9297);
   U9897 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_2_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_482_port, B2 => n2597, 
                           ZN => n14875);
   U9898 : INV_X1 port map( A => n14874, ZN => n9298);
   U9899 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_1_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_481_port, B2 => n2597, 
                           ZN => n14874);
   U9900 : INV_X1 port map( A => n14871, ZN => n9299);
   U9901 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_0_0_port, 
                           A2 => n2596, B1 => 
                           DataPath_RF_bus_reg_dataout_480_port, B2 => n2597, 
                           ZN => n14871);
   U9902 : INV_X1 port map( A => n14938, ZN => n9300);
   U9903 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_543_port, B2 => n2605, 
                           ZN => n14938);
   U9904 : INV_X1 port map( A => n14937, ZN => n9301);
   U9905 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_542_port, B2 => n2605, 
                           ZN => n14937);
   U9906 : INV_X1 port map( A => n14936, ZN => n9302);
   U9907 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_541_port, B2 => n2605, 
                           ZN => n14936);
   U9908 : INV_X1 port map( A => n14935, ZN => n9303);
   U9909 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_540_port, B2 => n2605, 
                           ZN => n14935);
   U9910 : INV_X1 port map( A => n14934, ZN => n9304);
   U9911 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_539_port, B2 => n2605, 
                           ZN => n14934);
   U9912 : INV_X1 port map( A => n14933, ZN => n9305);
   U9913 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_538_port, B2 => n2605, 
                           ZN => n14933);
   U9914 : INV_X1 port map( A => n14932, ZN => n9306);
   U9915 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_537_port, B2 => n2605, 
                           ZN => n14932);
   U9916 : INV_X1 port map( A => n14931, ZN => n9307);
   U9917 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_536_port, B2 => n2605, 
                           ZN => n14931);
   U9918 : INV_X1 port map( A => n14930, ZN => n9308);
   U9919 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_535_port, B2 => n2604, 
                           ZN => n14930);
   U9920 : INV_X1 port map( A => n14929, ZN => n9309);
   U9921 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_534_port, B2 => n2604, 
                           ZN => n14929);
   U9922 : INV_X1 port map( A => n14928, ZN => n9310);
   U9923 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_533_port, B2 => n2604, 
                           ZN => n14928);
   U9924 : INV_X1 port map( A => n14927, ZN => n9311);
   U9925 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port, 
                           A2 => n2600, B1 => 
                           DataPath_RF_bus_reg_dataout_532_port, B2 => n2604, 
                           ZN => n14927);
   U9926 : INV_X1 port map( A => n14926, ZN => n9312);
   U9927 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_531_port, B2 => n2604, 
                           ZN => n14926);
   U9928 : INV_X1 port map( A => n14925, ZN => n9313);
   U9929 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_530_port, B2 => n2604, 
                           ZN => n14925);
   U9930 : INV_X1 port map( A => n14924, ZN => n9314);
   U9931 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_529_port, B2 => n2604, 
                           ZN => n14924);
   U9932 : INV_X1 port map( A => n14923, ZN => n9315);
   U9933 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_528_port, B2 => n2604, 
                           ZN => n14923);
   U9934 : INV_X1 port map( A => n14922, ZN => n9316);
   U9935 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_527_port, B2 => n2604, 
                           ZN => n14922);
   U9936 : INV_X1 port map( A => n14921, ZN => n9317);
   U9937 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_526_port, B2 => n2604, 
                           ZN => n14921);
   U9938 : INV_X1 port map( A => n14920, ZN => n9318);
   U9939 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_525_port, B2 => n2604, 
                           ZN => n14920);
   U9940 : INV_X1 port map( A => n14919, ZN => n9319);
   U9941 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_524_port, B2 => n2604, 
                           ZN => n14919);
   U9942 : INV_X1 port map( A => n14918, ZN => n9320);
   U9943 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_523_port, B2 => n2603, 
                           ZN => n14918);
   U9944 : INV_X1 port map( A => n14917, ZN => n9321);
   U9945 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_522_port, B2 => n2603, 
                           ZN => n14917);
   U9946 : INV_X1 port map( A => n14916, ZN => n9322);
   U9947 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_521_port, B2 => n2603, 
                           ZN => n14916);
   U9948 : INV_X1 port map( A => n14915, ZN => n9323);
   U9949 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2601, B1 => 
                           DataPath_RF_bus_reg_dataout_520_port, B2 => n2603, 
                           ZN => n14915);
   U9950 : INV_X1 port map( A => n14914, ZN => n9324);
   U9951 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_519_port, B2 => n2603, 
                           ZN => n14914);
   U9952 : INV_X1 port map( A => n14913, ZN => n9325);
   U9953 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_518_port, B2 => n2603, 
                           ZN => n14913);
   U9954 : INV_X1 port map( A => n14912, ZN => n9326);
   U9955 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_517_port, B2 => n2603, 
                           ZN => n14912);
   U9956 : INV_X1 port map( A => n14911, ZN => n9327);
   U9957 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_516_port, B2 => n2603, 
                           ZN => n14911);
   U9958 : INV_X1 port map( A => n14910, ZN => n9328);
   U9959 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_515_port, B2 => n2603, 
                           ZN => n14910);
   U9960 : INV_X1 port map( A => n14909, ZN => n9329);
   U9961 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_514_port, B2 => n2603, 
                           ZN => n14909);
   U9962 : INV_X1 port map( A => n14908, ZN => n9330);
   U9963 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_513_port, B2 => n2603, 
                           ZN => n14908);
   U9964 : INV_X1 port map( A => n14905, ZN => n9331);
   U9965 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2602, B1 => 
                           DataPath_RF_bus_reg_dataout_512_port, B2 => n2603, 
                           ZN => n14905);
   U9966 : INV_X1 port map( A => n14972, ZN => n9332);
   U9967 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_575_port, B2 => n2611, 
                           ZN => n14972);
   U9968 : INV_X1 port map( A => n14971, ZN => n9333);
   U9969 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_574_port, B2 => n2611, 
                           ZN => n14971);
   U9970 : INV_X1 port map( A => n14970, ZN => n9334);
   U9971 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_573_port, B2 => n2611, 
                           ZN => n14970);
   U9972 : INV_X1 port map( A => n14969, ZN => n9335);
   U9973 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_572_port, B2 => n2611, 
                           ZN => n14969);
   U9974 : INV_X1 port map( A => n14968, ZN => n9336);
   U9975 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_571_port, B2 => n2611, 
                           ZN => n14968);
   U9976 : INV_X1 port map( A => n14967, ZN => n9337);
   U9977 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_570_port, B2 => n2611, 
                           ZN => n14967);
   U9978 : INV_X1 port map( A => n14966, ZN => n9338);
   U9979 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_569_port, B2 => n2611, 
                           ZN => n14966);
   U9980 : INV_X1 port map( A => n14965, ZN => n9339);
   U9981 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_568_port, B2 => n2611, 
                           ZN => n14965);
   U9982 : INV_X1 port map( A => n14964, ZN => n9340);
   U9983 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_567_port, B2 => n2610, 
                           ZN => n14964);
   U9984 : INV_X1 port map( A => n14963, ZN => n9341);
   U9985 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_566_port, B2 => n2610, 
                           ZN => n14963);
   U9986 : INV_X1 port map( A => n14962, ZN => n9342);
   U9987 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_565_port, B2 => n2610, 
                           ZN => n14962);
   U9988 : INV_X1 port map( A => n14961, ZN => n9343);
   U9989 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port, 
                           A2 => n2606, B1 => 
                           DataPath_RF_bus_reg_dataout_564_port, B2 => n2610, 
                           ZN => n14961);
   U9990 : INV_X1 port map( A => n14960, ZN => n9344);
   U9991 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port, 
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_563_port, B2 => n2610, 
                           ZN => n14960);
   U9992 : INV_X1 port map( A => n14959, ZN => n9345);
   U9993 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port, 
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_562_port, B2 => n2610, 
                           ZN => n14959);
   U9994 : INV_X1 port map( A => n14958, ZN => n9346);
   U9995 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port, 
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_561_port, B2 => n2610, 
                           ZN => n14958);
   U9996 : INV_X1 port map( A => n14957, ZN => n9347);
   U9997 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port, 
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_560_port, B2 => n2610, 
                           ZN => n14957);
   U9998 : INV_X1 port map( A => n14956, ZN => n9348);
   U9999 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port, 
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_559_port, B2 => n2610, 
                           ZN => n14956);
   U10000 : INV_X1 port map( A => n14955, ZN => n9349);
   U10001 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_558_port, B2 => n2610, 
                           ZN => n14955);
   U10002 : INV_X1 port map( A => n14954, ZN => n9350);
   U10003 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_557_port, B2 => n2610, 
                           ZN => n14954);
   U10004 : INV_X1 port map( A => n14953, ZN => n9351);
   U10005 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_556_port, B2 => n2610, 
                           ZN => n14953);
   U10006 : INV_X1 port map( A => n14952, ZN => n9352);
   U10007 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_555_port, B2 => n2609, 
                           ZN => n14952);
   U10008 : INV_X1 port map( A => n14951, ZN => n9353);
   U10009 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_554_port, B2 => n2609, 
                           ZN => n14951);
   U10010 : INV_X1 port map( A => n14950, ZN => n9354);
   U10011 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_553_port, B2 => n2609, 
                           ZN => n14950);
   U10012 : INV_X1 port map( A => n14949, ZN => n9355);
   U10013 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2607, B1 => 
                           DataPath_RF_bus_reg_dataout_552_port, B2 => n2609, 
                           ZN => n14949);
   U10014 : INV_X1 port map( A => n14948, ZN => n9356);
   U10015 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_551_port, B2 => n2609, 
                           ZN => n14948);
   U10016 : INV_X1 port map( A => n14947, ZN => n9357);
   U10017 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_550_port, B2 => n2609, 
                           ZN => n14947);
   U10018 : INV_X1 port map( A => n14946, ZN => n9358);
   U10019 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_549_port, B2 => n2609, 
                           ZN => n14946);
   U10020 : INV_X1 port map( A => n14945, ZN => n9359);
   U10021 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_548_port, B2 => n2609, 
                           ZN => n14945);
   U10022 : INV_X1 port map( A => n14944, ZN => n9360);
   U10023 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_547_port, B2 => n2609, 
                           ZN => n14944);
   U10024 : INV_X1 port map( A => n14943, ZN => n9361);
   U10025 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_546_port, B2 => n2609, 
                           ZN => n14943);
   U10026 : INV_X1 port map( A => n14942, ZN => n9362);
   U10027 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_545_port, B2 => n2609, 
                           ZN => n14942);
   U10028 : INV_X1 port map( A => n14939, ZN => n9363);
   U10029 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2608, B1 => 
                           DataPath_RF_bus_reg_dataout_544_port, B2 => n2609, 
                           ZN => n14939);
   U10030 : INV_X1 port map( A => n15006, ZN => n9364);
   U10031 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_607_port, B2 => n2617, 
                           ZN => n15006);
   U10032 : INV_X1 port map( A => n15005, ZN => n9365);
   U10033 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_606_port, B2 => n2617, 
                           ZN => n15005);
   U10034 : INV_X1 port map( A => n15004, ZN => n9366);
   U10035 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_605_port, B2 => n2617, 
                           ZN => n15004);
   U10036 : INV_X1 port map( A => n15003, ZN => n9367);
   U10037 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_604_port, B2 => n2617, 
                           ZN => n15003);
   U10038 : INV_X1 port map( A => n15002, ZN => n9368);
   U10039 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_603_port, B2 => n2617, 
                           ZN => n15002);
   U10040 : INV_X1 port map( A => n15001, ZN => n9369);
   U10041 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_602_port, B2 => n2617, 
                           ZN => n15001);
   U10042 : INV_X1 port map( A => n15000, ZN => n9370);
   U10043 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_601_port, B2 => n2617, 
                           ZN => n15000);
   U10044 : INV_X1 port map( A => n14999, ZN => n9371);
   U10045 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_600_port, B2 => n2617, 
                           ZN => n14999);
   U10046 : INV_X1 port map( A => n14998, ZN => n9372);
   U10047 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_599_port, B2 => n2616, 
                           ZN => n14998);
   U10048 : INV_X1 port map( A => n14997, ZN => n9373);
   U10049 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_598_port, B2 => n2616, 
                           ZN => n14997);
   U10050 : INV_X1 port map( A => n14996, ZN => n9374);
   U10051 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_597_port, B2 => n2616, 
                           ZN => n14996);
   U10052 : INV_X1 port map( A => n14995, ZN => n9375);
   U10053 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2612, B1 => 
                           DataPath_RF_bus_reg_dataout_596_port, B2 => n2616, 
                           ZN => n14995);
   U10054 : INV_X1 port map( A => n14994, ZN => n9376);
   U10055 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_595_port, B2 => n2616, 
                           ZN => n14994);
   U10056 : INV_X1 port map( A => n14993, ZN => n9377);
   U10057 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_594_port, B2 => n2616, 
                           ZN => n14993);
   U10058 : INV_X1 port map( A => n14992, ZN => n9378);
   U10059 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_593_port, B2 => n2616, 
                           ZN => n14992);
   U10060 : INV_X1 port map( A => n14991, ZN => n9379);
   U10061 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_592_port, B2 => n2616, 
                           ZN => n14991);
   U10062 : INV_X1 port map( A => n14990, ZN => n9380);
   U10063 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_591_port, B2 => n2616, 
                           ZN => n14990);
   U10064 : INV_X1 port map( A => n14989, ZN => n9381);
   U10065 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_590_port, B2 => n2616, 
                           ZN => n14989);
   U10066 : INV_X1 port map( A => n14988, ZN => n9382);
   U10067 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_589_port, B2 => n2616, 
                           ZN => n14988);
   U10068 : INV_X1 port map( A => n14987, ZN => n9383);
   U10069 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_588_port, B2 => n2616, 
                           ZN => n14987);
   U10070 : INV_X1 port map( A => n14986, ZN => n9384);
   U10071 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_587_port, B2 => n2615, 
                           ZN => n14986);
   U10072 : INV_X1 port map( A => n14985, ZN => n9385);
   U10073 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_586_port, B2 => n2615, 
                           ZN => n14985);
   U10074 : INV_X1 port map( A => n14984, ZN => n9386);
   U10075 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_585_port, B2 => n2615, 
                           ZN => n14984);
   U10076 : INV_X1 port map( A => n14983, ZN => n9387);
   U10077 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2613, B1 => 
                           DataPath_RF_bus_reg_dataout_584_port, B2 => n2615, 
                           ZN => n14983);
   U10078 : INV_X1 port map( A => n14982, ZN => n9388);
   U10079 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_583_port, B2 => n2615, 
                           ZN => n14982);
   U10080 : INV_X1 port map( A => n14981, ZN => n9389);
   U10081 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_582_port, B2 => n2615, 
                           ZN => n14981);
   U10082 : INV_X1 port map( A => n14980, ZN => n9390);
   U10083 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_581_port, B2 => n2615, 
                           ZN => n14980);
   U10084 : INV_X1 port map( A => n14979, ZN => n9391);
   U10085 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_580_port, B2 => n2615, 
                           ZN => n14979);
   U10086 : INV_X1 port map( A => n14978, ZN => n9392);
   U10087 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_579_port, B2 => n2615, 
                           ZN => n14978);
   U10088 : INV_X1 port map( A => n14977, ZN => n9393);
   U10089 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_578_port, B2 => n2615, 
                           ZN => n14977);
   U10090 : INV_X1 port map( A => n14976, ZN => n9394);
   U10091 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_577_port, B2 => n2615, 
                           ZN => n14976);
   U10092 : INV_X1 port map( A => n14973, ZN => n9395);
   U10093 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2614, B1 => 
                           DataPath_RF_bus_reg_dataout_576_port, B2 => n2615, 
                           ZN => n14973);
   U10094 : INV_X1 port map( A => n15040, ZN => n9396);
   U10095 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_639_port, B2 => n2623, 
                           ZN => n15040);
   U10096 : INV_X1 port map( A => n15039, ZN => n9397);
   U10097 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_638_port, B2 => n2623, 
                           ZN => n15039);
   U10098 : INV_X1 port map( A => n15038, ZN => n9398);
   U10099 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_637_port, B2 => n2623, 
                           ZN => n15038);
   U10100 : INV_X1 port map( A => n15037, ZN => n9399);
   U10101 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_636_port, B2 => n2623, 
                           ZN => n15037);
   U10102 : INV_X1 port map( A => n15036, ZN => n9400);
   U10103 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_635_port, B2 => n2623, 
                           ZN => n15036);
   U10104 : INV_X1 port map( A => n15035, ZN => n9401);
   U10105 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_634_port, B2 => n2623, 
                           ZN => n15035);
   U10106 : INV_X1 port map( A => n15034, ZN => n9402);
   U10107 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_633_port, B2 => n2623, 
                           ZN => n15034);
   U10108 : INV_X1 port map( A => n15033, ZN => n9403);
   U10109 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_632_port, B2 => n2623, 
                           ZN => n15033);
   U10110 : INV_X1 port map( A => n15032, ZN => n9404);
   U10111 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_631_port, B2 => n2622, 
                           ZN => n15032);
   U10112 : INV_X1 port map( A => n15031, ZN => n9405);
   U10113 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_630_port, B2 => n2622, 
                           ZN => n15031);
   U10114 : INV_X1 port map( A => n15030, ZN => n9406);
   U10115 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_629_port, B2 => n2622, 
                           ZN => n15030);
   U10116 : INV_X1 port map( A => n15029, ZN => n9407);
   U10117 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2618, B1 => 
                           DataPath_RF_bus_reg_dataout_628_port, B2 => n2622, 
                           ZN => n15029);
   U10118 : INV_X1 port map( A => n15028, ZN => n9408);
   U10119 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_627_port, B2 => n2622, 
                           ZN => n15028);
   U10120 : INV_X1 port map( A => n15027, ZN => n9409);
   U10121 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_626_port, B2 => n2622, 
                           ZN => n15027);
   U10122 : INV_X1 port map( A => n15026, ZN => n9410);
   U10123 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_625_port, B2 => n2622, 
                           ZN => n15026);
   U10124 : INV_X1 port map( A => n15025, ZN => n9411);
   U10125 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_624_port, B2 => n2622, 
                           ZN => n15025);
   U10126 : INV_X1 port map( A => n15024, ZN => n9412);
   U10127 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_623_port, B2 => n2622, 
                           ZN => n15024);
   U10128 : INV_X1 port map( A => n15023, ZN => n9413);
   U10129 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_622_port, B2 => n2622, 
                           ZN => n15023);
   U10130 : INV_X1 port map( A => n15022, ZN => n9414);
   U10131 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_621_port, B2 => n2622, 
                           ZN => n15022);
   U10132 : INV_X1 port map( A => n15021, ZN => n9415);
   U10133 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_620_port, B2 => n2622, 
                           ZN => n15021);
   U10134 : INV_X1 port map( A => n15020, ZN => n9416);
   U10135 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_619_port, B2 => n2621, 
                           ZN => n15020);
   U10136 : INV_X1 port map( A => n15019, ZN => n9417);
   U10137 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_618_port, B2 => n2621, 
                           ZN => n15019);
   U10138 : INV_X1 port map( A => n15018, ZN => n9418);
   U10139 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_617_port, B2 => n2621, 
                           ZN => n15018);
   U10140 : INV_X1 port map( A => n15017, ZN => n9419);
   U10141 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2619, B1 => 
                           DataPath_RF_bus_reg_dataout_616_port, B2 => n2621, 
                           ZN => n15017);
   U10142 : INV_X1 port map( A => n15016, ZN => n9420);
   U10143 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_615_port, B2 => n2621, 
                           ZN => n15016);
   U10144 : INV_X1 port map( A => n15015, ZN => n9421);
   U10145 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_614_port, B2 => n2621, 
                           ZN => n15015);
   U10146 : INV_X1 port map( A => n15014, ZN => n9422);
   U10147 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_613_port, B2 => n2621, 
                           ZN => n15014);
   U10148 : INV_X1 port map( A => n15013, ZN => n9423);
   U10149 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_612_port, B2 => n2621, 
                           ZN => n15013);
   U10150 : INV_X1 port map( A => n15012, ZN => n9424);
   U10151 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_611_port, B2 => n2621, 
                           ZN => n15012);
   U10152 : INV_X1 port map( A => n15011, ZN => n9425);
   U10153 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_610_port, B2 => n2621, 
                           ZN => n15011);
   U10154 : INV_X1 port map( A => n15010, ZN => n9426);
   U10155 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_609_port, B2 => n2621, 
                           ZN => n15010);
   U10156 : INV_X1 port map( A => n15007, ZN => n9427);
   U10157 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2620, B1 => 
                           DataPath_RF_bus_reg_dataout_608_port, B2 => n2621, 
                           ZN => n15007);
   U10158 : INV_X1 port map( A => n15074, ZN => n9428);
   U10159 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_671_port, B2 => n2629, 
                           ZN => n15074);
   U10160 : INV_X1 port map( A => n15073, ZN => n9429);
   U10161 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_670_port, B2 => n2629, 
                           ZN => n15073);
   U10162 : INV_X1 port map( A => n15072, ZN => n9430);
   U10163 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_669_port, B2 => n2629, 
                           ZN => n15072);
   U10164 : INV_X1 port map( A => n15071, ZN => n9431);
   U10165 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_668_port, B2 => n2629, 
                           ZN => n15071);
   U10166 : INV_X1 port map( A => n15070, ZN => n9432);
   U10167 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_667_port, B2 => n2629, 
                           ZN => n15070);
   U10168 : INV_X1 port map( A => n15069, ZN => n9433);
   U10169 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_666_port, B2 => n2629, 
                           ZN => n15069);
   U10170 : INV_X1 port map( A => n15068, ZN => n9434);
   U10171 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_665_port, B2 => n2629, 
                           ZN => n15068);
   U10172 : INV_X1 port map( A => n15067, ZN => n9435);
   U10173 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_664_port, B2 => n2629, 
                           ZN => n15067);
   U10174 : INV_X1 port map( A => n15066, ZN => n9436);
   U10175 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_663_port, B2 => n2628, 
                           ZN => n15066);
   U10176 : INV_X1 port map( A => n15065, ZN => n9437);
   U10177 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_662_port, B2 => n2628, 
                           ZN => n15065);
   U10178 : INV_X1 port map( A => n15064, ZN => n9438);
   U10179 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_661_port, B2 => n2628, 
                           ZN => n15064);
   U10180 : INV_X1 port map( A => n15063, ZN => n9439);
   U10181 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2624, B1 => 
                           DataPath_RF_bus_reg_dataout_660_port, B2 => n2628, 
                           ZN => n15063);
   U10182 : INV_X1 port map( A => n15062, ZN => n9440);
   U10183 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_659_port, B2 => n2628, 
                           ZN => n15062);
   U10184 : INV_X1 port map( A => n15061, ZN => n9441);
   U10185 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_658_port, B2 => n2628, 
                           ZN => n15061);
   U10186 : INV_X1 port map( A => n15060, ZN => n9442);
   U10187 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_657_port, B2 => n2628, 
                           ZN => n15060);
   U10188 : INV_X1 port map( A => n15059, ZN => n9443);
   U10189 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_656_port, B2 => n2628, 
                           ZN => n15059);
   U10190 : INV_X1 port map( A => n15058, ZN => n9444);
   U10191 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_655_port, B2 => n2628, 
                           ZN => n15058);
   U10192 : INV_X1 port map( A => n15057, ZN => n9445);
   U10193 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_654_port, B2 => n2628, 
                           ZN => n15057);
   U10194 : INV_X1 port map( A => n15056, ZN => n9446);
   U10195 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_653_port, B2 => n2628, 
                           ZN => n15056);
   U10196 : INV_X1 port map( A => n15055, ZN => n9447);
   U10197 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_652_port, B2 => n2628, 
                           ZN => n15055);
   U10198 : INV_X1 port map( A => n15054, ZN => n9448);
   U10199 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_651_port, B2 => n2627, 
                           ZN => n15054);
   U10200 : INV_X1 port map( A => n15053, ZN => n9449);
   U10201 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_650_port, B2 => n2627, 
                           ZN => n15053);
   U10202 : INV_X1 port map( A => n15052, ZN => n9450);
   U10203 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_649_port, B2 => n2627, 
                           ZN => n15052);
   U10204 : INV_X1 port map( A => n15051, ZN => n9451);
   U10205 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2625, B1 => 
                           DataPath_RF_bus_reg_dataout_648_port, B2 => n2627, 
                           ZN => n15051);
   U10206 : INV_X1 port map( A => n15050, ZN => n9452);
   U10207 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_647_port, B2 => n2627, 
                           ZN => n15050);
   U10208 : INV_X1 port map( A => n15049, ZN => n9453);
   U10209 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_646_port, B2 => n2627, 
                           ZN => n15049);
   U10210 : INV_X1 port map( A => n15048, ZN => n9454);
   U10211 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_645_port, B2 => n2627, 
                           ZN => n15048);
   U10212 : INV_X1 port map( A => n15047, ZN => n9455);
   U10213 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_644_port, B2 => n2627, 
                           ZN => n15047);
   U10214 : INV_X1 port map( A => n15046, ZN => n9456);
   U10215 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_643_port, B2 => n2627, 
                           ZN => n15046);
   U10216 : INV_X1 port map( A => n15045, ZN => n9457);
   U10217 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_642_port, B2 => n2627, 
                           ZN => n15045);
   U10218 : INV_X1 port map( A => n15044, ZN => n9458);
   U10219 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_641_port, B2 => n2627, 
                           ZN => n15044);
   U10220 : INV_X1 port map( A => n15041, ZN => n9459);
   U10221 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2626, B1 => 
                           DataPath_RF_bus_reg_dataout_640_port, B2 => n2627, 
                           ZN => n15041);
   U10222 : INV_X1 port map( A => n15108, ZN => n9460);
   U10223 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_703_port, B2 => n2635, 
                           ZN => n15108);
   U10224 : INV_X1 port map( A => n15107, ZN => n9461);
   U10225 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_702_port, B2 => n2635, 
                           ZN => n15107);
   U10226 : INV_X1 port map( A => n15106, ZN => n9462);
   U10227 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_701_port, B2 => n2635, 
                           ZN => n15106);
   U10228 : INV_X1 port map( A => n15105, ZN => n9463);
   U10229 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_700_port, B2 => n2635, 
                           ZN => n15105);
   U10230 : INV_X1 port map( A => n15104, ZN => n9464);
   U10231 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_699_port, B2 => n2635, 
                           ZN => n15104);
   U10232 : INV_X1 port map( A => n15103, ZN => n9465);
   U10233 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_698_port, B2 => n2635, 
                           ZN => n15103);
   U10234 : INV_X1 port map( A => n15102, ZN => n9466);
   U10235 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_697_port, B2 => n2635, 
                           ZN => n15102);
   U10236 : INV_X1 port map( A => n15101, ZN => n9467);
   U10237 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_696_port, B2 => n2635, 
                           ZN => n15101);
   U10238 : INV_X1 port map( A => n15100, ZN => n9468);
   U10239 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_695_port, B2 => n2634, 
                           ZN => n15100);
   U10240 : INV_X1 port map( A => n15099, ZN => n9469);
   U10241 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_694_port, B2 => n2634, 
                           ZN => n15099);
   U10242 : INV_X1 port map( A => n15098, ZN => n9470);
   U10243 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_693_port, B2 => n2634, 
                           ZN => n15098);
   U10244 : INV_X1 port map( A => n15097, ZN => n9471);
   U10245 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2630, B1 => 
                           DataPath_RF_bus_reg_dataout_692_port, B2 => n2634, 
                           ZN => n15097);
   U10246 : INV_X1 port map( A => n15096, ZN => n9472);
   U10247 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_691_port, B2 => n2634, 
                           ZN => n15096);
   U10248 : INV_X1 port map( A => n15095, ZN => n9473);
   U10249 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_690_port, B2 => n2634, 
                           ZN => n15095);
   U10250 : INV_X1 port map( A => n15094, ZN => n9474);
   U10251 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_689_port, B2 => n2634, 
                           ZN => n15094);
   U10252 : INV_X1 port map( A => n15093, ZN => n9475);
   U10253 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_688_port, B2 => n2634, 
                           ZN => n15093);
   U10254 : INV_X1 port map( A => n15092, ZN => n9476);
   U10255 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_687_port, B2 => n2634, 
                           ZN => n15092);
   U10256 : INV_X1 port map( A => n15091, ZN => n9477);
   U10257 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_686_port, B2 => n2634, 
                           ZN => n15091);
   U10258 : INV_X1 port map( A => n15090, ZN => n9478);
   U10259 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_685_port, B2 => n2634, 
                           ZN => n15090);
   U10260 : INV_X1 port map( A => n15089, ZN => n9479);
   U10261 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_684_port, B2 => n2634, 
                           ZN => n15089);
   U10262 : INV_X1 port map( A => n15088, ZN => n9480);
   U10263 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_683_port, B2 => n2633, 
                           ZN => n15088);
   U10264 : INV_X1 port map( A => n15087, ZN => n9481);
   U10265 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_682_port, B2 => n2633, 
                           ZN => n15087);
   U10266 : INV_X1 port map( A => n15086, ZN => n9482);
   U10267 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_681_port, B2 => n2633, 
                           ZN => n15086);
   U10268 : INV_X1 port map( A => n15085, ZN => n9483);
   U10269 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2631, B1 => 
                           DataPath_RF_bus_reg_dataout_680_port, B2 => n2633, 
                           ZN => n15085);
   U10270 : INV_X1 port map( A => n15084, ZN => n9484);
   U10271 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_679_port, B2 => n2633, 
                           ZN => n15084);
   U10272 : INV_X1 port map( A => n15083, ZN => n9485);
   U10273 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_678_port, B2 => n2633, 
                           ZN => n15083);
   U10274 : INV_X1 port map( A => n15082, ZN => n9486);
   U10275 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_677_port, B2 => n2633, 
                           ZN => n15082);
   U10276 : INV_X1 port map( A => n15081, ZN => n9487);
   U10277 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_676_port, B2 => n2633, 
                           ZN => n15081);
   U10278 : INV_X1 port map( A => n15080, ZN => n9488);
   U10279 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_675_port, B2 => n2633, 
                           ZN => n15080);
   U10280 : INV_X1 port map( A => n15079, ZN => n9489);
   U10281 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_674_port, B2 => n2633, 
                           ZN => n15079);
   U10282 : INV_X1 port map( A => n15078, ZN => n9490);
   U10283 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_673_port, B2 => n2633, 
                           ZN => n15078);
   U10284 : INV_X1 port map( A => n15075, ZN => n9491);
   U10285 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2632, B1 => 
                           DataPath_RF_bus_reg_dataout_672_port, B2 => n2633, 
                           ZN => n15075);
   U10286 : INV_X1 port map( A => n15142, ZN => n9492);
   U10287 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_735_port, B2 => n2641, 
                           ZN => n15142);
   U10288 : INV_X1 port map( A => n15141, ZN => n9493);
   U10289 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_734_port, B2 => n2641, 
                           ZN => n15141);
   U10290 : INV_X1 port map( A => n15140, ZN => n9494);
   U10291 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_733_port, B2 => n2641, 
                           ZN => n15140);
   U10292 : INV_X1 port map( A => n15139, ZN => n9495);
   U10293 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_732_port, B2 => n2641, 
                           ZN => n15139);
   U10294 : INV_X1 port map( A => n15138, ZN => n9496);
   U10295 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_731_port, B2 => n2641, 
                           ZN => n15138);
   U10296 : INV_X1 port map( A => n15137, ZN => n9497);
   U10297 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_730_port, B2 => n2641, 
                           ZN => n15137);
   U10298 : INV_X1 port map( A => n15136, ZN => n9498);
   U10299 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_729_port, B2 => n2641, 
                           ZN => n15136);
   U10300 : INV_X1 port map( A => n15135, ZN => n9499);
   U10301 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_728_port, B2 => n2641, 
                           ZN => n15135);
   U10302 : INV_X1 port map( A => n15134, ZN => n9500);
   U10303 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_727_port, B2 => n2640, 
                           ZN => n15134);
   U10304 : INV_X1 port map( A => n15133, ZN => n9501);
   U10305 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_726_port, B2 => n2640, 
                           ZN => n15133);
   U10306 : INV_X1 port map( A => n15132, ZN => n9502);
   U10307 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_725_port, B2 => n2640, 
                           ZN => n15132);
   U10308 : INV_X1 port map( A => n15131, ZN => n9503);
   U10309 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2636, B1 => 
                           DataPath_RF_bus_reg_dataout_724_port, B2 => n2640, 
                           ZN => n15131);
   U10310 : INV_X1 port map( A => n15130, ZN => n9504);
   U10311 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_723_port, B2 => n2640, 
                           ZN => n15130);
   U10312 : INV_X1 port map( A => n15129, ZN => n9505);
   U10313 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_722_port, B2 => n2640, 
                           ZN => n15129);
   U10314 : INV_X1 port map( A => n15128, ZN => n9506);
   U10315 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_721_port, B2 => n2640, 
                           ZN => n15128);
   U10316 : INV_X1 port map( A => n15127, ZN => n9507);
   U10317 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_720_port, B2 => n2640, 
                           ZN => n15127);
   U10318 : INV_X1 port map( A => n15126, ZN => n9508);
   U10319 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_719_port, B2 => n2640, 
                           ZN => n15126);
   U10320 : INV_X1 port map( A => n15125, ZN => n9509);
   U10321 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_718_port, B2 => n2640, 
                           ZN => n15125);
   U10322 : INV_X1 port map( A => n15124, ZN => n9510);
   U10323 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_717_port, B2 => n2640, 
                           ZN => n15124);
   U10324 : INV_X1 port map( A => n15123, ZN => n9511);
   U10325 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_716_port, B2 => n2640, 
                           ZN => n15123);
   U10326 : INV_X1 port map( A => n15122, ZN => n9512);
   U10327 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_715_port, B2 => n2639, 
                           ZN => n15122);
   U10328 : INV_X1 port map( A => n15121, ZN => n9513);
   U10329 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_714_port, B2 => n2639, 
                           ZN => n15121);
   U10330 : INV_X1 port map( A => n15120, ZN => n9514);
   U10331 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_713_port, B2 => n2639, 
                           ZN => n15120);
   U10332 : INV_X1 port map( A => n15119, ZN => n9515);
   U10333 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2637, B1 => 
                           DataPath_RF_bus_reg_dataout_712_port, B2 => n2639, 
                           ZN => n15119);
   U10334 : INV_X1 port map( A => n15118, ZN => n9516);
   U10335 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_711_port, B2 => n2639, 
                           ZN => n15118);
   U10336 : INV_X1 port map( A => n15117, ZN => n9517);
   U10337 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_710_port, B2 => n2639, 
                           ZN => n15117);
   U10338 : INV_X1 port map( A => n15116, ZN => n9518);
   U10339 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_709_port, B2 => n2639, 
                           ZN => n15116);
   U10340 : INV_X1 port map( A => n15115, ZN => n9519);
   U10341 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_708_port, B2 => n2639, 
                           ZN => n15115);
   U10342 : INV_X1 port map( A => n15114, ZN => n9520);
   U10343 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_707_port, B2 => n2639, 
                           ZN => n15114);
   U10344 : INV_X1 port map( A => n15113, ZN => n9521);
   U10345 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_706_port, B2 => n2639, 
                           ZN => n15113);
   U10346 : INV_X1 port map( A => n15112, ZN => n9522);
   U10347 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_705_port, B2 => n2639, 
                           ZN => n15112);
   U10348 : INV_X1 port map( A => n15109, ZN => n9523);
   U10349 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2638, B1 => 
                           DataPath_RF_bus_reg_dataout_704_port, B2 => n2639, 
                           ZN => n15109);
   U10350 : INV_X1 port map( A => n15176, ZN => n9524);
   U10351 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_767_port, B2 => n2647, 
                           ZN => n15176);
   U10352 : INV_X1 port map( A => n15175, ZN => n9525);
   U10353 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_766_port, B2 => n2647, 
                           ZN => n15175);
   U10354 : INV_X1 port map( A => n15174, ZN => n9526);
   U10355 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_765_port, B2 => n2647, 
                           ZN => n15174);
   U10356 : INV_X1 port map( A => n15173, ZN => n9527);
   U10357 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_764_port, B2 => n2647, 
                           ZN => n15173);
   U10358 : INV_X1 port map( A => n15172, ZN => n9528);
   U10359 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_763_port, B2 => n2647, 
                           ZN => n15172);
   U10360 : INV_X1 port map( A => n15171, ZN => n9529);
   U10361 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_762_port, B2 => n2647, 
                           ZN => n15171);
   U10362 : INV_X1 port map( A => n15170, ZN => n9530);
   U10363 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_761_port, B2 => n2647, 
                           ZN => n15170);
   U10364 : INV_X1 port map( A => n15169, ZN => n9531);
   U10365 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_760_port, B2 => n2647, 
                           ZN => n15169);
   U10366 : INV_X1 port map( A => n15168, ZN => n9532);
   U10367 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_759_port, B2 => n2646, 
                           ZN => n15168);
   U10368 : INV_X1 port map( A => n15167, ZN => n9533);
   U10369 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_758_port, B2 => n2646, 
                           ZN => n15167);
   U10370 : INV_X1 port map( A => n15166, ZN => n9534);
   U10371 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_757_port, B2 => n2646, 
                           ZN => n15166);
   U10372 : INV_X1 port map( A => n15165, ZN => n9535);
   U10373 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2642, B1 => 
                           DataPath_RF_bus_reg_dataout_756_port, B2 => n2646, 
                           ZN => n15165);
   U10374 : INV_X1 port map( A => n15164, ZN => n9536);
   U10375 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_755_port, B2 => n2646, 
                           ZN => n15164);
   U10376 : INV_X1 port map( A => n15163, ZN => n9537);
   U10377 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_754_port, B2 => n2646, 
                           ZN => n15163);
   U10378 : INV_X1 port map( A => n15162, ZN => n9538);
   U10379 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_753_port, B2 => n2646, 
                           ZN => n15162);
   U10380 : INV_X1 port map( A => n15161, ZN => n9539);
   U10381 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_752_port, B2 => n2646, 
                           ZN => n15161);
   U10382 : INV_X1 port map( A => n15160, ZN => n9540);
   U10383 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_751_port, B2 => n2646, 
                           ZN => n15160);
   U10384 : INV_X1 port map( A => n15159, ZN => n9541);
   U10385 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_750_port, B2 => n2646, 
                           ZN => n15159);
   U10386 : INV_X1 port map( A => n15158, ZN => n9542);
   U10387 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_749_port, B2 => n2646, 
                           ZN => n15158);
   U10388 : INV_X1 port map( A => n15157, ZN => n9543);
   U10389 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_748_port, B2 => n2646, 
                           ZN => n15157);
   U10390 : INV_X1 port map( A => n15156, ZN => n9544);
   U10391 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_747_port, B2 => n2645, 
                           ZN => n15156);
   U10392 : INV_X1 port map( A => n15155, ZN => n9545);
   U10393 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_746_port, B2 => n2645, 
                           ZN => n15155);
   U10394 : INV_X1 port map( A => n15154, ZN => n9546);
   U10395 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_745_port, B2 => n2645, 
                           ZN => n15154);
   U10396 : INV_X1 port map( A => n15153, ZN => n9547);
   U10397 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2643, B1 => 
                           DataPath_RF_bus_reg_dataout_744_port, B2 => n2645, 
                           ZN => n15153);
   U10398 : INV_X1 port map( A => n15152, ZN => n9548);
   U10399 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_743_port, B2 => n2645, 
                           ZN => n15152);
   U10400 : INV_X1 port map( A => n15151, ZN => n9549);
   U10401 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_742_port, B2 => n2645, 
                           ZN => n15151);
   U10402 : INV_X1 port map( A => n15150, ZN => n9550);
   U10403 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_741_port, B2 => n2645, 
                           ZN => n15150);
   U10404 : INV_X1 port map( A => n15149, ZN => n9551);
   U10405 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_740_port, B2 => n2645, 
                           ZN => n15149);
   U10406 : INV_X1 port map( A => n15148, ZN => n9552);
   U10407 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_739_port, B2 => n2645, 
                           ZN => n15148);
   U10408 : INV_X1 port map( A => n15147, ZN => n9553);
   U10409 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_738_port, B2 => n2645, 
                           ZN => n15147);
   U10410 : INV_X1 port map( A => n15146, ZN => n9554);
   U10411 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_737_port, B2 => n2645, 
                           ZN => n15146);
   U10412 : INV_X1 port map( A => n15143, ZN => n9555);
   U10413 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2644, B1 => 
                           DataPath_RF_bus_reg_dataout_736_port, B2 => n2645, 
                           ZN => n15143);
   U10414 : INV_X1 port map( A => n15210, ZN => n9556);
   U10415 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_799_port, B2 => n2653, 
                           ZN => n15210);
   U10416 : INV_X1 port map( A => n15209, ZN => n9557);
   U10417 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_798_port, B2 => n2653, 
                           ZN => n15209);
   U10418 : INV_X1 port map( A => n15208, ZN => n9558);
   U10419 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_797_port, B2 => n2653, 
                           ZN => n15208);
   U10420 : INV_X1 port map( A => n15207, ZN => n9559);
   U10421 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_796_port, B2 => n2653, 
                           ZN => n15207);
   U10422 : INV_X1 port map( A => n15206, ZN => n9560);
   U10423 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_795_port, B2 => n2653, 
                           ZN => n15206);
   U10424 : INV_X1 port map( A => n15205, ZN => n9561);
   U10425 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_794_port, B2 => n2653, 
                           ZN => n15205);
   U10426 : INV_X1 port map( A => n15204, ZN => n9562);
   U10427 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_793_port, B2 => n2653, 
                           ZN => n15204);
   U10428 : INV_X1 port map( A => n15203, ZN => n9563);
   U10429 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_792_port, B2 => n2653, 
                           ZN => n15203);
   U10430 : INV_X1 port map( A => n15202, ZN => n9564);
   U10431 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_791_port, B2 => n2652, 
                           ZN => n15202);
   U10432 : INV_X1 port map( A => n15201, ZN => n9565);
   U10433 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_790_port, B2 => n2652, 
                           ZN => n15201);
   U10434 : INV_X1 port map( A => n15200, ZN => n9566);
   U10435 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_789_port, B2 => n2652, 
                           ZN => n15200);
   U10436 : INV_X1 port map( A => n15199, ZN => n9567);
   U10437 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2648, B1 => 
                           DataPath_RF_bus_reg_dataout_788_port, B2 => n2652, 
                           ZN => n15199);
   U10438 : INV_X1 port map( A => n15198, ZN => n9568);
   U10439 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_787_port, B2 => n2652, 
                           ZN => n15198);
   U10440 : INV_X1 port map( A => n15197, ZN => n9569);
   U10441 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_786_port, B2 => n2652, 
                           ZN => n15197);
   U10442 : INV_X1 port map( A => n15196, ZN => n9570);
   U10443 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_785_port, B2 => n2652, 
                           ZN => n15196);
   U10444 : INV_X1 port map( A => n15195, ZN => n9571);
   U10445 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_784_port, B2 => n2652, 
                           ZN => n15195);
   U10446 : INV_X1 port map( A => n15194, ZN => n9572);
   U10447 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_783_port, B2 => n2652, 
                           ZN => n15194);
   U10448 : INV_X1 port map( A => n15193, ZN => n9573);
   U10449 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_782_port, B2 => n2652, 
                           ZN => n15193);
   U10450 : INV_X1 port map( A => n15192, ZN => n9574);
   U10451 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_781_port, B2 => n2652, 
                           ZN => n15192);
   U10452 : INV_X1 port map( A => n15191, ZN => n9575);
   U10453 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_780_port, B2 => n2652, 
                           ZN => n15191);
   U10454 : INV_X1 port map( A => n15190, ZN => n9576);
   U10455 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_779_port, B2 => n2651, 
                           ZN => n15190);
   U10456 : INV_X1 port map( A => n15189, ZN => n9577);
   U10457 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_778_port, B2 => n2651, 
                           ZN => n15189);
   U10458 : INV_X1 port map( A => n15188, ZN => n9578);
   U10459 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_777_port, B2 => n2651, 
                           ZN => n15188);
   U10460 : INV_X1 port map( A => n15187, ZN => n9579);
   U10461 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2649, B1 => 
                           DataPath_RF_bus_reg_dataout_776_port, B2 => n2651, 
                           ZN => n15187);
   U10462 : INV_X1 port map( A => n15186, ZN => n9580);
   U10463 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_775_port, B2 => n2651, 
                           ZN => n15186);
   U10464 : INV_X1 port map( A => n15185, ZN => n9581);
   U10465 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_774_port, B2 => n2651, 
                           ZN => n15185);
   U10466 : INV_X1 port map( A => n15184, ZN => n9582);
   U10467 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_773_port, B2 => n2651, 
                           ZN => n15184);
   U10468 : INV_X1 port map( A => n15183, ZN => n9583);
   U10469 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_772_port, B2 => n2651, 
                           ZN => n15183);
   U10470 : INV_X1 port map( A => n15182, ZN => n9584);
   U10471 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_771_port, B2 => n2651, 
                           ZN => n15182);
   U10472 : INV_X1 port map( A => n15181, ZN => n9585);
   U10473 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_770_port, B2 => n2651, 
                           ZN => n15181);
   U10474 : INV_X1 port map( A => n15180, ZN => n9586);
   U10475 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_769_port, B2 => n2651, 
                           ZN => n15180);
   U10476 : INV_X1 port map( A => n15177, ZN => n9587);
   U10477 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2650, B1 => 
                           DataPath_RF_bus_reg_dataout_768_port, B2 => n2651, 
                           ZN => n15177);
   U10478 : INV_X1 port map( A => n15244, ZN => n9588);
   U10479 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_831_port, B2 => n2659, 
                           ZN => n15244);
   U10480 : INV_X1 port map( A => n15243, ZN => n9589);
   U10481 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_830_port, B2 => n2659, 
                           ZN => n15243);
   U10482 : INV_X1 port map( A => n15242, ZN => n9590);
   U10483 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_829_port, B2 => n2659, 
                           ZN => n15242);
   U10484 : INV_X1 port map( A => n15241, ZN => n9591);
   U10485 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_828_port, B2 => n2659, 
                           ZN => n15241);
   U10486 : INV_X1 port map( A => n15240, ZN => n9592);
   U10487 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_827_port, B2 => n2659, 
                           ZN => n15240);
   U10488 : INV_X1 port map( A => n15239, ZN => n9593);
   U10489 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_826_port, B2 => n2659, 
                           ZN => n15239);
   U10490 : INV_X1 port map( A => n15238, ZN => n9594);
   U10491 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_825_port, B2 => n2659, 
                           ZN => n15238);
   U10492 : INV_X1 port map( A => n15237, ZN => n9595);
   U10493 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_824_port, B2 => n2659, 
                           ZN => n15237);
   U10494 : INV_X1 port map( A => n15236, ZN => n9596);
   U10495 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_823_port, B2 => n2658, 
                           ZN => n15236);
   U10496 : INV_X1 port map( A => n15235, ZN => n9597);
   U10497 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_822_port, B2 => n2658, 
                           ZN => n15235);
   U10498 : INV_X1 port map( A => n15234, ZN => n9598);
   U10499 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_821_port, B2 => n2658, 
                           ZN => n15234);
   U10500 : INV_X1 port map( A => n15233, ZN => n9599);
   U10501 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2654, B1 => 
                           DataPath_RF_bus_reg_dataout_820_port, B2 => n2658, 
                           ZN => n15233);
   U10502 : INV_X1 port map( A => n15232, ZN => n9600);
   U10503 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_819_port, B2 => n2658, 
                           ZN => n15232);
   U10504 : INV_X1 port map( A => n15231, ZN => n9601);
   U10505 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_818_port, B2 => n2658, 
                           ZN => n15231);
   U10506 : INV_X1 port map( A => n15230, ZN => n9602);
   U10507 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_817_port, B2 => n2658, 
                           ZN => n15230);
   U10508 : INV_X1 port map( A => n15229, ZN => n9603);
   U10509 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_816_port, B2 => n2658, 
                           ZN => n15229);
   U10510 : INV_X1 port map( A => n15228, ZN => n9604);
   U10511 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_815_port, B2 => n2658, 
                           ZN => n15228);
   U10512 : INV_X1 port map( A => n15227, ZN => n9605);
   U10513 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_814_port, B2 => n2658, 
                           ZN => n15227);
   U10514 : INV_X1 port map( A => n15226, ZN => n9606);
   U10515 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_813_port, B2 => n2658, 
                           ZN => n15226);
   U10516 : INV_X1 port map( A => n15225, ZN => n9607);
   U10517 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_812_port, B2 => n2658, 
                           ZN => n15225);
   U10518 : INV_X1 port map( A => n15224, ZN => n9608);
   U10519 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_811_port, B2 => n2657, 
                           ZN => n15224);
   U10520 : INV_X1 port map( A => n15223, ZN => n9609);
   U10521 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_810_port, B2 => n2657, 
                           ZN => n15223);
   U10522 : INV_X1 port map( A => n15222, ZN => n9610);
   U10523 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_809_port, B2 => n2657, 
                           ZN => n15222);
   U10524 : INV_X1 port map( A => n15221, ZN => n9611);
   U10525 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2655, B1 => 
                           DataPath_RF_bus_reg_dataout_808_port, B2 => n2657, 
                           ZN => n15221);
   U10526 : INV_X1 port map( A => n15220, ZN => n9612);
   U10527 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_807_port, B2 => n2657, 
                           ZN => n15220);
   U10528 : INV_X1 port map( A => n15219, ZN => n9613);
   U10529 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_806_port, B2 => n2657, 
                           ZN => n15219);
   U10530 : INV_X1 port map( A => n15218, ZN => n9614);
   U10531 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_805_port, B2 => n2657, 
                           ZN => n15218);
   U10532 : INV_X1 port map( A => n15217, ZN => n9615);
   U10533 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_804_port, B2 => n2657, 
                           ZN => n15217);
   U10534 : INV_X1 port map( A => n15216, ZN => n9616);
   U10535 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_803_port, B2 => n2657, 
                           ZN => n15216);
   U10536 : INV_X1 port map( A => n15215, ZN => n9617);
   U10537 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_802_port, B2 => n2657, 
                           ZN => n15215);
   U10538 : INV_X1 port map( A => n15214, ZN => n9618);
   U10539 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_801_port, B2 => n2657, 
                           ZN => n15214);
   U10540 : INV_X1 port map( A => n15211, ZN => n9619);
   U10541 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2656, B1 => 
                           DataPath_RF_bus_reg_dataout_800_port, B2 => n2657, 
                           ZN => n15211);
   U10542 : INV_X1 port map( A => n15278, ZN => n9620);
   U10543 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_863_port, B2 => n2665, 
                           ZN => n15278);
   U10544 : INV_X1 port map( A => n15277, ZN => n9621);
   U10545 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_862_port, B2 => n2665, 
                           ZN => n15277);
   U10546 : INV_X1 port map( A => n15276, ZN => n9622);
   U10547 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_861_port, B2 => n2665, 
                           ZN => n15276);
   U10548 : INV_X1 port map( A => n15275, ZN => n9623);
   U10549 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_860_port, B2 => n2665, 
                           ZN => n15275);
   U10550 : INV_X1 port map( A => n15274, ZN => n9624);
   U10551 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_859_port, B2 => n2665, 
                           ZN => n15274);
   U10552 : INV_X1 port map( A => n15273, ZN => n9625);
   U10553 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_858_port, B2 => n2665, 
                           ZN => n15273);
   U10554 : INV_X1 port map( A => n15272, ZN => n9626);
   U10555 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_857_port, B2 => n2665, 
                           ZN => n15272);
   U10556 : INV_X1 port map( A => n15271, ZN => n9627);
   U10557 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_856_port, B2 => n2665, 
                           ZN => n15271);
   U10558 : INV_X1 port map( A => n15270, ZN => n9628);
   U10559 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_855_port, B2 => n2664, 
                           ZN => n15270);
   U10560 : INV_X1 port map( A => n15269, ZN => n9629);
   U10561 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_854_port, B2 => n2664, 
                           ZN => n15269);
   U10562 : INV_X1 port map( A => n15268, ZN => n9630);
   U10563 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_853_port, B2 => n2664, 
                           ZN => n15268);
   U10564 : INV_X1 port map( A => n15267, ZN => n9631);
   U10565 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2660, B1 => 
                           DataPath_RF_bus_reg_dataout_852_port, B2 => n2664, 
                           ZN => n15267);
   U10566 : INV_X1 port map( A => n15266, ZN => n9632);
   U10567 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_851_port, B2 => n2664, 
                           ZN => n15266);
   U10568 : INV_X1 port map( A => n15265, ZN => n9633);
   U10569 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_850_port, B2 => n2664, 
                           ZN => n15265);
   U10570 : INV_X1 port map( A => n15264, ZN => n9634);
   U10571 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_849_port, B2 => n2664, 
                           ZN => n15264);
   U10572 : INV_X1 port map( A => n15263, ZN => n9635);
   U10573 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_848_port, B2 => n2664, 
                           ZN => n15263);
   U10574 : INV_X1 port map( A => n15262, ZN => n9636);
   U10575 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_847_port, B2 => n2664, 
                           ZN => n15262);
   U10576 : INV_X1 port map( A => n15261, ZN => n9637);
   U10577 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_846_port, B2 => n2664, 
                           ZN => n15261);
   U10578 : INV_X1 port map( A => n15260, ZN => n9638);
   U10579 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_845_port, B2 => n2664, 
                           ZN => n15260);
   U10580 : INV_X1 port map( A => n15259, ZN => n9639);
   U10581 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_844_port, B2 => n2664, 
                           ZN => n15259);
   U10582 : INV_X1 port map( A => n15258, ZN => n9640);
   U10583 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_843_port, B2 => n2663, 
                           ZN => n15258);
   U10584 : INV_X1 port map( A => n15257, ZN => n9641);
   U10585 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_842_port, B2 => n2663, 
                           ZN => n15257);
   U10586 : INV_X1 port map( A => n15256, ZN => n9642);
   U10587 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_841_port, B2 => n2663, 
                           ZN => n15256);
   U10588 : INV_X1 port map( A => n15255, ZN => n9643);
   U10589 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2661, B1 => 
                           DataPath_RF_bus_reg_dataout_840_port, B2 => n2663, 
                           ZN => n15255);
   U10590 : INV_X1 port map( A => n15254, ZN => n9644);
   U10591 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_839_port, B2 => n2663, 
                           ZN => n15254);
   U10592 : INV_X1 port map( A => n15253, ZN => n9645);
   U10593 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_838_port, B2 => n2663, 
                           ZN => n15253);
   U10594 : INV_X1 port map( A => n15252, ZN => n9646);
   U10595 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_837_port, B2 => n2663, 
                           ZN => n15252);
   U10596 : INV_X1 port map( A => n15251, ZN => n9647);
   U10597 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_836_port, B2 => n2663, 
                           ZN => n15251);
   U10598 : INV_X1 port map( A => n15250, ZN => n9648);
   U10599 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_835_port, B2 => n2663, 
                           ZN => n15250);
   U10600 : INV_X1 port map( A => n15249, ZN => n9649);
   U10601 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_834_port, B2 => n2663, 
                           ZN => n15249);
   U10602 : INV_X1 port map( A => n15248, ZN => n9650);
   U10603 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_833_port, B2 => n2663, 
                           ZN => n15248);
   U10604 : INV_X1 port map( A => n15245, ZN => n9651);
   U10605 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2662, B1 => 
                           DataPath_RF_bus_reg_dataout_832_port, B2 => n2663, 
                           ZN => n15245);
   U10606 : INV_X1 port map( A => n15312, ZN => n9652);
   U10607 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_895_port, B2 => n2671, 
                           ZN => n15312);
   U10608 : INV_X1 port map( A => n15311, ZN => n9653);
   U10609 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_894_port, B2 => n2671, 
                           ZN => n15311);
   U10610 : INV_X1 port map( A => n15310, ZN => n9654);
   U10611 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_893_port, B2 => n2671, 
                           ZN => n15310);
   U10612 : INV_X1 port map( A => n15309, ZN => n9655);
   U10613 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_892_port, B2 => n2671, 
                           ZN => n15309);
   U10614 : INV_X1 port map( A => n15308, ZN => n9656);
   U10615 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_891_port, B2 => n2671, 
                           ZN => n15308);
   U10616 : INV_X1 port map( A => n15307, ZN => n9657);
   U10617 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_890_port, B2 => n2671, 
                           ZN => n15307);
   U10618 : INV_X1 port map( A => n15306, ZN => n9658);
   U10619 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_889_port, B2 => n2671, 
                           ZN => n15306);
   U10620 : INV_X1 port map( A => n15305, ZN => n9659);
   U10621 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_888_port, B2 => n2671, 
                           ZN => n15305);
   U10622 : INV_X1 port map( A => n15304, ZN => n9660);
   U10623 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_887_port, B2 => n2670, 
                           ZN => n15304);
   U10624 : INV_X1 port map( A => n15303, ZN => n9661);
   U10625 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_886_port, B2 => n2670, 
                           ZN => n15303);
   U10626 : INV_X1 port map( A => n15302, ZN => n9662);
   U10627 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_885_port, B2 => n2670, 
                           ZN => n15302);
   U10628 : INV_X1 port map( A => n15301, ZN => n9663);
   U10629 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2666, B1 => 
                           DataPath_RF_bus_reg_dataout_884_port, B2 => n2670, 
                           ZN => n15301);
   U10630 : INV_X1 port map( A => n15300, ZN => n9664);
   U10631 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_883_port, B2 => n2670, 
                           ZN => n15300);
   U10632 : INV_X1 port map( A => n15299, ZN => n9665);
   U10633 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_882_port, B2 => n2670, 
                           ZN => n15299);
   U10634 : INV_X1 port map( A => n15298, ZN => n9666);
   U10635 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_881_port, B2 => n2670, 
                           ZN => n15298);
   U10636 : INV_X1 port map( A => n15297, ZN => n9667);
   U10637 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_880_port, B2 => n2670, 
                           ZN => n15297);
   U10638 : INV_X1 port map( A => n15296, ZN => n9668);
   U10639 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_879_port, B2 => n2670, 
                           ZN => n15296);
   U10640 : INV_X1 port map( A => n15295, ZN => n9669);
   U10641 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_878_port, B2 => n2670, 
                           ZN => n15295);
   U10642 : INV_X1 port map( A => n15294, ZN => n9670);
   U10643 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_877_port, B2 => n2670, 
                           ZN => n15294);
   U10644 : INV_X1 port map( A => n15293, ZN => n9671);
   U10645 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_876_port, B2 => n2670, 
                           ZN => n15293);
   U10646 : INV_X1 port map( A => n15292, ZN => n9672);
   U10647 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_875_port, B2 => n2669, 
                           ZN => n15292);
   U10648 : INV_X1 port map( A => n15291, ZN => n9673);
   U10649 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_874_port, B2 => n2669, 
                           ZN => n15291);
   U10650 : INV_X1 port map( A => n15290, ZN => n9674);
   U10651 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_873_port, B2 => n2669, 
                           ZN => n15290);
   U10652 : INV_X1 port map( A => n15289, ZN => n9675);
   U10653 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2667, B1 => 
                           DataPath_RF_bus_reg_dataout_872_port, B2 => n2669, 
                           ZN => n15289);
   U10654 : INV_X1 port map( A => n15288, ZN => n9676);
   U10655 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_871_port, B2 => n2669, 
                           ZN => n15288);
   U10656 : INV_X1 port map( A => n15287, ZN => n9677);
   U10657 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_870_port, B2 => n2669, 
                           ZN => n15287);
   U10658 : INV_X1 port map( A => n15286, ZN => n9678);
   U10659 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_869_port, B2 => n2669, 
                           ZN => n15286);
   U10660 : INV_X1 port map( A => n15285, ZN => n9679);
   U10661 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_868_port, B2 => n2669, 
                           ZN => n15285);
   U10662 : INV_X1 port map( A => n15284, ZN => n9680);
   U10663 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_867_port, B2 => n2669, 
                           ZN => n15284);
   U10664 : INV_X1 port map( A => n15283, ZN => n9681);
   U10665 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_866_port, B2 => n2669, 
                           ZN => n15283);
   U10666 : INV_X1 port map( A => n15282, ZN => n9682);
   U10667 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_865_port, B2 => n2669, 
                           ZN => n15282);
   U10668 : INV_X1 port map( A => n15279, ZN => n9683);
   U10669 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2668, B1 => 
                           DataPath_RF_bus_reg_dataout_864_port, B2 => n2669, 
                           ZN => n15279);
   U10670 : INV_X1 port map( A => n15346, ZN => n9684);
   U10671 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_927_port, B2 => n2677, 
                           ZN => n15346);
   U10672 : INV_X1 port map( A => n15345, ZN => n9685);
   U10673 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_926_port, B2 => n2677, 
                           ZN => n15345);
   U10674 : INV_X1 port map( A => n15344, ZN => n9686);
   U10675 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_925_port, B2 => n2677, 
                           ZN => n15344);
   U10676 : INV_X1 port map( A => n15343, ZN => n9687);
   U10677 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_924_port, B2 => n2677, 
                           ZN => n15343);
   U10678 : INV_X1 port map( A => n15342, ZN => n9688);
   U10679 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_923_port, B2 => n2677, 
                           ZN => n15342);
   U10680 : INV_X1 port map( A => n15341, ZN => n9689);
   U10681 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_922_port, B2 => n2677, 
                           ZN => n15341);
   U10682 : INV_X1 port map( A => n15340, ZN => n9690);
   U10683 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_921_port, B2 => n2677, 
                           ZN => n15340);
   U10684 : INV_X1 port map( A => n15339, ZN => n9691);
   U10685 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_920_port, B2 => n2677, 
                           ZN => n15339);
   U10686 : INV_X1 port map( A => n15338, ZN => n9692);
   U10687 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_919_port, B2 => n2676, 
                           ZN => n15338);
   U10688 : INV_X1 port map( A => n15337, ZN => n9693);
   U10689 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_918_port, B2 => n2676, 
                           ZN => n15337);
   U10690 : INV_X1 port map( A => n15336, ZN => n9694);
   U10691 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_917_port, B2 => n2676, 
                           ZN => n15336);
   U10692 : INV_X1 port map( A => n15335, ZN => n9695);
   U10693 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2672, B1 => 
                           DataPath_RF_bus_reg_dataout_916_port, B2 => n2676, 
                           ZN => n15335);
   U10694 : INV_X1 port map( A => n15334, ZN => n9696);
   U10695 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_915_port, B2 => n2676, 
                           ZN => n15334);
   U10696 : INV_X1 port map( A => n15333, ZN => n9697);
   U10697 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_914_port, B2 => n2676, 
                           ZN => n15333);
   U10698 : INV_X1 port map( A => n15332, ZN => n9698);
   U10699 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_913_port, B2 => n2676, 
                           ZN => n15332);
   U10700 : INV_X1 port map( A => n15331, ZN => n9699);
   U10701 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_912_port, B2 => n2676, 
                           ZN => n15331);
   U10702 : INV_X1 port map( A => n15330, ZN => n9700);
   U10703 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_911_port, B2 => n2676, 
                           ZN => n15330);
   U10704 : INV_X1 port map( A => n15329, ZN => n9701);
   U10705 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_910_port, B2 => n2676, 
                           ZN => n15329);
   U10706 : INV_X1 port map( A => n15328, ZN => n9702);
   U10707 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_909_port, B2 => n2676, 
                           ZN => n15328);
   U10708 : INV_X1 port map( A => n15327, ZN => n9703);
   U10709 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_908_port, B2 => n2676, 
                           ZN => n15327);
   U10710 : INV_X1 port map( A => n15326, ZN => n9704);
   U10711 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_907_port, B2 => n2675, 
                           ZN => n15326);
   U10712 : INV_X1 port map( A => n15325, ZN => n9705);
   U10713 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_906_port, B2 => n2675, 
                           ZN => n15325);
   U10714 : INV_X1 port map( A => n15324, ZN => n9706);
   U10715 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_905_port, B2 => n2675, 
                           ZN => n15324);
   U10716 : INV_X1 port map( A => n15323, ZN => n9707);
   U10717 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2673, B1 => 
                           DataPath_RF_bus_reg_dataout_904_port, B2 => n2675, 
                           ZN => n15323);
   U10718 : INV_X1 port map( A => n15322, ZN => n9708);
   U10719 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_903_port, B2 => n2675, 
                           ZN => n15322);
   U10720 : INV_X1 port map( A => n15321, ZN => n9709);
   U10721 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_902_port, B2 => n2675, 
                           ZN => n15321);
   U10722 : INV_X1 port map( A => n15320, ZN => n9710);
   U10723 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_901_port, B2 => n2675, 
                           ZN => n15320);
   U10724 : INV_X1 port map( A => n15319, ZN => n9711);
   U10725 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_900_port, B2 => n2675, 
                           ZN => n15319);
   U10726 : INV_X1 port map( A => n15318, ZN => n9712);
   U10727 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_899_port, B2 => n2675, 
                           ZN => n15318);
   U10728 : INV_X1 port map( A => n15317, ZN => n9713);
   U10729 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_898_port, B2 => n2675, 
                           ZN => n15317);
   U10730 : INV_X1 port map( A => n15316, ZN => n9714);
   U10731 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_897_port, B2 => n2675, 
                           ZN => n15316);
   U10732 : INV_X1 port map( A => n15313, ZN => n9715);
   U10733 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2674, B1 => 
                           DataPath_RF_bus_reg_dataout_896_port, B2 => n2675, 
                           ZN => n15313);
   U10734 : INV_X1 port map( A => n15380, ZN => n9716);
   U10735 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_959_port, B2 => n2683, 
                           ZN => n15380);
   U10736 : INV_X1 port map( A => n15379, ZN => n9717);
   U10737 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_958_port, B2 => n2683, 
                           ZN => n15379);
   U10738 : INV_X1 port map( A => n15378, ZN => n9718);
   U10739 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_957_port, B2 => n2683, 
                           ZN => n15378);
   U10740 : INV_X1 port map( A => n15377, ZN => n9719);
   U10741 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_956_port, B2 => n2683, 
                           ZN => n15377);
   U10742 : INV_X1 port map( A => n15376, ZN => n9720);
   U10743 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_955_port, B2 => n2683, 
                           ZN => n15376);
   U10744 : INV_X1 port map( A => n15375, ZN => n9721);
   U10745 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_954_port, B2 => n2683, 
                           ZN => n15375);
   U10746 : INV_X1 port map( A => n15374, ZN => n9722);
   U10747 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_953_port, B2 => n2683, 
                           ZN => n15374);
   U10748 : INV_X1 port map( A => n15373, ZN => n9723);
   U10749 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_952_port, B2 => n2683, 
                           ZN => n15373);
   U10750 : INV_X1 port map( A => n15372, ZN => n9724);
   U10751 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_951_port, B2 => n2682, 
                           ZN => n15372);
   U10752 : INV_X1 port map( A => n15371, ZN => n9725);
   U10753 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_950_port, B2 => n2682, 
                           ZN => n15371);
   U10754 : INV_X1 port map( A => n15370, ZN => n9726);
   U10755 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_949_port, B2 => n2682, 
                           ZN => n15370);
   U10756 : INV_X1 port map( A => n15369, ZN => n9727);
   U10757 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2678, B1 => 
                           DataPath_RF_bus_reg_dataout_948_port, B2 => n2682, 
                           ZN => n15369);
   U10758 : INV_X1 port map( A => n15368, ZN => n9728);
   U10759 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_947_port, B2 => n2682, 
                           ZN => n15368);
   U10760 : INV_X1 port map( A => n15367, ZN => n9729);
   U10761 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_946_port, B2 => n2682, 
                           ZN => n15367);
   U10762 : INV_X1 port map( A => n15366, ZN => n9730);
   U10763 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_945_port, B2 => n2682, 
                           ZN => n15366);
   U10764 : INV_X1 port map( A => n15365, ZN => n9731);
   U10765 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_944_port, B2 => n2682, 
                           ZN => n15365);
   U10766 : INV_X1 port map( A => n15364, ZN => n9732);
   U10767 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_943_port, B2 => n2682, 
                           ZN => n15364);
   U10768 : INV_X1 port map( A => n15363, ZN => n9733);
   U10769 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_942_port, B2 => n2682, 
                           ZN => n15363);
   U10770 : INV_X1 port map( A => n15362, ZN => n9734);
   U10771 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_941_port, B2 => n2682, 
                           ZN => n15362);
   U10772 : INV_X1 port map( A => n15361, ZN => n9735);
   U10773 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_940_port, B2 => n2682, 
                           ZN => n15361);
   U10774 : INV_X1 port map( A => n15360, ZN => n9736);
   U10775 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_939_port, B2 => n2681, 
                           ZN => n15360);
   U10776 : INV_X1 port map( A => n15359, ZN => n9737);
   U10777 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_938_port, B2 => n2681, 
                           ZN => n15359);
   U10778 : INV_X1 port map( A => n15358, ZN => n9738);
   U10779 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_937_port, B2 => n2681, 
                           ZN => n15358);
   U10780 : INV_X1 port map( A => n15357, ZN => n9739);
   U10781 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2679, B1 => 
                           DataPath_RF_bus_reg_dataout_936_port, B2 => n2681, 
                           ZN => n15357);
   U10782 : INV_X1 port map( A => n15356, ZN => n9740);
   U10783 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_935_port, B2 => n2681, 
                           ZN => n15356);
   U10784 : INV_X1 port map( A => n15355, ZN => n9741);
   U10785 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_934_port, B2 => n2681, 
                           ZN => n15355);
   U10786 : INV_X1 port map( A => n15354, ZN => n9742);
   U10787 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_933_port, B2 => n2681, 
                           ZN => n15354);
   U10788 : INV_X1 port map( A => n15353, ZN => n9743);
   U10789 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_932_port, B2 => n2681, 
                           ZN => n15353);
   U10790 : INV_X1 port map( A => n15352, ZN => n9744);
   U10791 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_931_port, B2 => n2681, 
                           ZN => n15352);
   U10792 : INV_X1 port map( A => n15351, ZN => n9745);
   U10793 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_930_port, B2 => n2681, 
                           ZN => n15351);
   U10794 : INV_X1 port map( A => n15350, ZN => n9746);
   U10795 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_929_port, B2 => n2681, 
                           ZN => n15350);
   U10796 : INV_X1 port map( A => n15347, ZN => n9747);
   U10797 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2680, B1 => 
                           DataPath_RF_bus_reg_dataout_928_port, B2 => n2681, 
                           ZN => n15347);
   U10798 : INV_X1 port map( A => n15414, ZN => n9748);
   U10799 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_991_port, B2 => n2689, 
                           ZN => n15414);
   U10800 : INV_X1 port map( A => n15413, ZN => n9749);
   U10801 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_990_port, B2 => n2689, 
                           ZN => n15413);
   U10802 : INV_X1 port map( A => n15412, ZN => n9750);
   U10803 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_989_port, B2 => n2689, 
                           ZN => n15412);
   U10804 : INV_X1 port map( A => n15411, ZN => n9751);
   U10805 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_988_port, B2 => n2689, 
                           ZN => n15411);
   U10806 : INV_X1 port map( A => n15410, ZN => n9752);
   U10807 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_987_port, B2 => n2689, 
                           ZN => n15410);
   U10808 : INV_X1 port map( A => n15409, ZN => n9753);
   U10809 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_986_port, B2 => n2689, 
                           ZN => n15409);
   U10810 : INV_X1 port map( A => n15408, ZN => n9754);
   U10811 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_985_port, B2 => n2689, 
                           ZN => n15408);
   U10812 : INV_X1 port map( A => n15407, ZN => n9755);
   U10813 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_984_port, B2 => n2689, 
                           ZN => n15407);
   U10814 : INV_X1 port map( A => n15406, ZN => n9756);
   U10815 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_983_port, B2 => n2688, 
                           ZN => n15406);
   U10816 : INV_X1 port map( A => n15405, ZN => n9757);
   U10817 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_982_port, B2 => n2688, 
                           ZN => n15405);
   U10818 : INV_X1 port map( A => n15404, ZN => n9758);
   U10819 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_981_port, B2 => n2688, 
                           ZN => n15404);
   U10820 : INV_X1 port map( A => n15403, ZN => n9759);
   U10821 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2684, B1 => 
                           DataPath_RF_bus_reg_dataout_980_port, B2 => n2688, 
                           ZN => n15403);
   U10822 : INV_X1 port map( A => n15402, ZN => n9760);
   U10823 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_979_port, B2 => n2688, 
                           ZN => n15402);
   U10824 : INV_X1 port map( A => n15401, ZN => n9761);
   U10825 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_978_port, B2 => n2688, 
                           ZN => n15401);
   U10826 : INV_X1 port map( A => n15400, ZN => n9762);
   U10827 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_977_port, B2 => n2688, 
                           ZN => n15400);
   U10828 : INV_X1 port map( A => n15399, ZN => n9763);
   U10829 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_976_port, B2 => n2688, 
                           ZN => n15399);
   U10830 : INV_X1 port map( A => n15398, ZN => n9764);
   U10831 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_975_port, B2 => n2688, 
                           ZN => n15398);
   U10832 : INV_X1 port map( A => n15397, ZN => n9765);
   U10833 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_974_port, B2 => n2688, 
                           ZN => n15397);
   U10834 : INV_X1 port map( A => n15396, ZN => n9766);
   U10835 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_973_port, B2 => n2688, 
                           ZN => n15396);
   U10836 : INV_X1 port map( A => n15395, ZN => n9767);
   U10837 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_972_port, B2 => n2688, 
                           ZN => n15395);
   U10838 : INV_X1 port map( A => n15394, ZN => n9768);
   U10839 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_971_port, B2 => n2687, 
                           ZN => n15394);
   U10840 : INV_X1 port map( A => n15393, ZN => n9769);
   U10841 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_970_port, B2 => n2687, 
                           ZN => n15393);
   U10842 : INV_X1 port map( A => n15392, ZN => n9770);
   U10843 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_969_port, B2 => n2687, 
                           ZN => n15392);
   U10844 : INV_X1 port map( A => n15391, ZN => n9771);
   U10845 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2685, B1 => 
                           DataPath_RF_bus_reg_dataout_968_port, B2 => n2687, 
                           ZN => n15391);
   U10846 : INV_X1 port map( A => n15390, ZN => n9772);
   U10847 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_967_port, B2 => n2687, 
                           ZN => n15390);
   U10848 : INV_X1 port map( A => n15389, ZN => n9773);
   U10849 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_966_port, B2 => n2687, 
                           ZN => n15389);
   U10850 : INV_X1 port map( A => n15388, ZN => n9774);
   U10851 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_965_port, B2 => n2687, 
                           ZN => n15388);
   U10852 : INV_X1 port map( A => n15387, ZN => n9775);
   U10853 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_964_port, B2 => n2687, 
                           ZN => n15387);
   U10854 : INV_X1 port map( A => n15386, ZN => n9776);
   U10855 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_963_port, B2 => n2687, 
                           ZN => n15386);
   U10856 : INV_X1 port map( A => n15385, ZN => n9777);
   U10857 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_962_port, B2 => n2687, 
                           ZN => n15385);
   U10858 : INV_X1 port map( A => n15384, ZN => n9778);
   U10859 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_961_port, B2 => n2687, 
                           ZN => n15384);
   U10860 : INV_X1 port map( A => n15381, ZN => n9779);
   U10861 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2686, B1 => 
                           DataPath_RF_bus_reg_dataout_960_port, B2 => n2687, 
                           ZN => n15381);
   U10862 : INV_X1 port map( A => n15448, ZN => n9780);
   U10863 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_31_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1023_port, B2 => n2695, 
                           ZN => n15448);
   U10864 : INV_X1 port map( A => n15447, ZN => n9781);
   U10865 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_30_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1022_port, B2 => n2695, 
                           ZN => n15447);
   U10866 : INV_X1 port map( A => n15446, ZN => n9782);
   U10867 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_29_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1021_port, B2 => n2695, 
                           ZN => n15446);
   U10868 : INV_X1 port map( A => n15445, ZN => n9783);
   U10869 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_28_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1020_port, B2 => n2695, 
                           ZN => n15445);
   U10870 : INV_X1 port map( A => n15444, ZN => n9784);
   U10871 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_27_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1019_port, B2 => n2695, 
                           ZN => n15444);
   U10872 : INV_X1 port map( A => n15443, ZN => n9785);
   U10873 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_26_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1018_port, B2 => n2695, 
                           ZN => n15443);
   U10874 : INV_X1 port map( A => n15442, ZN => n9786);
   U10875 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_25_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1017_port, B2 => n2695, 
                           ZN => n15442);
   U10876 : INV_X1 port map( A => n15441, ZN => n9787);
   U10877 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_24_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1016_port, B2 => n2695, 
                           ZN => n15441);
   U10878 : INV_X1 port map( A => n15440, ZN => n9788);
   U10879 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_23_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1015_port, B2 => n2694, 
                           ZN => n15440);
   U10880 : INV_X1 port map( A => n15439, ZN => n9789);
   U10881 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_22_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1014_port, B2 => n2694, 
                           ZN => n15439);
   U10882 : INV_X1 port map( A => n15438, ZN => n9790);
   U10883 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_21_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1013_port, B2 => n2694, 
                           ZN => n15438);
   U10884 : INV_X1 port map( A => n15437, ZN => n9791);
   U10885 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_20_port,
                           A2 => n2690, B1 => 
                           DataPath_RF_bus_reg_dataout_1012_port, B2 => n2694, 
                           ZN => n15437);
   U10886 : INV_X1 port map( A => n15436, ZN => n9792);
   U10887 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_19_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1011_port, B2 => n2694, 
                           ZN => n15436);
   U10888 : INV_X1 port map( A => n15435, ZN => n9793);
   U10889 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_18_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1010_port, B2 => n2694, 
                           ZN => n15435);
   U10890 : INV_X1 port map( A => n15434, ZN => n9794);
   U10891 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_17_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1009_port, B2 => n2694, 
                           ZN => n15434);
   U10892 : INV_X1 port map( A => n15433, ZN => n9795);
   U10893 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_16_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1008_port, B2 => n2694, 
                           ZN => n15433);
   U10894 : INV_X1 port map( A => n15432, ZN => n9796);
   U10895 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_15_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1007_port, B2 => n2694, 
                           ZN => n15432);
   U10896 : INV_X1 port map( A => n15431, ZN => n9797);
   U10897 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_14_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1006_port, B2 => n2694, 
                           ZN => n15431);
   U10898 : INV_X1 port map( A => n15430, ZN => n9798);
   U10899 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_13_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1005_port, B2 => n2694, 
                           ZN => n15430);
   U10900 : INV_X1 port map( A => n15429, ZN => n9799);
   U10901 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_12_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1004_port, B2 => n2694, 
                           ZN => n15429);
   U10902 : INV_X1 port map( A => n15428, ZN => n9800);
   U10903 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_11_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1003_port, B2 => n2693, 
                           ZN => n15428);
   U10904 : INV_X1 port map( A => n15427, ZN => n9801);
   U10905 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_10_port,
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1002_port, B2 => n2693, 
                           ZN => n15427);
   U10906 : INV_X1 port map( A => n15426, ZN => n9802);
   U10907 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_9_port, 
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1001_port, B2 => n2693, 
                           ZN => n15426);
   U10908 : INV_X1 port map( A => n15425, ZN => n9803);
   U10909 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_8_port, 
                           A2 => n2691, B1 => 
                           DataPath_RF_bus_reg_dataout_1000_port, B2 => n2693, 
                           ZN => n15425);
   U10910 : INV_X1 port map( A => n15424, ZN => n9804);
   U10911 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_7_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_999_port, B2 => n2693, 
                           ZN => n15424);
   U10912 : INV_X1 port map( A => n15423, ZN => n9805);
   U10913 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_6_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_998_port, B2 => n2693, 
                           ZN => n15423);
   U10914 : INV_X1 port map( A => n15422, ZN => n9806);
   U10915 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_5_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_997_port, B2 => n2693, 
                           ZN => n15422);
   U10916 : INV_X1 port map( A => n15421, ZN => n9807);
   U10917 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_4_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_996_port, B2 => n2693, 
                           ZN => n15421);
   U10918 : INV_X1 port map( A => n15420, ZN => n9808);
   U10919 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_3_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_995_port, B2 => n2693, 
                           ZN => n15420);
   U10920 : INV_X1 port map( A => n15419, ZN => n9809);
   U10921 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_2_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_994_port, B2 => n2693, 
                           ZN => n15419);
   U10922 : INV_X1 port map( A => n15418, ZN => n9810);
   U10923 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_1_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_993_port, B2 => n2693, 
                           ZN => n15418);
   U10924 : INV_X1 port map( A => n15415, ZN => n9811);
   U10925 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_1_0_port, 
                           A2 => n2692, B1 => 
                           DataPath_RF_bus_reg_dataout_992_port, B2 => n2693, 
                           ZN => n15415);
   U10926 : INV_X1 port map( A => n15482, ZN => n9812);
   U10927 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1055_port, B2 => n2701, 
                           ZN => n15482);
   U10928 : INV_X1 port map( A => n15481, ZN => n9813);
   U10929 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1054_port, B2 => n2701, 
                           ZN => n15481);
   U10930 : INV_X1 port map( A => n15480, ZN => n9814);
   U10931 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1053_port, B2 => n2701, 
                           ZN => n15480);
   U10932 : INV_X1 port map( A => n15479, ZN => n9815);
   U10933 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1052_port, B2 => n2701, 
                           ZN => n15479);
   U10934 : INV_X1 port map( A => n15478, ZN => n9816);
   U10935 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1051_port, B2 => n2701, 
                           ZN => n15478);
   U10936 : INV_X1 port map( A => n15477, ZN => n9817);
   U10937 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1050_port, B2 => n2701, 
                           ZN => n15477);
   U10938 : INV_X1 port map( A => n15476, ZN => n9818);
   U10939 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1049_port, B2 => n2701, 
                           ZN => n15476);
   U10940 : INV_X1 port map( A => n15475, ZN => n9819);
   U10941 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1048_port, B2 => n2701, 
                           ZN => n15475);
   U10942 : INV_X1 port map( A => n15474, ZN => n9820);
   U10943 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1047_port, B2 => n2700, 
                           ZN => n15474);
   U10944 : INV_X1 port map( A => n15473, ZN => n9821);
   U10945 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1046_port, B2 => n2700, 
                           ZN => n15473);
   U10946 : INV_X1 port map( A => n15472, ZN => n9822);
   U10947 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1045_port, B2 => n2700, 
                           ZN => n15472);
   U10948 : INV_X1 port map( A => n15471, ZN => n9823);
   U10949 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2696, B1 => 
                           DataPath_RF_bus_reg_dataout_1044_port, B2 => n2700, 
                           ZN => n15471);
   U10950 : INV_X1 port map( A => n15470, ZN => n9824);
   U10951 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1043_port, B2 => n2700, 
                           ZN => n15470);
   U10952 : INV_X1 port map( A => n15469, ZN => n9825);
   U10953 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1042_port, B2 => n2700, 
                           ZN => n15469);
   U10954 : INV_X1 port map( A => n15468, ZN => n9826);
   U10955 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1041_port, B2 => n2700, 
                           ZN => n15468);
   U10956 : INV_X1 port map( A => n15467, ZN => n9827);
   U10957 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1040_port, B2 => n2700, 
                           ZN => n15467);
   U10958 : INV_X1 port map( A => n15466, ZN => n9828);
   U10959 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1039_port, B2 => n2700, 
                           ZN => n15466);
   U10960 : INV_X1 port map( A => n15465, ZN => n9829);
   U10961 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1038_port, B2 => n2700, 
                           ZN => n15465);
   U10962 : INV_X1 port map( A => n15464, ZN => n9830);
   U10963 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1037_port, B2 => n2700, 
                           ZN => n15464);
   U10964 : INV_X1 port map( A => n15463, ZN => n9831);
   U10965 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1036_port, B2 => n2700, 
                           ZN => n15463);
   U10966 : INV_X1 port map( A => n15462, ZN => n9832);
   U10967 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1035_port, B2 => n2699, 
                           ZN => n15462);
   U10968 : INV_X1 port map( A => n15461, ZN => n9833);
   U10969 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1034_port, B2 => n2699, 
                           ZN => n15461);
   U10970 : INV_X1 port map( A => n15460, ZN => n9834);
   U10971 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1033_port, B2 => n2699, 
                           ZN => n15460);
   U10972 : INV_X1 port map( A => n15459, ZN => n9835);
   U10973 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2697, B1 => 
                           DataPath_RF_bus_reg_dataout_1032_port, B2 => n2699, 
                           ZN => n15459);
   U10974 : INV_X1 port map( A => n15458, ZN => n9836);
   U10975 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1031_port, B2 => n2699, 
                           ZN => n15458);
   U10976 : INV_X1 port map( A => n15457, ZN => n9837);
   U10977 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1030_port, B2 => n2699, 
                           ZN => n15457);
   U10978 : INV_X1 port map( A => n15456, ZN => n9838);
   U10979 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1029_port, B2 => n2699, 
                           ZN => n15456);
   U10980 : INV_X1 port map( A => n15455, ZN => n9839);
   U10981 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1028_port, B2 => n2699, 
                           ZN => n15455);
   U10982 : INV_X1 port map( A => n15454, ZN => n9840);
   U10983 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1027_port, B2 => n2699, 
                           ZN => n15454);
   U10984 : INV_X1 port map( A => n15453, ZN => n9841);
   U10985 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1026_port, B2 => n2699, 
                           ZN => n15453);
   U10986 : INV_X1 port map( A => n15452, ZN => n9842);
   U10987 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1025_port, B2 => n2699, 
                           ZN => n15452);
   U10988 : INV_X1 port map( A => n15449, ZN => n9843);
   U10989 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2698, B1 => 
                           DataPath_RF_bus_reg_dataout_1024_port, B2 => n2699, 
                           ZN => n15449);
   U10990 : INV_X1 port map( A => n15516, ZN => n9844);
   U10991 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1087_port, B2 => n2707, 
                           ZN => n15516);
   U10992 : INV_X1 port map( A => n15515, ZN => n9845);
   U10993 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1086_port, B2 => n2707, 
                           ZN => n15515);
   U10994 : INV_X1 port map( A => n15514, ZN => n9846);
   U10995 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1085_port, B2 => n2707, 
                           ZN => n15514);
   U10996 : INV_X1 port map( A => n15513, ZN => n9847);
   U10997 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1084_port, B2 => n2707, 
                           ZN => n15513);
   U10998 : INV_X1 port map( A => n15512, ZN => n9848);
   U10999 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1083_port, B2 => n2707, 
                           ZN => n15512);
   U11000 : INV_X1 port map( A => n15511, ZN => n9849);
   U11001 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1082_port, B2 => n2707, 
                           ZN => n15511);
   U11002 : INV_X1 port map( A => n15510, ZN => n9850);
   U11003 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1081_port, B2 => n2707, 
                           ZN => n15510);
   U11004 : INV_X1 port map( A => n15509, ZN => n9851);
   U11005 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1080_port, B2 => n2707, 
                           ZN => n15509);
   U11006 : INV_X1 port map( A => n15508, ZN => n9852);
   U11007 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1079_port, B2 => n2706, 
                           ZN => n15508);
   U11008 : INV_X1 port map( A => n15507, ZN => n9853);
   U11009 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1078_port, B2 => n2706, 
                           ZN => n15507);
   U11010 : INV_X1 port map( A => n15506, ZN => n9854);
   U11011 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1077_port, B2 => n2706, 
                           ZN => n15506);
   U11012 : INV_X1 port map( A => n15505, ZN => n9855);
   U11013 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2702, B1 => 
                           DataPath_RF_bus_reg_dataout_1076_port, B2 => n2706, 
                           ZN => n15505);
   U11014 : INV_X1 port map( A => n15504, ZN => n9856);
   U11015 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1075_port, B2 => n2706, 
                           ZN => n15504);
   U11016 : INV_X1 port map( A => n15503, ZN => n9857);
   U11017 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1074_port, B2 => n2706, 
                           ZN => n15503);
   U11018 : INV_X1 port map( A => n15502, ZN => n9858);
   U11019 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1073_port, B2 => n2706, 
                           ZN => n15502);
   U11020 : INV_X1 port map( A => n15501, ZN => n9859);
   U11021 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1072_port, B2 => n2706, 
                           ZN => n15501);
   U11022 : INV_X1 port map( A => n15500, ZN => n9860);
   U11023 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1071_port, B2 => n2706, 
                           ZN => n15500);
   U11024 : INV_X1 port map( A => n15499, ZN => n9861);
   U11025 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1070_port, B2 => n2706, 
                           ZN => n15499);
   U11026 : INV_X1 port map( A => n15498, ZN => n9862);
   U11027 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1069_port, B2 => n2706, 
                           ZN => n15498);
   U11028 : INV_X1 port map( A => n15497, ZN => n9863);
   U11029 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1068_port, B2 => n2706, 
                           ZN => n15497);
   U11030 : INV_X1 port map( A => n15496, ZN => n9864);
   U11031 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1067_port, B2 => n2705, 
                           ZN => n15496);
   U11032 : INV_X1 port map( A => n15495, ZN => n9865);
   U11033 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1066_port, B2 => n2705, 
                           ZN => n15495);
   U11034 : INV_X1 port map( A => n15494, ZN => n9866);
   U11035 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1065_port, B2 => n2705, 
                           ZN => n15494);
   U11036 : INV_X1 port map( A => n15493, ZN => n9867);
   U11037 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2703, B1 => 
                           DataPath_RF_bus_reg_dataout_1064_port, B2 => n2705, 
                           ZN => n15493);
   U11038 : INV_X1 port map( A => n15492, ZN => n9868);
   U11039 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1063_port, B2 => n2705, 
                           ZN => n15492);
   U11040 : INV_X1 port map( A => n15491, ZN => n9869);
   U11041 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1062_port, B2 => n2705, 
                           ZN => n15491);
   U11042 : INV_X1 port map( A => n15490, ZN => n9870);
   U11043 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1061_port, B2 => n2705, 
                           ZN => n15490);
   U11044 : INV_X1 port map( A => n15489, ZN => n9871);
   U11045 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1060_port, B2 => n2705, 
                           ZN => n15489);
   U11046 : INV_X1 port map( A => n15488, ZN => n9872);
   U11047 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1059_port, B2 => n2705, 
                           ZN => n15488);
   U11048 : INV_X1 port map( A => n15487, ZN => n9873);
   U11049 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1058_port, B2 => n2705, 
                           ZN => n15487);
   U11050 : INV_X1 port map( A => n15486, ZN => n9874);
   U11051 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1057_port, B2 => n2705, 
                           ZN => n15486);
   U11052 : INV_X1 port map( A => n15483, ZN => n9875);
   U11053 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2704, B1 => 
                           DataPath_RF_bus_reg_dataout_1056_port, B2 => n2705, 
                           ZN => n15483);
   U11054 : INV_X1 port map( A => n15550, ZN => n9876);
   U11055 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1119_port, B2 => n2713, 
                           ZN => n15550);
   U11056 : INV_X1 port map( A => n15549, ZN => n9877);
   U11057 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1118_port, B2 => n2713, 
                           ZN => n15549);
   U11058 : INV_X1 port map( A => n15548, ZN => n9878);
   U11059 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1117_port, B2 => n2713, 
                           ZN => n15548);
   U11060 : INV_X1 port map( A => n15547, ZN => n9879);
   U11061 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1116_port, B2 => n2713, 
                           ZN => n15547);
   U11062 : INV_X1 port map( A => n15546, ZN => n9880);
   U11063 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1115_port, B2 => n2713, 
                           ZN => n15546);
   U11064 : INV_X1 port map( A => n15545, ZN => n9881);
   U11065 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1114_port, B2 => n2713, 
                           ZN => n15545);
   U11066 : INV_X1 port map( A => n15544, ZN => n9882);
   U11067 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1113_port, B2 => n2713, 
                           ZN => n15544);
   U11068 : INV_X1 port map( A => n15543, ZN => n9883);
   U11069 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1112_port, B2 => n2713, 
                           ZN => n15543);
   U11070 : INV_X1 port map( A => n15542, ZN => n9884);
   U11071 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1111_port, B2 => n2712, 
                           ZN => n15542);
   U11072 : INV_X1 port map( A => n15541, ZN => n9885);
   U11073 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1110_port, B2 => n2712, 
                           ZN => n15541);
   U11074 : INV_X1 port map( A => n15540, ZN => n9886);
   U11075 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1109_port, B2 => n2712, 
                           ZN => n15540);
   U11076 : INV_X1 port map( A => n15539, ZN => n9887);
   U11077 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2708, B1 => 
                           DataPath_RF_bus_reg_dataout_1108_port, B2 => n2712, 
                           ZN => n15539);
   U11078 : INV_X1 port map( A => n15538, ZN => n9888);
   U11079 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1107_port, B2 => n2712, 
                           ZN => n15538);
   U11080 : INV_X1 port map( A => n15537, ZN => n9889);
   U11081 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1106_port, B2 => n2712, 
                           ZN => n15537);
   U11082 : INV_X1 port map( A => n15536, ZN => n9890);
   U11083 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1105_port, B2 => n2712, 
                           ZN => n15536);
   U11084 : INV_X1 port map( A => n15535, ZN => n9891);
   U11085 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1104_port, B2 => n2712, 
                           ZN => n15535);
   U11086 : INV_X1 port map( A => n15534, ZN => n9892);
   U11087 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1103_port, B2 => n2712, 
                           ZN => n15534);
   U11088 : INV_X1 port map( A => n15533, ZN => n9893);
   U11089 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1102_port, B2 => n2712, 
                           ZN => n15533);
   U11090 : INV_X1 port map( A => n15532, ZN => n9894);
   U11091 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1101_port, B2 => n2712, 
                           ZN => n15532);
   U11092 : INV_X1 port map( A => n15531, ZN => n9895);
   U11093 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1100_port, B2 => n2712, 
                           ZN => n15531);
   U11094 : INV_X1 port map( A => n15530, ZN => n9896);
   U11095 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1099_port, B2 => n2711, 
                           ZN => n15530);
   U11096 : INV_X1 port map( A => n15529, ZN => n9897);
   U11097 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1098_port, B2 => n2711, 
                           ZN => n15529);
   U11098 : INV_X1 port map( A => n15528, ZN => n9898);
   U11099 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1097_port, B2 => n2711, 
                           ZN => n15528);
   U11100 : INV_X1 port map( A => n15527, ZN => n9899);
   U11101 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2709, B1 => 
                           DataPath_RF_bus_reg_dataout_1096_port, B2 => n2711, 
                           ZN => n15527);
   U11102 : INV_X1 port map( A => n15526, ZN => n9900);
   U11103 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1095_port, B2 => n2711, 
                           ZN => n15526);
   U11104 : INV_X1 port map( A => n15525, ZN => n9901);
   U11105 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1094_port, B2 => n2711, 
                           ZN => n15525);
   U11106 : INV_X1 port map( A => n15524, ZN => n9902);
   U11107 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1093_port, B2 => n2711, 
                           ZN => n15524);
   U11108 : INV_X1 port map( A => n15523, ZN => n9903);
   U11109 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1092_port, B2 => n2711, 
                           ZN => n15523);
   U11110 : INV_X1 port map( A => n15522, ZN => n9904);
   U11111 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1091_port, B2 => n2711, 
                           ZN => n15522);
   U11112 : INV_X1 port map( A => n15521, ZN => n9905);
   U11113 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1090_port, B2 => n2711, 
                           ZN => n15521);
   U11114 : INV_X1 port map( A => n15520, ZN => n9906);
   U11115 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1089_port, B2 => n2711, 
                           ZN => n15520);
   U11116 : INV_X1 port map( A => n15517, ZN => n9907);
   U11117 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2710, B1 => 
                           DataPath_RF_bus_reg_dataout_1088_port, B2 => n2711, 
                           ZN => n15517);
   U11118 : INV_X1 port map( A => n15584, ZN => n9908);
   U11119 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1151_port, B2 => n2719, 
                           ZN => n15584);
   U11120 : INV_X1 port map( A => n15583, ZN => n9909);
   U11121 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1150_port, B2 => n2719, 
                           ZN => n15583);
   U11122 : INV_X1 port map( A => n15582, ZN => n9910);
   U11123 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1149_port, B2 => n2719, 
                           ZN => n15582);
   U11124 : INV_X1 port map( A => n15581, ZN => n9911);
   U11125 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1148_port, B2 => n2719, 
                           ZN => n15581);
   U11126 : INV_X1 port map( A => n15580, ZN => n9912);
   U11127 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1147_port, B2 => n2719, 
                           ZN => n15580);
   U11128 : INV_X1 port map( A => n15579, ZN => n9913);
   U11129 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1146_port, B2 => n2719, 
                           ZN => n15579);
   U11130 : INV_X1 port map( A => n15578, ZN => n9914);
   U11131 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1145_port, B2 => n2719, 
                           ZN => n15578);
   U11132 : INV_X1 port map( A => n15577, ZN => n9915);
   U11133 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1144_port, B2 => n2719, 
                           ZN => n15577);
   U11134 : INV_X1 port map( A => n15576, ZN => n9916);
   U11135 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1143_port, B2 => n2718, 
                           ZN => n15576);
   U11136 : INV_X1 port map( A => n15575, ZN => n9917);
   U11137 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1142_port, B2 => n2718, 
                           ZN => n15575);
   U11138 : INV_X1 port map( A => n15574, ZN => n9918);
   U11139 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1141_port, B2 => n2718, 
                           ZN => n15574);
   U11140 : INV_X1 port map( A => n15573, ZN => n9919);
   U11141 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2714, B1 => 
                           DataPath_RF_bus_reg_dataout_1140_port, B2 => n2718, 
                           ZN => n15573);
   U11142 : INV_X1 port map( A => n15572, ZN => n9920);
   U11143 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1139_port, B2 => n2718, 
                           ZN => n15572);
   U11144 : INV_X1 port map( A => n15571, ZN => n9921);
   U11145 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1138_port, B2 => n2718, 
                           ZN => n15571);
   U11146 : INV_X1 port map( A => n15570, ZN => n9922);
   U11147 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1137_port, B2 => n2718, 
                           ZN => n15570);
   U11148 : INV_X1 port map( A => n15569, ZN => n9923);
   U11149 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1136_port, B2 => n2718, 
                           ZN => n15569);
   U11150 : INV_X1 port map( A => n15568, ZN => n9924);
   U11151 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1135_port, B2 => n2718, 
                           ZN => n15568);
   U11152 : INV_X1 port map( A => n15567, ZN => n9925);
   U11153 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1134_port, B2 => n2718, 
                           ZN => n15567);
   U11154 : INV_X1 port map( A => n15566, ZN => n9926);
   U11155 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1133_port, B2 => n2718, 
                           ZN => n15566);
   U11156 : INV_X1 port map( A => n15565, ZN => n9927);
   U11157 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1132_port, B2 => n2718, 
                           ZN => n15565);
   U11158 : INV_X1 port map( A => n15564, ZN => n9928);
   U11159 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1131_port, B2 => n2717, 
                           ZN => n15564);
   U11160 : INV_X1 port map( A => n15563, ZN => n9929);
   U11161 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1130_port, B2 => n2717, 
                           ZN => n15563);
   U11162 : INV_X1 port map( A => n15562, ZN => n9930);
   U11163 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1129_port, B2 => n2717, 
                           ZN => n15562);
   U11164 : INV_X1 port map( A => n15561, ZN => n9931);
   U11165 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2715, B1 => 
                           DataPath_RF_bus_reg_dataout_1128_port, B2 => n2717, 
                           ZN => n15561);
   U11166 : INV_X1 port map( A => n15560, ZN => n9932);
   U11167 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1127_port, B2 => n2717, 
                           ZN => n15560);
   U11168 : INV_X1 port map( A => n15559, ZN => n9933);
   U11169 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1126_port, B2 => n2717, 
                           ZN => n15559);
   U11170 : INV_X1 port map( A => n15558, ZN => n9934);
   U11171 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1125_port, B2 => n2717, 
                           ZN => n15558);
   U11172 : INV_X1 port map( A => n15557, ZN => n9935);
   U11173 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1124_port, B2 => n2717, 
                           ZN => n15557);
   U11174 : INV_X1 port map( A => n15556, ZN => n9936);
   U11175 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1123_port, B2 => n2717, 
                           ZN => n15556);
   U11176 : INV_X1 port map( A => n15555, ZN => n9937);
   U11177 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1122_port, B2 => n2717, 
                           ZN => n15555);
   U11178 : INV_X1 port map( A => n15554, ZN => n9938);
   U11179 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1121_port, B2 => n2717, 
                           ZN => n15554);
   U11180 : INV_X1 port map( A => n15551, ZN => n9939);
   U11181 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2716, B1 => 
                           DataPath_RF_bus_reg_dataout_1120_port, B2 => n2717, 
                           ZN => n15551);
   U11182 : INV_X1 port map( A => n15618, ZN => n9940);
   U11183 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1183_port, B2 => n2725, 
                           ZN => n15618);
   U11184 : INV_X1 port map( A => n15617, ZN => n9941);
   U11185 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1182_port, B2 => n2725, 
                           ZN => n15617);
   U11186 : INV_X1 port map( A => n15616, ZN => n9942);
   U11187 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1181_port, B2 => n2725, 
                           ZN => n15616);
   U11188 : INV_X1 port map( A => n15615, ZN => n9943);
   U11189 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1180_port, B2 => n2725, 
                           ZN => n15615);
   U11190 : INV_X1 port map( A => n15614, ZN => n9944);
   U11191 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1179_port, B2 => n2725, 
                           ZN => n15614);
   U11192 : INV_X1 port map( A => n15613, ZN => n9945);
   U11193 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1178_port, B2 => n2725, 
                           ZN => n15613);
   U11194 : INV_X1 port map( A => n15612, ZN => n9946);
   U11195 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1177_port, B2 => n2725, 
                           ZN => n15612);
   U11196 : INV_X1 port map( A => n15611, ZN => n9947);
   U11197 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1176_port, B2 => n2725, 
                           ZN => n15611);
   U11198 : INV_X1 port map( A => n15610, ZN => n9948);
   U11199 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1175_port, B2 => n2724, 
                           ZN => n15610);
   U11200 : INV_X1 port map( A => n15609, ZN => n9949);
   U11201 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1174_port, B2 => n2724, 
                           ZN => n15609);
   U11202 : INV_X1 port map( A => n15608, ZN => n9950);
   U11203 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1173_port, B2 => n2724, 
                           ZN => n15608);
   U11204 : INV_X1 port map( A => n15607, ZN => n9951);
   U11205 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2720, B1 => 
                           DataPath_RF_bus_reg_dataout_1172_port, B2 => n2724, 
                           ZN => n15607);
   U11206 : INV_X1 port map( A => n15606, ZN => n9952);
   U11207 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1171_port, B2 => n2724, 
                           ZN => n15606);
   U11208 : INV_X1 port map( A => n15605, ZN => n9953);
   U11209 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1170_port, B2 => n2724, 
                           ZN => n15605);
   U11210 : INV_X1 port map( A => n15604, ZN => n9954);
   U11211 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1169_port, B2 => n2724, 
                           ZN => n15604);
   U11212 : INV_X1 port map( A => n15603, ZN => n9955);
   U11213 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1168_port, B2 => n2724, 
                           ZN => n15603);
   U11214 : INV_X1 port map( A => n15602, ZN => n9956);
   U11215 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1167_port, B2 => n2724, 
                           ZN => n15602);
   U11216 : INV_X1 port map( A => n15601, ZN => n9957);
   U11217 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1166_port, B2 => n2724, 
                           ZN => n15601);
   U11218 : INV_X1 port map( A => n15600, ZN => n9958);
   U11219 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1165_port, B2 => n2724, 
                           ZN => n15600);
   U11220 : INV_X1 port map( A => n15599, ZN => n9959);
   U11221 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1164_port, B2 => n2724, 
                           ZN => n15599);
   U11222 : INV_X1 port map( A => n15598, ZN => n9960);
   U11223 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1163_port, B2 => n2723, 
                           ZN => n15598);
   U11224 : INV_X1 port map( A => n15597, ZN => n9961);
   U11225 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1162_port, B2 => n2723, 
                           ZN => n15597);
   U11226 : INV_X1 port map( A => n15596, ZN => n9962);
   U11227 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1161_port, B2 => n2723, 
                           ZN => n15596);
   U11228 : INV_X1 port map( A => n15595, ZN => n9963);
   U11229 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2721, B1 => 
                           DataPath_RF_bus_reg_dataout_1160_port, B2 => n2723, 
                           ZN => n15595);
   U11230 : INV_X1 port map( A => n15594, ZN => n9964);
   U11231 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1159_port, B2 => n2723, 
                           ZN => n15594);
   U11232 : INV_X1 port map( A => n15593, ZN => n9965);
   U11233 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1158_port, B2 => n2723, 
                           ZN => n15593);
   U11234 : INV_X1 port map( A => n15592, ZN => n9966);
   U11235 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1157_port, B2 => n2723, 
                           ZN => n15592);
   U11236 : INV_X1 port map( A => n15591, ZN => n9967);
   U11237 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1156_port, B2 => n2723, 
                           ZN => n15591);
   U11238 : INV_X1 port map( A => n15590, ZN => n9968);
   U11239 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1155_port, B2 => n2723, 
                           ZN => n15590);
   U11240 : INV_X1 port map( A => n15589, ZN => n9969);
   U11241 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1154_port, B2 => n2723, 
                           ZN => n15589);
   U11242 : INV_X1 port map( A => n15588, ZN => n9970);
   U11243 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1153_port, B2 => n2723, 
                           ZN => n15588);
   U11244 : INV_X1 port map( A => n15585, ZN => n9971);
   U11245 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2722, B1 => 
                           DataPath_RF_bus_reg_dataout_1152_port, B2 => n2723, 
                           ZN => n15585);
   U11246 : INV_X1 port map( A => n15652, ZN => n9972);
   U11247 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1215_port, B2 => n2731, 
                           ZN => n15652);
   U11248 : INV_X1 port map( A => n15651, ZN => n9973);
   U11249 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1214_port, B2 => n2731, 
                           ZN => n15651);
   U11250 : INV_X1 port map( A => n15650, ZN => n9974);
   U11251 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1213_port, B2 => n2731, 
                           ZN => n15650);
   U11252 : INV_X1 port map( A => n15649, ZN => n9975);
   U11253 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1212_port, B2 => n2731, 
                           ZN => n15649);
   U11254 : INV_X1 port map( A => n15648, ZN => n9976);
   U11255 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1211_port, B2 => n2731, 
                           ZN => n15648);
   U11256 : INV_X1 port map( A => n15647, ZN => n9977);
   U11257 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1210_port, B2 => n2731, 
                           ZN => n15647);
   U11258 : INV_X1 port map( A => n15646, ZN => n9978);
   U11259 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1209_port, B2 => n2731, 
                           ZN => n15646);
   U11260 : INV_X1 port map( A => n15645, ZN => n9979);
   U11261 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1208_port, B2 => n2731, 
                           ZN => n15645);
   U11262 : INV_X1 port map( A => n15644, ZN => n9980);
   U11263 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1207_port, B2 => n2730, 
                           ZN => n15644);
   U11264 : INV_X1 port map( A => n15643, ZN => n9981);
   U11265 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1206_port, B2 => n2730, 
                           ZN => n15643);
   U11266 : INV_X1 port map( A => n15642, ZN => n9982);
   U11267 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1205_port, B2 => n2730, 
                           ZN => n15642);
   U11268 : INV_X1 port map( A => n15641, ZN => n9983);
   U11269 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2726, B1 => 
                           DataPath_RF_bus_reg_dataout_1204_port, B2 => n2730, 
                           ZN => n15641);
   U11270 : INV_X1 port map( A => n15640, ZN => n9984);
   U11271 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1203_port, B2 => n2730, 
                           ZN => n15640);
   U11272 : INV_X1 port map( A => n15639, ZN => n9985);
   U11273 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1202_port, B2 => n2730, 
                           ZN => n15639);
   U11274 : INV_X1 port map( A => n15638, ZN => n9986);
   U11275 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1201_port, B2 => n2730, 
                           ZN => n15638);
   U11276 : INV_X1 port map( A => n15637, ZN => n9987);
   U11277 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1200_port, B2 => n2730, 
                           ZN => n15637);
   U11278 : INV_X1 port map( A => n15636, ZN => n9988);
   U11279 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1199_port, B2 => n2730, 
                           ZN => n15636);
   U11280 : INV_X1 port map( A => n15635, ZN => n9989);
   U11281 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1198_port, B2 => n2730, 
                           ZN => n15635);
   U11282 : INV_X1 port map( A => n15634, ZN => n9990);
   U11283 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1197_port, B2 => n2730, 
                           ZN => n15634);
   U11284 : INV_X1 port map( A => n15633, ZN => n9991);
   U11285 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1196_port, B2 => n2730, 
                           ZN => n15633);
   U11286 : INV_X1 port map( A => n15632, ZN => n9992);
   U11287 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1195_port, B2 => n2729, 
                           ZN => n15632);
   U11288 : INV_X1 port map( A => n15631, ZN => n9993);
   U11289 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1194_port, B2 => n2729, 
                           ZN => n15631);
   U11290 : INV_X1 port map( A => n15630, ZN => n9994);
   U11291 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1193_port, B2 => n2729, 
                           ZN => n15630);
   U11292 : INV_X1 port map( A => n15629, ZN => n9995);
   U11293 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2727, B1 => 
                           DataPath_RF_bus_reg_dataout_1192_port, B2 => n2729, 
                           ZN => n15629);
   U11294 : INV_X1 port map( A => n15628, ZN => n9996);
   U11295 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1191_port, B2 => n2729, 
                           ZN => n15628);
   U11296 : INV_X1 port map( A => n15627, ZN => n9997);
   U11297 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1190_port, B2 => n2729, 
                           ZN => n15627);
   U11298 : INV_X1 port map( A => n15626, ZN => n9998);
   U11299 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1189_port, B2 => n2729, 
                           ZN => n15626);
   U11300 : INV_X1 port map( A => n15625, ZN => n9999);
   U11301 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1188_port, B2 => n2729, 
                           ZN => n15625);
   U11302 : INV_X1 port map( A => n15624, ZN => n10000);
   U11303 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1187_port, B2 => n2729, 
                           ZN => n15624);
   U11304 : INV_X1 port map( A => n15623, ZN => n10001);
   U11305 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1186_port, B2 => n2729, 
                           ZN => n15623);
   U11306 : INV_X1 port map( A => n15622, ZN => n10002);
   U11307 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1185_port, B2 => n2729, 
                           ZN => n15622);
   U11308 : INV_X1 port map( A => n15619, ZN => n10003);
   U11309 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2728, B1 => 
                           DataPath_RF_bus_reg_dataout_1184_port, B2 => n2729, 
                           ZN => n15619);
   U11310 : INV_X1 port map( A => n15686, ZN => n10004);
   U11311 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1247_port, B2 => n2737, 
                           ZN => n15686);
   U11312 : INV_X1 port map( A => n15685, ZN => n10005);
   U11313 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1246_port, B2 => n2737, 
                           ZN => n15685);
   U11314 : INV_X1 port map( A => n15684, ZN => n10006);
   U11315 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1245_port, B2 => n2737, 
                           ZN => n15684);
   U11316 : INV_X1 port map( A => n15683, ZN => n10007);
   U11317 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1244_port, B2 => n2737, 
                           ZN => n15683);
   U11318 : INV_X1 port map( A => n15682, ZN => n10008);
   U11319 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1243_port, B2 => n2737, 
                           ZN => n15682);
   U11320 : INV_X1 port map( A => n15681, ZN => n10009);
   U11321 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1242_port, B2 => n2737, 
                           ZN => n15681);
   U11322 : INV_X1 port map( A => n15680, ZN => n10010);
   U11323 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1241_port, B2 => n2737, 
                           ZN => n15680);
   U11324 : INV_X1 port map( A => n15679, ZN => n10011);
   U11325 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1240_port, B2 => n2737, 
                           ZN => n15679);
   U11326 : INV_X1 port map( A => n15678, ZN => n10012);
   U11327 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1239_port, B2 => n2736, 
                           ZN => n15678);
   U11328 : INV_X1 port map( A => n15677, ZN => n10013);
   U11329 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1238_port, B2 => n2736, 
                           ZN => n15677);
   U11330 : INV_X1 port map( A => n15676, ZN => n10014);
   U11331 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1237_port, B2 => n2736, 
                           ZN => n15676);
   U11332 : INV_X1 port map( A => n15675, ZN => n10015);
   U11333 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2732, B1 => 
                           DataPath_RF_bus_reg_dataout_1236_port, B2 => n2736, 
                           ZN => n15675);
   U11334 : INV_X1 port map( A => n15674, ZN => n10016);
   U11335 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1235_port, B2 => n2736, 
                           ZN => n15674);
   U11336 : INV_X1 port map( A => n15673, ZN => n10017);
   U11337 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1234_port, B2 => n2736, 
                           ZN => n15673);
   U11338 : INV_X1 port map( A => n15672, ZN => n10018);
   U11339 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1233_port, B2 => n2736, 
                           ZN => n15672);
   U11340 : INV_X1 port map( A => n15671, ZN => n10019);
   U11341 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1232_port, B2 => n2736, 
                           ZN => n15671);
   U11342 : INV_X1 port map( A => n15670, ZN => n10020);
   U11343 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1231_port, B2 => n2736, 
                           ZN => n15670);
   U11344 : INV_X1 port map( A => n15669, ZN => n10021);
   U11345 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1230_port, B2 => n2736, 
                           ZN => n15669);
   U11346 : INV_X1 port map( A => n15668, ZN => n10022);
   U11347 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1229_port, B2 => n2736, 
                           ZN => n15668);
   U11348 : INV_X1 port map( A => n15667, ZN => n10023);
   U11349 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1228_port, B2 => n2736, 
                           ZN => n15667);
   U11350 : INV_X1 port map( A => n15666, ZN => n10024);
   U11351 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1227_port, B2 => n2735, 
                           ZN => n15666);
   U11352 : INV_X1 port map( A => n15665, ZN => n10025);
   U11353 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1226_port, B2 => n2735, 
                           ZN => n15665);
   U11354 : INV_X1 port map( A => n15664, ZN => n10026);
   U11355 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1225_port, B2 => n2735, 
                           ZN => n15664);
   U11356 : INV_X1 port map( A => n15663, ZN => n10027);
   U11357 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2733, B1 => 
                           DataPath_RF_bus_reg_dataout_1224_port, B2 => n2735, 
                           ZN => n15663);
   U11358 : INV_X1 port map( A => n15662, ZN => n10028);
   U11359 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1223_port, B2 => n2735, 
                           ZN => n15662);
   U11360 : INV_X1 port map( A => n15661, ZN => n10029);
   U11361 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1222_port, B2 => n2735, 
                           ZN => n15661);
   U11362 : INV_X1 port map( A => n15660, ZN => n10030);
   U11363 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1221_port, B2 => n2735, 
                           ZN => n15660);
   U11364 : INV_X1 port map( A => n15659, ZN => n10031);
   U11365 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1220_port, B2 => n2735, 
                           ZN => n15659);
   U11366 : INV_X1 port map( A => n15658, ZN => n10032);
   U11367 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1219_port, B2 => n2735, 
                           ZN => n15658);
   U11368 : INV_X1 port map( A => n15657, ZN => n10033);
   U11369 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1218_port, B2 => n2735, 
                           ZN => n15657);
   U11370 : INV_X1 port map( A => n15656, ZN => n10034);
   U11371 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1217_port, B2 => n2735, 
                           ZN => n15656);
   U11372 : INV_X1 port map( A => n15653, ZN => n10035);
   U11373 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2734, B1 => 
                           DataPath_RF_bus_reg_dataout_1216_port, B2 => n2735, 
                           ZN => n15653);
   U11374 : INV_X1 port map( A => n15720, ZN => n10036);
   U11375 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1279_port, B2 => n2743, 
                           ZN => n15720);
   U11376 : INV_X1 port map( A => n15719, ZN => n10037);
   U11377 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1278_port, B2 => n2743, 
                           ZN => n15719);
   U11378 : INV_X1 port map( A => n15718, ZN => n10038);
   U11379 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1277_port, B2 => n2743, 
                           ZN => n15718);
   U11380 : INV_X1 port map( A => n15717, ZN => n10039);
   U11381 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1276_port, B2 => n2743, 
                           ZN => n15717);
   U11382 : INV_X1 port map( A => n15716, ZN => n10040);
   U11383 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1275_port, B2 => n2743, 
                           ZN => n15716);
   U11384 : INV_X1 port map( A => n15715, ZN => n10041);
   U11385 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1274_port, B2 => n2743, 
                           ZN => n15715);
   U11386 : INV_X1 port map( A => n15714, ZN => n10042);
   U11387 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1273_port, B2 => n2743, 
                           ZN => n15714);
   U11388 : INV_X1 port map( A => n15713, ZN => n10043);
   U11389 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1272_port, B2 => n2743, 
                           ZN => n15713);
   U11390 : INV_X1 port map( A => n15712, ZN => n10044);
   U11391 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1271_port, B2 => n2742, 
                           ZN => n15712);
   U11392 : INV_X1 port map( A => n15711, ZN => n10045);
   U11393 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1270_port, B2 => n2742, 
                           ZN => n15711);
   U11394 : INV_X1 port map( A => n15710, ZN => n10046);
   U11395 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1269_port, B2 => n2742, 
                           ZN => n15710);
   U11396 : INV_X1 port map( A => n15709, ZN => n10047);
   U11397 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2738, B1 => 
                           DataPath_RF_bus_reg_dataout_1268_port, B2 => n2742, 
                           ZN => n15709);
   U11398 : INV_X1 port map( A => n15708, ZN => n10048);
   U11399 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1267_port, B2 => n2742, 
                           ZN => n15708);
   U11400 : INV_X1 port map( A => n15707, ZN => n10049);
   U11401 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1266_port, B2 => n2742, 
                           ZN => n15707);
   U11402 : INV_X1 port map( A => n15706, ZN => n10050);
   U11403 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1265_port, B2 => n2742, 
                           ZN => n15706);
   U11404 : INV_X1 port map( A => n15705, ZN => n10051);
   U11405 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1264_port, B2 => n2742, 
                           ZN => n15705);
   U11406 : INV_X1 port map( A => n15704, ZN => n10052);
   U11407 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1263_port, B2 => n2742, 
                           ZN => n15704);
   U11408 : INV_X1 port map( A => n15703, ZN => n10053);
   U11409 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1262_port, B2 => n2742, 
                           ZN => n15703);
   U11410 : INV_X1 port map( A => n15702, ZN => n10054);
   U11411 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1261_port, B2 => n2742, 
                           ZN => n15702);
   U11412 : INV_X1 port map( A => n15701, ZN => n10055);
   U11413 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1260_port, B2 => n2742, 
                           ZN => n15701);
   U11414 : INV_X1 port map( A => n15700, ZN => n10056);
   U11415 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1259_port, B2 => n2741, 
                           ZN => n15700);
   U11416 : INV_X1 port map( A => n15699, ZN => n10057);
   U11417 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1258_port, B2 => n2741, 
                           ZN => n15699);
   U11418 : INV_X1 port map( A => n15698, ZN => n10058);
   U11419 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1257_port, B2 => n2741, 
                           ZN => n15698);
   U11420 : INV_X1 port map( A => n15697, ZN => n10059);
   U11421 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2739, B1 => 
                           DataPath_RF_bus_reg_dataout_1256_port, B2 => n2741, 
                           ZN => n15697);
   U11422 : INV_X1 port map( A => n15696, ZN => n10060);
   U11423 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1255_port, B2 => n2741, 
                           ZN => n15696);
   U11424 : INV_X1 port map( A => n15695, ZN => n10061);
   U11425 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1254_port, B2 => n2741, 
                           ZN => n15695);
   U11426 : INV_X1 port map( A => n15694, ZN => n10062);
   U11427 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1253_port, B2 => n2741, 
                           ZN => n15694);
   U11428 : INV_X1 port map( A => n15693, ZN => n10063);
   U11429 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1252_port, B2 => n2741, 
                           ZN => n15693);
   U11430 : INV_X1 port map( A => n15692, ZN => n10064);
   U11431 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1251_port, B2 => n2741, 
                           ZN => n15692);
   U11432 : INV_X1 port map( A => n15691, ZN => n10065);
   U11433 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1250_port, B2 => n2741, 
                           ZN => n15691);
   U11434 : INV_X1 port map( A => n15690, ZN => n10066);
   U11435 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1249_port, B2 => n2741, 
                           ZN => n15690);
   U11436 : INV_X1 port map( A => n15687, ZN => n10067);
   U11437 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2740, B1 => 
                           DataPath_RF_bus_reg_dataout_1248_port, B2 => n2741, 
                           ZN => n15687);
   U11438 : INV_X1 port map( A => n15754, ZN => n10068);
   U11439 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1311_port, B2 => n2749, 
                           ZN => n15754);
   U11440 : INV_X1 port map( A => n15753, ZN => n10069);
   U11441 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1310_port, B2 => n2749, 
                           ZN => n15753);
   U11442 : INV_X1 port map( A => n15752, ZN => n10070);
   U11443 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1309_port, B2 => n2749, 
                           ZN => n15752);
   U11444 : INV_X1 port map( A => n15751, ZN => n10071);
   U11445 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1308_port, B2 => n2749, 
                           ZN => n15751);
   U11446 : INV_X1 port map( A => n15750, ZN => n10072);
   U11447 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1307_port, B2 => n2749, 
                           ZN => n15750);
   U11448 : INV_X1 port map( A => n15749, ZN => n10073);
   U11449 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1306_port, B2 => n2749, 
                           ZN => n15749);
   U11450 : INV_X1 port map( A => n15748, ZN => n10074);
   U11451 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1305_port, B2 => n2749, 
                           ZN => n15748);
   U11452 : INV_X1 port map( A => n15747, ZN => n10075);
   U11453 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1304_port, B2 => n2749, 
                           ZN => n15747);
   U11454 : INV_X1 port map( A => n15746, ZN => n10076);
   U11455 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1303_port, B2 => n2748, 
                           ZN => n15746);
   U11456 : INV_X1 port map( A => n15745, ZN => n10077);
   U11457 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1302_port, B2 => n2748, 
                           ZN => n15745);
   U11458 : INV_X1 port map( A => n15744, ZN => n10078);
   U11459 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1301_port, B2 => n2748, 
                           ZN => n15744);
   U11460 : INV_X1 port map( A => n15743, ZN => n10079);
   U11461 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2744, B1 => 
                           DataPath_RF_bus_reg_dataout_1300_port, B2 => n2748, 
                           ZN => n15743);
   U11462 : INV_X1 port map( A => n15742, ZN => n10080);
   U11463 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1299_port, B2 => n2748, 
                           ZN => n15742);
   U11464 : INV_X1 port map( A => n15741, ZN => n10081);
   U11465 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1298_port, B2 => n2748, 
                           ZN => n15741);
   U11466 : INV_X1 port map( A => n15740, ZN => n10082);
   U11467 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1297_port, B2 => n2748, 
                           ZN => n15740);
   U11468 : INV_X1 port map( A => n15739, ZN => n10083);
   U11469 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1296_port, B2 => n2748, 
                           ZN => n15739);
   U11470 : INV_X1 port map( A => n15738, ZN => n10084);
   U11471 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1295_port, B2 => n2748, 
                           ZN => n15738);
   U11472 : INV_X1 port map( A => n15737, ZN => n10085);
   U11473 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1294_port, B2 => n2748, 
                           ZN => n15737);
   U11474 : INV_X1 port map( A => n15736, ZN => n10086);
   U11475 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1293_port, B2 => n2748, 
                           ZN => n15736);
   U11476 : INV_X1 port map( A => n15735, ZN => n10087);
   U11477 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1292_port, B2 => n2748, 
                           ZN => n15735);
   U11478 : INV_X1 port map( A => n15734, ZN => n10088);
   U11479 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1291_port, B2 => n2747, 
                           ZN => n15734);
   U11480 : INV_X1 port map( A => n15733, ZN => n10089);
   U11481 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1290_port, B2 => n2747, 
                           ZN => n15733);
   U11482 : INV_X1 port map( A => n15732, ZN => n10090);
   U11483 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1289_port, B2 => n2747, 
                           ZN => n15732);
   U11484 : INV_X1 port map( A => n15731, ZN => n10091);
   U11485 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2745, B1 => 
                           DataPath_RF_bus_reg_dataout_1288_port, B2 => n2747, 
                           ZN => n15731);
   U11486 : INV_X1 port map( A => n15730, ZN => n10092);
   U11487 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1287_port, B2 => n2747, 
                           ZN => n15730);
   U11488 : INV_X1 port map( A => n15729, ZN => n10093);
   U11489 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1286_port, B2 => n2747, 
                           ZN => n15729);
   U11490 : INV_X1 port map( A => n15728, ZN => n10094);
   U11491 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1285_port, B2 => n2747, 
                           ZN => n15728);
   U11492 : INV_X1 port map( A => n15727, ZN => n10095);
   U11493 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1284_port, B2 => n2747, 
                           ZN => n15727);
   U11494 : INV_X1 port map( A => n15726, ZN => n10096);
   U11495 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1283_port, B2 => n2747, 
                           ZN => n15726);
   U11496 : INV_X1 port map( A => n15725, ZN => n10097);
   U11497 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1282_port, B2 => n2747, 
                           ZN => n15725);
   U11498 : INV_X1 port map( A => n15724, ZN => n10098);
   U11499 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1281_port, B2 => n2747, 
                           ZN => n15724);
   U11500 : INV_X1 port map( A => n15721, ZN => n10099);
   U11501 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2746, B1 => 
                           DataPath_RF_bus_reg_dataout_1280_port, B2 => n2747, 
                           ZN => n15721);
   U11502 : INV_X1 port map( A => n15788, ZN => n10100);
   U11503 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1343_port, B2 => n2755, 
                           ZN => n15788);
   U11504 : INV_X1 port map( A => n15787, ZN => n10101);
   U11505 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1342_port, B2 => n2755, 
                           ZN => n15787);
   U11506 : INV_X1 port map( A => n15786, ZN => n10102);
   U11507 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1341_port, B2 => n2755, 
                           ZN => n15786);
   U11508 : INV_X1 port map( A => n15785, ZN => n10103);
   U11509 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1340_port, B2 => n2755, 
                           ZN => n15785);
   U11510 : INV_X1 port map( A => n15784, ZN => n10104);
   U11511 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1339_port, B2 => n2755, 
                           ZN => n15784);
   U11512 : INV_X1 port map( A => n15783, ZN => n10105);
   U11513 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1338_port, B2 => n2755, 
                           ZN => n15783);
   U11514 : INV_X1 port map( A => n15782, ZN => n10106);
   U11515 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1337_port, B2 => n2755, 
                           ZN => n15782);
   U11516 : INV_X1 port map( A => n15781, ZN => n10107);
   U11517 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1336_port, B2 => n2755, 
                           ZN => n15781);
   U11518 : INV_X1 port map( A => n15780, ZN => n10108);
   U11519 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1335_port, B2 => n2754, 
                           ZN => n15780);
   U11520 : INV_X1 port map( A => n15779, ZN => n10109);
   U11521 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1334_port, B2 => n2754, 
                           ZN => n15779);
   U11522 : INV_X1 port map( A => n15778, ZN => n10110);
   U11523 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1333_port, B2 => n2754, 
                           ZN => n15778);
   U11524 : INV_X1 port map( A => n15777, ZN => n10111);
   U11525 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2750, B1 => 
                           DataPath_RF_bus_reg_dataout_1332_port, B2 => n2754, 
                           ZN => n15777);
   U11526 : INV_X1 port map( A => n15776, ZN => n10112);
   U11527 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1331_port, B2 => n2754, 
                           ZN => n15776);
   U11528 : INV_X1 port map( A => n15775, ZN => n10113);
   U11529 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1330_port, B2 => n2754, 
                           ZN => n15775);
   U11530 : INV_X1 port map( A => n15774, ZN => n10114);
   U11531 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1329_port, B2 => n2754, 
                           ZN => n15774);
   U11532 : INV_X1 port map( A => n15773, ZN => n10115);
   U11533 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1328_port, B2 => n2754, 
                           ZN => n15773);
   U11534 : INV_X1 port map( A => n15772, ZN => n10116);
   U11535 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1327_port, B2 => n2754, 
                           ZN => n15772);
   U11536 : INV_X1 port map( A => n15771, ZN => n10117);
   U11537 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1326_port, B2 => n2754, 
                           ZN => n15771);
   U11538 : INV_X1 port map( A => n15770, ZN => n10118);
   U11539 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1325_port, B2 => n2754, 
                           ZN => n15770);
   U11540 : INV_X1 port map( A => n15769, ZN => n10119);
   U11541 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1324_port, B2 => n2754, 
                           ZN => n15769);
   U11542 : INV_X1 port map( A => n15768, ZN => n10120);
   U11543 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1323_port, B2 => n2753, 
                           ZN => n15768);
   U11544 : INV_X1 port map( A => n15767, ZN => n10121);
   U11545 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1322_port, B2 => n2753, 
                           ZN => n15767);
   U11546 : INV_X1 port map( A => n15766, ZN => n10122);
   U11547 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1321_port, B2 => n2753, 
                           ZN => n15766);
   U11548 : INV_X1 port map( A => n15765, ZN => n10123);
   U11549 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2751, B1 => 
                           DataPath_RF_bus_reg_dataout_1320_port, B2 => n2753, 
                           ZN => n15765);
   U11550 : INV_X1 port map( A => n15764, ZN => n10124);
   U11551 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1319_port, B2 => n2753, 
                           ZN => n15764);
   U11552 : INV_X1 port map( A => n15763, ZN => n10125);
   U11553 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1318_port, B2 => n2753, 
                           ZN => n15763);
   U11554 : INV_X1 port map( A => n15762, ZN => n10126);
   U11555 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1317_port, B2 => n2753, 
                           ZN => n15762);
   U11556 : INV_X1 port map( A => n15761, ZN => n10127);
   U11557 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1316_port, B2 => n2753, 
                           ZN => n15761);
   U11558 : INV_X1 port map( A => n15760, ZN => n10128);
   U11559 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1315_port, B2 => n2753, 
                           ZN => n15760);
   U11560 : INV_X1 port map( A => n15759, ZN => n10129);
   U11561 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1314_port, B2 => n2753, 
                           ZN => n15759);
   U11562 : INV_X1 port map( A => n15758, ZN => n10130);
   U11563 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1313_port, B2 => n2753, 
                           ZN => n15758);
   U11564 : INV_X1 port map( A => n15755, ZN => n10131);
   U11565 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2752, B1 => 
                           DataPath_RF_bus_reg_dataout_1312_port, B2 => n2753, 
                           ZN => n15755);
   U11566 : INV_X1 port map( A => n15822, ZN => n10132);
   U11567 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1375_port, B2 => n2761, 
                           ZN => n15822);
   U11568 : INV_X1 port map( A => n15821, ZN => n10133);
   U11569 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1374_port, B2 => n2761, 
                           ZN => n15821);
   U11570 : INV_X1 port map( A => n15820, ZN => n10134);
   U11571 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1373_port, B2 => n2761, 
                           ZN => n15820);
   U11572 : INV_X1 port map( A => n15819, ZN => n10135);
   U11573 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1372_port, B2 => n2761, 
                           ZN => n15819);
   U11574 : INV_X1 port map( A => n15818, ZN => n10136);
   U11575 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1371_port, B2 => n2761, 
                           ZN => n15818);
   U11576 : INV_X1 port map( A => n15817, ZN => n10137);
   U11577 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1370_port, B2 => n2761, 
                           ZN => n15817);
   U11578 : INV_X1 port map( A => n15816, ZN => n10138);
   U11579 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1369_port, B2 => n2761, 
                           ZN => n15816);
   U11580 : INV_X1 port map( A => n15815, ZN => n10139);
   U11581 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1368_port, B2 => n2761, 
                           ZN => n15815);
   U11582 : INV_X1 port map( A => n15814, ZN => n10140);
   U11583 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1367_port, B2 => n2760, 
                           ZN => n15814);
   U11584 : INV_X1 port map( A => n15813, ZN => n10141);
   U11585 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1366_port, B2 => n2760, 
                           ZN => n15813);
   U11586 : INV_X1 port map( A => n15812, ZN => n10142);
   U11587 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1365_port, B2 => n2760, 
                           ZN => n15812);
   U11588 : INV_X1 port map( A => n15811, ZN => n10143);
   U11589 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2756, B1 => 
                           DataPath_RF_bus_reg_dataout_1364_port, B2 => n2760, 
                           ZN => n15811);
   U11590 : INV_X1 port map( A => n15810, ZN => n10144);
   U11591 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1363_port, B2 => n2760, 
                           ZN => n15810);
   U11592 : INV_X1 port map( A => n15809, ZN => n10145);
   U11593 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1362_port, B2 => n2760, 
                           ZN => n15809);
   U11594 : INV_X1 port map( A => n15808, ZN => n10146);
   U11595 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1361_port, B2 => n2760, 
                           ZN => n15808);
   U11596 : INV_X1 port map( A => n15807, ZN => n10147);
   U11597 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1360_port, B2 => n2760, 
                           ZN => n15807);
   U11598 : INV_X1 port map( A => n15806, ZN => n10148);
   U11599 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1359_port, B2 => n2760, 
                           ZN => n15806);
   U11600 : INV_X1 port map( A => n15805, ZN => n10149);
   U11601 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1358_port, B2 => n2760, 
                           ZN => n15805);
   U11602 : INV_X1 port map( A => n15804, ZN => n10150);
   U11603 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1357_port, B2 => n2760, 
                           ZN => n15804);
   U11604 : INV_X1 port map( A => n15803, ZN => n10151);
   U11605 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1356_port, B2 => n2760, 
                           ZN => n15803);
   U11606 : INV_X1 port map( A => n15802, ZN => n10152);
   U11607 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1355_port, B2 => n2759, 
                           ZN => n15802);
   U11608 : INV_X1 port map( A => n15801, ZN => n10153);
   U11609 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1354_port, B2 => n2759, 
                           ZN => n15801);
   U11610 : INV_X1 port map( A => n15800, ZN => n10154);
   U11611 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1353_port, B2 => n2759, 
                           ZN => n15800);
   U11612 : INV_X1 port map( A => n15799, ZN => n10155);
   U11613 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2757, B1 => 
                           DataPath_RF_bus_reg_dataout_1352_port, B2 => n2759, 
                           ZN => n15799);
   U11614 : INV_X1 port map( A => n15798, ZN => n10156);
   U11615 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1351_port, B2 => n2759, 
                           ZN => n15798);
   U11616 : INV_X1 port map( A => n15797, ZN => n10157);
   U11617 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1350_port, B2 => n2759, 
                           ZN => n15797);
   U11618 : INV_X1 port map( A => n15796, ZN => n10158);
   U11619 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1349_port, B2 => n2759, 
                           ZN => n15796);
   U11620 : INV_X1 port map( A => n15795, ZN => n10159);
   U11621 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1348_port, B2 => n2759, 
                           ZN => n15795);
   U11622 : INV_X1 port map( A => n15794, ZN => n10160);
   U11623 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1347_port, B2 => n2759, 
                           ZN => n15794);
   U11624 : INV_X1 port map( A => n15793, ZN => n10161);
   U11625 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1346_port, B2 => n2759, 
                           ZN => n15793);
   U11626 : INV_X1 port map( A => n15792, ZN => n10162);
   U11627 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1345_port, B2 => n2759, 
                           ZN => n15792);
   U11628 : INV_X1 port map( A => n15789, ZN => n10163);
   U11629 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2758, B1 => 
                           DataPath_RF_bus_reg_dataout_1344_port, B2 => n2759, 
                           ZN => n15789);
   U11630 : INV_X1 port map( A => n15856, ZN => n10164);
   U11631 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1407_port, B2 => n2767, 
                           ZN => n15856);
   U11632 : INV_X1 port map( A => n15855, ZN => n10165);
   U11633 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1406_port, B2 => n2767, 
                           ZN => n15855);
   U11634 : INV_X1 port map( A => n15854, ZN => n10166);
   U11635 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1405_port, B2 => n2767, 
                           ZN => n15854);
   U11636 : INV_X1 port map( A => n15853, ZN => n10167);
   U11637 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1404_port, B2 => n2767, 
                           ZN => n15853);
   U11638 : INV_X1 port map( A => n15852, ZN => n10168);
   U11639 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1403_port, B2 => n2767, 
                           ZN => n15852);
   U11640 : INV_X1 port map( A => n15851, ZN => n10169);
   U11641 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1402_port, B2 => n2767, 
                           ZN => n15851);
   U11642 : INV_X1 port map( A => n15850, ZN => n10170);
   U11643 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1401_port, B2 => n2767, 
                           ZN => n15850);
   U11644 : INV_X1 port map( A => n15849, ZN => n10171);
   U11645 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1400_port, B2 => n2767, 
                           ZN => n15849);
   U11646 : INV_X1 port map( A => n15848, ZN => n10172);
   U11647 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1399_port, B2 => n2766, 
                           ZN => n15848);
   U11648 : INV_X1 port map( A => n15847, ZN => n10173);
   U11649 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1398_port, B2 => n2766, 
                           ZN => n15847);
   U11650 : INV_X1 port map( A => n15846, ZN => n10174);
   U11651 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1397_port, B2 => n2766, 
                           ZN => n15846);
   U11652 : INV_X1 port map( A => n15845, ZN => n10175);
   U11653 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2762, B1 => 
                           DataPath_RF_bus_reg_dataout_1396_port, B2 => n2766, 
                           ZN => n15845);
   U11654 : INV_X1 port map( A => n15844, ZN => n10176);
   U11655 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1395_port, B2 => n2766, 
                           ZN => n15844);
   U11656 : INV_X1 port map( A => n15843, ZN => n10177);
   U11657 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1394_port, B2 => n2766, 
                           ZN => n15843);
   U11658 : INV_X1 port map( A => n15842, ZN => n10178);
   U11659 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1393_port, B2 => n2766, 
                           ZN => n15842);
   U11660 : INV_X1 port map( A => n15841, ZN => n10179);
   U11661 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1392_port, B2 => n2766, 
                           ZN => n15841);
   U11662 : INV_X1 port map( A => n15840, ZN => n10180);
   U11663 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1391_port, B2 => n2766, 
                           ZN => n15840);
   U11664 : INV_X1 port map( A => n15839, ZN => n10181);
   U11665 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1390_port, B2 => n2766, 
                           ZN => n15839);
   U11666 : INV_X1 port map( A => n15838, ZN => n10182);
   U11667 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1389_port, B2 => n2766, 
                           ZN => n15838);
   U11668 : INV_X1 port map( A => n15837, ZN => n10183);
   U11669 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1388_port, B2 => n2766, 
                           ZN => n15837);
   U11670 : INV_X1 port map( A => n15836, ZN => n10184);
   U11671 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1387_port, B2 => n2765, 
                           ZN => n15836);
   U11672 : INV_X1 port map( A => n15835, ZN => n10185);
   U11673 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1386_port, B2 => n2765, 
                           ZN => n15835);
   U11674 : INV_X1 port map( A => n15834, ZN => n10186);
   U11675 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1385_port, B2 => n2765, 
                           ZN => n15834);
   U11676 : INV_X1 port map( A => n15833, ZN => n10187);
   U11677 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2763, B1 => 
                           DataPath_RF_bus_reg_dataout_1384_port, B2 => n2765, 
                           ZN => n15833);
   U11678 : INV_X1 port map( A => n15832, ZN => n10188);
   U11679 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1383_port, B2 => n2765, 
                           ZN => n15832);
   U11680 : INV_X1 port map( A => n15831, ZN => n10189);
   U11681 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1382_port, B2 => n2765, 
                           ZN => n15831);
   U11682 : INV_X1 port map( A => n15830, ZN => n10190);
   U11683 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1381_port, B2 => n2765, 
                           ZN => n15830);
   U11684 : INV_X1 port map( A => n15829, ZN => n10191);
   U11685 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1380_port, B2 => n2765, 
                           ZN => n15829);
   U11686 : INV_X1 port map( A => n15828, ZN => n10192);
   U11687 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1379_port, B2 => n2765, 
                           ZN => n15828);
   U11688 : INV_X1 port map( A => n15827, ZN => n10193);
   U11689 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1378_port, B2 => n2765, 
                           ZN => n15827);
   U11690 : INV_X1 port map( A => n15826, ZN => n10194);
   U11691 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1377_port, B2 => n2765, 
                           ZN => n15826);
   U11692 : INV_X1 port map( A => n15823, ZN => n10195);
   U11693 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2764, B1 => 
                           DataPath_RF_bus_reg_dataout_1376_port, B2 => n2765, 
                           ZN => n15823);
   U11694 : INV_X1 port map( A => n15890, ZN => n10196);
   U11695 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1439_port, B2 => n2773, 
                           ZN => n15890);
   U11696 : INV_X1 port map( A => n15889, ZN => n10197);
   U11697 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1438_port, B2 => n2773, 
                           ZN => n15889);
   U11698 : INV_X1 port map( A => n15888, ZN => n10198);
   U11699 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1437_port, B2 => n2773, 
                           ZN => n15888);
   U11700 : INV_X1 port map( A => n15887, ZN => n10199);
   U11701 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1436_port, B2 => n2773, 
                           ZN => n15887);
   U11702 : INV_X1 port map( A => n15886, ZN => n10200);
   U11703 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1435_port, B2 => n2773, 
                           ZN => n15886);
   U11704 : INV_X1 port map( A => n15885, ZN => n10201);
   U11705 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1434_port, B2 => n2773, 
                           ZN => n15885);
   U11706 : INV_X1 port map( A => n15884, ZN => n10202);
   U11707 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1433_port, B2 => n2773, 
                           ZN => n15884);
   U11708 : INV_X1 port map( A => n15883, ZN => n10203);
   U11709 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1432_port, B2 => n2773, 
                           ZN => n15883);
   U11710 : INV_X1 port map( A => n15882, ZN => n10204);
   U11711 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1431_port, B2 => n2772, 
                           ZN => n15882);
   U11712 : INV_X1 port map( A => n15881, ZN => n10205);
   U11713 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1430_port, B2 => n2772, 
                           ZN => n15881);
   U11714 : INV_X1 port map( A => n15880, ZN => n10206);
   U11715 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1429_port, B2 => n2772, 
                           ZN => n15880);
   U11716 : INV_X1 port map( A => n15879, ZN => n10207);
   U11717 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2768, B1 => 
                           DataPath_RF_bus_reg_dataout_1428_port, B2 => n2772, 
                           ZN => n15879);
   U11718 : INV_X1 port map( A => n15878, ZN => n10208);
   U11719 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1427_port, B2 => n2772, 
                           ZN => n15878);
   U11720 : INV_X1 port map( A => n15877, ZN => n10209);
   U11721 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1426_port, B2 => n2772, 
                           ZN => n15877);
   U11722 : INV_X1 port map( A => n15876, ZN => n10210);
   U11723 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1425_port, B2 => n2772, 
                           ZN => n15876);
   U11724 : INV_X1 port map( A => n15875, ZN => n10211);
   U11725 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1424_port, B2 => n2772, 
                           ZN => n15875);
   U11726 : INV_X1 port map( A => n15874, ZN => n10212);
   U11727 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1423_port, B2 => n2772, 
                           ZN => n15874);
   U11728 : INV_X1 port map( A => n15873, ZN => n10213);
   U11729 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1422_port, B2 => n2772, 
                           ZN => n15873);
   U11730 : INV_X1 port map( A => n15872, ZN => n10214);
   U11731 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1421_port, B2 => n2772, 
                           ZN => n15872);
   U11732 : INV_X1 port map( A => n15871, ZN => n10215);
   U11733 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1420_port, B2 => n2772, 
                           ZN => n15871);
   U11734 : INV_X1 port map( A => n15870, ZN => n10216);
   U11735 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1419_port, B2 => n2771, 
                           ZN => n15870);
   U11736 : INV_X1 port map( A => n15869, ZN => n10217);
   U11737 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1418_port, B2 => n2771, 
                           ZN => n15869);
   U11738 : INV_X1 port map( A => n15868, ZN => n10218);
   U11739 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1417_port, B2 => n2771, 
                           ZN => n15868);
   U11740 : INV_X1 port map( A => n15867, ZN => n10219);
   U11741 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2769, B1 => 
                           DataPath_RF_bus_reg_dataout_1416_port, B2 => n2771, 
                           ZN => n15867);
   U11742 : INV_X1 port map( A => n15866, ZN => n10220);
   U11743 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1415_port, B2 => n2771, 
                           ZN => n15866);
   U11744 : INV_X1 port map( A => n15865, ZN => n10221);
   U11745 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1414_port, B2 => n2771, 
                           ZN => n15865);
   U11746 : INV_X1 port map( A => n15864, ZN => n10222);
   U11747 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1413_port, B2 => n2771, 
                           ZN => n15864);
   U11748 : INV_X1 port map( A => n15863, ZN => n10223);
   U11749 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1412_port, B2 => n2771, 
                           ZN => n15863);
   U11750 : INV_X1 port map( A => n15862, ZN => n10224);
   U11751 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1411_port, B2 => n2771, 
                           ZN => n15862);
   U11752 : INV_X1 port map( A => n15861, ZN => n10225);
   U11753 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1410_port, B2 => n2771, 
                           ZN => n15861);
   U11754 : INV_X1 port map( A => n15860, ZN => n10226);
   U11755 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1409_port, B2 => n2771, 
                           ZN => n15860);
   U11756 : INV_X1 port map( A => n15857, ZN => n10227);
   U11757 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2770, B1 => 
                           DataPath_RF_bus_reg_dataout_1408_port, B2 => n2771, 
                           ZN => n15857);
   U11758 : INV_X1 port map( A => n15924, ZN => n10228);
   U11759 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1471_port, B2 => n2779, 
                           ZN => n15924);
   U11760 : INV_X1 port map( A => n15923, ZN => n10229);
   U11761 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1470_port, B2 => n2779, 
                           ZN => n15923);
   U11762 : INV_X1 port map( A => n15922, ZN => n10230);
   U11763 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1469_port, B2 => n2779, 
                           ZN => n15922);
   U11764 : INV_X1 port map( A => n15921, ZN => n10231);
   U11765 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1468_port, B2 => n2779, 
                           ZN => n15921);
   U11766 : INV_X1 port map( A => n15920, ZN => n10232);
   U11767 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1467_port, B2 => n2779, 
                           ZN => n15920);
   U11768 : INV_X1 port map( A => n15919, ZN => n10233);
   U11769 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1466_port, B2 => n2779, 
                           ZN => n15919);
   U11770 : INV_X1 port map( A => n15918, ZN => n10234);
   U11771 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1465_port, B2 => n2779, 
                           ZN => n15918);
   U11772 : INV_X1 port map( A => n15917, ZN => n10235);
   U11773 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1464_port, B2 => n2779, 
                           ZN => n15917);
   U11774 : INV_X1 port map( A => n15916, ZN => n10236);
   U11775 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1463_port, B2 => n2778, 
                           ZN => n15916);
   U11776 : INV_X1 port map( A => n15915, ZN => n10237);
   U11777 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1462_port, B2 => n2778, 
                           ZN => n15915);
   U11778 : INV_X1 port map( A => n15914, ZN => n10238);
   U11779 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1461_port, B2 => n2778, 
                           ZN => n15914);
   U11780 : INV_X1 port map( A => n15913, ZN => n10239);
   U11781 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2774, B1 => 
                           DataPath_RF_bus_reg_dataout_1460_port, B2 => n2778, 
                           ZN => n15913);
   U11782 : INV_X1 port map( A => n15912, ZN => n10240);
   U11783 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1459_port, B2 => n2778, 
                           ZN => n15912);
   U11784 : INV_X1 port map( A => n15911, ZN => n10241);
   U11785 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1458_port, B2 => n2778, 
                           ZN => n15911);
   U11786 : INV_X1 port map( A => n15910, ZN => n10242);
   U11787 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1457_port, B2 => n2778, 
                           ZN => n15910);
   U11788 : INV_X1 port map( A => n15909, ZN => n10243);
   U11789 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1456_port, B2 => n2778, 
                           ZN => n15909);
   U11790 : INV_X1 port map( A => n15908, ZN => n10244);
   U11791 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1455_port, B2 => n2778, 
                           ZN => n15908);
   U11792 : INV_X1 port map( A => n15907, ZN => n10245);
   U11793 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1454_port, B2 => n2778, 
                           ZN => n15907);
   U11794 : INV_X1 port map( A => n15906, ZN => n10246);
   U11795 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1453_port, B2 => n2778, 
                           ZN => n15906);
   U11796 : INV_X1 port map( A => n15905, ZN => n10247);
   U11797 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1452_port, B2 => n2778, 
                           ZN => n15905);
   U11798 : INV_X1 port map( A => n15904, ZN => n10248);
   U11799 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1451_port, B2 => n2777, 
                           ZN => n15904);
   U11800 : INV_X1 port map( A => n15903, ZN => n10249);
   U11801 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1450_port, B2 => n2777, 
                           ZN => n15903);
   U11802 : INV_X1 port map( A => n15902, ZN => n10250);
   U11803 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1449_port, B2 => n2777, 
                           ZN => n15902);
   U11804 : INV_X1 port map( A => n15901, ZN => n10251);
   U11805 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2775, B1 => 
                           DataPath_RF_bus_reg_dataout_1448_port, B2 => n2777, 
                           ZN => n15901);
   U11806 : INV_X1 port map( A => n15900, ZN => n10252);
   U11807 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1447_port, B2 => n2777, 
                           ZN => n15900);
   U11808 : INV_X1 port map( A => n15899, ZN => n10253);
   U11809 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1446_port, B2 => n2777, 
                           ZN => n15899);
   U11810 : INV_X1 port map( A => n15898, ZN => n10254);
   U11811 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1445_port, B2 => n2777, 
                           ZN => n15898);
   U11812 : INV_X1 port map( A => n15897, ZN => n10255);
   U11813 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1444_port, B2 => n2777, 
                           ZN => n15897);
   U11814 : INV_X1 port map( A => n15896, ZN => n10256);
   U11815 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1443_port, B2 => n2777, 
                           ZN => n15896);
   U11816 : INV_X1 port map( A => n15895, ZN => n10257);
   U11817 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1442_port, B2 => n2777, 
                           ZN => n15895);
   U11818 : INV_X1 port map( A => n15894, ZN => n10258);
   U11819 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1441_port, B2 => n2777, 
                           ZN => n15894);
   U11820 : INV_X1 port map( A => n15891, ZN => n10259);
   U11821 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2776, B1 => 
                           DataPath_RF_bus_reg_dataout_1440_port, B2 => n2777, 
                           ZN => n15891);
   U11822 : INV_X1 port map( A => n15958, ZN => n10260);
   U11823 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1503_port, B2 => n2785, 
                           ZN => n15958);
   U11824 : INV_X1 port map( A => n15957, ZN => n10261);
   U11825 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1502_port, B2 => n2785, 
                           ZN => n15957);
   U11826 : INV_X1 port map( A => n15956, ZN => n10262);
   U11827 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1501_port, B2 => n2785, 
                           ZN => n15956);
   U11828 : INV_X1 port map( A => n15955, ZN => n10263);
   U11829 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1500_port, B2 => n2785, 
                           ZN => n15955);
   U11830 : INV_X1 port map( A => n15954, ZN => n10264);
   U11831 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1499_port, B2 => n2785, 
                           ZN => n15954);
   U11832 : INV_X1 port map( A => n15953, ZN => n10265);
   U11833 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1498_port, B2 => n2785, 
                           ZN => n15953);
   U11834 : INV_X1 port map( A => n15952, ZN => n10266);
   U11835 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1497_port, B2 => n2785, 
                           ZN => n15952);
   U11836 : INV_X1 port map( A => n15951, ZN => n10267);
   U11837 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1496_port, B2 => n2785, 
                           ZN => n15951);
   U11838 : INV_X1 port map( A => n15950, ZN => n10268);
   U11839 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1495_port, B2 => n2784, 
                           ZN => n15950);
   U11840 : INV_X1 port map( A => n15949, ZN => n10269);
   U11841 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1494_port, B2 => n2784, 
                           ZN => n15949);
   U11842 : INV_X1 port map( A => n15948, ZN => n10270);
   U11843 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1493_port, B2 => n2784, 
                           ZN => n15948);
   U11844 : INV_X1 port map( A => n15947, ZN => n10271);
   U11845 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2780, B1 => 
                           DataPath_RF_bus_reg_dataout_1492_port, B2 => n2784, 
                           ZN => n15947);
   U11846 : INV_X1 port map( A => n15946, ZN => n10272);
   U11847 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1491_port, B2 => n2784, 
                           ZN => n15946);
   U11848 : INV_X1 port map( A => n15945, ZN => n10273);
   U11849 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1490_port, B2 => n2784, 
                           ZN => n15945);
   U11850 : INV_X1 port map( A => n15944, ZN => n10274);
   U11851 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1489_port, B2 => n2784, 
                           ZN => n15944);
   U11852 : INV_X1 port map( A => n15943, ZN => n10275);
   U11853 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1488_port, B2 => n2784, 
                           ZN => n15943);
   U11854 : INV_X1 port map( A => n15942, ZN => n10276);
   U11855 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1487_port, B2 => n2784, 
                           ZN => n15942);
   U11856 : INV_X1 port map( A => n15941, ZN => n10277);
   U11857 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1486_port, B2 => n2784, 
                           ZN => n15941);
   U11858 : INV_X1 port map( A => n15940, ZN => n10278);
   U11859 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1485_port, B2 => n2784, 
                           ZN => n15940);
   U11860 : INV_X1 port map( A => n15939, ZN => n10279);
   U11861 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1484_port, B2 => n2784, 
                           ZN => n15939);
   U11862 : INV_X1 port map( A => n15938, ZN => n10280);
   U11863 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1483_port, B2 => n2783, 
                           ZN => n15938);
   U11864 : INV_X1 port map( A => n15937, ZN => n10281);
   U11865 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1482_port, B2 => n2783, 
                           ZN => n15937);
   U11866 : INV_X1 port map( A => n15936, ZN => n10282);
   U11867 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1481_port, B2 => n2783, 
                           ZN => n15936);
   U11868 : INV_X1 port map( A => n15935, ZN => n10283);
   U11869 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2781, B1 => 
                           DataPath_RF_bus_reg_dataout_1480_port, B2 => n2783, 
                           ZN => n15935);
   U11870 : INV_X1 port map( A => n15934, ZN => n10284);
   U11871 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1479_port, B2 => n2783, 
                           ZN => n15934);
   U11872 : INV_X1 port map( A => n15933, ZN => n10285);
   U11873 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1478_port, B2 => n2783, 
                           ZN => n15933);
   U11874 : INV_X1 port map( A => n15932, ZN => n10286);
   U11875 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1477_port, B2 => n2783, 
                           ZN => n15932);
   U11876 : INV_X1 port map( A => n15931, ZN => n10287);
   U11877 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1476_port, B2 => n2783, 
                           ZN => n15931);
   U11878 : INV_X1 port map( A => n15930, ZN => n10288);
   U11879 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1475_port, B2 => n2783, 
                           ZN => n15930);
   U11880 : INV_X1 port map( A => n15929, ZN => n10289);
   U11881 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1474_port, B2 => n2783, 
                           ZN => n15929);
   U11882 : INV_X1 port map( A => n15928, ZN => n10290);
   U11883 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1473_port, B2 => n2783, 
                           ZN => n15928);
   U11884 : INV_X1 port map( A => n15925, ZN => n10291);
   U11885 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2782, B1 => 
                           DataPath_RF_bus_reg_dataout_1472_port, B2 => n2783, 
                           ZN => n15925);
   U11886 : INV_X1 port map( A => n15992, ZN => n10292);
   U11887 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_31_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1535_port, B2 => n2791, 
                           ZN => n15992);
   U11888 : INV_X1 port map( A => n15991, ZN => n10293);
   U11889 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_30_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1534_port, B2 => n2791, 
                           ZN => n15991);
   U11890 : INV_X1 port map( A => n15990, ZN => n10294);
   U11891 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_29_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1533_port, B2 => n2791, 
                           ZN => n15990);
   U11892 : INV_X1 port map( A => n15989, ZN => n10295);
   U11893 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_28_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1532_port, B2 => n2791, 
                           ZN => n15989);
   U11894 : INV_X1 port map( A => n15988, ZN => n10296);
   U11895 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_27_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1531_port, B2 => n2791, 
                           ZN => n15988);
   U11896 : INV_X1 port map( A => n15987, ZN => n10297);
   U11897 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_26_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1530_port, B2 => n2791, 
                           ZN => n15987);
   U11898 : INV_X1 port map( A => n15986, ZN => n10298);
   U11899 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_25_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1529_port, B2 => n2791, 
                           ZN => n15986);
   U11900 : INV_X1 port map( A => n15985, ZN => n10299);
   U11901 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_24_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1528_port, B2 => n2791, 
                           ZN => n15985);
   U11902 : INV_X1 port map( A => n15984, ZN => n10300);
   U11903 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_23_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1527_port, B2 => n2790, 
                           ZN => n15984);
   U11904 : INV_X1 port map( A => n15983, ZN => n10301);
   U11905 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_22_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1526_port, B2 => n2790, 
                           ZN => n15983);
   U11906 : INV_X1 port map( A => n15982, ZN => n10302);
   U11907 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_21_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1525_port, B2 => n2790, 
                           ZN => n15982);
   U11908 : INV_X1 port map( A => n15981, ZN => n10303);
   U11909 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_20_port,
                           A2 => n2786, B1 => 
                           DataPath_RF_bus_reg_dataout_1524_port, B2 => n2790, 
                           ZN => n15981);
   U11910 : INV_X1 port map( A => n15980, ZN => n10304);
   U11911 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_19_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1523_port, B2 => n2790, 
                           ZN => n15980);
   U11912 : INV_X1 port map( A => n15979, ZN => n10305);
   U11913 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_18_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1522_port, B2 => n2790, 
                           ZN => n15979);
   U11914 : INV_X1 port map( A => n15978, ZN => n10306);
   U11915 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_17_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1521_port, B2 => n2790, 
                           ZN => n15978);
   U11916 : INV_X1 port map( A => n15977, ZN => n10307);
   U11917 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_16_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1520_port, B2 => n2790, 
                           ZN => n15977);
   U11918 : INV_X1 port map( A => n15976, ZN => n10308);
   U11919 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_15_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1519_port, B2 => n2790, 
                           ZN => n15976);
   U11920 : INV_X1 port map( A => n15975, ZN => n10309);
   U11921 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_14_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1518_port, B2 => n2790, 
                           ZN => n15975);
   U11922 : INV_X1 port map( A => n15974, ZN => n10310);
   U11923 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_13_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1517_port, B2 => n2790, 
                           ZN => n15974);
   U11924 : INV_X1 port map( A => n15973, ZN => n10311);
   U11925 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_12_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1516_port, B2 => n2790, 
                           ZN => n15973);
   U11926 : INV_X1 port map( A => n15972, ZN => n10312);
   U11927 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_11_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1515_port, B2 => n2789, 
                           ZN => n15972);
   U11928 : INV_X1 port map( A => n15971, ZN => n10313);
   U11929 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_10_port,
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1514_port, B2 => n2789, 
                           ZN => n15971);
   U11930 : INV_X1 port map( A => n15970, ZN => n10314);
   U11931 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_9_port, 
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1513_port, B2 => n2789, 
                           ZN => n15970);
   U11932 : INV_X1 port map( A => n15969, ZN => n10315);
   U11933 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_8_port, 
                           A2 => n2787, B1 => 
                           DataPath_RF_bus_reg_dataout_1512_port, B2 => n2789, 
                           ZN => n15969);
   U11934 : INV_X1 port map( A => n15968, ZN => n10316);
   U11935 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_7_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1511_port, B2 => n2789, 
                           ZN => n15968);
   U11936 : INV_X1 port map( A => n15967, ZN => n10317);
   U11937 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_6_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1510_port, B2 => n2789, 
                           ZN => n15967);
   U11938 : INV_X1 port map( A => n15966, ZN => n10318);
   U11939 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_5_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1509_port, B2 => n2789, 
                           ZN => n15966);
   U11940 : INV_X1 port map( A => n15965, ZN => n10319);
   U11941 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_4_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1508_port, B2 => n2789, 
                           ZN => n15965);
   U11942 : INV_X1 port map( A => n15964, ZN => n10320);
   U11943 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_3_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1507_port, B2 => n2789, 
                           ZN => n15964);
   U11944 : INV_X1 port map( A => n15963, ZN => n10321);
   U11945 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_2_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1506_port, B2 => n2789, 
                           ZN => n15963);
   U11946 : INV_X1 port map( A => n15962, ZN => n10322);
   U11947 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_1_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1505_port, B2 => n2789, 
                           ZN => n15962);
   U11948 : INV_X1 port map( A => n15959, ZN => n10323);
   U11949 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_2_0_port, 
                           A2 => n2788, B1 => 
                           DataPath_RF_bus_reg_dataout_1504_port, B2 => n2789, 
                           ZN => n15959);
   U11950 : INV_X1 port map( A => n16026, ZN => n10324);
   U11951 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1567_port, B2 => n2797, 
                           ZN => n16026);
   U11952 : INV_X1 port map( A => n16025, ZN => n10325);
   U11953 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1566_port, B2 => n2797, 
                           ZN => n16025);
   U11954 : INV_X1 port map( A => n16024, ZN => n10326);
   U11955 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1565_port, B2 => n2797, 
                           ZN => n16024);
   U11956 : INV_X1 port map( A => n16023, ZN => n10327);
   U11957 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1564_port, B2 => n2797, 
                           ZN => n16023);
   U11958 : INV_X1 port map( A => n16022, ZN => n10328);
   U11959 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1563_port, B2 => n2797, 
                           ZN => n16022);
   U11960 : INV_X1 port map( A => n16021, ZN => n10329);
   U11961 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1562_port, B2 => n2797, 
                           ZN => n16021);
   U11962 : INV_X1 port map( A => n16020, ZN => n10330);
   U11963 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1561_port, B2 => n2797, 
                           ZN => n16020);
   U11964 : INV_X1 port map( A => n16019, ZN => n10331);
   U11965 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1560_port, B2 => n2797, 
                           ZN => n16019);
   U11966 : INV_X1 port map( A => n16018, ZN => n10332);
   U11967 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1559_port, B2 => n2796, 
                           ZN => n16018);
   U11968 : INV_X1 port map( A => n16017, ZN => n10333);
   U11969 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1558_port, B2 => n2796, 
                           ZN => n16017);
   U11970 : INV_X1 port map( A => n16016, ZN => n10334);
   U11971 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1557_port, B2 => n2796, 
                           ZN => n16016);
   U11972 : INV_X1 port map( A => n16015, ZN => n10335);
   U11973 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2792, B1 => 
                           DataPath_RF_bus_reg_dataout_1556_port, B2 => n2796, 
                           ZN => n16015);
   U11974 : INV_X1 port map( A => n16014, ZN => n10336);
   U11975 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1555_port, B2 => n2796, 
                           ZN => n16014);
   U11976 : INV_X1 port map( A => n16013, ZN => n10337);
   U11977 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1554_port, B2 => n2796, 
                           ZN => n16013);
   U11978 : INV_X1 port map( A => n16012, ZN => n10338);
   U11979 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1553_port, B2 => n2796, 
                           ZN => n16012);
   U11980 : INV_X1 port map( A => n16011, ZN => n10339);
   U11981 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1552_port, B2 => n2796, 
                           ZN => n16011);
   U11982 : INV_X1 port map( A => n16010, ZN => n10340);
   U11983 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1551_port, B2 => n2796, 
                           ZN => n16010);
   U11984 : INV_X1 port map( A => n16009, ZN => n10341);
   U11985 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1550_port, B2 => n2796, 
                           ZN => n16009);
   U11986 : INV_X1 port map( A => n16008, ZN => n10342);
   U11987 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1549_port, B2 => n2796, 
                           ZN => n16008);
   U11988 : INV_X1 port map( A => n16007, ZN => n10343);
   U11989 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1548_port, B2 => n2796, 
                           ZN => n16007);
   U11990 : INV_X1 port map( A => n16006, ZN => n10344);
   U11991 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1547_port, B2 => n2795, 
                           ZN => n16006);
   U11992 : INV_X1 port map( A => n16005, ZN => n10345);
   U11993 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1546_port, B2 => n2795, 
                           ZN => n16005);
   U11994 : INV_X1 port map( A => n16004, ZN => n10346);
   U11995 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1545_port, B2 => n2795, 
                           ZN => n16004);
   U11996 : INV_X1 port map( A => n16003, ZN => n10347);
   U11997 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2793, B1 => 
                           DataPath_RF_bus_reg_dataout_1544_port, B2 => n2795, 
                           ZN => n16003);
   U11998 : INV_X1 port map( A => n16002, ZN => n10348);
   U11999 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1543_port, B2 => n2795, 
                           ZN => n16002);
   U12000 : INV_X1 port map( A => n16001, ZN => n10349);
   U12001 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1542_port, B2 => n2795, 
                           ZN => n16001);
   U12002 : INV_X1 port map( A => n16000, ZN => n10350);
   U12003 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1541_port, B2 => n2795, 
                           ZN => n16000);
   U12004 : INV_X1 port map( A => n15999, ZN => n10351);
   U12005 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1540_port, B2 => n2795, 
                           ZN => n15999);
   U12006 : INV_X1 port map( A => n15998, ZN => n10352);
   U12007 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1539_port, B2 => n2795, 
                           ZN => n15998);
   U12008 : INV_X1 port map( A => n15997, ZN => n10353);
   U12009 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1538_port, B2 => n2795, 
                           ZN => n15997);
   U12010 : INV_X1 port map( A => n15996, ZN => n10354);
   U12011 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1537_port, B2 => n2795, 
                           ZN => n15996);
   U12012 : INV_X1 port map( A => n15993, ZN => n10355);
   U12013 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2794, B1 => 
                           DataPath_RF_bus_reg_dataout_1536_port, B2 => n2795, 
                           ZN => n15993);
   U12014 : INV_X1 port map( A => n16060, ZN => n10356);
   U12015 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1599_port, B2 => n2803, 
                           ZN => n16060);
   U12016 : INV_X1 port map( A => n16059, ZN => n10357);
   U12017 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1598_port, B2 => n2803, 
                           ZN => n16059);
   U12018 : INV_X1 port map( A => n16058, ZN => n10358);
   U12019 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1597_port, B2 => n2803, 
                           ZN => n16058);
   U12020 : INV_X1 port map( A => n16057, ZN => n10359);
   U12021 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1596_port, B2 => n2803, 
                           ZN => n16057);
   U12022 : INV_X1 port map( A => n16056, ZN => n10360);
   U12023 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1595_port, B2 => n2803, 
                           ZN => n16056);
   U12024 : INV_X1 port map( A => n16055, ZN => n10361);
   U12025 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1594_port, B2 => n2803, 
                           ZN => n16055);
   U12026 : INV_X1 port map( A => n16054, ZN => n10362);
   U12027 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1593_port, B2 => n2803, 
                           ZN => n16054);
   U12028 : INV_X1 port map( A => n16053, ZN => n10363);
   U12029 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1592_port, B2 => n2803, 
                           ZN => n16053);
   U12030 : INV_X1 port map( A => n16052, ZN => n10364);
   U12031 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1591_port, B2 => n2802, 
                           ZN => n16052);
   U12032 : INV_X1 port map( A => n16051, ZN => n10365);
   U12033 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1590_port, B2 => n2802, 
                           ZN => n16051);
   U12034 : INV_X1 port map( A => n16050, ZN => n10366);
   U12035 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1589_port, B2 => n2802, 
                           ZN => n16050);
   U12036 : INV_X1 port map( A => n16049, ZN => n10367);
   U12037 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2798, B1 => 
                           DataPath_RF_bus_reg_dataout_1588_port, B2 => n2802, 
                           ZN => n16049);
   U12038 : INV_X1 port map( A => n16048, ZN => n10368);
   U12039 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1587_port, B2 => n2802, 
                           ZN => n16048);
   U12040 : INV_X1 port map( A => n16047, ZN => n10369);
   U12041 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1586_port, B2 => n2802, 
                           ZN => n16047);
   U12042 : INV_X1 port map( A => n16046, ZN => n10370);
   U12043 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1585_port, B2 => n2802, 
                           ZN => n16046);
   U12044 : INV_X1 port map( A => n16045, ZN => n10371);
   U12045 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1584_port, B2 => n2802, 
                           ZN => n16045);
   U12046 : INV_X1 port map( A => n16044, ZN => n10372);
   U12047 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1583_port, B2 => n2802, 
                           ZN => n16044);
   U12048 : INV_X1 port map( A => n16043, ZN => n10373);
   U12049 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1582_port, B2 => n2802, 
                           ZN => n16043);
   U12050 : INV_X1 port map( A => n16042, ZN => n10374);
   U12051 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1581_port, B2 => n2802, 
                           ZN => n16042);
   U12052 : INV_X1 port map( A => n16041, ZN => n10375);
   U12053 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1580_port, B2 => n2802, 
                           ZN => n16041);
   U12054 : INV_X1 port map( A => n16040, ZN => n10376);
   U12055 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1579_port, B2 => n2801, 
                           ZN => n16040);
   U12056 : INV_X1 port map( A => n16039, ZN => n10377);
   U12057 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1578_port, B2 => n2801, 
                           ZN => n16039);
   U12058 : INV_X1 port map( A => n16038, ZN => n10378);
   U12059 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1577_port, B2 => n2801, 
                           ZN => n16038);
   U12060 : INV_X1 port map( A => n16037, ZN => n10379);
   U12061 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2799, B1 => 
                           DataPath_RF_bus_reg_dataout_1576_port, B2 => n2801, 
                           ZN => n16037);
   U12062 : INV_X1 port map( A => n16036, ZN => n10380);
   U12063 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1575_port, B2 => n2801, 
                           ZN => n16036);
   U12064 : INV_X1 port map( A => n16035, ZN => n10381);
   U12065 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1574_port, B2 => n2801, 
                           ZN => n16035);
   U12066 : INV_X1 port map( A => n16034, ZN => n10382);
   U12067 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1573_port, B2 => n2801, 
                           ZN => n16034);
   U12068 : INV_X1 port map( A => n16033, ZN => n10383);
   U12069 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1572_port, B2 => n2801, 
                           ZN => n16033);
   U12070 : INV_X1 port map( A => n16032, ZN => n10384);
   U12071 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1571_port, B2 => n2801, 
                           ZN => n16032);
   U12072 : INV_X1 port map( A => n16031, ZN => n10385);
   U12073 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1570_port, B2 => n2801, 
                           ZN => n16031);
   U12074 : INV_X1 port map( A => n16030, ZN => n10386);
   U12075 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1569_port, B2 => n2801, 
                           ZN => n16030);
   U12076 : INV_X1 port map( A => n16027, ZN => n10387);
   U12077 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2800, B1 => 
                           DataPath_RF_bus_reg_dataout_1568_port, B2 => n2801, 
                           ZN => n16027);
   U12078 : INV_X1 port map( A => n16094, ZN => n10388);
   U12079 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1631_port, B2 => n2809, 
                           ZN => n16094);
   U12080 : INV_X1 port map( A => n16093, ZN => n10389);
   U12081 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1630_port, B2 => n2809, 
                           ZN => n16093);
   U12082 : INV_X1 port map( A => n16092, ZN => n10390);
   U12083 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1629_port, B2 => n2809, 
                           ZN => n16092);
   U12084 : INV_X1 port map( A => n16091, ZN => n10391);
   U12085 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1628_port, B2 => n2809, 
                           ZN => n16091);
   U12086 : INV_X1 port map( A => n16090, ZN => n10392);
   U12087 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1627_port, B2 => n2809, 
                           ZN => n16090);
   U12088 : INV_X1 port map( A => n16089, ZN => n10393);
   U12089 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1626_port, B2 => n2809, 
                           ZN => n16089);
   U12090 : INV_X1 port map( A => n16088, ZN => n10394);
   U12091 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1625_port, B2 => n2809, 
                           ZN => n16088);
   U12092 : INV_X1 port map( A => n16087, ZN => n10395);
   U12093 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1624_port, B2 => n2809, 
                           ZN => n16087);
   U12094 : INV_X1 port map( A => n16086, ZN => n10396);
   U12095 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1623_port, B2 => n2808, 
                           ZN => n16086);
   U12096 : INV_X1 port map( A => n16085, ZN => n10397);
   U12097 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1622_port, B2 => n2808, 
                           ZN => n16085);
   U12098 : INV_X1 port map( A => n16084, ZN => n10398);
   U12099 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1621_port, B2 => n2808, 
                           ZN => n16084);
   U12100 : INV_X1 port map( A => n16083, ZN => n10399);
   U12101 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2804, B1 => 
                           DataPath_RF_bus_reg_dataout_1620_port, B2 => n2808, 
                           ZN => n16083);
   U12102 : INV_X1 port map( A => n16082, ZN => n10400);
   U12103 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1619_port, B2 => n2808, 
                           ZN => n16082);
   U12104 : INV_X1 port map( A => n16081, ZN => n10401);
   U12105 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1618_port, B2 => n2808, 
                           ZN => n16081);
   U12106 : INV_X1 port map( A => n16080, ZN => n10402);
   U12107 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1617_port, B2 => n2808, 
                           ZN => n16080);
   U12108 : INV_X1 port map( A => n16079, ZN => n10403);
   U12109 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1616_port, B2 => n2808, 
                           ZN => n16079);
   U12110 : INV_X1 port map( A => n16078, ZN => n10404);
   U12111 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1615_port, B2 => n2808, 
                           ZN => n16078);
   U12112 : INV_X1 port map( A => n16077, ZN => n10405);
   U12113 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1614_port, B2 => n2808, 
                           ZN => n16077);
   U12114 : INV_X1 port map( A => n16076, ZN => n10406);
   U12115 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1613_port, B2 => n2808, 
                           ZN => n16076);
   U12116 : INV_X1 port map( A => n16075, ZN => n10407);
   U12117 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1612_port, B2 => n2808, 
                           ZN => n16075);
   U12118 : INV_X1 port map( A => n16074, ZN => n10408);
   U12119 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1611_port, B2 => n2807, 
                           ZN => n16074);
   U12120 : INV_X1 port map( A => n16073, ZN => n10409);
   U12121 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1610_port, B2 => n2807, 
                           ZN => n16073);
   U12122 : INV_X1 port map( A => n16072, ZN => n10410);
   U12123 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1609_port, B2 => n2807, 
                           ZN => n16072);
   U12124 : INV_X1 port map( A => n16071, ZN => n10411);
   U12125 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2805, B1 => 
                           DataPath_RF_bus_reg_dataout_1608_port, B2 => n2807, 
                           ZN => n16071);
   U12126 : INV_X1 port map( A => n16070, ZN => n10412);
   U12127 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1607_port, B2 => n2807, 
                           ZN => n16070);
   U12128 : INV_X1 port map( A => n16069, ZN => n10413);
   U12129 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1606_port, B2 => n2807, 
                           ZN => n16069);
   U12130 : INV_X1 port map( A => n16068, ZN => n10414);
   U12131 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1605_port, B2 => n2807, 
                           ZN => n16068);
   U12132 : INV_X1 port map( A => n16067, ZN => n10415);
   U12133 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1604_port, B2 => n2807, 
                           ZN => n16067);
   U12134 : INV_X1 port map( A => n16066, ZN => n10416);
   U12135 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1603_port, B2 => n2807, 
                           ZN => n16066);
   U12136 : INV_X1 port map( A => n16065, ZN => n10417);
   U12137 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1602_port, B2 => n2807, 
                           ZN => n16065);
   U12138 : INV_X1 port map( A => n16064, ZN => n10418);
   U12139 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1601_port, B2 => n2807, 
                           ZN => n16064);
   U12140 : INV_X1 port map( A => n16061, ZN => n10419);
   U12141 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2806, B1 => 
                           DataPath_RF_bus_reg_dataout_1600_port, B2 => n2807, 
                           ZN => n16061);
   U12142 : INV_X1 port map( A => n16128, ZN => n10420);
   U12143 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1663_port, B2 => n2815, 
                           ZN => n16128);
   U12144 : INV_X1 port map( A => n16127, ZN => n10421);
   U12145 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1662_port, B2 => n2815, 
                           ZN => n16127);
   U12146 : INV_X1 port map( A => n16126, ZN => n10422);
   U12147 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1661_port, B2 => n2815, 
                           ZN => n16126);
   U12148 : INV_X1 port map( A => n16125, ZN => n10423);
   U12149 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1660_port, B2 => n2815, 
                           ZN => n16125);
   U12150 : INV_X1 port map( A => n16124, ZN => n10424);
   U12151 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1659_port, B2 => n2815, 
                           ZN => n16124);
   U12152 : INV_X1 port map( A => n16123, ZN => n10425);
   U12153 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1658_port, B2 => n2815, 
                           ZN => n16123);
   U12154 : INV_X1 port map( A => n16122, ZN => n10426);
   U12155 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1657_port, B2 => n2815, 
                           ZN => n16122);
   U12156 : INV_X1 port map( A => n16121, ZN => n10427);
   U12157 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1656_port, B2 => n2815, 
                           ZN => n16121);
   U12158 : INV_X1 port map( A => n16120, ZN => n10428);
   U12159 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1655_port, B2 => n2814, 
                           ZN => n16120);
   U12160 : INV_X1 port map( A => n16119, ZN => n10429);
   U12161 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1654_port, B2 => n2814, 
                           ZN => n16119);
   U12162 : INV_X1 port map( A => n16118, ZN => n10430);
   U12163 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1653_port, B2 => n2814, 
                           ZN => n16118);
   U12164 : INV_X1 port map( A => n16117, ZN => n10431);
   U12165 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2810, B1 => 
                           DataPath_RF_bus_reg_dataout_1652_port, B2 => n2814, 
                           ZN => n16117);
   U12166 : INV_X1 port map( A => n16116, ZN => n10432);
   U12167 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1651_port, B2 => n2814, 
                           ZN => n16116);
   U12168 : INV_X1 port map( A => n16115, ZN => n10433);
   U12169 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1650_port, B2 => n2814, 
                           ZN => n16115);
   U12170 : INV_X1 port map( A => n16114, ZN => n10434);
   U12171 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1649_port, B2 => n2814, 
                           ZN => n16114);
   U12172 : INV_X1 port map( A => n16113, ZN => n10435);
   U12173 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1648_port, B2 => n2814, 
                           ZN => n16113);
   U12174 : INV_X1 port map( A => n16112, ZN => n10436);
   U12175 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1647_port, B2 => n2814, 
                           ZN => n16112);
   U12176 : INV_X1 port map( A => n16111, ZN => n10437);
   U12177 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1646_port, B2 => n2814, 
                           ZN => n16111);
   U12178 : INV_X1 port map( A => n16110, ZN => n10438);
   U12179 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1645_port, B2 => n2814, 
                           ZN => n16110);
   U12180 : INV_X1 port map( A => n16109, ZN => n10439);
   U12181 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1644_port, B2 => n2814, 
                           ZN => n16109);
   U12182 : INV_X1 port map( A => n16108, ZN => n10440);
   U12183 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1643_port, B2 => n2813, 
                           ZN => n16108);
   U12184 : INV_X1 port map( A => n16107, ZN => n10441);
   U12185 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1642_port, B2 => n2813, 
                           ZN => n16107);
   U12186 : INV_X1 port map( A => n16106, ZN => n10442);
   U12187 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1641_port, B2 => n2813, 
                           ZN => n16106);
   U12188 : INV_X1 port map( A => n16105, ZN => n10443);
   U12189 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2811, B1 => 
                           DataPath_RF_bus_reg_dataout_1640_port, B2 => n2813, 
                           ZN => n16105);
   U12190 : INV_X1 port map( A => n16104, ZN => n10444);
   U12191 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1639_port, B2 => n2813, 
                           ZN => n16104);
   U12192 : INV_X1 port map( A => n16103, ZN => n10445);
   U12193 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1638_port, B2 => n2813, 
                           ZN => n16103);
   U12194 : INV_X1 port map( A => n16102, ZN => n10446);
   U12195 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1637_port, B2 => n2813, 
                           ZN => n16102);
   U12196 : INV_X1 port map( A => n16101, ZN => n10447);
   U12197 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1636_port, B2 => n2813, 
                           ZN => n16101);
   U12198 : INV_X1 port map( A => n16100, ZN => n10448);
   U12199 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1635_port, B2 => n2813, 
                           ZN => n16100);
   U12200 : INV_X1 port map( A => n16099, ZN => n10449);
   U12201 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1634_port, B2 => n2813, 
                           ZN => n16099);
   U12202 : INV_X1 port map( A => n16098, ZN => n10450);
   U12203 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1633_port, B2 => n2813, 
                           ZN => n16098);
   U12204 : INV_X1 port map( A => n16095, ZN => n10451);
   U12205 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2812, B1 => 
                           DataPath_RF_bus_reg_dataout_1632_port, B2 => n2813, 
                           ZN => n16095);
   U12206 : INV_X1 port map( A => n16162, ZN => n10452);
   U12207 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1695_port, B2 => n2821, 
                           ZN => n16162);
   U12208 : INV_X1 port map( A => n16161, ZN => n10453);
   U12209 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1694_port, B2 => n2821, 
                           ZN => n16161);
   U12210 : INV_X1 port map( A => n16160, ZN => n10454);
   U12211 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1693_port, B2 => n2821, 
                           ZN => n16160);
   U12212 : INV_X1 port map( A => n16159, ZN => n10455);
   U12213 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1692_port, B2 => n2821, 
                           ZN => n16159);
   U12214 : INV_X1 port map( A => n16158, ZN => n10456);
   U12215 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1691_port, B2 => n2821, 
                           ZN => n16158);
   U12216 : INV_X1 port map( A => n16157, ZN => n10457);
   U12217 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1690_port, B2 => n2821, 
                           ZN => n16157);
   U12218 : INV_X1 port map( A => n16156, ZN => n10458);
   U12219 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1689_port, B2 => n2821, 
                           ZN => n16156);
   U12220 : INV_X1 port map( A => n16155, ZN => n10459);
   U12221 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1688_port, B2 => n2821, 
                           ZN => n16155);
   U12222 : INV_X1 port map( A => n16154, ZN => n10460);
   U12223 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1687_port, B2 => n2820, 
                           ZN => n16154);
   U12224 : INV_X1 port map( A => n16153, ZN => n10461);
   U12225 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1686_port, B2 => n2820, 
                           ZN => n16153);
   U12226 : INV_X1 port map( A => n16152, ZN => n10462);
   U12227 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1685_port, B2 => n2820, 
                           ZN => n16152);
   U12228 : INV_X1 port map( A => n16151, ZN => n10463);
   U12229 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2816, B1 => 
                           DataPath_RF_bus_reg_dataout_1684_port, B2 => n2820, 
                           ZN => n16151);
   U12230 : INV_X1 port map( A => n16150, ZN => n10464);
   U12231 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1683_port, B2 => n2820, 
                           ZN => n16150);
   U12232 : INV_X1 port map( A => n16149, ZN => n10465);
   U12233 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1682_port, B2 => n2820, 
                           ZN => n16149);
   U12234 : INV_X1 port map( A => n16148, ZN => n10466);
   U12235 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1681_port, B2 => n2820, 
                           ZN => n16148);
   U12236 : INV_X1 port map( A => n16147, ZN => n10467);
   U12237 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1680_port, B2 => n2820, 
                           ZN => n16147);
   U12238 : INV_X1 port map( A => n16146, ZN => n10468);
   U12239 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1679_port, B2 => n2820, 
                           ZN => n16146);
   U12240 : INV_X1 port map( A => n16145, ZN => n10469);
   U12241 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1678_port, B2 => n2820, 
                           ZN => n16145);
   U12242 : INV_X1 port map( A => n16144, ZN => n10470);
   U12243 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1677_port, B2 => n2820, 
                           ZN => n16144);
   U12244 : INV_X1 port map( A => n16143, ZN => n10471);
   U12245 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1676_port, B2 => n2820, 
                           ZN => n16143);
   U12246 : INV_X1 port map( A => n16142, ZN => n10472);
   U12247 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1675_port, B2 => n2819, 
                           ZN => n16142);
   U12248 : INV_X1 port map( A => n16141, ZN => n10473);
   U12249 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1674_port, B2 => n2819, 
                           ZN => n16141);
   U12250 : INV_X1 port map( A => n16140, ZN => n10474);
   U12251 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1673_port, B2 => n2819, 
                           ZN => n16140);
   U12252 : INV_X1 port map( A => n16139, ZN => n10475);
   U12253 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2817, B1 => 
                           DataPath_RF_bus_reg_dataout_1672_port, B2 => n2819, 
                           ZN => n16139);
   U12254 : INV_X1 port map( A => n16138, ZN => n10476);
   U12255 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1671_port, B2 => n2819, 
                           ZN => n16138);
   U12256 : INV_X1 port map( A => n16137, ZN => n10477);
   U12257 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1670_port, B2 => n2819, 
                           ZN => n16137);
   U12258 : INV_X1 port map( A => n16136, ZN => n10478);
   U12259 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1669_port, B2 => n2819, 
                           ZN => n16136);
   U12260 : INV_X1 port map( A => n16135, ZN => n10479);
   U12261 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1668_port, B2 => n2819, 
                           ZN => n16135);
   U12262 : INV_X1 port map( A => n16134, ZN => n10480);
   U12263 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1667_port, B2 => n2819, 
                           ZN => n16134);
   U12264 : INV_X1 port map( A => n16133, ZN => n10481);
   U12265 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1666_port, B2 => n2819, 
                           ZN => n16133);
   U12266 : INV_X1 port map( A => n16132, ZN => n10482);
   U12267 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1665_port, B2 => n2819, 
                           ZN => n16132);
   U12268 : INV_X1 port map( A => n16129, ZN => n10483);
   U12269 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2818, B1 => 
                           DataPath_RF_bus_reg_dataout_1664_port, B2 => n2819, 
                           ZN => n16129);
   U12270 : INV_X1 port map( A => n16196, ZN => n10484);
   U12271 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1727_port, B2 => n2827, 
                           ZN => n16196);
   U12272 : INV_X1 port map( A => n16195, ZN => n10485);
   U12273 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1726_port, B2 => n2827, 
                           ZN => n16195);
   U12274 : INV_X1 port map( A => n16194, ZN => n10486);
   U12275 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1725_port, B2 => n2827, 
                           ZN => n16194);
   U12276 : INV_X1 port map( A => n16193, ZN => n10487);
   U12277 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1724_port, B2 => n2827, 
                           ZN => n16193);
   U12278 : INV_X1 port map( A => n16192, ZN => n10488);
   U12279 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1723_port, B2 => n2827, 
                           ZN => n16192);
   U12280 : INV_X1 port map( A => n16191, ZN => n10489);
   U12281 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1722_port, B2 => n2827, 
                           ZN => n16191);
   U12282 : INV_X1 port map( A => n16190, ZN => n10490);
   U12283 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1721_port, B2 => n2827, 
                           ZN => n16190);
   U12284 : INV_X1 port map( A => n16189, ZN => n10491);
   U12285 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1720_port, B2 => n2827, 
                           ZN => n16189);
   U12286 : INV_X1 port map( A => n16188, ZN => n10492);
   U12287 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1719_port, B2 => n2826, 
                           ZN => n16188);
   U12288 : INV_X1 port map( A => n16187, ZN => n10493);
   U12289 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1718_port, B2 => n2826, 
                           ZN => n16187);
   U12290 : INV_X1 port map( A => n16186, ZN => n10494);
   U12291 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1717_port, B2 => n2826, 
                           ZN => n16186);
   U12292 : INV_X1 port map( A => n16185, ZN => n10495);
   U12293 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2822, B1 => 
                           DataPath_RF_bus_reg_dataout_1716_port, B2 => n2826, 
                           ZN => n16185);
   U12294 : INV_X1 port map( A => n16184, ZN => n10496);
   U12295 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1715_port, B2 => n2826, 
                           ZN => n16184);
   U12296 : INV_X1 port map( A => n16183, ZN => n10497);
   U12297 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1714_port, B2 => n2826, 
                           ZN => n16183);
   U12298 : INV_X1 port map( A => n16182, ZN => n10498);
   U12299 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1713_port, B2 => n2826, 
                           ZN => n16182);
   U12300 : INV_X1 port map( A => n16181, ZN => n10499);
   U12301 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1712_port, B2 => n2826, 
                           ZN => n16181);
   U12302 : INV_X1 port map( A => n16180, ZN => n10500);
   U12303 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1711_port, B2 => n2826, 
                           ZN => n16180);
   U12304 : INV_X1 port map( A => n16179, ZN => n10501);
   U12305 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1710_port, B2 => n2826, 
                           ZN => n16179);
   U12306 : INV_X1 port map( A => n16178, ZN => n10502);
   U12307 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1709_port, B2 => n2826, 
                           ZN => n16178);
   U12308 : INV_X1 port map( A => n16177, ZN => n10503);
   U12309 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1708_port, B2 => n2826, 
                           ZN => n16177);
   U12310 : INV_X1 port map( A => n16176, ZN => n10504);
   U12311 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1707_port, B2 => n2825, 
                           ZN => n16176);
   U12312 : INV_X1 port map( A => n16175, ZN => n10505);
   U12313 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1706_port, B2 => n2825, 
                           ZN => n16175);
   U12314 : INV_X1 port map( A => n16174, ZN => n10506);
   U12315 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1705_port, B2 => n2825, 
                           ZN => n16174);
   U12316 : INV_X1 port map( A => n16173, ZN => n10507);
   U12317 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2823, B1 => 
                           DataPath_RF_bus_reg_dataout_1704_port, B2 => n2825, 
                           ZN => n16173);
   U12318 : INV_X1 port map( A => n16172, ZN => n10508);
   U12319 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1703_port, B2 => n2825, 
                           ZN => n16172);
   U12320 : INV_X1 port map( A => n16171, ZN => n10509);
   U12321 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1702_port, B2 => n2825, 
                           ZN => n16171);
   U12322 : INV_X1 port map( A => n16170, ZN => n10510);
   U12323 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1701_port, B2 => n2825, 
                           ZN => n16170);
   U12324 : INV_X1 port map( A => n16169, ZN => n10511);
   U12325 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1700_port, B2 => n2825, 
                           ZN => n16169);
   U12326 : INV_X1 port map( A => n16168, ZN => n10512);
   U12327 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1699_port, B2 => n2825, 
                           ZN => n16168);
   U12328 : INV_X1 port map( A => n16167, ZN => n10513);
   U12329 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1698_port, B2 => n2825, 
                           ZN => n16167);
   U12330 : INV_X1 port map( A => n16166, ZN => n10514);
   U12331 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1697_port, B2 => n2825, 
                           ZN => n16166);
   U12332 : INV_X1 port map( A => n16163, ZN => n10515);
   U12333 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2824, B1 => 
                           DataPath_RF_bus_reg_dataout_1696_port, B2 => n2825, 
                           ZN => n16163);
   U12334 : INV_X1 port map( A => n16230, ZN => n10516);
   U12335 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1759_port, B2 => n2833, 
                           ZN => n16230);
   U12336 : INV_X1 port map( A => n16229, ZN => n10517);
   U12337 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1758_port, B2 => n2833, 
                           ZN => n16229);
   U12338 : INV_X1 port map( A => n16228, ZN => n10518);
   U12339 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1757_port, B2 => n2833, 
                           ZN => n16228);
   U12340 : INV_X1 port map( A => n16227, ZN => n10519);
   U12341 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1756_port, B2 => n2833, 
                           ZN => n16227);
   U12342 : INV_X1 port map( A => n16226, ZN => n10520);
   U12343 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1755_port, B2 => n2833, 
                           ZN => n16226);
   U12344 : INV_X1 port map( A => n16225, ZN => n10521);
   U12345 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1754_port, B2 => n2833, 
                           ZN => n16225);
   U12346 : INV_X1 port map( A => n16224, ZN => n10522);
   U12347 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1753_port, B2 => n2833, 
                           ZN => n16224);
   U12348 : INV_X1 port map( A => n16223, ZN => n10523);
   U12349 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1752_port, B2 => n2833, 
                           ZN => n16223);
   U12350 : INV_X1 port map( A => n16222, ZN => n10524);
   U12351 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1751_port, B2 => n2832, 
                           ZN => n16222);
   U12352 : INV_X1 port map( A => n16221, ZN => n10525);
   U12353 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1750_port, B2 => n2832, 
                           ZN => n16221);
   U12354 : INV_X1 port map( A => n16220, ZN => n10526);
   U12355 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1749_port, B2 => n2832, 
                           ZN => n16220);
   U12356 : INV_X1 port map( A => n16219, ZN => n10527);
   U12357 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2828, B1 => 
                           DataPath_RF_bus_reg_dataout_1748_port, B2 => n2832, 
                           ZN => n16219);
   U12358 : INV_X1 port map( A => n16218, ZN => n10528);
   U12359 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1747_port, B2 => n2832, 
                           ZN => n16218);
   U12360 : INV_X1 port map( A => n16217, ZN => n10529);
   U12361 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1746_port, B2 => n2832, 
                           ZN => n16217);
   U12362 : INV_X1 port map( A => n16216, ZN => n10530);
   U12363 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1745_port, B2 => n2832, 
                           ZN => n16216);
   U12364 : INV_X1 port map( A => n16215, ZN => n10531);
   U12365 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1744_port, B2 => n2832, 
                           ZN => n16215);
   U12366 : INV_X1 port map( A => n16214, ZN => n10532);
   U12367 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1743_port, B2 => n2832, 
                           ZN => n16214);
   U12368 : INV_X1 port map( A => n16213, ZN => n10533);
   U12369 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1742_port, B2 => n2832, 
                           ZN => n16213);
   U12370 : INV_X1 port map( A => n16212, ZN => n10534);
   U12371 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1741_port, B2 => n2832, 
                           ZN => n16212);
   U12372 : INV_X1 port map( A => n16211, ZN => n10535);
   U12373 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1740_port, B2 => n2832, 
                           ZN => n16211);
   U12374 : INV_X1 port map( A => n16210, ZN => n10536);
   U12375 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1739_port, B2 => n2831, 
                           ZN => n16210);
   U12376 : INV_X1 port map( A => n16209, ZN => n10537);
   U12377 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1738_port, B2 => n2831, 
                           ZN => n16209);
   U12378 : INV_X1 port map( A => n16208, ZN => n10538);
   U12379 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1737_port, B2 => n2831, 
                           ZN => n16208);
   U12380 : INV_X1 port map( A => n16207, ZN => n10539);
   U12381 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2829, B1 => 
                           DataPath_RF_bus_reg_dataout_1736_port, B2 => n2831, 
                           ZN => n16207);
   U12382 : INV_X1 port map( A => n16206, ZN => n10540);
   U12383 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1735_port, B2 => n2831, 
                           ZN => n16206);
   U12384 : INV_X1 port map( A => n16205, ZN => n10541);
   U12385 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1734_port, B2 => n2831, 
                           ZN => n16205);
   U12386 : INV_X1 port map( A => n16204, ZN => n10542);
   U12387 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1733_port, B2 => n2831, 
                           ZN => n16204);
   U12388 : INV_X1 port map( A => n16203, ZN => n10543);
   U12389 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1732_port, B2 => n2831, 
                           ZN => n16203);
   U12390 : INV_X1 port map( A => n16202, ZN => n10544);
   U12391 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1731_port, B2 => n2831, 
                           ZN => n16202);
   U12392 : INV_X1 port map( A => n16201, ZN => n10545);
   U12393 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1730_port, B2 => n2831, 
                           ZN => n16201);
   U12394 : INV_X1 port map( A => n16200, ZN => n10546);
   U12395 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1729_port, B2 => n2831, 
                           ZN => n16200);
   U12396 : INV_X1 port map( A => n16197, ZN => n10547);
   U12397 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2830, B1 => 
                           DataPath_RF_bus_reg_dataout_1728_port, B2 => n2831, 
                           ZN => n16197);
   U12398 : INV_X1 port map( A => n16264, ZN => n10548);
   U12399 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1791_port, B2 => n2839, 
                           ZN => n16264);
   U12400 : INV_X1 port map( A => n16263, ZN => n10549);
   U12401 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1790_port, B2 => n2839, 
                           ZN => n16263);
   U12402 : INV_X1 port map( A => n16262, ZN => n10550);
   U12403 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1789_port, B2 => n2839, 
                           ZN => n16262);
   U12404 : INV_X1 port map( A => n16261, ZN => n10551);
   U12405 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1788_port, B2 => n2839, 
                           ZN => n16261);
   U12406 : INV_X1 port map( A => n16260, ZN => n10552);
   U12407 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1787_port, B2 => n2839, 
                           ZN => n16260);
   U12408 : INV_X1 port map( A => n16259, ZN => n10553);
   U12409 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1786_port, B2 => n2839, 
                           ZN => n16259);
   U12410 : INV_X1 port map( A => n16258, ZN => n10554);
   U12411 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1785_port, B2 => n2839, 
                           ZN => n16258);
   U12412 : INV_X1 port map( A => n16257, ZN => n10555);
   U12413 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1784_port, B2 => n2839, 
                           ZN => n16257);
   U12414 : INV_X1 port map( A => n16256, ZN => n10556);
   U12415 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1783_port, B2 => n2838, 
                           ZN => n16256);
   U12416 : INV_X1 port map( A => n16255, ZN => n10557);
   U12417 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1782_port, B2 => n2838, 
                           ZN => n16255);
   U12418 : INV_X1 port map( A => n16254, ZN => n10558);
   U12419 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1781_port, B2 => n2838, 
                           ZN => n16254);
   U12420 : INV_X1 port map( A => n16253, ZN => n10559);
   U12421 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2834, B1 => 
                           DataPath_RF_bus_reg_dataout_1780_port, B2 => n2838, 
                           ZN => n16253);
   U12422 : INV_X1 port map( A => n16252, ZN => n10560);
   U12423 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1779_port, B2 => n2838, 
                           ZN => n16252);
   U12424 : INV_X1 port map( A => n16251, ZN => n10561);
   U12425 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1778_port, B2 => n2838, 
                           ZN => n16251);
   U12426 : INV_X1 port map( A => n16250, ZN => n10562);
   U12427 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1777_port, B2 => n2838, 
                           ZN => n16250);
   U12428 : INV_X1 port map( A => n16249, ZN => n10563);
   U12429 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1776_port, B2 => n2838, 
                           ZN => n16249);
   U12430 : INV_X1 port map( A => n16248, ZN => n10564);
   U12431 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1775_port, B2 => n2838, 
                           ZN => n16248);
   U12432 : INV_X1 port map( A => n16247, ZN => n10565);
   U12433 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1774_port, B2 => n2838, 
                           ZN => n16247);
   U12434 : INV_X1 port map( A => n16246, ZN => n10566);
   U12435 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1773_port, B2 => n2838, 
                           ZN => n16246);
   U12436 : INV_X1 port map( A => n16245, ZN => n10567);
   U12437 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1772_port, B2 => n2838, 
                           ZN => n16245);
   U12438 : INV_X1 port map( A => n16244, ZN => n10568);
   U12439 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1771_port, B2 => n2837, 
                           ZN => n16244);
   U12440 : INV_X1 port map( A => n16243, ZN => n10569);
   U12441 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1770_port, B2 => n2837, 
                           ZN => n16243);
   U12442 : INV_X1 port map( A => n16242, ZN => n10570);
   U12443 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1769_port, B2 => n2837, 
                           ZN => n16242);
   U12444 : INV_X1 port map( A => n16241, ZN => n10571);
   U12445 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2835, B1 => 
                           DataPath_RF_bus_reg_dataout_1768_port, B2 => n2837, 
                           ZN => n16241);
   U12446 : INV_X1 port map( A => n16240, ZN => n10572);
   U12447 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1767_port, B2 => n2837, 
                           ZN => n16240);
   U12448 : INV_X1 port map( A => n16239, ZN => n10573);
   U12449 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1766_port, B2 => n2837, 
                           ZN => n16239);
   U12450 : INV_X1 port map( A => n16238, ZN => n10574);
   U12451 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1765_port, B2 => n2837, 
                           ZN => n16238);
   U12452 : INV_X1 port map( A => n16237, ZN => n10575);
   U12453 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1764_port, B2 => n2837, 
                           ZN => n16237);
   U12454 : INV_X1 port map( A => n16236, ZN => n10576);
   U12455 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1763_port, B2 => n2837, 
                           ZN => n16236);
   U12456 : INV_X1 port map( A => n16235, ZN => n10577);
   U12457 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1762_port, B2 => n2837, 
                           ZN => n16235);
   U12458 : INV_X1 port map( A => n16234, ZN => n10578);
   U12459 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1761_port, B2 => n2837, 
                           ZN => n16234);
   U12460 : INV_X1 port map( A => n16231, ZN => n10579);
   U12461 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2836, B1 => 
                           DataPath_RF_bus_reg_dataout_1760_port, B2 => n2837, 
                           ZN => n16231);
   U12462 : INV_X1 port map( A => n16298, ZN => n10580);
   U12463 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1823_port, B2 => n2845, 
                           ZN => n16298);
   U12464 : INV_X1 port map( A => n16297, ZN => n10581);
   U12465 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1822_port, B2 => n2845, 
                           ZN => n16297);
   U12466 : INV_X1 port map( A => n16296, ZN => n10582);
   U12467 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1821_port, B2 => n2845, 
                           ZN => n16296);
   U12468 : INV_X1 port map( A => n16295, ZN => n10583);
   U12469 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1820_port, B2 => n2845, 
                           ZN => n16295);
   U12470 : INV_X1 port map( A => n16294, ZN => n10584);
   U12471 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1819_port, B2 => n2845, 
                           ZN => n16294);
   U12472 : INV_X1 port map( A => n16293, ZN => n10585);
   U12473 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1818_port, B2 => n2845, 
                           ZN => n16293);
   U12474 : INV_X1 port map( A => n16292, ZN => n10586);
   U12475 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1817_port, B2 => n2845, 
                           ZN => n16292);
   U12476 : INV_X1 port map( A => n16291, ZN => n10587);
   U12477 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1816_port, B2 => n2845, 
                           ZN => n16291);
   U12478 : INV_X1 port map( A => n16290, ZN => n10588);
   U12479 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1815_port, B2 => n2844, 
                           ZN => n16290);
   U12480 : INV_X1 port map( A => n16289, ZN => n10589);
   U12481 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1814_port, B2 => n2844, 
                           ZN => n16289);
   U12482 : INV_X1 port map( A => n16288, ZN => n10590);
   U12483 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1813_port, B2 => n2844, 
                           ZN => n16288);
   U12484 : INV_X1 port map( A => n16287, ZN => n10591);
   U12485 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2840, B1 => 
                           DataPath_RF_bus_reg_dataout_1812_port, B2 => n2844, 
                           ZN => n16287);
   U12486 : INV_X1 port map( A => n16286, ZN => n10592);
   U12487 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1811_port, B2 => n2844, 
                           ZN => n16286);
   U12488 : INV_X1 port map( A => n16285, ZN => n10593);
   U12489 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1810_port, B2 => n2844, 
                           ZN => n16285);
   U12490 : INV_X1 port map( A => n16284, ZN => n10594);
   U12491 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1809_port, B2 => n2844, 
                           ZN => n16284);
   U12492 : INV_X1 port map( A => n16283, ZN => n10595);
   U12493 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1808_port, B2 => n2844, 
                           ZN => n16283);
   U12494 : INV_X1 port map( A => n16282, ZN => n10596);
   U12495 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1807_port, B2 => n2844, 
                           ZN => n16282);
   U12496 : INV_X1 port map( A => n16281, ZN => n10597);
   U12497 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1806_port, B2 => n2844, 
                           ZN => n16281);
   U12498 : INV_X1 port map( A => n16280, ZN => n10598);
   U12499 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1805_port, B2 => n2844, 
                           ZN => n16280);
   U12500 : INV_X1 port map( A => n16279, ZN => n10599);
   U12501 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1804_port, B2 => n2844, 
                           ZN => n16279);
   U12502 : INV_X1 port map( A => n16278, ZN => n10600);
   U12503 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1803_port, B2 => n2843, 
                           ZN => n16278);
   U12504 : INV_X1 port map( A => n16277, ZN => n10601);
   U12505 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1802_port, B2 => n2843, 
                           ZN => n16277);
   U12506 : INV_X1 port map( A => n16276, ZN => n10602);
   U12507 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1801_port, B2 => n2843, 
                           ZN => n16276);
   U12508 : INV_X1 port map( A => n16275, ZN => n10603);
   U12509 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2841, B1 => 
                           DataPath_RF_bus_reg_dataout_1800_port, B2 => n2843, 
                           ZN => n16275);
   U12510 : INV_X1 port map( A => n16274, ZN => n10604);
   U12511 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1799_port, B2 => n2843, 
                           ZN => n16274);
   U12512 : INV_X1 port map( A => n16273, ZN => n10605);
   U12513 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1798_port, B2 => n2843, 
                           ZN => n16273);
   U12514 : INV_X1 port map( A => n16272, ZN => n10606);
   U12515 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1797_port, B2 => n2843, 
                           ZN => n16272);
   U12516 : INV_X1 port map( A => n16271, ZN => n10607);
   U12517 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1796_port, B2 => n2843, 
                           ZN => n16271);
   U12518 : INV_X1 port map( A => n16270, ZN => n10608);
   U12519 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1795_port, B2 => n2843, 
                           ZN => n16270);
   U12520 : INV_X1 port map( A => n16269, ZN => n10609);
   U12521 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1794_port, B2 => n2843, 
                           ZN => n16269);
   U12522 : INV_X1 port map( A => n16268, ZN => n10610);
   U12523 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1793_port, B2 => n2843, 
                           ZN => n16268);
   U12524 : INV_X1 port map( A => n16265, ZN => n10611);
   U12525 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2842, B1 => 
                           DataPath_RF_bus_reg_dataout_1792_port, B2 => n2843, 
                           ZN => n16265);
   U12526 : INV_X1 port map( A => n16332, ZN => n10612);
   U12527 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1855_port, B2 => n2851, 
                           ZN => n16332);
   U12528 : INV_X1 port map( A => n16331, ZN => n10613);
   U12529 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1854_port, B2 => n2851, 
                           ZN => n16331);
   U12530 : INV_X1 port map( A => n16330, ZN => n10614);
   U12531 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1853_port, B2 => n2851, 
                           ZN => n16330);
   U12532 : INV_X1 port map( A => n16329, ZN => n10615);
   U12533 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1852_port, B2 => n2851, 
                           ZN => n16329);
   U12534 : INV_X1 port map( A => n16328, ZN => n10616);
   U12535 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1851_port, B2 => n2851, 
                           ZN => n16328);
   U12536 : INV_X1 port map( A => n16327, ZN => n10617);
   U12537 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1850_port, B2 => n2851, 
                           ZN => n16327);
   U12538 : INV_X1 port map( A => n16326, ZN => n10618);
   U12539 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1849_port, B2 => n2851, 
                           ZN => n16326);
   U12540 : INV_X1 port map( A => n16325, ZN => n10619);
   U12541 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1848_port, B2 => n2851, 
                           ZN => n16325);
   U12542 : INV_X1 port map( A => n16324, ZN => n10620);
   U12543 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1847_port, B2 => n2850, 
                           ZN => n16324);
   U12544 : INV_X1 port map( A => n16323, ZN => n10621);
   U12545 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1846_port, B2 => n2850, 
                           ZN => n16323);
   U12546 : INV_X1 port map( A => n16322, ZN => n10622);
   U12547 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1845_port, B2 => n2850, 
                           ZN => n16322);
   U12548 : INV_X1 port map( A => n16321, ZN => n10623);
   U12549 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2846, B1 => 
                           DataPath_RF_bus_reg_dataout_1844_port, B2 => n2850, 
                           ZN => n16321);
   U12550 : INV_X1 port map( A => n16320, ZN => n10624);
   U12551 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1843_port, B2 => n2850, 
                           ZN => n16320);
   U12552 : INV_X1 port map( A => n16319, ZN => n10625);
   U12553 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1842_port, B2 => n2850, 
                           ZN => n16319);
   U12554 : INV_X1 port map( A => n16318, ZN => n10626);
   U12555 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1841_port, B2 => n2850, 
                           ZN => n16318);
   U12556 : INV_X1 port map( A => n16317, ZN => n10627);
   U12557 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1840_port, B2 => n2850, 
                           ZN => n16317);
   U12558 : INV_X1 port map( A => n16316, ZN => n10628);
   U12559 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1839_port, B2 => n2850, 
                           ZN => n16316);
   U12560 : INV_X1 port map( A => n16315, ZN => n10629);
   U12561 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1838_port, B2 => n2850, 
                           ZN => n16315);
   U12562 : INV_X1 port map( A => n16314, ZN => n10630);
   U12563 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1837_port, B2 => n2850, 
                           ZN => n16314);
   U12564 : INV_X1 port map( A => n16313, ZN => n10631);
   U12565 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1836_port, B2 => n2850, 
                           ZN => n16313);
   U12566 : INV_X1 port map( A => n16312, ZN => n10632);
   U12567 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1835_port, B2 => n2849, 
                           ZN => n16312);
   U12568 : INV_X1 port map( A => n16311, ZN => n10633);
   U12569 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1834_port, B2 => n2849, 
                           ZN => n16311);
   U12570 : INV_X1 port map( A => n16310, ZN => n10634);
   U12571 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1833_port, B2 => n2849, 
                           ZN => n16310);
   U12572 : INV_X1 port map( A => n16309, ZN => n10635);
   U12573 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2847, B1 => 
                           DataPath_RF_bus_reg_dataout_1832_port, B2 => n2849, 
                           ZN => n16309);
   U12574 : INV_X1 port map( A => n16308, ZN => n10636);
   U12575 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1831_port, B2 => n2849, 
                           ZN => n16308);
   U12576 : INV_X1 port map( A => n16307, ZN => n10637);
   U12577 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1830_port, B2 => n2849, 
                           ZN => n16307);
   U12578 : INV_X1 port map( A => n16306, ZN => n10638);
   U12579 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1829_port, B2 => n2849, 
                           ZN => n16306);
   U12580 : INV_X1 port map( A => n16305, ZN => n10639);
   U12581 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1828_port, B2 => n2849, 
                           ZN => n16305);
   U12582 : INV_X1 port map( A => n16304, ZN => n10640);
   U12583 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1827_port, B2 => n2849, 
                           ZN => n16304);
   U12584 : INV_X1 port map( A => n16303, ZN => n10641);
   U12585 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1826_port, B2 => n2849, 
                           ZN => n16303);
   U12586 : INV_X1 port map( A => n16302, ZN => n10642);
   U12587 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1825_port, B2 => n2849, 
                           ZN => n16302);
   U12588 : INV_X1 port map( A => n16299, ZN => n10643);
   U12589 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2848, B1 => 
                           DataPath_RF_bus_reg_dataout_1824_port, B2 => n2849, 
                           ZN => n16299);
   U12590 : INV_X1 port map( A => n16366, ZN => n10644);
   U12591 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1887_port, B2 => n2857, 
                           ZN => n16366);
   U12592 : INV_X1 port map( A => n16365, ZN => n10645);
   U12593 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1886_port, B2 => n2857, 
                           ZN => n16365);
   U12594 : INV_X1 port map( A => n16364, ZN => n10646);
   U12595 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1885_port, B2 => n2857, 
                           ZN => n16364);
   U12596 : INV_X1 port map( A => n16363, ZN => n10647);
   U12597 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1884_port, B2 => n2857, 
                           ZN => n16363);
   U12598 : INV_X1 port map( A => n16362, ZN => n10648);
   U12599 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1883_port, B2 => n2857, 
                           ZN => n16362);
   U12600 : INV_X1 port map( A => n16361, ZN => n10649);
   U12601 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1882_port, B2 => n2857, 
                           ZN => n16361);
   U12602 : INV_X1 port map( A => n16360, ZN => n10650);
   U12603 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1881_port, B2 => n2857, 
                           ZN => n16360);
   U12604 : INV_X1 port map( A => n16359, ZN => n10651);
   U12605 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1880_port, B2 => n2857, 
                           ZN => n16359);
   U12606 : INV_X1 port map( A => n16358, ZN => n10652);
   U12607 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1879_port, B2 => n2856, 
                           ZN => n16358);
   U12608 : INV_X1 port map( A => n16357, ZN => n10653);
   U12609 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1878_port, B2 => n2856, 
                           ZN => n16357);
   U12610 : INV_X1 port map( A => n16356, ZN => n10654);
   U12611 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1877_port, B2 => n2856, 
                           ZN => n16356);
   U12612 : INV_X1 port map( A => n16355, ZN => n10655);
   U12613 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2852, B1 => 
                           DataPath_RF_bus_reg_dataout_1876_port, B2 => n2856, 
                           ZN => n16355);
   U12614 : INV_X1 port map( A => n16354, ZN => n10656);
   U12615 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1875_port, B2 => n2856, 
                           ZN => n16354);
   U12616 : INV_X1 port map( A => n16353, ZN => n10657);
   U12617 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1874_port, B2 => n2856, 
                           ZN => n16353);
   U12618 : INV_X1 port map( A => n16352, ZN => n10658);
   U12619 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1873_port, B2 => n2856, 
                           ZN => n16352);
   U12620 : INV_X1 port map( A => n16351, ZN => n10659);
   U12621 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1872_port, B2 => n2856, 
                           ZN => n16351);
   U12622 : INV_X1 port map( A => n16350, ZN => n10660);
   U12623 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1871_port, B2 => n2856, 
                           ZN => n16350);
   U12624 : INV_X1 port map( A => n16349, ZN => n10661);
   U12625 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1870_port, B2 => n2856, 
                           ZN => n16349);
   U12626 : INV_X1 port map( A => n16348, ZN => n10662);
   U12627 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1869_port, B2 => n2856, 
                           ZN => n16348);
   U12628 : INV_X1 port map( A => n16347, ZN => n10663);
   U12629 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1868_port, B2 => n2856, 
                           ZN => n16347);
   U12630 : INV_X1 port map( A => n16346, ZN => n10664);
   U12631 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1867_port, B2 => n2855, 
                           ZN => n16346);
   U12632 : INV_X1 port map( A => n16345, ZN => n10665);
   U12633 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1866_port, B2 => n2855, 
                           ZN => n16345);
   U12634 : INV_X1 port map( A => n16344, ZN => n10666);
   U12635 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1865_port, B2 => n2855, 
                           ZN => n16344);
   U12636 : INV_X1 port map( A => n16343, ZN => n10667);
   U12637 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2853, B1 => 
                           DataPath_RF_bus_reg_dataout_1864_port, B2 => n2855, 
                           ZN => n16343);
   U12638 : INV_X1 port map( A => n16342, ZN => n10668);
   U12639 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1863_port, B2 => n2855, 
                           ZN => n16342);
   U12640 : INV_X1 port map( A => n16341, ZN => n10669);
   U12641 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1862_port, B2 => n2855, 
                           ZN => n16341);
   U12642 : INV_X1 port map( A => n16340, ZN => n10670);
   U12643 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1861_port, B2 => n2855, 
                           ZN => n16340);
   U12644 : INV_X1 port map( A => n16339, ZN => n10671);
   U12645 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1860_port, B2 => n2855, 
                           ZN => n16339);
   U12646 : INV_X1 port map( A => n16338, ZN => n10672);
   U12647 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1859_port, B2 => n2855, 
                           ZN => n16338);
   U12648 : INV_X1 port map( A => n16337, ZN => n10673);
   U12649 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1858_port, B2 => n2855, 
                           ZN => n16337);
   U12650 : INV_X1 port map( A => n16336, ZN => n10674);
   U12651 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1857_port, B2 => n2855, 
                           ZN => n16336);
   U12652 : INV_X1 port map( A => n16333, ZN => n10675);
   U12653 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2854, B1 => 
                           DataPath_RF_bus_reg_dataout_1856_port, B2 => n2855, 
                           ZN => n16333);
   U12654 : INV_X1 port map( A => n16400, ZN => n10676);
   U12655 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1919_port, B2 => n2863, 
                           ZN => n16400);
   U12656 : INV_X1 port map( A => n16399, ZN => n10677);
   U12657 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1918_port, B2 => n2863, 
                           ZN => n16399);
   U12658 : INV_X1 port map( A => n16398, ZN => n10678);
   U12659 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1917_port, B2 => n2863, 
                           ZN => n16398);
   U12660 : INV_X1 port map( A => n16397, ZN => n10679);
   U12661 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1916_port, B2 => n2863, 
                           ZN => n16397);
   U12662 : INV_X1 port map( A => n16396, ZN => n10680);
   U12663 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1915_port, B2 => n2863, 
                           ZN => n16396);
   U12664 : INV_X1 port map( A => n16395, ZN => n10681);
   U12665 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1914_port, B2 => n2863, 
                           ZN => n16395);
   U12666 : INV_X1 port map( A => n16394, ZN => n10682);
   U12667 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1913_port, B2 => n2863, 
                           ZN => n16394);
   U12668 : INV_X1 port map( A => n16393, ZN => n10683);
   U12669 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1912_port, B2 => n2863, 
                           ZN => n16393);
   U12670 : INV_X1 port map( A => n16392, ZN => n10684);
   U12671 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1911_port, B2 => n2862, 
                           ZN => n16392);
   U12672 : INV_X1 port map( A => n16391, ZN => n10685);
   U12673 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1910_port, B2 => n2862, 
                           ZN => n16391);
   U12674 : INV_X1 port map( A => n16390, ZN => n10686);
   U12675 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1909_port, B2 => n2862, 
                           ZN => n16390);
   U12676 : INV_X1 port map( A => n16389, ZN => n10687);
   U12677 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2858, B1 => 
                           DataPath_RF_bus_reg_dataout_1908_port, B2 => n2862, 
                           ZN => n16389);
   U12678 : INV_X1 port map( A => n16388, ZN => n10688);
   U12679 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1907_port, B2 => n2862, 
                           ZN => n16388);
   U12680 : INV_X1 port map( A => n16387, ZN => n10689);
   U12681 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1906_port, B2 => n2862, 
                           ZN => n16387);
   U12682 : INV_X1 port map( A => n16386, ZN => n10690);
   U12683 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1905_port, B2 => n2862, 
                           ZN => n16386);
   U12684 : INV_X1 port map( A => n16385, ZN => n10691);
   U12685 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1904_port, B2 => n2862, 
                           ZN => n16385);
   U12686 : INV_X1 port map( A => n16384, ZN => n10692);
   U12687 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1903_port, B2 => n2862, 
                           ZN => n16384);
   U12688 : INV_X1 port map( A => n16383, ZN => n10693);
   U12689 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1902_port, B2 => n2862, 
                           ZN => n16383);
   U12690 : INV_X1 port map( A => n16382, ZN => n10694);
   U12691 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1901_port, B2 => n2862, 
                           ZN => n16382);
   U12692 : INV_X1 port map( A => n16381, ZN => n10695);
   U12693 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1900_port, B2 => n2862, 
                           ZN => n16381);
   U12694 : INV_X1 port map( A => n16380, ZN => n10696);
   U12695 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1899_port, B2 => n2861, 
                           ZN => n16380);
   U12696 : INV_X1 port map( A => n16379, ZN => n10697);
   U12697 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1898_port, B2 => n2861, 
                           ZN => n16379);
   U12698 : INV_X1 port map( A => n16378, ZN => n10698);
   U12699 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1897_port, B2 => n2861, 
                           ZN => n16378);
   U12700 : INV_X1 port map( A => n16377, ZN => n10699);
   U12701 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2859, B1 => 
                           DataPath_RF_bus_reg_dataout_1896_port, B2 => n2861, 
                           ZN => n16377);
   U12702 : INV_X1 port map( A => n16376, ZN => n10700);
   U12703 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1895_port, B2 => n2861, 
                           ZN => n16376);
   U12704 : INV_X1 port map( A => n16375, ZN => n10701);
   U12705 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1894_port, B2 => n2861, 
                           ZN => n16375);
   U12706 : INV_X1 port map( A => n16374, ZN => n10702);
   U12707 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1893_port, B2 => n2861, 
                           ZN => n16374);
   U12708 : INV_X1 port map( A => n16373, ZN => n10703);
   U12709 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1892_port, B2 => n2861, 
                           ZN => n16373);
   U12710 : INV_X1 port map( A => n16372, ZN => n10704);
   U12711 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1891_port, B2 => n2861, 
                           ZN => n16372);
   U12712 : INV_X1 port map( A => n16371, ZN => n10705);
   U12713 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1890_port, B2 => n2861, 
                           ZN => n16371);
   U12714 : INV_X1 port map( A => n16370, ZN => n10706);
   U12715 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1889_port, B2 => n2861, 
                           ZN => n16370);
   U12716 : INV_X1 port map( A => n16367, ZN => n10707);
   U12717 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2860, B1 => 
                           DataPath_RF_bus_reg_dataout_1888_port, B2 => n2861, 
                           ZN => n16367);
   U12718 : INV_X1 port map( A => n16434, ZN => n10708);
   U12719 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1951_port, B2 => n2869, 
                           ZN => n16434);
   U12720 : INV_X1 port map( A => n16433, ZN => n10709);
   U12721 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1950_port, B2 => n2869, 
                           ZN => n16433);
   U12722 : INV_X1 port map( A => n16432, ZN => n10710);
   U12723 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1949_port, B2 => n2869, 
                           ZN => n16432);
   U12724 : INV_X1 port map( A => n16431, ZN => n10711);
   U12725 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1948_port, B2 => n2869, 
                           ZN => n16431);
   U12726 : INV_X1 port map( A => n16430, ZN => n10712);
   U12727 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1947_port, B2 => n2869, 
                           ZN => n16430);
   U12728 : INV_X1 port map( A => n16429, ZN => n10713);
   U12729 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1946_port, B2 => n2869, 
                           ZN => n16429);
   U12730 : INV_X1 port map( A => n16428, ZN => n10714);
   U12731 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1945_port, B2 => n2869, 
                           ZN => n16428);
   U12732 : INV_X1 port map( A => n16427, ZN => n10715);
   U12733 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1944_port, B2 => n2869, 
                           ZN => n16427);
   U12734 : INV_X1 port map( A => n16426, ZN => n10716);
   U12735 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1943_port, B2 => n2868, 
                           ZN => n16426);
   U12736 : INV_X1 port map( A => n16425, ZN => n10717);
   U12737 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1942_port, B2 => n2868, 
                           ZN => n16425);
   U12738 : INV_X1 port map( A => n16424, ZN => n10718);
   U12739 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1941_port, B2 => n2868, 
                           ZN => n16424);
   U12740 : INV_X1 port map( A => n16423, ZN => n10719);
   U12741 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2864, B1 => 
                           DataPath_RF_bus_reg_dataout_1940_port, B2 => n2868, 
                           ZN => n16423);
   U12742 : INV_X1 port map( A => n16422, ZN => n10720);
   U12743 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1939_port, B2 => n2868, 
                           ZN => n16422);
   U12744 : INV_X1 port map( A => n16421, ZN => n10721);
   U12745 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1938_port, B2 => n2868, 
                           ZN => n16421);
   U12746 : INV_X1 port map( A => n16420, ZN => n10722);
   U12747 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1937_port, B2 => n2868, 
                           ZN => n16420);
   U12748 : INV_X1 port map( A => n16419, ZN => n10723);
   U12749 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1936_port, B2 => n2868, 
                           ZN => n16419);
   U12750 : INV_X1 port map( A => n16418, ZN => n10724);
   U12751 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1935_port, B2 => n2868, 
                           ZN => n16418);
   U12752 : INV_X1 port map( A => n16417, ZN => n10725);
   U12753 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1934_port, B2 => n2868, 
                           ZN => n16417);
   U12754 : INV_X1 port map( A => n16416, ZN => n10726);
   U12755 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1933_port, B2 => n2868, 
                           ZN => n16416);
   U12756 : INV_X1 port map( A => n16415, ZN => n10727);
   U12757 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1932_port, B2 => n2868, 
                           ZN => n16415);
   U12758 : INV_X1 port map( A => n16414, ZN => n10728);
   U12759 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1931_port, B2 => n2867, 
                           ZN => n16414);
   U12760 : INV_X1 port map( A => n16413, ZN => n10729);
   U12761 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1930_port, B2 => n2867, 
                           ZN => n16413);
   U12762 : INV_X1 port map( A => n16412, ZN => n10730);
   U12763 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1929_port, B2 => n2867, 
                           ZN => n16412);
   U12764 : INV_X1 port map( A => n16411, ZN => n10731);
   U12765 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2865, B1 => 
                           DataPath_RF_bus_reg_dataout_1928_port, B2 => n2867, 
                           ZN => n16411);
   U12766 : INV_X1 port map( A => n16410, ZN => n10732);
   U12767 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1927_port, B2 => n2867, 
                           ZN => n16410);
   U12768 : INV_X1 port map( A => n16409, ZN => n10733);
   U12769 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1926_port, B2 => n2867, 
                           ZN => n16409);
   U12770 : INV_X1 port map( A => n16408, ZN => n10734);
   U12771 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1925_port, B2 => n2867, 
                           ZN => n16408);
   U12772 : INV_X1 port map( A => n16407, ZN => n10735);
   U12773 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1924_port, B2 => n2867, 
                           ZN => n16407);
   U12774 : INV_X1 port map( A => n16406, ZN => n10736);
   U12775 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1923_port, B2 => n2867, 
                           ZN => n16406);
   U12776 : INV_X1 port map( A => n16405, ZN => n10737);
   U12777 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1922_port, B2 => n2867, 
                           ZN => n16405);
   U12778 : INV_X1 port map( A => n16404, ZN => n10738);
   U12779 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1921_port, B2 => n2867, 
                           ZN => n16404);
   U12780 : INV_X1 port map( A => n16401, ZN => n10739);
   U12781 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2866, B1 => 
                           DataPath_RF_bus_reg_dataout_1920_port, B2 => n2867, 
                           ZN => n16401);
   U12782 : INV_X1 port map( A => n16468, ZN => n10740);
   U12783 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1983_port, B2 => n2875, 
                           ZN => n16468);
   U12784 : INV_X1 port map( A => n16467, ZN => n10741);
   U12785 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1982_port, B2 => n2875, 
                           ZN => n16467);
   U12786 : INV_X1 port map( A => n16466, ZN => n10742);
   U12787 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1981_port, B2 => n2875, 
                           ZN => n16466);
   U12788 : INV_X1 port map( A => n16465, ZN => n10743);
   U12789 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1980_port, B2 => n2875, 
                           ZN => n16465);
   U12790 : INV_X1 port map( A => n16464, ZN => n10744);
   U12791 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1979_port, B2 => n2875, 
                           ZN => n16464);
   U12792 : INV_X1 port map( A => n16463, ZN => n10745);
   U12793 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1978_port, B2 => n2875, 
                           ZN => n16463);
   U12794 : INV_X1 port map( A => n16462, ZN => n10746);
   U12795 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1977_port, B2 => n2875, 
                           ZN => n16462);
   U12796 : INV_X1 port map( A => n16461, ZN => n10747);
   U12797 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1976_port, B2 => n2875, 
                           ZN => n16461);
   U12798 : INV_X1 port map( A => n16460, ZN => n10748);
   U12799 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1975_port, B2 => n2874, 
                           ZN => n16460);
   U12800 : INV_X1 port map( A => n16459, ZN => n10749);
   U12801 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1974_port, B2 => n2874, 
                           ZN => n16459);
   U12802 : INV_X1 port map( A => n16458, ZN => n10750);
   U12803 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1973_port, B2 => n2874, 
                           ZN => n16458);
   U12804 : INV_X1 port map( A => n16457, ZN => n10751);
   U12805 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2870, B1 => 
                           DataPath_RF_bus_reg_dataout_1972_port, B2 => n2874, 
                           ZN => n16457);
   U12806 : INV_X1 port map( A => n16456, ZN => n10752);
   U12807 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1971_port, B2 => n2874, 
                           ZN => n16456);
   U12808 : INV_X1 port map( A => n16455, ZN => n10753);
   U12809 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1970_port, B2 => n2874, 
                           ZN => n16455);
   U12810 : INV_X1 port map( A => n16454, ZN => n10754);
   U12811 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1969_port, B2 => n2874, 
                           ZN => n16454);
   U12812 : INV_X1 port map( A => n16453, ZN => n10755);
   U12813 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1968_port, B2 => n2874, 
                           ZN => n16453);
   U12814 : INV_X1 port map( A => n16452, ZN => n10756);
   U12815 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1967_port, B2 => n2874, 
                           ZN => n16452);
   U12816 : INV_X1 port map( A => n16451, ZN => n10757);
   U12817 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1966_port, B2 => n2874, 
                           ZN => n16451);
   U12818 : INV_X1 port map( A => n16450, ZN => n10758);
   U12819 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1965_port, B2 => n2874, 
                           ZN => n16450);
   U12820 : INV_X1 port map( A => n16449, ZN => n10759);
   U12821 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1964_port, B2 => n2874, 
                           ZN => n16449);
   U12822 : INV_X1 port map( A => n16448, ZN => n10760);
   U12823 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1963_port, B2 => n2873, 
                           ZN => n16448);
   U12824 : INV_X1 port map( A => n16447, ZN => n10761);
   U12825 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1962_port, B2 => n2873, 
                           ZN => n16447);
   U12826 : INV_X1 port map( A => n16446, ZN => n10762);
   U12827 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1961_port, B2 => n2873, 
                           ZN => n16446);
   U12828 : INV_X1 port map( A => n16445, ZN => n10763);
   U12829 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2871, B1 => 
                           DataPath_RF_bus_reg_dataout_1960_port, B2 => n2873, 
                           ZN => n16445);
   U12830 : INV_X1 port map( A => n16444, ZN => n10764);
   U12831 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1959_port, B2 => n2873, 
                           ZN => n16444);
   U12832 : INV_X1 port map( A => n16443, ZN => n10765);
   U12833 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1958_port, B2 => n2873, 
                           ZN => n16443);
   U12834 : INV_X1 port map( A => n16442, ZN => n10766);
   U12835 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1957_port, B2 => n2873, 
                           ZN => n16442);
   U12836 : INV_X1 port map( A => n16441, ZN => n10767);
   U12837 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1956_port, B2 => n2873, 
                           ZN => n16441);
   U12838 : INV_X1 port map( A => n16440, ZN => n10768);
   U12839 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1955_port, B2 => n2873, 
                           ZN => n16440);
   U12840 : INV_X1 port map( A => n16439, ZN => n10769);
   U12841 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1954_port, B2 => n2873, 
                           ZN => n16439);
   U12842 : INV_X1 port map( A => n16438, ZN => n10770);
   U12843 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1953_port, B2 => n2873, 
                           ZN => n16438);
   U12844 : INV_X1 port map( A => n16435, ZN => n10771);
   U12845 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2872, B1 => 
                           DataPath_RF_bus_reg_dataout_1952_port, B2 => n2873, 
                           ZN => n16435);
   U12846 : INV_X1 port map( A => n16502, ZN => n10772);
   U12847 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2015_port, B2 => n2881, 
                           ZN => n16502);
   U12848 : INV_X1 port map( A => n16501, ZN => n10773);
   U12849 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2014_port, B2 => n2881, 
                           ZN => n16501);
   U12850 : INV_X1 port map( A => n16500, ZN => n10774);
   U12851 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2013_port, B2 => n2881, 
                           ZN => n16500);
   U12852 : INV_X1 port map( A => n16499, ZN => n10775);
   U12853 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2012_port, B2 => n2881, 
                           ZN => n16499);
   U12854 : INV_X1 port map( A => n16498, ZN => n10776);
   U12855 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2011_port, B2 => n2881, 
                           ZN => n16498);
   U12856 : INV_X1 port map( A => n16497, ZN => n10777);
   U12857 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2010_port, B2 => n2881, 
                           ZN => n16497);
   U12858 : INV_X1 port map( A => n16496, ZN => n10778);
   U12859 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2009_port, B2 => n2881, 
                           ZN => n16496);
   U12860 : INV_X1 port map( A => n16495, ZN => n10779);
   U12861 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2008_port, B2 => n2881, 
                           ZN => n16495);
   U12862 : INV_X1 port map( A => n16494, ZN => n10780);
   U12863 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2007_port, B2 => n2880, 
                           ZN => n16494);
   U12864 : INV_X1 port map( A => n16493, ZN => n10781);
   U12865 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2006_port, B2 => n2880, 
                           ZN => n16493);
   U12866 : INV_X1 port map( A => n16492, ZN => n10782);
   U12867 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2005_port, B2 => n2880, 
                           ZN => n16492);
   U12868 : INV_X1 port map( A => n16491, ZN => n10783);
   U12869 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2876, B1 => 
                           DataPath_RF_bus_reg_dataout_2004_port, B2 => n2880, 
                           ZN => n16491);
   U12870 : INV_X1 port map( A => n16490, ZN => n10784);
   U12871 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_2003_port, B2 => n2880, 
                           ZN => n16490);
   U12872 : INV_X1 port map( A => n16489, ZN => n10785);
   U12873 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_2002_port, B2 => n2880, 
                           ZN => n16489);
   U12874 : INV_X1 port map( A => n16488, ZN => n10786);
   U12875 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_2001_port, B2 => n2880, 
                           ZN => n16488);
   U12876 : INV_X1 port map( A => n16487, ZN => n10787);
   U12877 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_2000_port, B2 => n2880, 
                           ZN => n16487);
   U12878 : INV_X1 port map( A => n16486, ZN => n10788);
   U12879 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1999_port, B2 => n2880, 
                           ZN => n16486);
   U12880 : INV_X1 port map( A => n16485, ZN => n10789);
   U12881 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1998_port, B2 => n2880, 
                           ZN => n16485);
   U12882 : INV_X1 port map( A => n16484, ZN => n10790);
   U12883 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1997_port, B2 => n2880, 
                           ZN => n16484);
   U12884 : INV_X1 port map( A => n16483, ZN => n10791);
   U12885 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1996_port, B2 => n2880, 
                           ZN => n16483);
   U12886 : INV_X1 port map( A => n16482, ZN => n10792);
   U12887 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1995_port, B2 => n2879, 
                           ZN => n16482);
   U12888 : INV_X1 port map( A => n16481, ZN => n10793);
   U12889 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1994_port, B2 => n2879, 
                           ZN => n16481);
   U12890 : INV_X1 port map( A => n16480, ZN => n10794);
   U12891 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1993_port, B2 => n2879, 
                           ZN => n16480);
   U12892 : INV_X1 port map( A => n16479, ZN => n10795);
   U12893 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2877, B1 => 
                           DataPath_RF_bus_reg_dataout_1992_port, B2 => n2879, 
                           ZN => n16479);
   U12894 : INV_X1 port map( A => n16478, ZN => n10796);
   U12895 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1991_port, B2 => n2879, 
                           ZN => n16478);
   U12896 : INV_X1 port map( A => n16477, ZN => n10797);
   U12897 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1990_port, B2 => n2879, 
                           ZN => n16477);
   U12898 : INV_X1 port map( A => n16476, ZN => n10798);
   U12899 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1989_port, B2 => n2879, 
                           ZN => n16476);
   U12900 : INV_X1 port map( A => n16475, ZN => n10799);
   U12901 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1988_port, B2 => n2879, 
                           ZN => n16475);
   U12902 : INV_X1 port map( A => n16474, ZN => n10800);
   U12903 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1987_port, B2 => n2879, 
                           ZN => n16474);
   U12904 : INV_X1 port map( A => n16473, ZN => n10801);
   U12905 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1986_port, B2 => n2879, 
                           ZN => n16473);
   U12906 : INV_X1 port map( A => n16472, ZN => n10802);
   U12907 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1985_port, B2 => n2879, 
                           ZN => n16472);
   U12908 : INV_X1 port map( A => n16469, ZN => n10803);
   U12909 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2878, B1 => 
                           DataPath_RF_bus_reg_dataout_1984_port, B2 => n2879, 
                           ZN => n16469);
   U12910 : INV_X1 port map( A => n16536, ZN => n10804);
   U12911 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_31_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2047_port, B2 => n2887, 
                           ZN => n16536);
   U12912 : INV_X1 port map( A => n16535, ZN => n10805);
   U12913 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_30_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2046_port, B2 => n2887, 
                           ZN => n16535);
   U12914 : INV_X1 port map( A => n16534, ZN => n10806);
   U12915 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_29_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2045_port, B2 => n2887, 
                           ZN => n16534);
   U12916 : INV_X1 port map( A => n16533, ZN => n10807);
   U12917 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_28_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2044_port, B2 => n2887, 
                           ZN => n16533);
   U12918 : INV_X1 port map( A => n16532, ZN => n10808);
   U12919 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_27_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2043_port, B2 => n2887, 
                           ZN => n16532);
   U12920 : INV_X1 port map( A => n16531, ZN => n10809);
   U12921 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_26_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2042_port, B2 => n2887, 
                           ZN => n16531);
   U12922 : INV_X1 port map( A => n16530, ZN => n10810);
   U12923 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_25_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2041_port, B2 => n2887, 
                           ZN => n16530);
   U12924 : INV_X1 port map( A => n16529, ZN => n10811);
   U12925 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_24_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2040_port, B2 => n2887, 
                           ZN => n16529);
   U12926 : INV_X1 port map( A => n16528, ZN => n10812);
   U12927 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_23_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2039_port, B2 => n2886, 
                           ZN => n16528);
   U12928 : INV_X1 port map( A => n16527, ZN => n10813);
   U12929 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_22_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2038_port, B2 => n2886, 
                           ZN => n16527);
   U12930 : INV_X1 port map( A => n16526, ZN => n10814);
   U12931 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_21_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2037_port, B2 => n2886, 
                           ZN => n16526);
   U12932 : INV_X1 port map( A => n16525, ZN => n10815);
   U12933 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_20_port,
                           A2 => n2882, B1 => 
                           DataPath_RF_bus_reg_dataout_2036_port, B2 => n2886, 
                           ZN => n16525);
   U12934 : INV_X1 port map( A => n16524, ZN => n10816);
   U12935 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_19_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2035_port, B2 => n2886, 
                           ZN => n16524);
   U12936 : INV_X1 port map( A => n16523, ZN => n10817);
   U12937 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_18_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2034_port, B2 => n2886, 
                           ZN => n16523);
   U12938 : INV_X1 port map( A => n16522, ZN => n10818);
   U12939 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_17_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2033_port, B2 => n2886, 
                           ZN => n16522);
   U12940 : INV_X1 port map( A => n16521, ZN => n10819);
   U12941 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_16_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2032_port, B2 => n2886, 
                           ZN => n16521);
   U12942 : INV_X1 port map( A => n16520, ZN => n10820);
   U12943 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_15_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2031_port, B2 => n2886, 
                           ZN => n16520);
   U12944 : INV_X1 port map( A => n16519, ZN => n10821);
   U12945 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_14_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2030_port, B2 => n2886, 
                           ZN => n16519);
   U12946 : INV_X1 port map( A => n16518, ZN => n10822);
   U12947 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_13_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2029_port, B2 => n2886, 
                           ZN => n16518);
   U12948 : INV_X1 port map( A => n16517, ZN => n10823);
   U12949 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_12_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2028_port, B2 => n2886, 
                           ZN => n16517);
   U12950 : INV_X1 port map( A => n16516, ZN => n10824);
   U12951 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_11_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2027_port, B2 => n2885, 
                           ZN => n16516);
   U12952 : INV_X1 port map( A => n16515, ZN => n10825);
   U12953 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_10_port,
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2026_port, B2 => n2885, 
                           ZN => n16515);
   U12954 : INV_X1 port map( A => n16514, ZN => n10826);
   U12955 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_9_port, 
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2025_port, B2 => n2885, 
                           ZN => n16514);
   U12956 : INV_X1 port map( A => n16513, ZN => n10827);
   U12957 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_8_port, 
                           A2 => n2883, B1 => 
                           DataPath_RF_bus_reg_dataout_2024_port, B2 => n2885, 
                           ZN => n16513);
   U12958 : INV_X1 port map( A => n16512, ZN => n10828);
   U12959 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_7_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2023_port, B2 => n2885, 
                           ZN => n16512);
   U12960 : INV_X1 port map( A => n16511, ZN => n10829);
   U12961 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_6_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2022_port, B2 => n2885, 
                           ZN => n16511);
   U12962 : INV_X1 port map( A => n16510, ZN => n10830);
   U12963 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_5_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2021_port, B2 => n2885, 
                           ZN => n16510);
   U12964 : INV_X1 port map( A => n16509, ZN => n10831);
   U12965 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_4_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2020_port, B2 => n2885, 
                           ZN => n16509);
   U12966 : INV_X1 port map( A => n16508, ZN => n10832);
   U12967 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_3_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2019_port, B2 => n2885, 
                           ZN => n16508);
   U12968 : INV_X1 port map( A => n16507, ZN => n10833);
   U12969 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_2_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2018_port, B2 => n2885, 
                           ZN => n16507);
   U12970 : INV_X1 port map( A => n16506, ZN => n10834);
   U12971 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_1_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2017_port, B2 => n2885, 
                           ZN => n16506);
   U12972 : INV_X1 port map( A => n16503, ZN => n10835);
   U12973 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_3_0_port, 
                           A2 => n2884, B1 => 
                           DataPath_RF_bus_reg_dataout_2016_port, B2 => n2885, 
                           ZN => n16503);
   U12974 : INV_X1 port map( A => n16570, ZN => n10836);
   U12975 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2079_port, B2 => n2893, 
                           ZN => n16570);
   U12976 : INV_X1 port map( A => n16569, ZN => n10837);
   U12977 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2078_port, B2 => n2893, 
                           ZN => n16569);
   U12978 : INV_X1 port map( A => n16568, ZN => n10838);
   U12979 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2077_port, B2 => n2893, 
                           ZN => n16568);
   U12980 : INV_X1 port map( A => n16567, ZN => n10839);
   U12981 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2076_port, B2 => n2893, 
                           ZN => n16567);
   U12982 : INV_X1 port map( A => n16566, ZN => n10840);
   U12983 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2075_port, B2 => n2893, 
                           ZN => n16566);
   U12984 : INV_X1 port map( A => n16565, ZN => n10841);
   U12985 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2074_port, B2 => n2893, 
                           ZN => n16565);
   U12986 : INV_X1 port map( A => n16564, ZN => n10842);
   U12987 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2073_port, B2 => n2893, 
                           ZN => n16564);
   U12988 : INV_X1 port map( A => n16563, ZN => n10843);
   U12989 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2072_port, B2 => n2893, 
                           ZN => n16563);
   U12990 : INV_X1 port map( A => n16562, ZN => n10844);
   U12991 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2071_port, B2 => n2892, 
                           ZN => n16562);
   U12992 : INV_X1 port map( A => n16561, ZN => n10845);
   U12993 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2070_port, B2 => n2892, 
                           ZN => n16561);
   U12994 : INV_X1 port map( A => n16560, ZN => n10846);
   U12995 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2069_port, B2 => n2892, 
                           ZN => n16560);
   U12996 : INV_X1 port map( A => n16559, ZN => n10847);
   U12997 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2888, B1 => 
                           DataPath_RF_bus_reg_dataout_2068_port, B2 => n2892, 
                           ZN => n16559);
   U12998 : INV_X1 port map( A => n16558, ZN => n10848);
   U12999 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2067_port, B2 => n2892, 
                           ZN => n16558);
   U13000 : INV_X1 port map( A => n16557, ZN => n10849);
   U13001 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2066_port, B2 => n2892, 
                           ZN => n16557);
   U13002 : INV_X1 port map( A => n16556, ZN => n10850);
   U13003 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2065_port, B2 => n2892, 
                           ZN => n16556);
   U13004 : INV_X1 port map( A => n16555, ZN => n10851);
   U13005 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2064_port, B2 => n2892, 
                           ZN => n16555);
   U13006 : INV_X1 port map( A => n16554, ZN => n10852);
   U13007 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2063_port, B2 => n2892, 
                           ZN => n16554);
   U13008 : INV_X1 port map( A => n16553, ZN => n10853);
   U13009 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2062_port, B2 => n2892, 
                           ZN => n16553);
   U13010 : INV_X1 port map( A => n16552, ZN => n10854);
   U13011 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2061_port, B2 => n2892, 
                           ZN => n16552);
   U13012 : INV_X1 port map( A => n16551, ZN => n10855);
   U13013 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2060_port, B2 => n2892, 
                           ZN => n16551);
   U13014 : INV_X1 port map( A => n16550, ZN => n10856);
   U13015 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2059_port, B2 => n2891, 
                           ZN => n16550);
   U13016 : INV_X1 port map( A => n16549, ZN => n10857);
   U13017 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2058_port, B2 => n2891, 
                           ZN => n16549);
   U13018 : INV_X1 port map( A => n16548, ZN => n10858);
   U13019 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2057_port, B2 => n2891, 
                           ZN => n16548);
   U13020 : INV_X1 port map( A => n16547, ZN => n10859);
   U13021 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2889, B1 => 
                           DataPath_RF_bus_reg_dataout_2056_port, B2 => n2891, 
                           ZN => n16547);
   U13022 : INV_X1 port map( A => n16546, ZN => n10860);
   U13023 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2055_port, B2 => n2891, 
                           ZN => n16546);
   U13024 : INV_X1 port map( A => n16545, ZN => n10861);
   U13025 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2054_port, B2 => n2891, 
                           ZN => n16545);
   U13026 : INV_X1 port map( A => n16544, ZN => n10862);
   U13027 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2053_port, B2 => n2891, 
                           ZN => n16544);
   U13028 : INV_X1 port map( A => n16543, ZN => n10863);
   U13029 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2052_port, B2 => n2891, 
                           ZN => n16543);
   U13030 : INV_X1 port map( A => n16542, ZN => n10864);
   U13031 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2051_port, B2 => n2891, 
                           ZN => n16542);
   U13032 : INV_X1 port map( A => n16541, ZN => n10865);
   U13033 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2050_port, B2 => n2891, 
                           ZN => n16541);
   U13034 : INV_X1 port map( A => n16540, ZN => n10866);
   U13035 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2049_port, B2 => n2891, 
                           ZN => n16540);
   U13036 : INV_X1 port map( A => n16537, ZN => n10867);
   U13037 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2890, B1 => 
                           DataPath_RF_bus_reg_dataout_2048_port, B2 => n2891, 
                           ZN => n16537);
   U13038 : INV_X1 port map( A => n16604, ZN => n10868);
   U13039 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2111_port, B2 => n2899, 
                           ZN => n16604);
   U13040 : INV_X1 port map( A => n16603, ZN => n10869);
   U13041 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2110_port, B2 => n2899, 
                           ZN => n16603);
   U13042 : INV_X1 port map( A => n16602, ZN => n10870);
   U13043 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2109_port, B2 => n2899, 
                           ZN => n16602);
   U13044 : INV_X1 port map( A => n16601, ZN => n10871);
   U13045 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2108_port, B2 => n2899, 
                           ZN => n16601);
   U13046 : INV_X1 port map( A => n16600, ZN => n10872);
   U13047 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2107_port, B2 => n2899, 
                           ZN => n16600);
   U13048 : INV_X1 port map( A => n16599, ZN => n10873);
   U13049 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2106_port, B2 => n2899, 
                           ZN => n16599);
   U13050 : INV_X1 port map( A => n16598, ZN => n10874);
   U13051 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2105_port, B2 => n2899, 
                           ZN => n16598);
   U13052 : INV_X1 port map( A => n16597, ZN => n10875);
   U13053 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2104_port, B2 => n2899, 
                           ZN => n16597);
   U13054 : INV_X1 port map( A => n16596, ZN => n10876);
   U13055 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2103_port, B2 => n2898, 
                           ZN => n16596);
   U13056 : INV_X1 port map( A => n16595, ZN => n10877);
   U13057 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2102_port, B2 => n2898, 
                           ZN => n16595);
   U13058 : INV_X1 port map( A => n16594, ZN => n10878);
   U13059 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2101_port, B2 => n2898, 
                           ZN => n16594);
   U13060 : INV_X1 port map( A => n16593, ZN => n10879);
   U13061 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2894, B1 => 
                           DataPath_RF_bus_reg_dataout_2100_port, B2 => n2898, 
                           ZN => n16593);
   U13062 : INV_X1 port map( A => n16592, ZN => n10880);
   U13063 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2099_port, B2 => n2898, 
                           ZN => n16592);
   U13064 : INV_X1 port map( A => n16591, ZN => n10881);
   U13065 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2098_port, B2 => n2898, 
                           ZN => n16591);
   U13066 : INV_X1 port map( A => n16590, ZN => n10882);
   U13067 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2097_port, B2 => n2898, 
                           ZN => n16590);
   U13068 : INV_X1 port map( A => n16589, ZN => n10883);
   U13069 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2096_port, B2 => n2898, 
                           ZN => n16589);
   U13070 : INV_X1 port map( A => n16588, ZN => n10884);
   U13071 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2095_port, B2 => n2898, 
                           ZN => n16588);
   U13072 : INV_X1 port map( A => n16587, ZN => n10885);
   U13073 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2094_port, B2 => n2898, 
                           ZN => n16587);
   U13074 : INV_X1 port map( A => n16586, ZN => n10886);
   U13075 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2093_port, B2 => n2898, 
                           ZN => n16586);
   U13076 : INV_X1 port map( A => n16585, ZN => n10887);
   U13077 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2092_port, B2 => n2898, 
                           ZN => n16585);
   U13078 : INV_X1 port map( A => n16584, ZN => n10888);
   U13079 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2091_port, B2 => n2897, 
                           ZN => n16584);
   U13080 : INV_X1 port map( A => n16583, ZN => n10889);
   U13081 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2090_port, B2 => n2897, 
                           ZN => n16583);
   U13082 : INV_X1 port map( A => n16582, ZN => n10890);
   U13083 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2089_port, B2 => n2897, 
                           ZN => n16582);
   U13084 : INV_X1 port map( A => n16581, ZN => n10891);
   U13085 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2895, B1 => 
                           DataPath_RF_bus_reg_dataout_2088_port, B2 => n2897, 
                           ZN => n16581);
   U13086 : INV_X1 port map( A => n16580, ZN => n10892);
   U13087 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2087_port, B2 => n2897, 
                           ZN => n16580);
   U13088 : INV_X1 port map( A => n16579, ZN => n10893);
   U13089 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2086_port, B2 => n2897, 
                           ZN => n16579);
   U13090 : INV_X1 port map( A => n16578, ZN => n10894);
   U13091 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2085_port, B2 => n2897, 
                           ZN => n16578);
   U13092 : INV_X1 port map( A => n16577, ZN => n10895);
   U13093 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2084_port, B2 => n2897, 
                           ZN => n16577);
   U13094 : INV_X1 port map( A => n16576, ZN => n10896);
   U13095 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2083_port, B2 => n2897, 
                           ZN => n16576);
   U13096 : INV_X1 port map( A => n16575, ZN => n10897);
   U13097 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2082_port, B2 => n2897, 
                           ZN => n16575);
   U13098 : INV_X1 port map( A => n16574, ZN => n10898);
   U13099 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2081_port, B2 => n2897, 
                           ZN => n16574);
   U13100 : INV_X1 port map( A => n16571, ZN => n10899);
   U13101 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2896, B1 => 
                           DataPath_RF_bus_reg_dataout_2080_port, B2 => n2897, 
                           ZN => n16571);
   U13102 : INV_X1 port map( A => n16638, ZN => n10900);
   U13103 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2143_port, B2 => n2905, 
                           ZN => n16638);
   U13104 : INV_X1 port map( A => n16637, ZN => n10901);
   U13105 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2142_port, B2 => n2905, 
                           ZN => n16637);
   U13106 : INV_X1 port map( A => n16636, ZN => n10902);
   U13107 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2141_port, B2 => n2905, 
                           ZN => n16636);
   U13108 : INV_X1 port map( A => n16635, ZN => n10903);
   U13109 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2140_port, B2 => n2905, 
                           ZN => n16635);
   U13110 : INV_X1 port map( A => n16634, ZN => n10904);
   U13111 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2139_port, B2 => n2905, 
                           ZN => n16634);
   U13112 : INV_X1 port map( A => n16633, ZN => n10905);
   U13113 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2138_port, B2 => n2905, 
                           ZN => n16633);
   U13114 : INV_X1 port map( A => n16632, ZN => n10906);
   U13115 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2137_port, B2 => n2905, 
                           ZN => n16632);
   U13116 : INV_X1 port map( A => n16631, ZN => n10907);
   U13117 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2136_port, B2 => n2905, 
                           ZN => n16631);
   U13118 : INV_X1 port map( A => n16630, ZN => n10908);
   U13119 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2135_port, B2 => n2904, 
                           ZN => n16630);
   U13120 : INV_X1 port map( A => n16629, ZN => n10909);
   U13121 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2134_port, B2 => n2904, 
                           ZN => n16629);
   U13122 : INV_X1 port map( A => n16628, ZN => n10910);
   U13123 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2133_port, B2 => n2904, 
                           ZN => n16628);
   U13124 : INV_X1 port map( A => n16627, ZN => n10911);
   U13125 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2900, B1 => 
                           DataPath_RF_bus_reg_dataout_2132_port, B2 => n2904, 
                           ZN => n16627);
   U13126 : INV_X1 port map( A => n16626, ZN => n10912);
   U13127 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2131_port, B2 => n2904, 
                           ZN => n16626);
   U13128 : INV_X1 port map( A => n16625, ZN => n10913);
   U13129 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2130_port, B2 => n2904, 
                           ZN => n16625);
   U13130 : INV_X1 port map( A => n16624, ZN => n10914);
   U13131 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2129_port, B2 => n2904, 
                           ZN => n16624);
   U13132 : INV_X1 port map( A => n16623, ZN => n10915);
   U13133 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2128_port, B2 => n2904, 
                           ZN => n16623);
   U13134 : INV_X1 port map( A => n16622, ZN => n10916);
   U13135 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2127_port, B2 => n2904, 
                           ZN => n16622);
   U13136 : INV_X1 port map( A => n16621, ZN => n10917);
   U13137 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2126_port, B2 => n2904, 
                           ZN => n16621);
   U13138 : INV_X1 port map( A => n16620, ZN => n10918);
   U13139 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2125_port, B2 => n2904, 
                           ZN => n16620);
   U13140 : INV_X1 port map( A => n16619, ZN => n10919);
   U13141 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2124_port, B2 => n2904, 
                           ZN => n16619);
   U13142 : INV_X1 port map( A => n16618, ZN => n10920);
   U13143 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2123_port, B2 => n2903, 
                           ZN => n16618);
   U13144 : INV_X1 port map( A => n16617, ZN => n10921);
   U13145 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2122_port, B2 => n2903, 
                           ZN => n16617);
   U13146 : INV_X1 port map( A => n16616, ZN => n10922);
   U13147 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2121_port, B2 => n2903, 
                           ZN => n16616);
   U13148 : INV_X1 port map( A => n16615, ZN => n10923);
   U13149 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2901, B1 => 
                           DataPath_RF_bus_reg_dataout_2120_port, B2 => n2903, 
                           ZN => n16615);
   U13150 : INV_X1 port map( A => n16614, ZN => n10924);
   U13151 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2119_port, B2 => n2903, 
                           ZN => n16614);
   U13152 : INV_X1 port map( A => n16613, ZN => n10925);
   U13153 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2118_port, B2 => n2903, 
                           ZN => n16613);
   U13154 : INV_X1 port map( A => n16612, ZN => n10926);
   U13155 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2117_port, B2 => n2903, 
                           ZN => n16612);
   U13156 : INV_X1 port map( A => n16611, ZN => n10927);
   U13157 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2116_port, B2 => n2903, 
                           ZN => n16611);
   U13158 : INV_X1 port map( A => n16610, ZN => n10928);
   U13159 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2115_port, B2 => n2903, 
                           ZN => n16610);
   U13160 : INV_X1 port map( A => n16609, ZN => n10929);
   U13161 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2114_port, B2 => n2903, 
                           ZN => n16609);
   U13162 : INV_X1 port map( A => n16608, ZN => n10930);
   U13163 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2113_port, B2 => n2903, 
                           ZN => n16608);
   U13164 : INV_X1 port map( A => n16605, ZN => n10931);
   U13165 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2902, B1 => 
                           DataPath_RF_bus_reg_dataout_2112_port, B2 => n2903, 
                           ZN => n16605);
   U13166 : INV_X1 port map( A => n16672, ZN => n10932);
   U13167 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2175_port, B2 => n2911, 
                           ZN => n16672);
   U13168 : INV_X1 port map( A => n16671, ZN => n10933);
   U13169 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2174_port, B2 => n2911, 
                           ZN => n16671);
   U13170 : INV_X1 port map( A => n16670, ZN => n10934);
   U13171 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2173_port, B2 => n2911, 
                           ZN => n16670);
   U13172 : INV_X1 port map( A => n16669, ZN => n10935);
   U13173 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2172_port, B2 => n2911, 
                           ZN => n16669);
   U13174 : INV_X1 port map( A => n16668, ZN => n10936);
   U13175 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2171_port, B2 => n2911, 
                           ZN => n16668);
   U13176 : INV_X1 port map( A => n16667, ZN => n10937);
   U13177 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2170_port, B2 => n2911, 
                           ZN => n16667);
   U13178 : INV_X1 port map( A => n16666, ZN => n10938);
   U13179 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2169_port, B2 => n2911, 
                           ZN => n16666);
   U13180 : INV_X1 port map( A => n16665, ZN => n10939);
   U13181 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2168_port, B2 => n2911, 
                           ZN => n16665);
   U13182 : INV_X1 port map( A => n16664, ZN => n10940);
   U13183 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2167_port, B2 => n2910, 
                           ZN => n16664);
   U13184 : INV_X1 port map( A => n16663, ZN => n10941);
   U13185 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2166_port, B2 => n2910, 
                           ZN => n16663);
   U13186 : INV_X1 port map( A => n16662, ZN => n10942);
   U13187 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2165_port, B2 => n2910, 
                           ZN => n16662);
   U13188 : INV_X1 port map( A => n16661, ZN => n10943);
   U13189 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2906, B1 => 
                           DataPath_RF_bus_reg_dataout_2164_port, B2 => n2910, 
                           ZN => n16661);
   U13190 : INV_X1 port map( A => n16660, ZN => n10944);
   U13191 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2163_port, B2 => n2910, 
                           ZN => n16660);
   U13192 : INV_X1 port map( A => n16659, ZN => n10945);
   U13193 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2162_port, B2 => n2910, 
                           ZN => n16659);
   U13194 : INV_X1 port map( A => n16658, ZN => n10946);
   U13195 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2161_port, B2 => n2910, 
                           ZN => n16658);
   U13196 : INV_X1 port map( A => n16657, ZN => n10947);
   U13197 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2160_port, B2 => n2910, 
                           ZN => n16657);
   U13198 : INV_X1 port map( A => n16656, ZN => n10948);
   U13199 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2159_port, B2 => n2910, 
                           ZN => n16656);
   U13200 : INV_X1 port map( A => n16655, ZN => n10949);
   U13201 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2158_port, B2 => n2910, 
                           ZN => n16655);
   U13202 : INV_X1 port map( A => n16654, ZN => n10950);
   U13203 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2157_port, B2 => n2910, 
                           ZN => n16654);
   U13204 : INV_X1 port map( A => n16653, ZN => n10951);
   U13205 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2156_port, B2 => n2910, 
                           ZN => n16653);
   U13206 : INV_X1 port map( A => n16652, ZN => n10952);
   U13207 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2155_port, B2 => n2909, 
                           ZN => n16652);
   U13208 : INV_X1 port map( A => n16651, ZN => n10953);
   U13209 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2154_port, B2 => n2909, 
                           ZN => n16651);
   U13210 : INV_X1 port map( A => n16650, ZN => n10954);
   U13211 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2153_port, B2 => n2909, 
                           ZN => n16650);
   U13212 : INV_X1 port map( A => n16649, ZN => n10955);
   U13213 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2907, B1 => 
                           DataPath_RF_bus_reg_dataout_2152_port, B2 => n2909, 
                           ZN => n16649);
   U13214 : INV_X1 port map( A => n16648, ZN => n10956);
   U13215 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2151_port, B2 => n2909, 
                           ZN => n16648);
   U13216 : INV_X1 port map( A => n16647, ZN => n10957);
   U13217 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2150_port, B2 => n2909, 
                           ZN => n16647);
   U13218 : INV_X1 port map( A => n16646, ZN => n10958);
   U13219 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2149_port, B2 => n2909, 
                           ZN => n16646);
   U13220 : INV_X1 port map( A => n16645, ZN => n10959);
   U13221 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2148_port, B2 => n2909, 
                           ZN => n16645);
   U13222 : INV_X1 port map( A => n16644, ZN => n10960);
   U13223 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2147_port, B2 => n2909, 
                           ZN => n16644);
   U13224 : INV_X1 port map( A => n16643, ZN => n10961);
   U13225 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2146_port, B2 => n2909, 
                           ZN => n16643);
   U13226 : INV_X1 port map( A => n16642, ZN => n10962);
   U13227 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2145_port, B2 => n2909, 
                           ZN => n16642);
   U13228 : INV_X1 port map( A => n16639, ZN => n10963);
   U13229 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2908, B1 => 
                           DataPath_RF_bus_reg_dataout_2144_port, B2 => n2909, 
                           ZN => n16639);
   U13230 : INV_X1 port map( A => n16706, ZN => n10964);
   U13231 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2207_port, B2 => n2917, 
                           ZN => n16706);
   U13232 : INV_X1 port map( A => n16705, ZN => n10965);
   U13233 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2206_port, B2 => n2917, 
                           ZN => n16705);
   U13234 : INV_X1 port map( A => n16704, ZN => n10966);
   U13235 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2205_port, B2 => n2917, 
                           ZN => n16704);
   U13236 : INV_X1 port map( A => n16703, ZN => n10967);
   U13237 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2204_port, B2 => n2917, 
                           ZN => n16703);
   U13238 : INV_X1 port map( A => n16702, ZN => n10968);
   U13239 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2203_port, B2 => n2917, 
                           ZN => n16702);
   U13240 : INV_X1 port map( A => n16701, ZN => n10969);
   U13241 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2202_port, B2 => n2917, 
                           ZN => n16701);
   U13242 : INV_X1 port map( A => n16700, ZN => n10970);
   U13243 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2201_port, B2 => n2917, 
                           ZN => n16700);
   U13244 : INV_X1 port map( A => n16699, ZN => n10971);
   U13245 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2200_port, B2 => n2917, 
                           ZN => n16699);
   U13246 : INV_X1 port map( A => n16698, ZN => n10972);
   U13247 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2199_port, B2 => n2916, 
                           ZN => n16698);
   U13248 : INV_X1 port map( A => n16697, ZN => n10973);
   U13249 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2198_port, B2 => n2916, 
                           ZN => n16697);
   U13250 : INV_X1 port map( A => n16696, ZN => n10974);
   U13251 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2197_port, B2 => n2916, 
                           ZN => n16696);
   U13252 : INV_X1 port map( A => n16695, ZN => n10975);
   U13253 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2912, B1 => 
                           DataPath_RF_bus_reg_dataout_2196_port, B2 => n2916, 
                           ZN => n16695);
   U13254 : INV_X1 port map( A => n16694, ZN => n10976);
   U13255 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2195_port, B2 => n2916, 
                           ZN => n16694);
   U13256 : INV_X1 port map( A => n16693, ZN => n10977);
   U13257 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2194_port, B2 => n2916, 
                           ZN => n16693);
   U13258 : INV_X1 port map( A => n16692, ZN => n10978);
   U13259 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2193_port, B2 => n2916, 
                           ZN => n16692);
   U13260 : INV_X1 port map( A => n16691, ZN => n10979);
   U13261 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2192_port, B2 => n2916, 
                           ZN => n16691);
   U13262 : INV_X1 port map( A => n16690, ZN => n10980);
   U13263 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2191_port, B2 => n2916, 
                           ZN => n16690);
   U13264 : INV_X1 port map( A => n16689, ZN => n10981);
   U13265 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2190_port, B2 => n2916, 
                           ZN => n16689);
   U13266 : INV_X1 port map( A => n16688, ZN => n10982);
   U13267 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2189_port, B2 => n2916, 
                           ZN => n16688);
   U13268 : INV_X1 port map( A => n16687, ZN => n10983);
   U13269 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2188_port, B2 => n2916, 
                           ZN => n16687);
   U13270 : INV_X1 port map( A => n16686, ZN => n10984);
   U13271 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2187_port, B2 => n2915, 
                           ZN => n16686);
   U13272 : INV_X1 port map( A => n16685, ZN => n10985);
   U13273 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2186_port, B2 => n2915, 
                           ZN => n16685);
   U13274 : INV_X1 port map( A => n16684, ZN => n10986);
   U13275 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2185_port, B2 => n2915, 
                           ZN => n16684);
   U13276 : INV_X1 port map( A => n16683, ZN => n10987);
   U13277 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2913, B1 => 
                           DataPath_RF_bus_reg_dataout_2184_port, B2 => n2915, 
                           ZN => n16683);
   U13278 : INV_X1 port map( A => n16682, ZN => n10988);
   U13279 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2183_port, B2 => n2915, 
                           ZN => n16682);
   U13280 : INV_X1 port map( A => n16681, ZN => n10989);
   U13281 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2182_port, B2 => n2915, 
                           ZN => n16681);
   U13282 : INV_X1 port map( A => n16680, ZN => n10990);
   U13283 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2181_port, B2 => n2915, 
                           ZN => n16680);
   U13284 : INV_X1 port map( A => n16679, ZN => n10991);
   U13285 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2180_port, B2 => n2915, 
                           ZN => n16679);
   U13286 : INV_X1 port map( A => n16678, ZN => n10992);
   U13287 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2179_port, B2 => n2915, 
                           ZN => n16678);
   U13288 : INV_X1 port map( A => n16677, ZN => n10993);
   U13289 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2178_port, B2 => n2915, 
                           ZN => n16677);
   U13290 : INV_X1 port map( A => n16676, ZN => n10994);
   U13291 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2177_port, B2 => n2915, 
                           ZN => n16676);
   U13292 : INV_X1 port map( A => n16673, ZN => n10995);
   U13293 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2914, B1 => 
                           DataPath_RF_bus_reg_dataout_2176_port, B2 => n2915, 
                           ZN => n16673);
   U13294 : INV_X1 port map( A => n16740, ZN => n10996);
   U13295 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2239_port, B2 => n2923, 
                           ZN => n16740);
   U13296 : INV_X1 port map( A => n16739, ZN => n10997);
   U13297 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2238_port, B2 => n2923, 
                           ZN => n16739);
   U13298 : INV_X1 port map( A => n16738, ZN => n10998);
   U13299 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2237_port, B2 => n2923, 
                           ZN => n16738);
   U13300 : INV_X1 port map( A => n16737, ZN => n10999);
   U13301 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2236_port, B2 => n2923, 
                           ZN => n16737);
   U13302 : INV_X1 port map( A => n16736, ZN => n11000);
   U13303 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2235_port, B2 => n2923, 
                           ZN => n16736);
   U13304 : INV_X1 port map( A => n16735, ZN => n11001);
   U13305 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2234_port, B2 => n2923, 
                           ZN => n16735);
   U13306 : INV_X1 port map( A => n16734, ZN => n11002);
   U13307 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2233_port, B2 => n2923, 
                           ZN => n16734);
   U13308 : INV_X1 port map( A => n16733, ZN => n11003);
   U13309 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2232_port, B2 => n2923, 
                           ZN => n16733);
   U13310 : INV_X1 port map( A => n16732, ZN => n11004);
   U13311 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2231_port, B2 => n2922, 
                           ZN => n16732);
   U13312 : INV_X1 port map( A => n16731, ZN => n11005);
   U13313 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2230_port, B2 => n2922, 
                           ZN => n16731);
   U13314 : INV_X1 port map( A => n16730, ZN => n11006);
   U13315 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2229_port, B2 => n2922, 
                           ZN => n16730);
   U13316 : INV_X1 port map( A => n16729, ZN => n11007);
   U13317 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2918, B1 => 
                           DataPath_RF_bus_reg_dataout_2228_port, B2 => n2922, 
                           ZN => n16729);
   U13318 : INV_X1 port map( A => n16728, ZN => n11008);
   U13319 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2227_port, B2 => n2922, 
                           ZN => n16728);
   U13320 : INV_X1 port map( A => n16727, ZN => n11009);
   U13321 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2226_port, B2 => n2922, 
                           ZN => n16727);
   U13322 : INV_X1 port map( A => n16726, ZN => n11010);
   U13323 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2225_port, B2 => n2922, 
                           ZN => n16726);
   U13324 : INV_X1 port map( A => n16725, ZN => n11011);
   U13325 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2224_port, B2 => n2922, 
                           ZN => n16725);
   U13326 : INV_X1 port map( A => n16724, ZN => n11012);
   U13327 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2223_port, B2 => n2922, 
                           ZN => n16724);
   U13328 : INV_X1 port map( A => n16723, ZN => n11013);
   U13329 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2222_port, B2 => n2922, 
                           ZN => n16723);
   U13330 : INV_X1 port map( A => n16722, ZN => n11014);
   U13331 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2221_port, B2 => n2922, 
                           ZN => n16722);
   U13332 : INV_X1 port map( A => n16721, ZN => n11015);
   U13333 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2220_port, B2 => n2922, 
                           ZN => n16721);
   U13334 : INV_X1 port map( A => n16720, ZN => n11016);
   U13335 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2219_port, B2 => n2921, 
                           ZN => n16720);
   U13336 : INV_X1 port map( A => n16719, ZN => n11017);
   U13337 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2218_port, B2 => n2921, 
                           ZN => n16719);
   U13338 : INV_X1 port map( A => n16718, ZN => n11018);
   U13339 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2217_port, B2 => n2921, 
                           ZN => n16718);
   U13340 : INV_X1 port map( A => n16717, ZN => n11019);
   U13341 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2919, B1 => 
                           DataPath_RF_bus_reg_dataout_2216_port, B2 => n2921, 
                           ZN => n16717);
   U13342 : INV_X1 port map( A => n16716, ZN => n11020);
   U13343 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2215_port, B2 => n2921, 
                           ZN => n16716);
   U13344 : INV_X1 port map( A => n16715, ZN => n11021);
   U13345 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2214_port, B2 => n2921, 
                           ZN => n16715);
   U13346 : INV_X1 port map( A => n16714, ZN => n11022);
   U13347 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2213_port, B2 => n2921, 
                           ZN => n16714);
   U13348 : INV_X1 port map( A => n16713, ZN => n11023);
   U13349 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2212_port, B2 => n2921, 
                           ZN => n16713);
   U13350 : INV_X1 port map( A => n16712, ZN => n11024);
   U13351 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2211_port, B2 => n2921, 
                           ZN => n16712);
   U13352 : INV_X1 port map( A => n16711, ZN => n11025);
   U13353 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2210_port, B2 => n2921, 
                           ZN => n16711);
   U13354 : INV_X1 port map( A => n16710, ZN => n11026);
   U13355 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2209_port, B2 => n2921, 
                           ZN => n16710);
   U13356 : INV_X1 port map( A => n16707, ZN => n11027);
   U13357 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2920, B1 => 
                           DataPath_RF_bus_reg_dataout_2208_port, B2 => n2921, 
                           ZN => n16707);
   U13358 : INV_X1 port map( A => n16774, ZN => n11028);
   U13359 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2271_port, B2 => n2929, 
                           ZN => n16774);
   U13360 : INV_X1 port map( A => n16773, ZN => n11029);
   U13361 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2270_port, B2 => n2929, 
                           ZN => n16773);
   U13362 : INV_X1 port map( A => n16772, ZN => n11030);
   U13363 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2269_port, B2 => n2929, 
                           ZN => n16772);
   U13364 : INV_X1 port map( A => n16771, ZN => n11031);
   U13365 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2268_port, B2 => n2929, 
                           ZN => n16771);
   U13366 : INV_X1 port map( A => n16770, ZN => n11032);
   U13367 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2267_port, B2 => n2929, 
                           ZN => n16770);
   U13368 : INV_X1 port map( A => n16769, ZN => n11033);
   U13369 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2266_port, B2 => n2929, 
                           ZN => n16769);
   U13370 : INV_X1 port map( A => n16768, ZN => n11034);
   U13371 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2265_port, B2 => n2929, 
                           ZN => n16768);
   U13372 : INV_X1 port map( A => n16767, ZN => n11035);
   U13373 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2264_port, B2 => n2929, 
                           ZN => n16767);
   U13374 : INV_X1 port map( A => n16766, ZN => n11036);
   U13375 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2263_port, B2 => n2928, 
                           ZN => n16766);
   U13376 : INV_X1 port map( A => n16765, ZN => n11037);
   U13377 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2262_port, B2 => n2928, 
                           ZN => n16765);
   U13378 : INV_X1 port map( A => n16764, ZN => n11038);
   U13379 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2261_port, B2 => n2928, 
                           ZN => n16764);
   U13380 : INV_X1 port map( A => n16763, ZN => n11039);
   U13381 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2924, B1 => 
                           DataPath_RF_bus_reg_dataout_2260_port, B2 => n2928, 
                           ZN => n16763);
   U13382 : INV_X1 port map( A => n16762, ZN => n11040);
   U13383 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2259_port, B2 => n2928, 
                           ZN => n16762);
   U13384 : INV_X1 port map( A => n16761, ZN => n11041);
   U13385 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2258_port, B2 => n2928, 
                           ZN => n16761);
   U13386 : INV_X1 port map( A => n16760, ZN => n11042);
   U13387 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2257_port, B2 => n2928, 
                           ZN => n16760);
   U13388 : INV_X1 port map( A => n16759, ZN => n11043);
   U13389 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2256_port, B2 => n2928, 
                           ZN => n16759);
   U13390 : INV_X1 port map( A => n16758, ZN => n11044);
   U13391 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2255_port, B2 => n2928, 
                           ZN => n16758);
   U13392 : INV_X1 port map( A => n16757, ZN => n11045);
   U13393 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2254_port, B2 => n2928, 
                           ZN => n16757);
   U13394 : INV_X1 port map( A => n16756, ZN => n11046);
   U13395 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2253_port, B2 => n2928, 
                           ZN => n16756);
   U13396 : INV_X1 port map( A => n16755, ZN => n11047);
   U13397 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2252_port, B2 => n2928, 
                           ZN => n16755);
   U13398 : INV_X1 port map( A => n16754, ZN => n11048);
   U13399 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2251_port, B2 => n2927, 
                           ZN => n16754);
   U13400 : INV_X1 port map( A => n16753, ZN => n11049);
   U13401 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2250_port, B2 => n2927, 
                           ZN => n16753);
   U13402 : INV_X1 port map( A => n16752, ZN => n11050);
   U13403 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2249_port, B2 => n2927, 
                           ZN => n16752);
   U13404 : INV_X1 port map( A => n16751, ZN => n11051);
   U13405 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2925, B1 => 
                           DataPath_RF_bus_reg_dataout_2248_port, B2 => n2927, 
                           ZN => n16751);
   U13406 : INV_X1 port map( A => n16750, ZN => n11052);
   U13407 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2247_port, B2 => n2927, 
                           ZN => n16750);
   U13408 : INV_X1 port map( A => n16749, ZN => n11053);
   U13409 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2246_port, B2 => n2927, 
                           ZN => n16749);
   U13410 : INV_X1 port map( A => n16748, ZN => n11054);
   U13411 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2245_port, B2 => n2927, 
                           ZN => n16748);
   U13412 : INV_X1 port map( A => n16747, ZN => n11055);
   U13413 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2244_port, B2 => n2927, 
                           ZN => n16747);
   U13414 : INV_X1 port map( A => n16746, ZN => n11056);
   U13415 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2243_port, B2 => n2927, 
                           ZN => n16746);
   U13416 : INV_X1 port map( A => n16745, ZN => n11057);
   U13417 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2242_port, B2 => n2927, 
                           ZN => n16745);
   U13418 : INV_X1 port map( A => n16744, ZN => n11058);
   U13419 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2241_port, B2 => n2927, 
                           ZN => n16744);
   U13420 : INV_X1 port map( A => n16741, ZN => n11059);
   U13421 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2926, B1 => 
                           DataPath_RF_bus_reg_dataout_2240_port, B2 => n2927, 
                           ZN => n16741);
   U13422 : INV_X1 port map( A => n16808, ZN => n11060);
   U13423 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2303_port, B2 => n2935, 
                           ZN => n16808);
   U13424 : INV_X1 port map( A => n16807, ZN => n11061);
   U13425 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2302_port, B2 => n2935, 
                           ZN => n16807);
   U13426 : INV_X1 port map( A => n16806, ZN => n11062);
   U13427 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2301_port, B2 => n2935, 
                           ZN => n16806);
   U13428 : INV_X1 port map( A => n16805, ZN => n11063);
   U13429 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2300_port, B2 => n2935, 
                           ZN => n16805);
   U13430 : INV_X1 port map( A => n16804, ZN => n11064);
   U13431 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2299_port, B2 => n2935, 
                           ZN => n16804);
   U13432 : INV_X1 port map( A => n16803, ZN => n11065);
   U13433 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2298_port, B2 => n2935, 
                           ZN => n16803);
   U13434 : INV_X1 port map( A => n16802, ZN => n11066);
   U13435 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2297_port, B2 => n2935, 
                           ZN => n16802);
   U13436 : INV_X1 port map( A => n16801, ZN => n11067);
   U13437 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2296_port, B2 => n2935, 
                           ZN => n16801);
   U13438 : INV_X1 port map( A => n16800, ZN => n11068);
   U13439 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2295_port, B2 => n2934, 
                           ZN => n16800);
   U13440 : INV_X1 port map( A => n16799, ZN => n11069);
   U13441 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2294_port, B2 => n2934, 
                           ZN => n16799);
   U13442 : INV_X1 port map( A => n16798, ZN => n11070);
   U13443 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2293_port, B2 => n2934, 
                           ZN => n16798);
   U13444 : INV_X1 port map( A => n16797, ZN => n11071);
   U13445 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2930, B1 => 
                           DataPath_RF_bus_reg_dataout_2292_port, B2 => n2934, 
                           ZN => n16797);
   U13446 : INV_X1 port map( A => n16796, ZN => n11072);
   U13447 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2291_port, B2 => n2934, 
                           ZN => n16796);
   U13448 : INV_X1 port map( A => n16795, ZN => n11073);
   U13449 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2290_port, B2 => n2934, 
                           ZN => n16795);
   U13450 : INV_X1 port map( A => n16794, ZN => n11074);
   U13451 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2289_port, B2 => n2934, 
                           ZN => n16794);
   U13452 : INV_X1 port map( A => n16793, ZN => n11075);
   U13453 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2288_port, B2 => n2934, 
                           ZN => n16793);
   U13454 : INV_X1 port map( A => n16792, ZN => n11076);
   U13455 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2287_port, B2 => n2934, 
                           ZN => n16792);
   U13456 : INV_X1 port map( A => n16791, ZN => n11077);
   U13457 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2286_port, B2 => n2934, 
                           ZN => n16791);
   U13458 : INV_X1 port map( A => n16790, ZN => n11078);
   U13459 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2285_port, B2 => n2934, 
                           ZN => n16790);
   U13460 : INV_X1 port map( A => n16789, ZN => n11079);
   U13461 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2284_port, B2 => n2934, 
                           ZN => n16789);
   U13462 : INV_X1 port map( A => n16788, ZN => n11080);
   U13463 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2283_port, B2 => n2933, 
                           ZN => n16788);
   U13464 : INV_X1 port map( A => n16787, ZN => n11081);
   U13465 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2282_port, B2 => n2933, 
                           ZN => n16787);
   U13466 : INV_X1 port map( A => n16786, ZN => n11082);
   U13467 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2281_port, B2 => n2933, 
                           ZN => n16786);
   U13468 : INV_X1 port map( A => n16785, ZN => n11083);
   U13469 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2931, B1 => 
                           DataPath_RF_bus_reg_dataout_2280_port, B2 => n2933, 
                           ZN => n16785);
   U13470 : INV_X1 port map( A => n16784, ZN => n11084);
   U13471 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2279_port, B2 => n2933, 
                           ZN => n16784);
   U13472 : INV_X1 port map( A => n16783, ZN => n11085);
   U13473 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2278_port, B2 => n2933, 
                           ZN => n16783);
   U13474 : INV_X1 port map( A => n16782, ZN => n11086);
   U13475 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2277_port, B2 => n2933, 
                           ZN => n16782);
   U13476 : INV_X1 port map( A => n16781, ZN => n11087);
   U13477 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2276_port, B2 => n2933, 
                           ZN => n16781);
   U13478 : INV_X1 port map( A => n16780, ZN => n11088);
   U13479 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2275_port, B2 => n2933, 
                           ZN => n16780);
   U13480 : INV_X1 port map( A => n16779, ZN => n11089);
   U13481 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2274_port, B2 => n2933, 
                           ZN => n16779);
   U13482 : INV_X1 port map( A => n16778, ZN => n11090);
   U13483 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2273_port, B2 => n2933, 
                           ZN => n16778);
   U13484 : INV_X1 port map( A => n16775, ZN => n11091);
   U13485 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2932, B1 => 
                           DataPath_RF_bus_reg_dataout_2272_port, B2 => n2933, 
                           ZN => n16775);
   U13486 : INV_X1 port map( A => n16842, ZN => n11092);
   U13487 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2335_port, B2 => n2941, 
                           ZN => n16842);
   U13488 : INV_X1 port map( A => n16841, ZN => n11093);
   U13489 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2334_port, B2 => n2941, 
                           ZN => n16841);
   U13490 : INV_X1 port map( A => n16840, ZN => n11094);
   U13491 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2333_port, B2 => n2941, 
                           ZN => n16840);
   U13492 : INV_X1 port map( A => n16839, ZN => n11095);
   U13493 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2332_port, B2 => n2941, 
                           ZN => n16839);
   U13494 : INV_X1 port map( A => n16838, ZN => n11096);
   U13495 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2331_port, B2 => n2941, 
                           ZN => n16838);
   U13496 : INV_X1 port map( A => n16837, ZN => n11097);
   U13497 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2330_port, B2 => n2941, 
                           ZN => n16837);
   U13498 : INV_X1 port map( A => n16836, ZN => n11098);
   U13499 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2329_port, B2 => n2941, 
                           ZN => n16836);
   U13500 : INV_X1 port map( A => n16835, ZN => n11099);
   U13501 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2328_port, B2 => n2941, 
                           ZN => n16835);
   U13502 : INV_X1 port map( A => n16834, ZN => n11100);
   U13503 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2327_port, B2 => n2940, 
                           ZN => n16834);
   U13504 : INV_X1 port map( A => n16833, ZN => n11101);
   U13505 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2326_port, B2 => n2940, 
                           ZN => n16833);
   U13506 : INV_X1 port map( A => n16832, ZN => n11102);
   U13507 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2325_port, B2 => n2940, 
                           ZN => n16832);
   U13508 : INV_X1 port map( A => n16831, ZN => n11103);
   U13509 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2936, B1 => 
                           DataPath_RF_bus_reg_dataout_2324_port, B2 => n2940, 
                           ZN => n16831);
   U13510 : INV_X1 port map( A => n16830, ZN => n11104);
   U13511 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2323_port, B2 => n2940, 
                           ZN => n16830);
   U13512 : INV_X1 port map( A => n16829, ZN => n11105);
   U13513 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2322_port, B2 => n2940, 
                           ZN => n16829);
   U13514 : INV_X1 port map( A => n16828, ZN => n11106);
   U13515 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2321_port, B2 => n2940, 
                           ZN => n16828);
   U13516 : INV_X1 port map( A => n16827, ZN => n11107);
   U13517 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2320_port, B2 => n2940, 
                           ZN => n16827);
   U13518 : INV_X1 port map( A => n16826, ZN => n11108);
   U13519 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2319_port, B2 => n2940, 
                           ZN => n16826);
   U13520 : INV_X1 port map( A => n16825, ZN => n11109);
   U13521 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2318_port, B2 => n2940, 
                           ZN => n16825);
   U13522 : INV_X1 port map( A => n16824, ZN => n11110);
   U13523 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2317_port, B2 => n2940, 
                           ZN => n16824);
   U13524 : INV_X1 port map( A => n16823, ZN => n11111);
   U13525 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2316_port, B2 => n2940, 
                           ZN => n16823);
   U13526 : INV_X1 port map( A => n16822, ZN => n11112);
   U13527 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2315_port, B2 => n2939, 
                           ZN => n16822);
   U13528 : INV_X1 port map( A => n16821, ZN => n11113);
   U13529 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2314_port, B2 => n2939, 
                           ZN => n16821);
   U13530 : INV_X1 port map( A => n16820, ZN => n11114);
   U13531 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2313_port, B2 => n2939, 
                           ZN => n16820);
   U13532 : INV_X1 port map( A => n16819, ZN => n11115);
   U13533 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2937, B1 => 
                           DataPath_RF_bus_reg_dataout_2312_port, B2 => n2939, 
                           ZN => n16819);
   U13534 : INV_X1 port map( A => n16818, ZN => n11116);
   U13535 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2311_port, B2 => n2939, 
                           ZN => n16818);
   U13536 : INV_X1 port map( A => n16817, ZN => n11117);
   U13537 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2310_port, B2 => n2939, 
                           ZN => n16817);
   U13538 : INV_X1 port map( A => n16816, ZN => n11118);
   U13539 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2309_port, B2 => n2939, 
                           ZN => n16816);
   U13540 : INV_X1 port map( A => n16815, ZN => n11119);
   U13541 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2308_port, B2 => n2939, 
                           ZN => n16815);
   U13542 : INV_X1 port map( A => n16814, ZN => n11120);
   U13543 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2307_port, B2 => n2939, 
                           ZN => n16814);
   U13544 : INV_X1 port map( A => n16813, ZN => n11121);
   U13545 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2306_port, B2 => n2939, 
                           ZN => n16813);
   U13546 : INV_X1 port map( A => n16812, ZN => n11122);
   U13547 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2305_port, B2 => n2939, 
                           ZN => n16812);
   U13548 : INV_X1 port map( A => n16809, ZN => n11123);
   U13549 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2938, B1 => 
                           DataPath_RF_bus_reg_dataout_2304_port, B2 => n2939, 
                           ZN => n16809);
   U13550 : INV_X1 port map( A => n16876, ZN => n11124);
   U13551 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2367_port, B2 => n2947, 
                           ZN => n16876);
   U13552 : INV_X1 port map( A => n16875, ZN => n11125);
   U13553 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2366_port, B2 => n2947, 
                           ZN => n16875);
   U13554 : INV_X1 port map( A => n16874, ZN => n11126);
   U13555 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2365_port, B2 => n2947, 
                           ZN => n16874);
   U13556 : INV_X1 port map( A => n16873, ZN => n11127);
   U13557 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2364_port, B2 => n2947, 
                           ZN => n16873);
   U13558 : INV_X1 port map( A => n16872, ZN => n11128);
   U13559 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2363_port, B2 => n2947, 
                           ZN => n16872);
   U13560 : INV_X1 port map( A => n16871, ZN => n11129);
   U13561 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2362_port, B2 => n2947, 
                           ZN => n16871);
   U13562 : INV_X1 port map( A => n16870, ZN => n11130);
   U13563 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2361_port, B2 => n2947, 
                           ZN => n16870);
   U13564 : INV_X1 port map( A => n16869, ZN => n11131);
   U13565 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2360_port, B2 => n2947, 
                           ZN => n16869);
   U13566 : INV_X1 port map( A => n16868, ZN => n11132);
   U13567 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2359_port, B2 => n2946, 
                           ZN => n16868);
   U13568 : INV_X1 port map( A => n16867, ZN => n11133);
   U13569 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2358_port, B2 => n2946, 
                           ZN => n16867);
   U13570 : INV_X1 port map( A => n16866, ZN => n11134);
   U13571 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2357_port, B2 => n2946, 
                           ZN => n16866);
   U13572 : INV_X1 port map( A => n16865, ZN => n11135);
   U13573 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2942, B1 => 
                           DataPath_RF_bus_reg_dataout_2356_port, B2 => n2946, 
                           ZN => n16865);
   U13574 : INV_X1 port map( A => n16864, ZN => n11136);
   U13575 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2355_port, B2 => n2946, 
                           ZN => n16864);
   U13576 : INV_X1 port map( A => n16863, ZN => n11137);
   U13577 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2354_port, B2 => n2946, 
                           ZN => n16863);
   U13578 : INV_X1 port map( A => n16862, ZN => n11138);
   U13579 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2353_port, B2 => n2946, 
                           ZN => n16862);
   U13580 : INV_X1 port map( A => n16861, ZN => n11139);
   U13581 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2352_port, B2 => n2946, 
                           ZN => n16861);
   U13582 : INV_X1 port map( A => n16860, ZN => n11140);
   U13583 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2351_port, B2 => n2946, 
                           ZN => n16860);
   U13584 : INV_X1 port map( A => n16859, ZN => n11141);
   U13585 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2350_port, B2 => n2946, 
                           ZN => n16859);
   U13586 : INV_X1 port map( A => n16858, ZN => n11142);
   U13587 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2349_port, B2 => n2946, 
                           ZN => n16858);
   U13588 : INV_X1 port map( A => n16857, ZN => n11143);
   U13589 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2348_port, B2 => n2946, 
                           ZN => n16857);
   U13590 : INV_X1 port map( A => n16856, ZN => n11144);
   U13591 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2347_port, B2 => n2945, 
                           ZN => n16856);
   U13592 : INV_X1 port map( A => n16855, ZN => n11145);
   U13593 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2346_port, B2 => n2945, 
                           ZN => n16855);
   U13594 : INV_X1 port map( A => n16854, ZN => n11146);
   U13595 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2345_port, B2 => n2945, 
                           ZN => n16854);
   U13596 : INV_X1 port map( A => n16853, ZN => n11147);
   U13597 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2943, B1 => 
                           DataPath_RF_bus_reg_dataout_2344_port, B2 => n2945, 
                           ZN => n16853);
   U13598 : INV_X1 port map( A => n16852, ZN => n11148);
   U13599 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2343_port, B2 => n2945, 
                           ZN => n16852);
   U13600 : INV_X1 port map( A => n16851, ZN => n11149);
   U13601 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2342_port, B2 => n2945, 
                           ZN => n16851);
   U13602 : INV_X1 port map( A => n16850, ZN => n11150);
   U13603 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2341_port, B2 => n2945, 
                           ZN => n16850);
   U13604 : INV_X1 port map( A => n16849, ZN => n11151);
   U13605 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2340_port, B2 => n2945, 
                           ZN => n16849);
   U13606 : INV_X1 port map( A => n16848, ZN => n11152);
   U13607 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2339_port, B2 => n2945, 
                           ZN => n16848);
   U13608 : INV_X1 port map( A => n16847, ZN => n11153);
   U13609 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2338_port, B2 => n2945, 
                           ZN => n16847);
   U13610 : INV_X1 port map( A => n16846, ZN => n11154);
   U13611 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2337_port, B2 => n2945, 
                           ZN => n16846);
   U13612 : INV_X1 port map( A => n16843, ZN => n11155);
   U13613 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2944, B1 => 
                           DataPath_RF_bus_reg_dataout_2336_port, B2 => n2945, 
                           ZN => n16843);
   U13614 : INV_X1 port map( A => n16910, ZN => n11156);
   U13615 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2399_port, B2 => n2953, 
                           ZN => n16910);
   U13616 : INV_X1 port map( A => n16909, ZN => n11157);
   U13617 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2398_port, B2 => n2953, 
                           ZN => n16909);
   U13618 : INV_X1 port map( A => n16908, ZN => n11158);
   U13619 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2397_port, B2 => n2953, 
                           ZN => n16908);
   U13620 : INV_X1 port map( A => n16907, ZN => n11159);
   U13621 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2396_port, B2 => n2953, 
                           ZN => n16907);
   U13622 : INV_X1 port map( A => n16906, ZN => n11160);
   U13623 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2395_port, B2 => n2953, 
                           ZN => n16906);
   U13624 : INV_X1 port map( A => n16905, ZN => n11161);
   U13625 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2394_port, B2 => n2953, 
                           ZN => n16905);
   U13626 : INV_X1 port map( A => n16904, ZN => n11162);
   U13627 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2393_port, B2 => n2953, 
                           ZN => n16904);
   U13628 : INV_X1 port map( A => n16903, ZN => n11163);
   U13629 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2392_port, B2 => n2953, 
                           ZN => n16903);
   U13630 : INV_X1 port map( A => n16902, ZN => n11164);
   U13631 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2391_port, B2 => n2952, 
                           ZN => n16902);
   U13632 : INV_X1 port map( A => n16901, ZN => n11165);
   U13633 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2390_port, B2 => n2952, 
                           ZN => n16901);
   U13634 : INV_X1 port map( A => n16900, ZN => n11166);
   U13635 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2389_port, B2 => n2952, 
                           ZN => n16900);
   U13636 : INV_X1 port map( A => n16899, ZN => n11167);
   U13637 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2948, B1 => 
                           DataPath_RF_bus_reg_dataout_2388_port, B2 => n2952, 
                           ZN => n16899);
   U13638 : INV_X1 port map( A => n16898, ZN => n11168);
   U13639 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2387_port, B2 => n2952, 
                           ZN => n16898);
   U13640 : INV_X1 port map( A => n16897, ZN => n11169);
   U13641 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2386_port, B2 => n2952, 
                           ZN => n16897);
   U13642 : INV_X1 port map( A => n16896, ZN => n11170);
   U13643 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2385_port, B2 => n2952, 
                           ZN => n16896);
   U13644 : INV_X1 port map( A => n16895, ZN => n11171);
   U13645 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2384_port, B2 => n2952, 
                           ZN => n16895);
   U13646 : INV_X1 port map( A => n16894, ZN => n11172);
   U13647 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2383_port, B2 => n2952, 
                           ZN => n16894);
   U13648 : INV_X1 port map( A => n16893, ZN => n11173);
   U13649 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2382_port, B2 => n2952, 
                           ZN => n16893);
   U13650 : INV_X1 port map( A => n16892, ZN => n11174);
   U13651 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2381_port, B2 => n2952, 
                           ZN => n16892);
   U13652 : INV_X1 port map( A => n16891, ZN => n11175);
   U13653 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2380_port, B2 => n2952, 
                           ZN => n16891);
   U13654 : INV_X1 port map( A => n16890, ZN => n11176);
   U13655 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2379_port, B2 => n2951, 
                           ZN => n16890);
   U13656 : INV_X1 port map( A => n16889, ZN => n11177);
   U13657 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2378_port, B2 => n2951, 
                           ZN => n16889);
   U13658 : INV_X1 port map( A => n16888, ZN => n11178);
   U13659 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2377_port, B2 => n2951, 
                           ZN => n16888);
   U13660 : INV_X1 port map( A => n16887, ZN => n11179);
   U13661 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2949, B1 => 
                           DataPath_RF_bus_reg_dataout_2376_port, B2 => n2951, 
                           ZN => n16887);
   U13662 : INV_X1 port map( A => n16886, ZN => n11180);
   U13663 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2375_port, B2 => n2951, 
                           ZN => n16886);
   U13664 : INV_X1 port map( A => n16885, ZN => n11181);
   U13665 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2374_port, B2 => n2951, 
                           ZN => n16885);
   U13666 : INV_X1 port map( A => n16884, ZN => n11182);
   U13667 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2373_port, B2 => n2951, 
                           ZN => n16884);
   U13668 : INV_X1 port map( A => n16883, ZN => n11183);
   U13669 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2372_port, B2 => n2951, 
                           ZN => n16883);
   U13670 : INV_X1 port map( A => n16882, ZN => n11184);
   U13671 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2371_port, B2 => n2951, 
                           ZN => n16882);
   U13672 : INV_X1 port map( A => n16881, ZN => n11185);
   U13673 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2370_port, B2 => n2951, 
                           ZN => n16881);
   U13674 : INV_X1 port map( A => n16880, ZN => n11186);
   U13675 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2369_port, B2 => n2951, 
                           ZN => n16880);
   U13676 : INV_X1 port map( A => n16877, ZN => n11187);
   U13677 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2950, B1 => 
                           DataPath_RF_bus_reg_dataout_2368_port, B2 => n2951, 
                           ZN => n16877);
   U13678 : INV_X1 port map( A => n16944, ZN => n11188);
   U13679 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2431_port, B2 => n2959, 
                           ZN => n16944);
   U13680 : INV_X1 port map( A => n16943, ZN => n11189);
   U13681 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2430_port, B2 => n2959, 
                           ZN => n16943);
   U13682 : INV_X1 port map( A => n16942, ZN => n11190);
   U13683 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2429_port, B2 => n2959, 
                           ZN => n16942);
   U13684 : INV_X1 port map( A => n16941, ZN => n11191);
   U13685 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2428_port, B2 => n2959, 
                           ZN => n16941);
   U13686 : INV_X1 port map( A => n16940, ZN => n11192);
   U13687 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2427_port, B2 => n2959, 
                           ZN => n16940);
   U13688 : INV_X1 port map( A => n16939, ZN => n11193);
   U13689 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2426_port, B2 => n2959, 
                           ZN => n16939);
   U13690 : INV_X1 port map( A => n16938, ZN => n11194);
   U13691 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2425_port, B2 => n2959, 
                           ZN => n16938);
   U13692 : INV_X1 port map( A => n16937, ZN => n11195);
   U13693 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2424_port, B2 => n2959, 
                           ZN => n16937);
   U13694 : INV_X1 port map( A => n16936, ZN => n11196);
   U13695 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2423_port, B2 => n2958, 
                           ZN => n16936);
   U13696 : INV_X1 port map( A => n16935, ZN => n11197);
   U13697 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2422_port, B2 => n2958, 
                           ZN => n16935);
   U13698 : INV_X1 port map( A => n16934, ZN => n11198);
   U13699 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2421_port, B2 => n2958, 
                           ZN => n16934);
   U13700 : INV_X1 port map( A => n16933, ZN => n11199);
   U13701 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2954, B1 => 
                           DataPath_RF_bus_reg_dataout_2420_port, B2 => n2958, 
                           ZN => n16933);
   U13702 : INV_X1 port map( A => n16932, ZN => n11200);
   U13703 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2419_port, B2 => n2958, 
                           ZN => n16932);
   U13704 : INV_X1 port map( A => n16931, ZN => n11201);
   U13705 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2418_port, B2 => n2958, 
                           ZN => n16931);
   U13706 : INV_X1 port map( A => n16930, ZN => n11202);
   U13707 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2417_port, B2 => n2958, 
                           ZN => n16930);
   U13708 : INV_X1 port map( A => n16929, ZN => n11203);
   U13709 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2416_port, B2 => n2958, 
                           ZN => n16929);
   U13710 : INV_X1 port map( A => n16928, ZN => n11204);
   U13711 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2415_port, B2 => n2958, 
                           ZN => n16928);
   U13712 : INV_X1 port map( A => n16927, ZN => n11205);
   U13713 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2414_port, B2 => n2958, 
                           ZN => n16927);
   U13714 : INV_X1 port map( A => n16926, ZN => n11206);
   U13715 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2413_port, B2 => n2958, 
                           ZN => n16926);
   U13716 : INV_X1 port map( A => n16925, ZN => n11207);
   U13717 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2412_port, B2 => n2958, 
                           ZN => n16925);
   U13718 : INV_X1 port map( A => n16924, ZN => n11208);
   U13719 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2411_port, B2 => n2957, 
                           ZN => n16924);
   U13720 : INV_X1 port map( A => n16923, ZN => n11209);
   U13721 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2410_port, B2 => n2957, 
                           ZN => n16923);
   U13722 : INV_X1 port map( A => n16922, ZN => n11210);
   U13723 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2409_port, B2 => n2957, 
                           ZN => n16922);
   U13724 : INV_X1 port map( A => n16921, ZN => n11211);
   U13725 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2955, B1 => 
                           DataPath_RF_bus_reg_dataout_2408_port, B2 => n2957, 
                           ZN => n16921);
   U13726 : INV_X1 port map( A => n16920, ZN => n11212);
   U13727 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2407_port, B2 => n2957, 
                           ZN => n16920);
   U13728 : INV_X1 port map( A => n16919, ZN => n11213);
   U13729 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2406_port, B2 => n2957, 
                           ZN => n16919);
   U13730 : INV_X1 port map( A => n16918, ZN => n11214);
   U13731 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2405_port, B2 => n2957, 
                           ZN => n16918);
   U13732 : INV_X1 port map( A => n16917, ZN => n11215);
   U13733 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2404_port, B2 => n2957, 
                           ZN => n16917);
   U13734 : INV_X1 port map( A => n16916, ZN => n11216);
   U13735 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2403_port, B2 => n2957, 
                           ZN => n16916);
   U13736 : INV_X1 port map( A => n16915, ZN => n11217);
   U13737 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2402_port, B2 => n2957, 
                           ZN => n16915);
   U13738 : INV_X1 port map( A => n16914, ZN => n11218);
   U13739 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2401_port, B2 => n2957, 
                           ZN => n16914);
   U13740 : INV_X1 port map( A => n16911, ZN => n11219);
   U13741 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2956, B1 => 
                           DataPath_RF_bus_reg_dataout_2400_port, B2 => n2957, 
                           ZN => n16911);
   U13742 : INV_X1 port map( A => n16978, ZN => n11220);
   U13743 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2463_port, B2 => n2965, 
                           ZN => n16978);
   U13744 : INV_X1 port map( A => n16977, ZN => n11221);
   U13745 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2462_port, B2 => n2965, 
                           ZN => n16977);
   U13746 : INV_X1 port map( A => n16976, ZN => n11222);
   U13747 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2461_port, B2 => n2965, 
                           ZN => n16976);
   U13748 : INV_X1 port map( A => n16975, ZN => n11223);
   U13749 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2460_port, B2 => n2965, 
                           ZN => n16975);
   U13750 : INV_X1 port map( A => n16974, ZN => n11224);
   U13751 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2459_port, B2 => n2965, 
                           ZN => n16974);
   U13752 : INV_X1 port map( A => n16973, ZN => n11225);
   U13753 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2458_port, B2 => n2965, 
                           ZN => n16973);
   U13754 : INV_X1 port map( A => n16972, ZN => n11226);
   U13755 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2457_port, B2 => n2965, 
                           ZN => n16972);
   U13756 : INV_X1 port map( A => n16971, ZN => n11227);
   U13757 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2456_port, B2 => n2965, 
                           ZN => n16971);
   U13758 : INV_X1 port map( A => n16970, ZN => n11228);
   U13759 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2455_port, B2 => n2964, 
                           ZN => n16970);
   U13760 : INV_X1 port map( A => n16969, ZN => n11229);
   U13761 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2454_port, B2 => n2964, 
                           ZN => n16969);
   U13762 : INV_X1 port map( A => n16968, ZN => n11230);
   U13763 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2453_port, B2 => n2964, 
                           ZN => n16968);
   U13764 : INV_X1 port map( A => n16967, ZN => n11231);
   U13765 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2960, B1 => 
                           DataPath_RF_bus_reg_dataout_2452_port, B2 => n2964, 
                           ZN => n16967);
   U13766 : INV_X1 port map( A => n16966, ZN => n11232);
   U13767 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2451_port, B2 => n2964, 
                           ZN => n16966);
   U13768 : INV_X1 port map( A => n16965, ZN => n11233);
   U13769 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2450_port, B2 => n2964, 
                           ZN => n16965);
   U13770 : INV_X1 port map( A => n16964, ZN => n11234);
   U13771 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2449_port, B2 => n2964, 
                           ZN => n16964);
   U13772 : INV_X1 port map( A => n16963, ZN => n11235);
   U13773 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2448_port, B2 => n2964, 
                           ZN => n16963);
   U13774 : INV_X1 port map( A => n16962, ZN => n11236);
   U13775 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2447_port, B2 => n2964, 
                           ZN => n16962);
   U13776 : INV_X1 port map( A => n16961, ZN => n11237);
   U13777 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2446_port, B2 => n2964, 
                           ZN => n16961);
   U13778 : INV_X1 port map( A => n16960, ZN => n11238);
   U13779 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2445_port, B2 => n2964, 
                           ZN => n16960);
   U13780 : INV_X1 port map( A => n16959, ZN => n11239);
   U13781 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2444_port, B2 => n2964, 
                           ZN => n16959);
   U13782 : INV_X1 port map( A => n16958, ZN => n11240);
   U13783 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2443_port, B2 => n2963, 
                           ZN => n16958);
   U13784 : INV_X1 port map( A => n16957, ZN => n11241);
   U13785 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2442_port, B2 => n2963, 
                           ZN => n16957);
   U13786 : INV_X1 port map( A => n16956, ZN => n11242);
   U13787 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2441_port, B2 => n2963, 
                           ZN => n16956);
   U13788 : INV_X1 port map( A => n16955, ZN => n11243);
   U13789 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2961, B1 => 
                           DataPath_RF_bus_reg_dataout_2440_port, B2 => n2963, 
                           ZN => n16955);
   U13790 : INV_X1 port map( A => n16954, ZN => n11244);
   U13791 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2439_port, B2 => n2963, 
                           ZN => n16954);
   U13792 : INV_X1 port map( A => n16953, ZN => n11245);
   U13793 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2438_port, B2 => n2963, 
                           ZN => n16953);
   U13794 : INV_X1 port map( A => n16952, ZN => n11246);
   U13795 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2437_port, B2 => n2963, 
                           ZN => n16952);
   U13796 : INV_X1 port map( A => n16951, ZN => n11247);
   U13797 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2436_port, B2 => n2963, 
                           ZN => n16951);
   U13798 : INV_X1 port map( A => n16950, ZN => n11248);
   U13799 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2435_port, B2 => n2963, 
                           ZN => n16950);
   U13800 : INV_X1 port map( A => n16949, ZN => n11249);
   U13801 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2434_port, B2 => n2963, 
                           ZN => n16949);
   U13802 : INV_X1 port map( A => n16948, ZN => n11250);
   U13803 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2433_port, B2 => n2963, 
                           ZN => n16948);
   U13804 : INV_X1 port map( A => n16945, ZN => n11251);
   U13805 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2962, B1 => 
                           DataPath_RF_bus_reg_dataout_2432_port, B2 => n2963, 
                           ZN => n16945);
   U13806 : INV_X1 port map( A => n17012, ZN => n11252);
   U13807 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2495_port, B2 => n2971, 
                           ZN => n17012);
   U13808 : INV_X1 port map( A => n17011, ZN => n11253);
   U13809 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2494_port, B2 => n2971, 
                           ZN => n17011);
   U13810 : INV_X1 port map( A => n17010, ZN => n11254);
   U13811 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2493_port, B2 => n2971, 
                           ZN => n17010);
   U13812 : INV_X1 port map( A => n17009, ZN => n11255);
   U13813 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2492_port, B2 => n2971, 
                           ZN => n17009);
   U13814 : INV_X1 port map( A => n17008, ZN => n11256);
   U13815 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2491_port, B2 => n2971, 
                           ZN => n17008);
   U13816 : INV_X1 port map( A => n17007, ZN => n11257);
   U13817 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2490_port, B2 => n2971, 
                           ZN => n17007);
   U13818 : INV_X1 port map( A => n17006, ZN => n11258);
   U13819 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2489_port, B2 => n2971, 
                           ZN => n17006);
   U13820 : INV_X1 port map( A => n17005, ZN => n11259);
   U13821 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2488_port, B2 => n2971, 
                           ZN => n17005);
   U13822 : INV_X1 port map( A => n17004, ZN => n11260);
   U13823 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2487_port, B2 => n2970, 
                           ZN => n17004);
   U13824 : INV_X1 port map( A => n17003, ZN => n11261);
   U13825 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2486_port, B2 => n2970, 
                           ZN => n17003);
   U13826 : INV_X1 port map( A => n17002, ZN => n11262);
   U13827 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2485_port, B2 => n2970, 
                           ZN => n17002);
   U13828 : INV_X1 port map( A => n17001, ZN => n11263);
   U13829 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2966, B1 => 
                           DataPath_RF_bus_reg_dataout_2484_port, B2 => n2970, 
                           ZN => n17001);
   U13830 : INV_X1 port map( A => n17000, ZN => n11264);
   U13831 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2483_port, B2 => n2970, 
                           ZN => n17000);
   U13832 : INV_X1 port map( A => n16999, ZN => n11265);
   U13833 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2482_port, B2 => n2970, 
                           ZN => n16999);
   U13834 : INV_X1 port map( A => n16998, ZN => n11266);
   U13835 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2481_port, B2 => n2970, 
                           ZN => n16998);
   U13836 : INV_X1 port map( A => n16997, ZN => n11267);
   U13837 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2480_port, B2 => n2970, 
                           ZN => n16997);
   U13838 : INV_X1 port map( A => n16996, ZN => n11268);
   U13839 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2479_port, B2 => n2970, 
                           ZN => n16996);
   U13840 : INV_X1 port map( A => n16995, ZN => n11269);
   U13841 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2478_port, B2 => n2970, 
                           ZN => n16995);
   U13842 : INV_X1 port map( A => n16994, ZN => n11270);
   U13843 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2477_port, B2 => n2970, 
                           ZN => n16994);
   U13844 : INV_X1 port map( A => n16993, ZN => n11271);
   U13845 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2476_port, B2 => n2970, 
                           ZN => n16993);
   U13846 : INV_X1 port map( A => n16992, ZN => n11272);
   U13847 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2475_port, B2 => n2969, 
                           ZN => n16992);
   U13848 : INV_X1 port map( A => n16991, ZN => n11273);
   U13849 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2474_port, B2 => n2969, 
                           ZN => n16991);
   U13850 : INV_X1 port map( A => n16990, ZN => n11274);
   U13851 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2473_port, B2 => n2969, 
                           ZN => n16990);
   U13852 : INV_X1 port map( A => n16989, ZN => n11275);
   U13853 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2967, B1 => 
                           DataPath_RF_bus_reg_dataout_2472_port, B2 => n2969, 
                           ZN => n16989);
   U13854 : INV_X1 port map( A => n16988, ZN => n11276);
   U13855 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2471_port, B2 => n2969, 
                           ZN => n16988);
   U13856 : INV_X1 port map( A => n16987, ZN => n11277);
   U13857 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2470_port, B2 => n2969, 
                           ZN => n16987);
   U13858 : INV_X1 port map( A => n16986, ZN => n11278);
   U13859 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2469_port, B2 => n2969, 
                           ZN => n16986);
   U13860 : INV_X1 port map( A => n16985, ZN => n11279);
   U13861 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2468_port, B2 => n2969, 
                           ZN => n16985);
   U13862 : INV_X1 port map( A => n16984, ZN => n11280);
   U13863 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2467_port, B2 => n2969, 
                           ZN => n16984);
   U13864 : INV_X1 port map( A => n16983, ZN => n11281);
   U13865 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2466_port, B2 => n2969, 
                           ZN => n16983);
   U13866 : INV_X1 port map( A => n16982, ZN => n11282);
   U13867 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2465_port, B2 => n2969, 
                           ZN => n16982);
   U13868 : INV_X1 port map( A => n16979, ZN => n11283);
   U13869 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2968, B1 => 
                           DataPath_RF_bus_reg_dataout_2464_port, B2 => n2969, 
                           ZN => n16979);
   U13870 : INV_X1 port map( A => n17046, ZN => n11284);
   U13871 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2527_port, B2 => n2977, 
                           ZN => n17046);
   U13872 : INV_X1 port map( A => n17045, ZN => n11285);
   U13873 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2526_port, B2 => n2977, 
                           ZN => n17045);
   U13874 : INV_X1 port map( A => n17044, ZN => n11286);
   U13875 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2525_port, B2 => n2977, 
                           ZN => n17044);
   U13876 : INV_X1 port map( A => n17043, ZN => n11287);
   U13877 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2524_port, B2 => n2977, 
                           ZN => n17043);
   U13878 : INV_X1 port map( A => n17042, ZN => n11288);
   U13879 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2523_port, B2 => n2977, 
                           ZN => n17042);
   U13880 : INV_X1 port map( A => n17041, ZN => n11289);
   U13881 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2522_port, B2 => n2977, 
                           ZN => n17041);
   U13882 : INV_X1 port map( A => n17040, ZN => n11290);
   U13883 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2521_port, B2 => n2977, 
                           ZN => n17040);
   U13884 : INV_X1 port map( A => n17039, ZN => n11291);
   U13885 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2520_port, B2 => n2977, 
                           ZN => n17039);
   U13886 : INV_X1 port map( A => n17038, ZN => n11292);
   U13887 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2519_port, B2 => n2976, 
                           ZN => n17038);
   U13888 : INV_X1 port map( A => n17037, ZN => n11293);
   U13889 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2518_port, B2 => n2976, 
                           ZN => n17037);
   U13890 : INV_X1 port map( A => n17036, ZN => n11294);
   U13891 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2517_port, B2 => n2976, 
                           ZN => n17036);
   U13892 : INV_X1 port map( A => n17035, ZN => n11295);
   U13893 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2972, B1 => 
                           DataPath_RF_bus_reg_dataout_2516_port, B2 => n2976, 
                           ZN => n17035);
   U13894 : INV_X1 port map( A => n17034, ZN => n11296);
   U13895 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2515_port, B2 => n2976, 
                           ZN => n17034);
   U13896 : INV_X1 port map( A => n17033, ZN => n11297);
   U13897 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2514_port, B2 => n2976, 
                           ZN => n17033);
   U13898 : INV_X1 port map( A => n17032, ZN => n11298);
   U13899 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2513_port, B2 => n2976, 
                           ZN => n17032);
   U13900 : INV_X1 port map( A => n17031, ZN => n11299);
   U13901 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2512_port, B2 => n2976, 
                           ZN => n17031);
   U13902 : INV_X1 port map( A => n17030, ZN => n11300);
   U13903 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2511_port, B2 => n2976, 
                           ZN => n17030);
   U13904 : INV_X1 port map( A => n17029, ZN => n11301);
   U13905 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2510_port, B2 => n2976, 
                           ZN => n17029);
   U13906 : INV_X1 port map( A => n17028, ZN => n11302);
   U13907 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2509_port, B2 => n2976, 
                           ZN => n17028);
   U13908 : INV_X1 port map( A => n17027, ZN => n11303);
   U13909 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2508_port, B2 => n2976, 
                           ZN => n17027);
   U13910 : INV_X1 port map( A => n17026, ZN => n11304);
   U13911 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2507_port, B2 => n2975, 
                           ZN => n17026);
   U13912 : INV_X1 port map( A => n17025, ZN => n11305);
   U13913 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2506_port, B2 => n2975, 
                           ZN => n17025);
   U13914 : INV_X1 port map( A => n17024, ZN => n11306);
   U13915 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2505_port, B2 => n2975, 
                           ZN => n17024);
   U13916 : INV_X1 port map( A => n17023, ZN => n11307);
   U13917 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2973, B1 => 
                           DataPath_RF_bus_reg_dataout_2504_port, B2 => n2975, 
                           ZN => n17023);
   U13918 : INV_X1 port map( A => n17022, ZN => n11308);
   U13919 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2503_port, B2 => n2975, 
                           ZN => n17022);
   U13920 : INV_X1 port map( A => n17021, ZN => n11309);
   U13921 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2502_port, B2 => n2975, 
                           ZN => n17021);
   U13922 : INV_X1 port map( A => n17020, ZN => n11310);
   U13923 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2501_port, B2 => n2975, 
                           ZN => n17020);
   U13924 : INV_X1 port map( A => n17019, ZN => n11311);
   U13925 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2500_port, B2 => n2975, 
                           ZN => n17019);
   U13926 : INV_X1 port map( A => n17018, ZN => n11312);
   U13927 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2499_port, B2 => n2975, 
                           ZN => n17018);
   U13928 : INV_X1 port map( A => n17017, ZN => n11313);
   U13929 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2498_port, B2 => n2975, 
                           ZN => n17017);
   U13930 : INV_X1 port map( A => n17016, ZN => n11314);
   U13931 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2497_port, B2 => n2975, 
                           ZN => n17016);
   U13932 : INV_X1 port map( A => n17013, ZN => n11315);
   U13933 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2974, B1 => 
                           DataPath_RF_bus_reg_dataout_2496_port, B2 => n2975, 
                           ZN => n17013);
   U13934 : INV_X1 port map( A => n17080, ZN => n11316);
   U13935 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_31_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2559_port, B2 => n2983, 
                           ZN => n17080);
   U13936 : INV_X1 port map( A => n17079, ZN => n11317);
   U13937 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_30_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2558_port, B2 => n2983, 
                           ZN => n17079);
   U13938 : INV_X1 port map( A => n17078, ZN => n11318);
   U13939 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_29_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2557_port, B2 => n2983, 
                           ZN => n17078);
   U13940 : INV_X1 port map( A => n17077, ZN => n11319);
   U13941 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_28_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2556_port, B2 => n2983, 
                           ZN => n17077);
   U13942 : INV_X1 port map( A => n17076, ZN => n11320);
   U13943 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_27_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2555_port, B2 => n2983, 
                           ZN => n17076);
   U13944 : INV_X1 port map( A => n17075, ZN => n11321);
   U13945 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_26_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2554_port, B2 => n2983, 
                           ZN => n17075);
   U13946 : INV_X1 port map( A => n17074, ZN => n11322);
   U13947 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_25_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2553_port, B2 => n2983, 
                           ZN => n17074);
   U13948 : INV_X1 port map( A => n17073, ZN => n11323);
   U13949 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_24_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2552_port, B2 => n2983, 
                           ZN => n17073);
   U13950 : INV_X1 port map( A => n17072, ZN => n11324);
   U13951 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_23_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2551_port, B2 => n2982, 
                           ZN => n17072);
   U13952 : INV_X1 port map( A => n17071, ZN => n11325);
   U13953 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_22_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2550_port, B2 => n2982, 
                           ZN => n17071);
   U13954 : INV_X1 port map( A => n17070, ZN => n11326);
   U13955 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_21_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2549_port, B2 => n2982, 
                           ZN => n17070);
   U13956 : INV_X1 port map( A => n17069, ZN => n11327);
   U13957 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_20_port,
                           A2 => n2978, B1 => 
                           DataPath_RF_bus_reg_dataout_2548_port, B2 => n2982, 
                           ZN => n17069);
   U13958 : INV_X1 port map( A => n17068, ZN => n11328);
   U13959 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_19_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2547_port, B2 => n2982, 
                           ZN => n17068);
   U13960 : INV_X1 port map( A => n17067, ZN => n11329);
   U13961 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_18_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2546_port, B2 => n2982, 
                           ZN => n17067);
   U13962 : INV_X1 port map( A => n17066, ZN => n11330);
   U13963 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_17_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2545_port, B2 => n2982, 
                           ZN => n17066);
   U13964 : INV_X1 port map( A => n17065, ZN => n11331);
   U13965 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_16_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2544_port, B2 => n2982, 
                           ZN => n17065);
   U13966 : INV_X1 port map( A => n17064, ZN => n11332);
   U13967 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_15_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2543_port, B2 => n2982, 
                           ZN => n17064);
   U13968 : INV_X1 port map( A => n17063, ZN => n11333);
   U13969 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_14_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2542_port, B2 => n2982, 
                           ZN => n17063);
   U13970 : INV_X1 port map( A => n17062, ZN => n11334);
   U13971 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_13_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2541_port, B2 => n2982, 
                           ZN => n17062);
   U13972 : INV_X1 port map( A => n17061, ZN => n11335);
   U13973 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_12_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2540_port, B2 => n2982, 
                           ZN => n17061);
   U13974 : INV_X1 port map( A => n17060, ZN => n11336);
   U13975 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_11_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2539_port, B2 => n2981, 
                           ZN => n17060);
   U13976 : INV_X1 port map( A => n17059, ZN => n11337);
   U13977 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_10_port,
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2538_port, B2 => n2981, 
                           ZN => n17059);
   U13978 : INV_X1 port map( A => n17058, ZN => n11338);
   U13979 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_9_port, 
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2537_port, B2 => n2981, 
                           ZN => n17058);
   U13980 : INV_X1 port map( A => n17057, ZN => n11339);
   U13981 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_8_port, 
                           A2 => n2979, B1 => 
                           DataPath_RF_bus_reg_dataout_2536_port, B2 => n2981, 
                           ZN => n17057);
   U13982 : INV_X1 port map( A => n17056, ZN => n11340);
   U13983 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_7_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2535_port, B2 => n2981, 
                           ZN => n17056);
   U13984 : INV_X1 port map( A => n17055, ZN => n11341);
   U13985 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_6_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2534_port, B2 => n2981, 
                           ZN => n17055);
   U13986 : INV_X1 port map( A => n17054, ZN => n11342);
   U13987 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_5_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2533_port, B2 => n2981, 
                           ZN => n17054);
   U13988 : INV_X1 port map( A => n17053, ZN => n11343);
   U13989 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_4_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2532_port, B2 => n2981, 
                           ZN => n17053);
   U13990 : INV_X1 port map( A => n17052, ZN => n11344);
   U13991 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_3_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2531_port, B2 => n2981, 
                           ZN => n17052);
   U13992 : INV_X1 port map( A => n17051, ZN => n11345);
   U13993 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_2_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2530_port, B2 => n2981, 
                           ZN => n17051);
   U13994 : INV_X1 port map( A => n17050, ZN => n11346);
   U13995 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_1_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2529_port, B2 => n2981, 
                           ZN => n17050);
   U13996 : INV_X1 port map( A => n17047, ZN => n11347);
   U13997 : AOI22_X1 port map( A1 => DataPath_RF_internal_inloc_data_4_0_port, 
                           A2 => n2980, B1 => 
                           DataPath_RF_bus_reg_dataout_2528_port, B2 => n2981, 
                           ZN => n17047);
   U13998 : INV_X1 port map( A => n17122, ZN => n11550);
   U13999 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_30_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_30_port, B2 
                           => n4111, ZN => n17122);
   U14000 : INV_X1 port map( A => n17124, ZN => n11552);
   U14001 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_29_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_29_port, B2 
                           => n4111, ZN => n17124);
   U14002 : INV_X1 port map( A => n17125, ZN => n11553);
   U14003 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_28_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_28_port, B2 
                           => n4111, ZN => n17125);
   U14004 : INV_X1 port map( A => n17126, ZN => n11554);
   U14005 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_27_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_27_port, B2 
                           => n4112, ZN => n17126);
   U14006 : INV_X1 port map( A => n17127, ZN => n11555);
   U14007 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_26_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_26_port, B2 
                           => n4112, ZN => n17127);
   U14008 : INV_X1 port map( A => n17128, ZN => n11556);
   U14009 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_25_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_25_port, B2 
                           => n4112, ZN => n17128);
   U14010 : INV_X1 port map( A => n17129, ZN => n11557);
   U14011 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_24_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_24_port, B2 
                           => n4112, ZN => n17129);
   U14012 : INV_X1 port map( A => n17130, ZN => n11558);
   U14013 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_23_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_23_port, B2 
                           => n4113, ZN => n17130);
   U14014 : INV_X1 port map( A => n17131, ZN => n11559);
   U14015 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_22_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_22_port, B2 
                           => n4113, ZN => n17131);
   U14016 : INV_X1 port map( A => n17132, ZN => n11560);
   U14017 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_21_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_21_port, B2 
                           => n4113, ZN => n17132);
   U14018 : INV_X1 port map( A => n17133, ZN => n11561);
   U14019 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_20_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_20_port, B2 
                           => n4113, ZN => n17133);
   U14020 : INV_X1 port map( A => n17135, ZN => n11563);
   U14021 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_19_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_19_port, B2 =>
                           n4114, ZN => n17135);
   U14022 : INV_X1 port map( A => n17136, ZN => n11564);
   U14023 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_18_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_18_port, B2 =>
                           n4114, ZN => n17136);
   U14024 : INV_X1 port map( A => n17137, ZN => n11565);
   U14025 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_17_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_17_port, B2 =>
                           n4114, ZN => n17137);
   U14026 : INV_X1 port map( A => n17138, ZN => n11566);
   U14027 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_16_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_16_port, B2 =>
                           n4115, ZN => n17138);
   U14028 : INV_X1 port map( A => n17139, ZN => n11567);
   U14029 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_15_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_15_port, B2 =>
                           n4115, ZN => n17139);
   U14030 : INV_X1 port map( A => n17140, ZN => n11568);
   U14031 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_14_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_14_port, B2 =>
                           n4115, ZN => n17140);
   U14032 : INV_X1 port map( A => n17141, ZN => n11569);
   U14033 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_13_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_13_port, B2 =>
                           n4115, ZN => n17141);
   U14034 : INV_X1 port map( A => n17142, ZN => n11570);
   U14035 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_12_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_12_port, B2 =>
                           n4116, ZN => n17142);
   U14036 : INV_X1 port map( A => n17143, ZN => n11571);
   U14037 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_11_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_11_port, B2 =>
                           n4116, ZN => n17143);
   U14038 : INV_X1 port map( A => n17144, ZN => n11572);
   U14039 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_10_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_10_port, B2 =>
                           n4116, ZN => n17144);
   U14040 : INV_X1 port map( A => n17123, ZN => n11551);
   U14041 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_2_port, A2 => 
                           n4108, B1 => DataPath_i_REG_MEM_ALUOUT_2_port, B2 =>
                           n4111, ZN => n17123);
   U14042 : INV_X1 port map( A => n17134, ZN => n11562);
   U14043 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_1_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_1_port, B2 => 
                           n4114, ZN => n17134);
   U14044 : INV_X1 port map( A => n17145, ZN => n11573);
   U14045 : AOI22_X1 port map( A1 => DataPath_i_REG_LDSTR_OUT_0_port, A2 => 
                           n256, B1 => DataPath_i_REG_MEM_ALUOUT_0_port, B2 => 
                           n4116, ZN => n17145);
   U14046 : INV_X1 port map( A => n14302, ZN => n8748);
   U14047 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_7_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_7_port, B2 => n2495, ZN => 
                           n14302);
   U14048 : INV_X1 port map( A => n14301, ZN => n8749);
   U14049 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_6_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_6_port, B2 => n2495, ZN => 
                           n14301);
   U14050 : INV_X1 port map( A => n14300, ZN => n8750);
   U14051 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_5_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_5_port, B2 => n2495, ZN => 
                           n14300);
   U14052 : INV_X1 port map( A => n14299, ZN => n8751);
   U14053 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_4_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_4_port, B2 => n2495, ZN => 
                           n14299);
   U14054 : INV_X1 port map( A => n14298, ZN => n8752);
   U14055 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_3_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_3_port, B2 => n2495, ZN => 
                           n14298);
   U14056 : INV_X1 port map( A => n14297, ZN => n8753);
   U14057 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_2_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_2_port, B2 => n2495, ZN => 
                           n14297);
   U14058 : INV_X1 port map( A => n14296, ZN => n8754);
   U14059 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_1_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_1_port, B2 => n2495, ZN => 
                           n14296);
   U14060 : INV_X1 port map( A => n14293, ZN => n8755);
   U14061 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_0_port, A2 => n2494, B1 => 
                           DataPath_i_REG_LDSTR_OUT_0_port, B2 => n2495, ZN => 
                           n14293);
   U14062 : INV_X1 port map( A => n14310, ZN => n8740);
   U14063 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_15_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_15_port, B2 => n2496, ZN =>
                           n14310);
   U14064 : INV_X1 port map( A => n14309, ZN => n8741);
   U14065 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_14_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_14_port, B2 => n2496, ZN =>
                           n14309);
   U14066 : INV_X1 port map( A => n14308, ZN => n8742);
   U14067 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_13_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_13_port, B2 => n2496, ZN =>
                           n14308);
   U14068 : INV_X1 port map( A => n14307, ZN => n8743);
   U14069 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_12_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_12_port, B2 => n2496, ZN =>
                           n14307);
   U14070 : INV_X1 port map( A => n14306, ZN => n8744);
   U14071 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_11_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_11_port, B2 => n2495, ZN =>
                           n14306);
   U14072 : INV_X1 port map( A => n14305, ZN => n8745);
   U14073 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_10_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_10_port, B2 => n2495, ZN =>
                           n14305);
   U14074 : INV_X1 port map( A => n14304, ZN => n8746);
   U14075 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_9_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_9_port, B2 => n2495, ZN => 
                           n14304);
   U14076 : INV_X1 port map( A => n14303, ZN => n8747);
   U14077 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_8_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_8_port, B2 => n2495, ZN => 
                           n14303);
   U14078 : INV_X1 port map( A => n14317, ZN => n8733);
   U14079 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_22_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_22_port, B2 => n2496, ZN =>
                           n14317);
   U14080 : INV_X1 port map( A => n14316, ZN => n8734);
   U14081 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_21_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_21_port, B2 => n2496, ZN =>
                           n14316);
   U14082 : INV_X1 port map( A => n14315, ZN => n8735);
   U14083 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_20_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_20_port, B2 => n2496, ZN =>
                           n14315);
   U14084 : INV_X1 port map( A => n14314, ZN => n8736);
   U14085 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_19_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_19_port, B2 => n2496, ZN =>
                           n14314);
   U14086 : INV_X1 port map( A => n14313, ZN => n8737);
   U14087 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_18_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_18_port, B2 => n2496, ZN =>
                           n14313);
   U14088 : INV_X1 port map( A => n14312, ZN => n8738);
   U14089 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_17_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_17_port, B2 => n2496, ZN =>
                           n14312);
   U14090 : INV_X1 port map( A => n14311, ZN => n8739);
   U14091 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_16_port, A2 => n2493, B1 => 
                           DataPath_i_REG_LDSTR_OUT_16_port, B2 => n2496, ZN =>
                           n14311);
   U14092 : INV_X1 port map( A => n14326, ZN => n8724);
   U14093 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_31_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_31_port, B2 => n2497, ZN =>
                           n14326);
   U14094 : INV_X1 port map( A => n14325, ZN => n8725);
   U14095 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_30_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_30_port, B2 => n2497, ZN =>
                           n14325);
   U14096 : INV_X1 port map( A => n14324, ZN => n8726);
   U14097 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_29_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_29_port, B2 => n2497, ZN =>
                           n14324);
   U14098 : INV_X1 port map( A => n14323, ZN => n8727);
   U14099 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_28_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_28_port, B2 => n2497, ZN =>
                           n14323);
   U14100 : INV_X1 port map( A => n14322, ZN => n8728);
   U14101 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_27_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_27_port, B2 => n2497, ZN =>
                           n14322);
   U14102 : INV_X1 port map( A => n14321, ZN => n8729);
   U14103 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_26_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_26_port, B2 => n2497, ZN =>
                           n14321);
   U14104 : INV_X1 port map( A => n14320, ZN => n8730);
   U14105 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_25_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_25_port, B2 => n2497, ZN =>
                           n14320);
   U14106 : INV_X1 port map( A => n14319, ZN => n8731);
   U14107 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_24_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_24_port, B2 => n2497, ZN =>
                           n14319);
   U14108 : INV_X1 port map( A => n14318, ZN => n8732);
   U14109 : AOI22_X1 port map( A1 => DRAM_DATA_OUT_23_port, A2 => n2492, B1 => 
                           DataPath_i_REG_LDSTR_OUT_23_port, B2 => n2496, ZN =>
                           n14318);
   U14110 : AOI222_X1 port map( A1 => DataPath_WRF_CUhw_N109, A2 => n3265, B1 
                           => DataPath_WRF_CUhw_N109, B2 => n3262, C1 => 
                           DataPath_WRF_CUhw_N109, C2 => n2475, ZN => 
                           DataPath_WRF_CUhw_n145);
   U14111 : AOI222_X1 port map( A1 => DataPath_WRF_CUhw_curr_addr_1_port, A2 =>
                           n3266, B1 => DataPath_WRF_CUhw_curr_addr_1_port, B2 
                           => n3263, C1 => DataPath_WRF_CUhw_curr_addr_1_port, 
                           C2 => n2475, ZN => DataPath_WRF_CUhw_n144);
   U14112 : AOI222_X1 port map( A1 => n304, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N111, B2 => n3262, C1 => n412, C2 
                           => n2476, ZN => DataPath_WRF_CUhw_n143);
   U14113 : XNOR2_X1 port map( A => n1855, B => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => 
                           DataPath_WRF_CUhw_N111);
   U14114 : NAND2_X1 port map( A1 => i_ALU_OP_0_port, A2 => i_ALU_OP_1_port, ZN
                           => n8140);
   U14115 : NAND2_X1 port map( A1 => i_ADD_WB_4_port, A2 => i_ADD_WB_3_port, ZN
                           => DataPath_RF_DEC_n17);
   U14116 : NAND2_X1 port map( A1 => i_ADD_WB_4_port, A2 => n11601, ZN => 
                           DataPath_RF_DEC_n16);
   U14117 : NAND2_X1 port map( A1 => i_ADD_WB_3_port, A2 => n11602, ZN => 
                           DataPath_RF_DEC_n15);
   U14118 : OAI221_X1 port map( B1 => DataPath_i_LGET_0_port, B2 => 
                           DataPath_SETCMP_n4, C1 => DataPath_i_LGET_0_port, C2
                           => DataPath_SETCMP_n5, A => DataPath_SETCMP_n6, ZN 
                           => DataPath_i_SETCMP_OUT_0_port);
   U14119 : OR2_X1 port map( A1 => i_SEL_LGET_0_port, A2 => i_SEL_LGET_1_port, 
                           ZN => DataPath_SETCMP_n5);
   U14120 : AOI21_X1 port map( B1 => DataPath_i_LGET_1_port, B2 => 
                           DataPath_SETCMP_n7, A => DataPath_SETCMP_n8, ZN => 
                           DataPath_SETCMP_n6);
   U14121 : AOI22_X1 port map( A1 => DRAM_DATA_IN(18), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_18_port, B2 => 
                           n4124, ZN => n17104);
   U14122 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n46);
   U14123 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n49);
   U14124 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n47);
   U14125 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n48);
   U14126 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n36);
   U14127 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n37);
   U14128 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n40);
   U14129 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n39);
   U14130 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n38);
   U14131 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n41);
   U14132 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n43);
   U14133 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n42);
   U14134 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n44);
   U14135 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n50);
   U14136 : AOI22_X1 port map( A1 => DRAM_DATA_IN(23), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_23_port, B2 => 
                           n4123, ZN => n17098);
   U14137 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_n52, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, B1 => 
                           n11446, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n45);
   U14138 : AOI22_X1 port map( A1 => DRAM_DATA_IN(31), A2 => n4118, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_31_port, B2 => n4120,
                           ZN => n17089);
   U14139 : AOI22_X1 port map( A1 => DRAM_DATA_IN(15), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_15_port, B2 => 
                           n4125, ZN => n17107);
   U14140 : AOI22_X1 port map( A1 => DRAM_DATA_IN(10), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_10_port, B2 => 
                           n4126, ZN => n17112);
   U14141 : AOI22_X1 port map( A1 => DRAM_DATA_IN(11), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_11_port, B2 => 
                           n4126, ZN => n17111);
   U14142 : AOI22_X1 port map( A1 => DRAM_DATA_IN(12), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_12_port, B2 => 
                           n4126, ZN => n17110);
   U14143 : AOI22_X1 port map( A1 => DRAM_DATA_IN(14), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_14_port, B2 => 
                           n4125, ZN => n17108);
   U14144 : AOI22_X1 port map( A1 => DRAM_DATA_IN(8), A2 => n4118, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_8_port, B2 => n4119, 
                           ZN => n17083);
   U14145 : AOI22_X1 port map( A1 => n4118, A2 => DRAM_DATA_IN(9), B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_9_port, B2 => n4124, 
                           ZN => n17082);
   U14146 : AOI22_X1 port map( A1 => DRAM_DATA_IN(13), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_13_port, B2 => 
                           n4126, ZN => n17109);
   U14147 : AOI22_X1 port map( A1 => DRAM_DATA_IN(16), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_16_port, B2 => 
                           n4125, ZN => n17106);
   U14148 : AOI22_X1 port map( A1 => DRAM_DATA_IN(17), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_17_port, B2 => 
                           n4125, ZN => n17105);
   U14149 : AOI22_X1 port map( A1 => DRAM_DATA_IN(19), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_19_port, B2 => 
                           n4124, ZN => n17103);
   U14150 : AOI22_X1 port map( A1 => DRAM_DATA_IN(20), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_20_port, B2 => 
                           n4123, ZN => n17101);
   U14151 : NOR2_X1 port map( A1 => CU_I_n98, A2 => CU_I_n71, ZN => i_EN3);
   U14152 : AOI22_X1 port map( A1 => DRAM_DATA_IN(21), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_21_port, B2 => 
                           n4123, ZN => n17100);
   U14153 : AOI22_X1 port map( A1 => DRAM_DATA_IN(22), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_22_port, B2 => 
                           n4123, ZN => n17099);
   U14154 : OAI221_X1 port map( B1 => n12952, B2 => n12953, C1 => n8647, C2 => 
                           n12950, A => n12954, ZN => n12979);
   U14155 : NAND4_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_N61, A2 => n11607,
                           A3 => n4143, A4 => n12955, ZN => n12954);
   U14156 : OAI221_X1 port map( B1 => DataPath_RF_PUSH_ADDRGEN_n27, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_n28, C1 => n8648, C2 => 
                           DataPath_RF_PUSH_ADDRGEN_n22, A => 
                           DataPath_RF_PUSH_ADDRGEN_n29, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n54);
   U14157 : NAND4_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_N61, A2 => n11597
                           , A3 => n4143, A4 => DataPath_RF_PUSH_ADDRGEN_n30, 
                           ZN => DataPath_RF_PUSH_ADDRGEN_n29);
   U14158 : OAI22_X1 port map( A1 => n4151, A2 => DataPath_WRF_CUhw_n28, B1 => 
                           n11468, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_10_port);
   U14159 : OAI22_X1 port map( A1 => n4143, A2 => DataPath_WRF_CUhw_n29, B1 => 
                           n11469, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_9_port);
   U14160 : OAI22_X1 port map( A1 => n4144, A2 => DataPath_WRF_CUhw_n30, B1 => 
                           n11470, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_8_port);
   U14161 : OAI22_X1 port map( A1 => n4147, A2 => DataPath_WRF_CUhw_n31, B1 => 
                           n11471, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_7_port);
   U14162 : OAI22_X1 port map( A1 => n4144, A2 => DataPath_WRF_CUhw_n32, B1 => 
                           n11472, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_6_port);
   U14163 : OAI22_X1 port map( A1 => n4144, A2 => DataPath_WRF_CUhw_n33, B1 => 
                           n11473, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_5_port);
   U14164 : OAI22_X1 port map( A1 => n4144, A2 => DataPath_WRF_CUhw_n34, B1 => 
                           n11474, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_4_port);
   U14165 : OAI22_X1 port map( A1 => n4145, A2 => DataPath_WRF_CUhw_n7, B1 => 
                           n11447, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_31_port);
   U14166 : OAI22_X1 port map( A1 => n4145, A2 => DataPath_WRF_CUhw_n8, B1 => 
                           n11448, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_30_port);
   U14167 : OAI22_X1 port map( A1 => n4146, A2 => DataPath_WRF_CUhw_n9, B1 => 
                           n11449, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_29_port);
   U14168 : OAI22_X1 port map( A1 => n4146, A2 => DataPath_WRF_CUhw_n10, B1 => 
                           n11450, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_28_port);
   U14169 : OAI22_X1 port map( A1 => n4146, A2 => DataPath_WRF_CUhw_n11, B1 => 
                           n11451, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_27_port);
   U14170 : OAI22_X1 port map( A1 => n4146, A2 => DataPath_WRF_CUhw_n12, B1 => 
                           n11452, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_26_port);
   U14171 : OAI22_X1 port map( A1 => n4147, A2 => DataPath_WRF_CUhw_n13, B1 => 
                           n11453, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_25_port);
   U14172 : OAI22_X1 port map( A1 => n4147, A2 => DataPath_WRF_CUhw_n14, B1 => 
                           n11454, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_24_port);
   U14173 : OAI22_X1 port map( A1 => n4147, A2 => DataPath_WRF_CUhw_n15, B1 => 
                           n11455, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_23_port);
   U14174 : OAI22_X1 port map( A1 => n4148, A2 => DataPath_WRF_CUhw_n16, B1 => 
                           n11456, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_22_port);
   U14175 : OAI22_X1 port map( A1 => n4148, A2 => DataPath_WRF_CUhw_n17, B1 => 
                           n11457, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_21_port);
   U14176 : OAI22_X1 port map( A1 => n4148, A2 => DataPath_WRF_CUhw_n18, B1 => 
                           n11458, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_20_port);
   U14177 : OAI22_X1 port map( A1 => n4149, A2 => DataPath_WRF_CUhw_n19, B1 => 
                           n11459, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_19_port);
   U14178 : OAI22_X1 port map( A1 => n4149, A2 => DataPath_WRF_CUhw_n20, B1 => 
                           n11460, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_18_port);
   U14179 : OAI22_X1 port map( A1 => n4149, A2 => DataPath_WRF_CUhw_n21, B1 => 
                           n11461, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_17_port);
   U14180 : OAI22_X1 port map( A1 => n4149, A2 => DataPath_WRF_CUhw_n22, B1 => 
                           n11462, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_16_port);
   U14181 : OAI22_X1 port map( A1 => n4150, A2 => DataPath_WRF_CUhw_n23, B1 => 
                           n11463, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_15_port);
   U14182 : OAI22_X1 port map( A1 => n4150, A2 => DataPath_WRF_CUhw_n24, B1 => 
                           n11464, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_14_port);
   U14183 : OAI22_X1 port map( A1 => n4150, A2 => DataPath_WRF_CUhw_n25, B1 => 
                           n11465, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_13_port);
   U14184 : OAI22_X1 port map( A1 => n4151, A2 => DataPath_WRF_CUhw_n26, B1 => 
                           n11466, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_12_port);
   U14185 : OAI22_X1 port map( A1 => n4145, A2 => DataPath_WRF_CUhw_n35, B1 => 
                           n11475, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_3_port);
   U14186 : OAI22_X1 port map( A1 => n4145, A2 => DataPath_WRF_CUhw_n36, B1 => 
                           n11476, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_2_port);
   U14187 : OAI22_X1 port map( A1 => n4148, A2 => DataPath_WRF_CUhw_n37, B1 => 
                           n11477, B2 => n4155, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_1_port);
   U14188 : OAI22_X1 port map( A1 => n4143, A2 => DataPath_WRF_CUhw_n38, B1 => 
                           n11478, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_0_port);
   U14189 : OAI22_X1 port map( A1 => n4150, A2 => DataPath_WRF_CUhw_n27, B1 => 
                           n11467, B2 => n4156, ZN => 
                           DataPath_i_RF_BUS_FROM_RF_CU_11_port);
   U14190 : AOI21_X1 port map( B1 => DataPath_RF_PUSH_ADDRGEN_n52, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, A => 
                           n11596, ZN => DataPath_RF_PUSH_ADDRGEN_n51);
   U14191 : INV_X1 port map( A => DataPath_RF_PUSH_ADDRGEN_n28, ZN => n11596);
   U14192 : XNOR2_X1 port map( A => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port,
                           B => DataPath_RF_PUSH_ADDRGEN_n20, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n28);
   U14193 : XNOR2_X1 port map( A => DataPath_RF_POP_ADDRGEN_curr_state_0_port, 
                           B => n12949, ZN => n12953);
   U14194 : OAI22_X1 port map( A1 => n11480, A2 => n4106, B1 => CU_I_n22, B2 =>
                           n11481, ZN => CU_I_n148);
   U14195 : AOI21_X1 port map( B1 => DataPath_n2, B2 => DataPath_n3, A => n2282
                           , ZN => DataPath_i_WF);
   U14196 : NOR2_X1 port map( A1 => i_ADD_WB_1_port, A2 => i_ADD_WB_0_port, ZN 
                           => DataPath_n2);
   U14197 : NOR3_X1 port map( A1 => i_ADD_WB_2_port, A2 => i_ADD_WB_4_port, A3 
                           => i_ADD_WB_3_port, ZN => DataPath_n3);
   U14198 : OAI22_X1 port map( A1 => DRAM_READNOTWRITE_port, A2 => n4106, B1 =>
                           CU_I_n105, B2 => CU_I_n22, ZN => CU_I_n136);
   U14199 : OAI22_X1 port map( A1 => CU_I_n104, A2 => n4106, B1 => CU_I_n103, 
                           B2 => CU_I_n22, ZN => CU_I_n137);
   U14200 : OAI22_X1 port map( A1 => CU_I_n102, A2 => n4106, B1 => CU_I_n101, 
                           B2 => CU_I_n22, ZN => CU_I_n138);
   U14201 : OAI22_X1 port map( A1 => n11579, A2 => n4106, B1 => CU_I_n99, B2 =>
                           CU_I_n22, ZN => CU_I_n139);
   U14202 : OAI22_X1 port map( A1 => CU_I_n111, A2 => n4106, B1 => CU_I_n110, 
                           B2 => CU_I_n22, ZN => CU_I_n141);
   U14203 : OAI22_X1 port map( A1 => CU_I_n113, A2 => n4106, B1 => CU_I_n112, 
                           B2 => CU_I_n22, ZN => CU_I_n142);
   U14204 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n31, B1 => 
                           n3261, B2 => n11471, ZN => DataPath_WRF_CUhw_n163);
   U14205 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n32, B1 => 
                           n3261, B2 => n11472, ZN => DataPath_WRF_CUhw_n162);
   U14206 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n33, B1 => 
                           n3261, B2 => n11473, ZN => DataPath_WRF_CUhw_n161);
   U14207 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n34, B1 => 
                           n3261, B2 => n11474, ZN => DataPath_WRF_CUhw_n160);
   U14208 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n35, B1 => 
                           n3261, B2 => n11475, ZN => DataPath_WRF_CUhw_n159);
   U14209 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n36, B1 => 
                           n3261, B2 => n11476, ZN => DataPath_WRF_CUhw_n158);
   U14210 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n37, B1 => 
                           n3261, B2 => n11477, ZN => DataPath_WRF_CUhw_n157);
   U14211 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n38, B1 => 
                           n3261, B2 => n11478, ZN => DataPath_WRF_CUhw_n156);
   U14212 : OAI22_X1 port map( A1 => n8647, A2 => n12949, B1 => n12951, B2 => 
                           n12952, ZN => n12978);
   U14213 : OAI22_X1 port map( A1 => n8648, A2 => DataPath_RF_PUSH_ADDRGEN_n20,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n26, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_n27, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n53);
   U14214 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n12905, 
                           B1 => DataPath_RF_c_swin_3_port, B2 => n12906, ZN =>
                           n12907);
   U14215 : AOI22_X1 port map( A1 => DataPath_RF_c_win_3_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n6, B1 => 
                           DataPath_RF_c_win_3_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n8);
   U14216 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_2_port, A2 => n12905, 
                           B1 => DataPath_RF_c_swin_2_port, B2 => n12906, ZN =>
                           n12909);
   U14217 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_1_port, A2 => n12905, 
                           B1 => DataPath_RF_c_swin_1_port, B2 => n12906, ZN =>
                           n12911);
   U14218 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_0_port, A2 => n12905, 
                           B1 => DataPath_RF_c_swin_0_port, B2 => n12906, ZN =>
                           n12913);
   U14219 : AOI22_X1 port map( A1 => DataPath_RF_c_win_2_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n6, B1 => 
                           DataPath_RF_c_win_2_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n10);
   U14220 : AOI22_X1 port map( A1 => DataPath_RF_c_win_1_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n6, B1 => 
                           DataPath_RF_c_win_1_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n12);
   U14221 : AOI22_X1 port map( A1 => DataPath_RF_c_win_0_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n6, B1 => 
                           DataPath_RF_c_win_0_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n7, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n14);
   U14222 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n7, B1 => 
                           n3259, B2 => n11447, ZN => DataPath_WRF_CUhw_n187);
   U14223 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n8, B1 => 
                           n3259, B2 => n11448, ZN => DataPath_WRF_CUhw_n186);
   U14224 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n9, B1 => 
                           n3259, B2 => n11449, ZN => DataPath_WRF_CUhw_n185);
   U14225 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n10, B1 => 
                           n3259, B2 => n11450, ZN => DataPath_WRF_CUhw_n184);
   U14226 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n11, B1 => 
                           n3259, B2 => n11451, ZN => DataPath_WRF_CUhw_n183);
   U14227 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n12, B1 => 
                           n3259, B2 => n11452, ZN => DataPath_WRF_CUhw_n182);
   U14228 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n13, B1 => 
                           n3259, B2 => n11453, ZN => DataPath_WRF_CUhw_n181);
   U14229 : OAI22_X1 port map( A1 => n3258, A2 => DataPath_WRF_CUhw_n14, B1 => 
                           n3259, B2 => n11454, ZN => DataPath_WRF_CUhw_n180);
   U14230 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n15, B1 => 
                           n3259, B2 => n11455, ZN => DataPath_WRF_CUhw_n179);
   U14231 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n16, B1 => 
                           n3259, B2 => n11456, ZN => DataPath_WRF_CUhw_n178);
   U14232 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n17, B1 => 
                           n3259, B2 => n11457, ZN => DataPath_WRF_CUhw_n177);
   U14233 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n18, B1 => 
                           n3259, B2 => n11458, ZN => DataPath_WRF_CUhw_n176);
   U14234 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n19, B1 => 
                           n3260, B2 => n11459, ZN => DataPath_WRF_CUhw_n175);
   U14235 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n20, B1 => 
                           n3260, B2 => n11460, ZN => DataPath_WRF_CUhw_n174);
   U14236 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n21, B1 => 
                           n3260, B2 => n11461, ZN => DataPath_WRF_CUhw_n173);
   U14237 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n22, B1 => 
                           n3260, B2 => n11462, ZN => DataPath_WRF_CUhw_n172);
   U14238 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n23, B1 => 
                           n3260, B2 => n11463, ZN => DataPath_WRF_CUhw_n171);
   U14239 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n24, B1 => 
                           n3260, B2 => n11464, ZN => DataPath_WRF_CUhw_n170);
   U14240 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n25, B1 => 
                           n3260, B2 => n11465, ZN => DataPath_WRF_CUhw_n169);
   U14241 : OAI22_X1 port map( A1 => n3257, A2 => DataPath_WRF_CUhw_n26, B1 => 
                           n3260, B2 => n11466, ZN => DataPath_WRF_CUhw_n168);
   U14242 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n27, B1 => 
                           n3260, B2 => n11467, ZN => DataPath_WRF_CUhw_n167);
   U14243 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n28, B1 => 
                           n3260, B2 => n11468, ZN => DataPath_WRF_CUhw_n166);
   U14244 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n29, B1 => 
                           n3260, B2 => n11469, ZN => DataPath_WRF_CUhw_n165);
   U14245 : OAI22_X1 port map( A1 => n3256, A2 => DataPath_WRF_CUhw_n30, B1 => 
                           n3260, B2 => n11470, ZN => DataPath_WRF_CUhw_n164);
   U14246 : NAND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_state_1_port, A2 =>
                           DataPath_WRF_CUhw_n73, ZN => DataPath_WRF_CUhw_n150)
                           ;
   U14247 : NAND2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port
                           , A2 => DataPath_RF_PUSH_ADDRGEN_n20, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_n26);
   U14248 : NAND2_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_state_0_port,
                           A2 => n12949, ZN => n12951);
   U14249 : AOI21_X1 port map( B1 => DataPath_SETCMP_n4, B2 => 
                           DataPath_SETCMP_n9, A => DataPath_i_LGET_1_port, ZN 
                           => DataPath_SETCMP_n8);
   U14250 : NOR3_X1 port map( A1 => CU_I_n71, A2 => CU_I_n111, A3 => n4157, ZN 
                           => CU_I_N50);
   U14251 : NOR3_X1 port map( A1 => CU_I_n71, A2 => CU_I_n113, A3 => n4157, ZN 
                           => CU_I_N49);
   U14252 : AND2_X1 port map( A1 => DataPath_WRF_CUhw_curr_state_1_port, A2 => 
                           DataPath_WRF_CUhw_curr_state_0_port, ZN => 
                           DataPath_WRF_CUhw_n148);
   U14253 : OAI21_X1 port map( B1 => CU_I_n140, B2 => CU_I_n22, A => n4107, ZN 
                           => CU_I_n157);
   U14254 : INV_X1 port map( A => n17097, ZN => n11364);
   U14255 : AOI22_X1 port map( A1 => DRAM_DATA_IN(24), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_24_port, B2 => 
                           n4122, ZN => n17097);
   U14256 : INV_X1 port map( A => n17094, ZN => n11358);
   U14257 : AOI22_X1 port map( A1 => DRAM_DATA_IN(27), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_27_port, B2 => 
                           n4122, ZN => n17094);
   U14258 : INV_X1 port map( A => n17093, ZN => n11356);
   U14259 : AOI22_X1 port map( A1 => DRAM_DATA_IN(28), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_28_port, B2 => 
                           n4121, ZN => n17093);
   U14260 : INV_X1 port map( A => n17092, ZN => n11354);
   U14261 : AOI22_X1 port map( A1 => DRAM_DATA_IN(29), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_29_port, B2 => 
                           n4121, ZN => n17092);
   U14262 : INV_X1 port map( A => n17090, ZN => n11352);
   U14263 : AOI22_X1 port map( A1 => DRAM_DATA_IN(30), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_30_port, B2 => 
                           n4121, ZN => n17090);
   U14264 : INV_X1 port map( A => n17095, ZN => n11360);
   U14265 : AOI22_X1 port map( A1 => DRAM_DATA_IN(26), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_26_port, B2 => 
                           n4122, ZN => n17095);
   U14266 : INV_X1 port map( A => n17096, ZN => n11362);
   U14267 : AOI22_X1 port map( A1 => DRAM_DATA_IN(25), A2 => i_DATAMEM_RM, B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_25_port, B2 => 
                           n4122, ZN => n17096);
   U14268 : BUF_X1 port map( A => DataPath_RF_c_win_4_port, Z => n3267);
   U14269 : BUF_X1 port map( A => DataPath_RF_c_win_4_port, Z => n3268);
   U14270 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_29_port, A2 => n4265,
                           ZN => n1992);
   U14271 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_28_port, A2 => n4260,
                           ZN => n1993);
   U14272 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_27_port, A2 => n4258,
                           ZN => n1994);
   U14273 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_26_port, A2 => n4259,
                           ZN => n1995);
   U14274 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_25_port, A2 => n4263,
                           ZN => n1996);
   U14275 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_24_port, A2 => n4263,
                           ZN => n1997);
   U14276 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_23_port, A2 => n4264,
                           ZN => n1998);
   U14277 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_22_port, A2 => n4265,
                           ZN => n1999);
   U14278 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_21_port, A2 => n4264,
                           ZN => n2000);
   U14279 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_20_port, A2 => n4261,
                           ZN => n2001);
   U14280 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_19_port, A2 => n4262,
                           ZN => n2002);
   U14281 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_18_port, A2 => n4263,
                           ZN => n2003);
   U14282 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_17_port, A2 => n4261,
                           ZN => n2004);
   U14283 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_16_port, A2 => n4265,
                           ZN => n2005);
   U14284 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_15_port, A2 => n4264,
                           ZN => n2006);
   U14285 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_14_port, A2 => n4261,
                           ZN => n2007);
   U14286 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_13_port, A2 => n4262,
                           ZN => n2008);
   U14287 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_12_port, A2 => n4257,
                           ZN => n2009);
   U14288 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_11_port, A2 => n4264,
                           ZN => n2010);
   U14289 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_10_port, A2 => n4260,
                           ZN => n2011);
   U14290 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_9_port, A2 => n4258, 
                           ZN => n2012);
   U14291 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_8_port, A2 => n4259, 
                           ZN => n2013);
   U14292 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_7_port, A2 => n4263, 
                           ZN => n2014);
   U14293 : NOR2_X1 port map( A1 => CU_I_n109, A2 => n4107, ZN => CU_I_n126);
   U14294 : NOR2_X1 port map( A1 => CU_I_n105, A2 => n4107, ZN => CU_I_n129);
   U14295 : NOR2_X1 port map( A1 => CU_I_n103, A2 => n4107, ZN => CU_I_n130);
   U14296 : NOR2_X1 port map( A1 => CU_I_n101, A2 => n4107, ZN => CU_I_n131);
   U14297 : NOR2_X1 port map( A1 => CU_I_n99, A2 => n4107, ZN => CU_I_n132);
   U14298 : NOR2_X1 port map( A1 => CU_I_n140, A2 => n4107, ZN => CU_I_n133);
   U14299 : NOR2_X1 port map( A1 => CU_I_n110, A2 => n4107, ZN => CU_I_n134);
   U14300 : NOR2_X1 port map( A1 => CU_I_n112, A2 => n4107, ZN => CU_I_n135);
   U14301 : NOR2_X1 port map( A1 => n4202, A2 => DataPath_WRF_CUhw_n152, ZN => 
                           DataPath_WRF_CUhw_N144_port);
   U14302 : AOI221_X1 port map( B1 => n3264, B2 => DataPath_RF_n10, C1 => 
                           DataPath_WRF_CUhw_n153, C2 => DataPath_WRF_CUhw_n154
                           , A => DataPath_WRF_CUhw_n155, ZN => 
                           DataPath_WRF_CUhw_n152);
   U14303 : NAND2_X1 port map( A1 => DataPath_WRF_CUhw_n73, A2 => n12957, ZN =>
                           DataPath_WRF_CUhw_n153);
   U14304 : OAI22_X1 port map( A1 => DataPath_WRF_CUhw_curr_state_1_port, A2 =>
                           DataPath_WRF_CUhw_curr_state_0_port, B1 => 
                           DataPath_WRF_CUhw_n150, B2 => n11400, ZN => 
                           DataPath_WRF_CUhw_n155);
   U14305 : AOI222_X1 port map( A1 => n309, A2 => n3265, B1 => 
                           DataPath_WRF_CUhw_N112_port, B2 => n3262, C1 => n420
                           , C2 => n2477, ZN => DataPath_WRF_CUhw_n142);
   U14306 : XNOR2_X1 port map( A => DataPath_WRF_CUhw_curr_addr_3_port, B => 
                           DataPath_WRF_CUhw_sub_85_aco_carry_3_port, ZN => 
                           DataPath_WRF_CUhw_N112_port);
   U14307 : INV_X1 port map( A => n14240, ZN => n8656);
   U14308 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB2_3_port, A2 => 
                           n14236, B1 => i_ADD_WB_3_port, B2 => n14237, ZN => 
                           n14240);
   U14309 : INV_X1 port map( A => n14264, ZN => n8720);
   U14310 : INV_X1 port map( A => n14262, ZN => n8722);
   U14311 : INV_X1 port map( A => n14259, ZN => n8723);
   U14312 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_26_port, A2 => n4259,
                           ZN => n2015);
   U14313 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_25_port, A2 => n4258,
                           ZN => n2016);
   U14314 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_24_port, A2 => n4261,
                           ZN => n2017);
   U14315 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_23_port, A2 => n4262,
                           ZN => n2018);
   U14316 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_22_port, A2 => n4257,
                           ZN => n2019);
   U14317 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_21_port, A2 => n4259,
                           ZN => n2020);
   U14318 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_20_port, A2 => n4258,
                           ZN => n2021);
   U14319 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_19_port, A2 => n4261,
                           ZN => n2022);
   U14320 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_18_port, A2 => n4262,
                           ZN => n2023);
   U14321 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_17_port, A2 => n4257,
                           ZN => n2024);
   U14322 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_16_port, A2 => n4264,
                           ZN => n2025);
   U14323 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_15_port, A2 => n4263,
                           ZN => n2026);
   U14324 : INV_X1 port map( A => n14239, ZN => n8657);
   U14325 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB2_2_port, A2 => 
                           n14236, B1 => i_ADD_WB_2_port, B2 => n14237, ZN => 
                           n14239);
   U14326 : INV_X1 port map( A => n14235, ZN => n8659);
   U14327 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB2_0_port, A2 => 
                           n14236, B1 => i_ADD_WB_0_port, B2 => n14237, ZN => 
                           n14235);
   U14328 : INV_X1 port map( A => n14238, ZN => n8658);
   U14329 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB2_1_port, A2 => 
                           n14236, B1 => i_ADD_WB_1_port, B2 => n14237, ZN => 
                           n14238);
   U14330 : INV_X1 port map( A => n14330, ZN => n8786);
   U14331 : AOI22_X1 port map( A1 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_1_port, A2 =>
                           n2500, B1 => DataPath_i_REG_MEM_ALUOUT_1_port, B2 =>
                           n2501, ZN => n14330);
   U14332 : INV_X1 port map( A => n14234, ZN => n8650);
   U14333 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_4_port, A2 => 
                           n14229, B1 => DataPath_i_PIPLIN_WRB2_4_port, B2 => 
                           n14230, ZN => n14234);
   U14334 : INV_X1 port map( A => n14233, ZN => n8651);
   U14335 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_3_port, A2 => 
                           n14229, B1 => DataPath_i_PIPLIN_WRB2_3_port, B2 => 
                           n14230, ZN => n14233);
   U14336 : INV_X1 port map( A => n14232, ZN => n8652);
   U14337 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_2_port, A2 => 
                           n14229, B1 => DataPath_i_PIPLIN_WRB2_2_port, B2 => 
                           n14230, ZN => n14232);
   U14338 : INV_X1 port map( A => n14231, ZN => n8653);
   U14339 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_1_port, A2 => 
                           n14229, B1 => DataPath_i_PIPLIN_WRB2_1_port, B2 => 
                           n14230, ZN => n14231);
   U14340 : INV_X1 port map( A => n14228, ZN => n8654);
   U14341 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_0_port, A2 => 
                           n14229, B1 => DataPath_i_PIPLIN_WRB2_0_port, B2 => 
                           n14230, ZN => n14228);
   U14342 : INV_X1 port map( A => n14241, ZN => n8655);
   U14343 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_WRB2_4_port, A2 => 
                           n14236, B1 => i_ADD_WB_4_port, B2 => n14237, ZN => 
                           n14241);
   U14344 : INV_X1 port map( A => n14327, ZN => n8787);
   U14345 : AOI22_X1 port map( A1 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_0_port, A2 =>
                           n2500, B1 => DataPath_i_REG_MEM_ALUOUT_0_port, B2 =>
                           n2501, ZN => n14327);
   U14346 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_1_port, A2 => n4263, 
                           ZN => n2027);
   U14347 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_0_port, A2 => n4264, 
                           ZN => n2028);
   U14348 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_3_port, A2 => n4266, ZN
                           => n2029);
   U14349 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_1_port, A2 => n4265, ZN
                           => n2030);
   U14350 : AND2_X1 port map( A1 => n1266, A2 => n4260, ZN => n2031);
   U14351 : INV_X1 port map( A => n14292, ZN => n8692);
   U14352 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_31_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_31_port, B2 => 
                           n2491, ZN => n14292);
   U14353 : INV_X1 port map( A => n14291, ZN => n8693);
   U14354 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_30_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_30_port, B2 => 
                           n2491, ZN => n14291);
   U14355 : INV_X1 port map( A => n14290, ZN => n8694);
   U14356 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_29_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_29_port, B2 => 
                           n2491, ZN => n14290);
   U14357 : INV_X1 port map( A => n14289, ZN => n8695);
   U14358 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_28_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_28_port, B2 => 
                           n2491, ZN => n14289);
   U14359 : INV_X1 port map( A => n14288, ZN => n8696);
   U14360 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_27_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_27_port, B2 => 
                           n2491, ZN => n14288);
   U14361 : INV_X1 port map( A => n14287, ZN => n8697);
   U14362 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_26_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_26_port, B2 => 
                           n2491, ZN => n14287);
   U14363 : INV_X1 port map( A => n14286, ZN => n8698);
   U14364 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_25_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_25_port, B2 => 
                           n2491, ZN => n14286);
   U14365 : INV_X1 port map( A => n14285, ZN => n8699);
   U14366 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_24_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_24_port, B2 => 
                           n2491, ZN => n14285);
   U14367 : INV_X1 port map( A => n14360, ZN => n8756);
   U14368 : AOI22_X1 port map( A1 => DRAM_ADDRESS_31_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_31_port, B2 => n2503, ZN 
                           => n14360);
   U14369 : INV_X1 port map( A => n14359, ZN => n8757);
   U14370 : AOI22_X1 port map( A1 => DRAM_ADDRESS_30_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_30_port, B2 => n2503, ZN 
                           => n14359);
   U14371 : INV_X1 port map( A => n14358, ZN => n8758);
   U14372 : AOI22_X1 port map( A1 => DRAM_ADDRESS_29_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_29_port, B2 => n2503, ZN 
                           => n14358);
   U14373 : INV_X1 port map( A => n14357, ZN => n8759);
   U14374 : AOI22_X1 port map( A1 => DRAM_ADDRESS_28_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_28_port, B2 => n2503, ZN 
                           => n14357);
   U14375 : INV_X1 port map( A => n14356, ZN => n8760);
   U14376 : AOI22_X1 port map( A1 => DRAM_ADDRESS_27_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_27_port, B2 => n2503, ZN 
                           => n14356);
   U14377 : INV_X1 port map( A => n14355, ZN => n8761);
   U14378 : AOI22_X1 port map( A1 => DRAM_ADDRESS_26_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_26_port, B2 => n2503, ZN 
                           => n14355);
   U14379 : INV_X1 port map( A => n14354, ZN => n8762);
   U14380 : AOI22_X1 port map( A1 => DRAM_ADDRESS_25_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_25_port, B2 => n2503, ZN 
                           => n14354);
   U14381 : INV_X1 port map( A => n14353, ZN => n8763);
   U14382 : AOI22_X1 port map( A1 => DRAM_ADDRESS_24_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_24_port, B2 => n2503, ZN 
                           => n14353);
   U14383 : INV_X1 port map( A => n14284, ZN => n8700);
   U14384 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_23_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_23_port, B2 => 
                           n2490, ZN => n14284);
   U14385 : INV_X1 port map( A => n14283, ZN => n8701);
   U14386 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_22_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_22_port, B2 => 
                           n2490, ZN => n14283);
   U14387 : INV_X1 port map( A => n14282, ZN => n8702);
   U14388 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_21_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_21_port, B2 => 
                           n2490, ZN => n14282);
   U14389 : INV_X1 port map( A => n14281, ZN => n8703);
   U14390 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_20_port, A2 => n2486, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_20_port, B2 => 
                           n2490, ZN => n14281);
   U14391 : INV_X1 port map( A => n14280, ZN => n8704);
   U14392 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_19_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_19_port, B2 => 
                           n2490, ZN => n14280);
   U14393 : INV_X1 port map( A => n14279, ZN => n8705);
   U14394 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_18_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_18_port, B2 => 
                           n2490, ZN => n14279);
   U14395 : INV_X1 port map( A => n14278, ZN => n8706);
   U14396 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_17_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_17_port, B2 => 
                           n2490, ZN => n14278);
   U14397 : INV_X1 port map( A => n14277, ZN => n8707);
   U14398 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_16_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_16_port, B2 => 
                           n2490, ZN => n14277);
   U14399 : INV_X1 port map( A => n14276, ZN => n8708);
   U14400 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_15_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_15_port, B2 => 
                           n2490, ZN => n14276);
   U14401 : INV_X1 port map( A => n14275, ZN => n8709);
   U14402 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_14_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_14_port, B2 => 
                           n2490, ZN => n14275);
   U14403 : INV_X1 port map( A => n14274, ZN => n8710);
   U14404 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_13_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_13_port, B2 => 
                           n2490, ZN => n14274);
   U14405 : INV_X1 port map( A => n14273, ZN => n8711);
   U14406 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_12_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_12_port, B2 => 
                           n2490, ZN => n14273);
   U14407 : INV_X1 port map( A => n14352, ZN => n8764);
   U14408 : AOI22_X1 port map( A1 => DRAM_ADDRESS_23_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_23_port, B2 => n2502, ZN 
                           => n14352);
   U14409 : INV_X1 port map( A => n14351, ZN => n8765);
   U14410 : AOI22_X1 port map( A1 => DRAM_ADDRESS_22_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_22_port, B2 => n2502, ZN 
                           => n14351);
   U14411 : INV_X1 port map( A => n14350, ZN => n8766);
   U14412 : AOI22_X1 port map( A1 => DRAM_ADDRESS_21_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_21_port, B2 => n2502, ZN 
                           => n14350);
   U14413 : INV_X1 port map( A => n14349, ZN => n8767);
   U14414 : AOI22_X1 port map( A1 => DRAM_ADDRESS_20_port, A2 => n2498, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_20_port, B2 => n2502, ZN 
                           => n14349);
   U14415 : INV_X1 port map( A => n14348, ZN => n8768);
   U14416 : AOI22_X1 port map( A1 => DRAM_ADDRESS_19_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_19_port, B2 => n2502, ZN 
                           => n14348);
   U14417 : INV_X1 port map( A => n14347, ZN => n8769);
   U14418 : AOI22_X1 port map( A1 => DRAM_ADDRESS_18_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_18_port, B2 => n2502, ZN 
                           => n14347);
   U14419 : INV_X1 port map( A => n14346, ZN => n8770);
   U14420 : AOI22_X1 port map( A1 => DRAM_ADDRESS_17_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_17_port, B2 => n2502, ZN 
                           => n14346);
   U14421 : INV_X1 port map( A => n14345, ZN => n8771);
   U14422 : AOI22_X1 port map( A1 => DRAM_ADDRESS_16_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_16_port, B2 => n2502, ZN 
                           => n14345);
   U14423 : INV_X1 port map( A => n14344, ZN => n8772);
   U14424 : AOI22_X1 port map( A1 => DRAM_ADDRESS_15_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_15_port, B2 => n2502, ZN 
                           => n14344);
   U14425 : INV_X1 port map( A => n14343, ZN => n8773);
   U14426 : AOI22_X1 port map( A1 => DRAM_ADDRESS_14_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_14_port, B2 => n2502, ZN 
                           => n14343);
   U14427 : INV_X1 port map( A => n14342, ZN => n8774);
   U14428 : AOI22_X1 port map( A1 => DRAM_ADDRESS_13_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_13_port, B2 => n2502, ZN 
                           => n14342);
   U14429 : INV_X1 port map( A => n14341, ZN => n8775);
   U14430 : AOI22_X1 port map( A1 => DRAM_ADDRESS_12_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_12_port, B2 => n2502, ZN 
                           => n14341);
   U14431 : INV_X1 port map( A => n14340, ZN => n8776);
   U14432 : AOI22_X1 port map( A1 => DRAM_ADDRESS_11_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_11_port, B2 => n2501, ZN 
                           => n14340);
   U14433 : INV_X1 port map( A => n14339, ZN => n8777);
   U14434 : AOI22_X1 port map( A1 => DRAM_ADDRESS_10_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_10_port, B2 => n2501, ZN 
                           => n14339);
   U14435 : INV_X1 port map( A => n14338, ZN => n8778);
   U14436 : AOI22_X1 port map( A1 => DRAM_ADDRESS_9_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_9_port, B2 => n2501, ZN =>
                           n14338);
   U14437 : INV_X1 port map( A => n14337, ZN => n8779);
   U14438 : AOI22_X1 port map( A1 => DRAM_ADDRESS_8_port, A2 => n2499, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_8_port, B2 => n2501, ZN =>
                           n14337);
   U14439 : INV_X1 port map( A => n14336, ZN => n8780);
   U14440 : AOI22_X1 port map( A1 => DRAM_ADDRESS_7_port, A2 => n2500, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_7_port, B2 => n2501, ZN =>
                           n14336);
   U14441 : INV_X1 port map( A => n14335, ZN => n8781);
   U14442 : AOI22_X1 port map( A1 => DRAM_ADDRESS_6_port, A2 => n2500, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_6_port, B2 => n2501, ZN =>
                           n14335);
   U14443 : INV_X1 port map( A => n14334, ZN => n8782);
   U14444 : AOI22_X1 port map( A1 => DRAM_ADDRESS_5_port, A2 => n2500, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_5_port, B2 => n2501, ZN =>
                           n14334);
   U14445 : INV_X1 port map( A => n14333, ZN => n8783);
   U14446 : AOI22_X1 port map( A1 => DRAM_ADDRESS_4_port, A2 => n2500, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_4_port, B2 => n2501, ZN =>
                           n14333);
   U14447 : INV_X1 port map( A => n14332, ZN => n8784);
   U14448 : AOI22_X1 port map( A1 => DRAM_ADDRESS_3_port, A2 => n2500, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_3_port, B2 => n2501, ZN =>
                           n14332);
   U14449 : INV_X1 port map( A => n14331, ZN => n8785);
   U14450 : AOI22_X1 port map( A1 => DRAM_ADDRESS_2_port, A2 => n2500, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_2_port, B2 => n2501, ZN =>
                           n14331);
   U14451 : INV_X1 port map( A => n14272, ZN => n8712);
   U14452 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_11_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_11_port, B2 => 
                           n2489, ZN => n14272);
   U14453 : INV_X1 port map( A => n14271, ZN => n8713);
   U14454 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_10_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_10_port, B2 => 
                           n2489, ZN => n14271);
   U14455 : INV_X1 port map( A => n14270, ZN => n8714);
   U14456 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_9_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_9_port, B2 => 
                           n2489, ZN => n14270);
   U14457 : INV_X1 port map( A => n14269, ZN => n8715);
   U14458 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_8_port, A2 => n2487, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_8_port, B2 => 
                           n2489, ZN => n14269);
   U14459 : INV_X1 port map( A => n14268, ZN => n8716);
   U14460 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_7_port, A2 => n2488, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_7_port, B2 => 
                           n2489, ZN => n14268);
   U14461 : INV_X1 port map( A => n14267, ZN => n8717);
   U14462 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_6_port, A2 => n2488, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_6_port, B2 => 
                           n2489, ZN => n14267);
   U14463 : INV_X1 port map( A => n14266, ZN => n8718);
   U14464 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_5_port, A2 => n2488, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_5_port, B2 => 
                           n2489, ZN => n14266);
   U14465 : INV_X1 port map( A => n14265, ZN => n8719);
   U14466 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_4_port, A2 => n2488, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_4_port, B2 => 
                           n2489, ZN => n14265);
   U14467 : INV_X1 port map( A => n14263, ZN => n8721);
   U14468 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_2_port, A2 => n2488, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_2_port, B2 => 
                           n2489, ZN => n14263);
   U14469 : AND2_X1 port map( A1 => DataPath_i_LGET_0_port, A2 => n4260, ZN => 
                           n2032);
   U14470 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_23_port, A2 => n4263, 
                           ZN => n2033);
   U14471 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_22_port, A2 => n4259, 
                           ZN => n2034);
   U14472 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_21_port, A2 => n4258, 
                           ZN => n2035);
   U14473 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_20_port, A2 => n4261, 
                           ZN => n2036);
   U14474 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_19_port, A2 => n4262, 
                           ZN => n2037);
   U14475 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_18_port, A2 => n4257, 
                           ZN => n2038);
   U14476 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_17_port, A2 => n4264, 
                           ZN => n2039);
   U14477 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_16_port, A2 => n4263, 
                           ZN => n2040);
   U14478 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_15_port, A2 => n4259, 
                           ZN => n2041);
   U14479 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_14_port, A2 => n4258, 
                           ZN => n2042);
   U14480 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_13_port, A2 => n4261, 
                           ZN => n2043);
   U14481 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_12_port, A2 => n4262, 
                           ZN => n2044);
   U14482 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_14_port, A2 => n4258,
                           ZN => n2045);
   U14483 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_13_port, A2 => n4261,
                           ZN => n2046);
   U14484 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_12_port, A2 => n4262,
                           ZN => n2047);
   U14485 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_11_port, A2 => n4257,
                           ZN => n2048);
   U14486 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_10_port, A2 => n4264,
                           ZN => n2049);
   U14487 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_9_port, A2 => n4263, 
                           ZN => n2050);
   U14488 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_8_port, A2 => n4259, 
                           ZN => n2051);
   U14489 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_7_port, A2 => n4258, 
                           ZN => n2052);
   U14490 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_6_port, A2 => n4261, 
                           ZN => n2053);
   U14491 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_5_port, A2 => n4262, 
                           ZN => n2054);
   U14492 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_4_port, A2 => n4257, 
                           ZN => n2055);
   U14493 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_30_port, A2 => n4264,
                           ZN => n2056);
   U14494 : INV_X1 port map( A => DataPath_RF_CWP_n13, ZN => n8649);
   U14495 : NAND2_X1 port map( A1 => DataPath_RF_next_cwp_4_port, A2 => n4258, 
                           ZN => DataPath_RF_CWP_n13);
   U14496 : NAND2_X1 port map( A1 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n2, A2 
                           => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n3, ZN => 
                           DataPath_RF_next_cwp_4_port);
   U14497 : AOI22_X1 port map( A1 => DataPath_RF_c_win_0_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4, B1 => 
                           DataPath_RF_c_win_3_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n3);
   U14498 : NAND2_X1 port map( A1 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n10, A2 
                           => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n11, ZN => 
                           DataPath_RF_next_cwp_2_port);
   U14499 : AOI22_X1 port map( A1 => DataPath_RF_c_win_3_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4, B1 => 
                           DataPath_RF_c_win_1_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n11);
   U14500 : NAND2_X1 port map( A1 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n12, A2 
                           => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n13, ZN => 
                           DataPath_RF_next_cwp_1_port);
   U14501 : AOI22_X1 port map( A1 => DataPath_RF_c_win_2_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4, B1 => 
                           DataPath_RF_c_win_0_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n13);
   U14502 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_30_port, A2 => n4264, 
                           ZN => n2057);
   U14503 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_29_port, A2 => n4263, 
                           ZN => n2058);
   U14504 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_28_port, A2 => n4259, 
                           ZN => n2059);
   U14505 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_27_port, A2 => n4258, 
                           ZN => n2060);
   U14506 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_26_port, A2 => n4261, 
                           ZN => n2061);
   U14507 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_25_port, A2 => n4262, 
                           ZN => n2062);
   U14508 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_24_port, A2 => n4257, 
                           ZN => n2063);
   U14509 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_23_port, A2 => n4264, 
                           ZN => n2064);
   U14510 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_22_port, A2 => n4263, 
                           ZN => n2065);
   U14511 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_21_port, A2 => n4259, 
                           ZN => n2066);
   U14512 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_20_port, A2 => n4258, 
                           ZN => n2067);
   U14513 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_19_port, A2 => n4261, 
                           ZN => n2068);
   U14514 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_18_port, A2 => n4259, 
                           ZN => n2069);
   U14515 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_17_port, A2 => n4258, 
                           ZN => n2070);
   U14516 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_16_port, A2 => n4261, 
                           ZN => n2071);
   U14517 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_15_port, A2 => n4262, 
                           ZN => n2072);
   U14518 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_14_port, A2 => n4257, 
                           ZN => n2073);
   U14519 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_13_port, A2 => n4264, 
                           ZN => n2074);
   U14520 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_12_port, A2 => n4263, 
                           ZN => n2075);
   U14521 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_11_port, A2 => n4259, 
                           ZN => n2076);
   U14522 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_10_port, A2 => n4258, 
                           ZN => n2077);
   U14523 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_9_port, A2 => n4261, ZN
                           => n2078);
   U14524 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_8_port, A2 => n4262, ZN
                           => n2079);
   U14525 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_7_port, A2 => n4257, ZN
                           => n2080);
   U14526 : NAND2_X1 port map( A1 => n12901, A2 => n12902, ZN => 
                           DataPath_RF_next_swp_4_port);
   U14527 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_0_port, A2 => n12903, 
                           B1 => DataPath_RF_c_swin_3_port, B2 => n12904, ZN =>
                           n12902);
   U14528 : NAND2_X1 port map( A1 => n12909, A2 => n12910, ZN => 
                           DataPath_RF_next_swp_2_port);
   U14529 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n12903, 
                           B1 => DataPath_RF_c_swin_1_port, B2 => n12904, ZN =>
                           n12910);
   U14530 : NAND2_X1 port map( A1 => n12911, A2 => n12912, ZN => 
                           DataPath_RF_next_swp_1_port);
   U14531 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_2_port, A2 => n12903, 
                           B1 => DataPath_RF_c_swin_0_port, B2 => n12904, ZN =>
                           n12912);
   U14532 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_31_port, A2 => n4260, 
                           ZN => n2081);
   U14533 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_30_port, A2 => n4259, 
                           ZN => n2082);
   U14534 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_29_port, A2 => n4263, 
                           ZN => n2083);
   U14535 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_28_port, A2 => n4266, 
                           ZN => n2084);
   U14536 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_27_port, A2 => n4265, 
                           ZN => n2085);
   U14537 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_26_port, A2 => n4262, 
                           ZN => n2086);
   U14538 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_25_port, A2 => n4265, 
                           ZN => n2087);
   U14539 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_24_port, A2 => n4264, 
                           ZN => n2088);
   U14540 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_3_port, A2 => n4261, 
                           ZN => n2089);
   U14541 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_2_port, A2 => n4262, 
                           ZN => n2090);
   U14542 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_1_port, A2 => n4257, 
                           ZN => n2091);
   U14543 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_0_port, A2 => n4259, 
                           ZN => n2092);
   U14544 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_4_port, A2 => n4264,
                           ZN => n2093);
   U14545 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_3_port, A2 => n4266,
                           ZN => n2094);
   U14546 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_2_port, A2 => n4265,
                           ZN => n2095);
   U14547 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_1_port, A2 => n4265,
                           ZN => n2096);
   U14548 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_WRB1_0_port, A2 => n4260,
                           ZN => n2097);
   U14549 : AND2_X1 port map( A1 => DataPath_i_LGET_1_port, A2 => n4260, ZN => 
                           n2098);
   U14550 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_31_port, A2 => n4260, 
                           ZN => n2099);
   U14551 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_6_port, A2 => n4259, ZN
                           => n2100);
   U14552 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_5_port, A2 => n4265, ZN
                           => n2101);
   U14553 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_4_port, A2 => n4260, ZN
                           => n2102);
   U14554 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_3_port, A2 => n4263, ZN
                           => n2103);
   U14555 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_2_port, A2 => n4260, ZN
                           => n2104);
   U14556 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_1_port, A2 => n4261, ZN
                           => n2105);
   U14557 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_A_0_port, A2 => n4266, ZN
                           => n2106);
   U14558 : NAND2_X1 port map( A1 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n8, A2 
                           => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n9, ZN => 
                           DataPath_RF_next_cwp_3_port);
   U14559 : AOI22_X1 port map( A1 => n3269, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4, B1 => 
                           DataPath_RF_c_win_2_port, B2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n9);
   U14560 : NAND2_X1 port map( A1 => n12907, A2 => n12908, ZN => 
                           DataPath_RF_next_swp_3_port);
   U14561 : AOI22_X1 port map( A1 => n3889, A2 => n12903, B1 => 
                           DataPath_RF_c_swin_2_port, B2 => n12904, ZN => 
                           n12908);
   U14562 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_31_port, A2 => n4265,
                           ZN => n2107);
   U14563 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_31_port, A2 => n4260,
                           ZN => n2108);
   U14564 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_30_port, A2 => n4257,
                           ZN => n2109);
   U14565 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_29_port, A2 => n4264,
                           ZN => n2110);
   U14566 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_28_port, A2 => n4258,
                           ZN => n2111);
   U14567 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN1_27_port, A2 => n4258,
                           ZN => n2112);
   U14568 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_6_port, A2 => n4261, 
                           ZN => n2113);
   U14569 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_5_port, A2 => n4260, 
                           ZN => n2114);
   U14570 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_4_port, A2 => n4262, 
                           ZN => n2115);
   U14571 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_3_port, A2 => n4263, 
                           ZN => n2116);
   U14572 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_IN2_2_port, A2 => n4257, 
                           ZN => n2117);
   U14573 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_11_port, A2 => n4262, 
                           ZN => n2118);
   U14574 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_10_port, A2 => n4260, 
                           ZN => n2119);
   U14575 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_9_port, A2 => n4260, ZN
                           => n2120);
   U14576 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_8_port, A2 => n4265, ZN
                           => n2121);
   U14577 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_7_port, A2 => n4258, ZN
                           => n2122);
   U14578 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_6_port, A2 => n4266, ZN
                           => n2123);
   U14579 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_5_port, A2 => n4257, ZN
                           => n2124);
   U14580 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_4_port, A2 => n4260, ZN
                           => n2125);
   U14581 : AND2_X1 port map( A1 => DataPath_i_PIPLIN_B_2_port, A2 => n4259, ZN
                           => n2126);
   U14582 : NAND2_X1 port map( A1 => n12913, A2 => n12914, ZN => 
                           DataPath_RF_next_swp_0_port);
   U14583 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_1_port, A2 => n12903, 
                           B1 => n3890, B2 => n12904, ZN => n12914);
   U14584 : NAND2_X1 port map( A1 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n14, A2 
                           => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n15, ZN => 
                           DataPath_RF_next_cwp_0_port);
   U14585 : AOI22_X1 port map( A1 => DataPath_RF_c_win_1_port, A2 => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n4, B1 => n3270, 
                           B2 => DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n5, ZN => 
                           DataPath_RF_CWP_NEXT_CALC_MUX_SEL_n15);
   U14586 : OAI22_X1 port map( A1 => n3904, A2 => DataPath_RF_PUSH_ADDRGEN_n13,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n40, B2 => 
                           DataPath_RF_n10, ZN => 
                           DataPath_RF_spill_address_ext_5_port);
   U14587 : OAI22_X1 port map( A1 => n3904, A2 => DataPath_RF_PUSH_ADDRGEN_n14,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n41, B2 => 
                           DataPath_RF_n10, ZN => 
                           DataPath_RF_spill_address_ext_4_port);
   U14588 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_96_port, A2 
                           => n3090, B1 => DataPath_RF_bus_reg_dataout_608_port
                           , B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1632_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n17);
   U14589 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_97_port, A2 
                           => n3090, B1 => DataPath_RF_bus_reg_dataout_609_port
                           , B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1633_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n15);
   U14590 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_98_port, A2 
                           => n3090, B1 => DataPath_RF_bus_reg_dataout_610_port
                           , B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1634_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n13);
   U14591 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_99_port, A2 
                           => n3090, B1 => DataPath_RF_bus_reg_dataout_611_port
                           , B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1635_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n11);
   U14592 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_9_port, A2 =>
                           n3090, B1 => DataPath_RF_bus_reg_dataout_521_port, 
                           B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1545_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n5);
   U14593 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_93_port, A2 
                           => n3090, B1 => DataPath_RF_bus_reg_dataout_605_port
                           , B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1629_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n23);
   U14594 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_94_port, A2 
                           => n3090, B1 => DataPath_RF_bus_reg_dataout_606_port
                           , B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1630_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n21);
   U14595 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_95_port, A2 
                           => n3090, B1 => DataPath_RF_bus_reg_dataout_607_port
                           , B2 => n3145, C1 => 
                           DataPath_RF_bus_reg_dataout_1631_port, C2 => n3191, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n19);
   U14596 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_192_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_704_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1728_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n827);
   U14597 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_32_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_544_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1568_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n521);
   U14598 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_160_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_672_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1696_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n897);
   U14599 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_64_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_576_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1600_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n87);
   U14600 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_0_port, A2 =>
                           n3048, B1 => DataPath_RF_bus_reg_dataout_512_port, 
                           B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1536_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1031);
   U14601 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_128_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_640_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1664_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n969);
   U14602 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_224_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_736_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1760_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n755);
   U14603 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_416_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_928_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1952_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n329);
   U14604 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_320_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_832_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1856_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n541);
   U14605 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_256_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_768_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1792_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n685);
   U14606 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_384_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_896_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1920_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n401);
   U14607 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_288_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_800_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1824_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n615);
   U14608 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_352_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_864_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1888_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n471);
   U14609 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_193_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_705_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1729_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n825);
   U14610 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_33_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_545_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1569_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n499);
   U14611 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_161_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_673_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1697_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n895);
   U14612 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_65_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_577_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1601_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n85);
   U14613 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1_port, A2 =>
                           n3057, B1 => DataPath_RF_bus_reg_dataout_513_port, 
                           B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1537_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n809);
   U14614 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_129_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_641_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1665_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n967);
   U14615 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_225_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_737_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1761_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n753);
   U14616 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_417_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_929_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1953_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n327);
   U14617 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_321_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_833_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1857_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n539);
   U14618 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_257_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_769_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1793_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n683);
   U14619 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_385_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_897_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1921_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n399);
   U14620 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_289_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_801_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1825_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n613);
   U14621 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_353_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_865_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1889_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n469);
   U14622 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_194_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_706_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1730_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n823);
   U14623 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_34_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_546_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1570_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n477);
   U14624 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_162_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_674_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1698_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n893);
   U14625 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_66_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_578_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1602_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n83);
   U14626 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2_port, A2 =>
                           n3066, B1 => DataPath_RF_bus_reg_dataout_514_port, 
                           B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1538_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n587);
   U14627 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_130_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_642_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1666_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n963);
   U14628 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_226_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_738_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1762_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n751);
   U14629 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_418_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_930_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1954_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n325);
   U14630 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_322_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_834_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1858_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n537);
   U14631 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_258_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_770_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1794_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n681);
   U14632 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_386_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_898_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1922_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n397);
   U14633 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_290_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_802_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1826_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n609);
   U14634 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_354_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_866_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1890_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n467);
   U14635 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_195_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_707_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1731_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n821);
   U14636 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_35_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_547_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1571_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n455);
   U14637 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_163_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_675_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1699_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n891);
   U14638 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_67_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_579_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1603_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n81);
   U14639 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_3_port, A2 =>
                           n3075, B1 => DataPath_RF_bus_reg_dataout_515_port, 
                           B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1539_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n365);
   U14640 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_131_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_643_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1667_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n961);
   U14641 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_227_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_739_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1763_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n749);
   U14642 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_419_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_931_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1955_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n323);
   U14643 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_323_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_835_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1859_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n535);
   U14644 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_259_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_771_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1795_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n679);
   U14645 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_387_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_899_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1923_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n395);
   U14646 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_291_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_803_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1827_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n607);
   U14647 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_355_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_867_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1891_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n465);
   U14648 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_196_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_708_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1732_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n819);
   U14649 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_100_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_612_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1636_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1029);
   U14650 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_36_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_548_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1572_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n433);
   U14651 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_164_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_676_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1700_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n889);
   U14652 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_68_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_580_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1604_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n79);
   U14653 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_4_port, A2 =>
                           n3085, B1 => DataPath_RF_bus_reg_dataout_516_port, 
                           B2 => n3140, C1 => 
                           DataPath_RF_bus_reg_dataout_1540_port, C2 => n3186, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n143);
   U14654 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_132_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_644_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1668_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n959);
   U14655 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_228_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_740_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1764_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n747);
   U14656 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_420_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_932_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1956_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n319);
   U14657 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_324_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_836_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1860_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n533);
   U14658 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_260_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_772_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1796_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n675);
   U14659 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_388_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_900_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1924_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n393);
   U14660 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_292_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_804_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1828_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n605);
   U14661 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_356_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_868_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1892_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n463);
   U14662 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_197_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_709_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1733_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n817);
   U14663 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_101_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_613_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1637_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1027);
   U14664 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_37_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_549_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1573_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n411);
   U14665 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_165_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_677_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1701_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n887);
   U14666 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_69_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_581_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1605_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n77);
   U14667 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_5_port, A2 =>
                           n3086, B1 => DataPath_RF_bus_reg_dataout_517_port, 
                           B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1541_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n97);
   U14668 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_133_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_645_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1669_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n957);
   U14669 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_229_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_741_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1765_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n745);
   U14670 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_421_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_933_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1957_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n317);
   U14671 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_325_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_837_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1861_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n531);
   U14672 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_261_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_773_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1797_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n673);
   U14673 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_389_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_901_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1925_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n391);
   U14674 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_293_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_805_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1829_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n603);
   U14675 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_357_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_869_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1893_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n461);
   U14676 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_198_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_710_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1734_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n815);
   U14677 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_102_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_614_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1638_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1025);
   U14678 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_38_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_550_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1574_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n389);
   U14679 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_166_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_678_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1702_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n885);
   U14680 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_70_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_582_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1606_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n73);
   U14681 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_6_port, A2 =>
                           n3087, B1 => DataPath_RF_bus_reg_dataout_518_port, 
                           B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1542_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n75);
   U14682 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_134_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_646_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1670_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n955);
   U14683 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_230_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_742_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1766_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n741);
   U14684 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_422_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_934_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1958_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n315);
   U14685 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_326_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_838_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1862_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n529);
   U14686 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_262_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_774_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1798_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n671);
   U14687 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_390_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_902_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1926_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n387);
   U14688 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_294_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_806_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1830_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n601);
   U14689 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_358_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_870_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1894_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n459);
   U14690 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_199_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_711_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1735_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n813);
   U14691 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_103_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_615_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1639_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1023);
   U14692 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_39_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_551_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1575_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n367);
   U14693 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_167_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_679_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1703_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n883);
   U14694 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_71_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_583_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1607_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n71);
   U14695 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_7_port, A2 =>
                           n3088, B1 => DataPath_RF_bus_reg_dataout_519_port, 
                           B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1543_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n53);
   U14696 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_135_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_647_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1671_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n953);
   U14697 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_231_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_743_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1767_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n739);
   U14698 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_423_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_935_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1959_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n313);
   U14699 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_327_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_839_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1863_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n527);
   U14700 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_263_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_775_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1799_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n669);
   U14701 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_391_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_903_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1927_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n385);
   U14702 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_295_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_807_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1831_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n599);
   U14703 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_359_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_871_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1895_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n457);
   U14704 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_200_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_712_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1736_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n807);
   U14705 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_104_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_616_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1640_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1021);
   U14706 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_40_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_552_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1576_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n343);
   U14707 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_168_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_680_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1704_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n881);
   U14708 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_72_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_584_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1608_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n69);
   U14709 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_8_port, A2 =>
                           n3089, B1 => DataPath_RF_bus_reg_dataout_520_port, 
                           B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1544_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n31);
   U14710 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_136_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_648_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1672_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n951);
   U14711 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_232_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_744_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1768_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n737);
   U14712 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_424_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_936_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1960_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n311);
   U14713 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_328_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_840_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1864_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n525);
   U14714 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_264_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_776_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1800_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n667);
   U14715 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_392_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_904_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1928_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n383);
   U14716 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_296_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_808_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1832_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n597);
   U14717 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_360_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_872_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1896_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n453);
   U14718 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_201_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_713_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1737_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n805);
   U14719 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_105_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_617_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1641_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1019);
   U14720 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_41_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_553_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1577_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n321);
   U14721 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_169_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_681_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1705_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n879);
   U14722 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_73_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_585_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1609_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n67);
   U14723 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_137_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_649_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1673_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n949);
   U14724 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_233_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_745_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1769_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n735);
   U14725 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_425_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_937_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1961_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n309);
   U14726 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_329_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_841_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1865_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n523);
   U14727 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_265_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_777_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1801_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n665);
   U14728 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_393_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_905_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1929_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n381);
   U14729 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_297_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_809_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1833_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n595);
   U14730 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_361_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_873_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1897_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n451);
   U14731 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_202_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_714_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1738_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n803);
   U14732 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_106_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_618_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1642_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1017);
   U14733 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_42_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_554_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1578_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n299);
   U14734 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_170_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_682_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1706_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n875);
   U14735 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_74_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_586_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1610_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n65);
   U14736 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_10_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_522_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1546_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1009);
   U14737 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_138_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_650_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1674_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n947);
   U14738 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_234_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_746_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1770_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n733);
   U14739 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_426_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_938_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1962_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n307);
   U14740 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_330_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_842_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1866_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n519);
   U14741 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_266_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_778_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1802_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n663);
   U14742 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_394_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_906_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1930_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n379);
   U14743 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_298_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_810_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1834_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n593);
   U14744 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_362_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_874_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1898_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n449);
   U14745 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_203_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_715_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1739_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n801);
   U14746 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_107_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_619_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1643_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1015);
   U14747 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_43_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_555_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1579_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n277);
   U14748 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_171_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_683_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1707_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n873);
   U14749 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_75_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_587_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1611_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n63);
   U14750 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_11_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_523_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1547_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n987);
   U14751 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_139_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_651_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1675_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n945);
   U14752 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_235_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_747_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1771_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n731);
   U14753 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_427_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_939_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1963_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n305);
   U14754 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_331_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_843_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1867_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n517);
   U14755 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_267_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_779_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1803_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n661);
   U14756 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_395_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_907_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1931_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n377);
   U14757 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_299_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_811_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1835_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n591);
   U14758 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_363_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_875_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1899_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n447);
   U14759 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_204_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_716_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1740_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n799);
   U14760 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_108_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_620_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1644_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1013);
   U14761 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_44_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_556_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1580_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n255);
   U14762 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_172_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_684_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1708_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n871);
   U14763 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_76_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_588_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1612_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n61);
   U14764 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_12_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_524_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1548_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n965);
   U14765 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_140_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_652_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1676_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n941);
   U14766 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_236_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_748_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1772_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n729);
   U14767 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_428_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_940_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1964_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n303);
   U14768 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_332_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_844_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1868_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n515);
   U14769 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_268_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_780_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1804_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n659);
   U14770 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_396_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_908_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1932_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n375);
   U14771 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_300_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_812_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1836_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n585);
   U14772 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_364_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_876_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1900_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n445);
   U14773 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_205_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_717_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1741_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n797);
   U14774 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_109_port, A2 
                           => n3048, B1 => DataPath_RF_bus_reg_dataout_621_port
                           , B2 => n3103, C1 => 
                           DataPath_RF_bus_reg_dataout_1645_port, C2 => n3149, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1011);
   U14775 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_45_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_557_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1581_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n233);
   U14776 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_173_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_685_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1709_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n869);
   U14777 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_77_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_589_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1613_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n59);
   U14778 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_13_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_525_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1549_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n943);
   U14779 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_141_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_653_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1677_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n939);
   U14780 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_237_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_749_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1773_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n727);
   U14781 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_429_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_941_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1965_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n301);
   U14782 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_333_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_845_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1869_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n513);
   U14783 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_269_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_781_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1805_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n657);
   U14784 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_397_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_909_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1933_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n373);
   U14785 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_301_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_813_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1837_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n583);
   U14786 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_365_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_877_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1901_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n443);
   U14787 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_206_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_718_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1742_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n795);
   U14788 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_110_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_622_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1646_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1007);
   U14789 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_46_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_558_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_1582_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n211);
   U14790 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_174_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_686_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1710_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n867);
   U14791 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_78_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_590_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1614_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n57);
   U14792 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_14_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_526_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1550_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n921);
   U14793 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_142_port, A2 
                           => n3051, B1 => DataPath_RF_bus_reg_dataout_654_port
                           , B2 => n3106, C1 => 
                           DataPath_RF_bus_reg_dataout_1678_port, C2 => n3152, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n937);
   U14794 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_238_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_750_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1774_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n725);
   U14795 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_430_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_942_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1966_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n297);
   U14796 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_334_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_846_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1870_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n511);
   U14797 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_270_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_782_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1806_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n653);
   U14798 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_398_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_910_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1934_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n371);
   U14799 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_302_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_814_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1838_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n581);
   U14800 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_366_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_878_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1902_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n441);
   U14801 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_207_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_719_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1743_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n793);
   U14802 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_111_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_623_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1647_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1005);
   U14803 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_47_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_559_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_1583_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n189);
   U14804 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_175_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_687_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1711_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n865);
   U14805 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_79_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_591_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1615_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n55);
   U14806 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_15_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_527_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1551_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n899);
   U14807 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_143_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_655_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1679_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n935);
   U14808 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_239_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_751_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1775_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n723);
   U14809 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_431_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_943_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1967_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n295);
   U14810 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_335_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_847_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1871_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n509);
   U14811 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_271_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_783_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1807_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n651);
   U14812 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_399_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_911_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1935_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n369);
   U14813 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_303_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_815_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1839_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n579);
   U14814 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_367_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_879_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1903_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n439);
   U14815 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_208_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_720_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1744_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n791);
   U14816 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_112_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_624_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1648_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1003);
   U14817 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_48_port, A2 
                           => n3084, B1 => DataPath_RF_bus_reg_dataout_560_port
                           , B2 => n3139, C1 => 
                           DataPath_RF_bus_reg_dataout_1584_port, C2 => n3185, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n167);
   U14818 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_176_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_688_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1712_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n863);
   U14819 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_80_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_592_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1616_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n51);
   U14820 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_16_port, A2 
                           => n3054, B1 => DataPath_RF_bus_reg_dataout_528_port
                           , B2 => n3109, C1 => 
                           DataPath_RF_bus_reg_dataout_1552_port, C2 => n3155, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n877);
   U14821 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_144_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_656_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1680_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n933);
   U14822 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_240_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_752_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1776_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n719);
   U14823 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_432_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_944_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1968_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n293);
   U14824 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_336_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_848_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1872_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n507);
   U14825 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_272_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_784_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1808_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n649);
   U14826 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_400_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_912_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1936_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n363);
   U14827 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_304_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_816_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1840_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n577);
   U14828 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_368_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_880_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1904_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n437);
   U14829 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_209_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_721_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1745_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n789);
   U14830 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_113_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_625_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1649_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1001);
   U14831 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_49_port, A2 
                           => n3084, B1 => DataPath_RF_bus_reg_dataout_561_port
                           , B2 => n3139, C1 => 
                           DataPath_RF_bus_reg_dataout_1585_port, C2 => n3185, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n145);
   U14832 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_177_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_689_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1713_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n861);
   U14833 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_81_port, A2 
                           => n3088, B1 => DataPath_RF_bus_reg_dataout_593_port
                           , B2 => n3143, C1 => 
                           DataPath_RF_bus_reg_dataout_1617_port, C2 => n3189, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n49);
   U14834 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_17_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_529_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1553_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n855);
   U14835 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_145_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_657_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1681_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n931);
   U14836 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_241_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_753_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1777_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n717);
   U14837 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_433_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_945_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1969_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n291);
   U14838 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_337_port, A2 
                           => n3069, B1 => DataPath_RF_bus_reg_dataout_849_port
                           , B2 => n3124, C1 => 
                           DataPath_RF_bus_reg_dataout_1873_port, C2 => n3170, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n505);
   U14839 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_273_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_785_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1809_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n647);
   U14840 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_401_port, A2 
                           => n3075, B1 => DataPath_RF_bus_reg_dataout_913_port
                           , B2 => n3130, C1 => 
                           DataPath_RF_bus_reg_dataout_1937_port, C2 => n3176, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n361);
   U14841 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_305_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_817_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1841_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n575);
   U14842 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_369_port, A2 
                           => n3072, B1 => DataPath_RF_bus_reg_dataout_881_port
                           , B2 => n3127, C1 => 
                           DataPath_RF_bus_reg_dataout_1905_port, C2 => n3173, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n435);
   U14843 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_210_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_722_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1746_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n785);
   U14844 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_114_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_626_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1650_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n999);
   U14845 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_50_port, A2 
                           => n3085, B1 => DataPath_RF_bus_reg_dataout_562_port
                           , B2 => n3140, C1 => 
                           DataPath_RF_bus_reg_dataout_1586_port, C2 => n3186, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n121);
   U14846 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_178_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_690_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1714_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n859);
   U14847 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_82_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_594_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1618_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n47);
   U14848 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_18_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_530_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1554_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n833);
   U14849 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_146_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_658_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1682_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n929);
   U14850 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_242_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_754_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1778_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n715);
   U14851 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_434_port, A2 
                           => n3078, B1 => DataPath_RF_bus_reg_dataout_946_port
                           , B2 => n3133, C1 => 
                           DataPath_RF_bus_reg_dataout_1970_port, C2 => n3179, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n289);
   U14852 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_338_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_850_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1874_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n503);
   U14853 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_274_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_786_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1810_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n645);
   U14854 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_402_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_914_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1938_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n359);
   U14855 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_306_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_818_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1842_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n573);
   U14856 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_370_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_882_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1906_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n431);
   U14857 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_211_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_723_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1747_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n783);
   U14858 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_115_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_627_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1651_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n997);
   U14859 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_51_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_563_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1587_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n115);
   U14860 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_179_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_691_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1715_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n857);
   U14861 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_83_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_595_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1619_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n45);
   U14862 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_19_port, A2 
                           => n3057, B1 => DataPath_RF_bus_reg_dataout_531_port
                           , B2 => n3112, C1 => 
                           DataPath_RF_bus_reg_dataout_1555_port, C2 => n3158, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n811);
   U14863 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_147_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_659_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1683_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n927);
   U14864 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_243_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_755_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1779_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n713);
   U14865 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_435_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_947_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1971_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n287);
   U14866 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_339_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_851_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1875_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n501);
   U14867 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_275_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_787_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1811_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n643);
   U14868 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_403_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_915_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1939_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n357);
   U14869 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_307_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_819_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1843_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n571);
   U14870 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_371_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_883_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1907_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n429);
   U14871 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_212_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_724_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1748_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n781);
   U14872 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_116_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_628_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1652_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n995);
   U14873 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_52_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_564_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1588_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n113);
   U14874 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_180_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_692_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1716_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n853);
   U14875 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_84_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_596_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1620_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n43);
   U14876 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_20_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_532_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1556_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n787);
   U14877 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_148_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_660_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1684_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n925);
   U14878 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_244_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_756_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1780_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n711);
   U14879 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_436_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_948_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1972_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n285);
   U14880 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_340_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_852_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1876_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n497);
   U14881 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_276_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_788_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1812_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n641);
   U14882 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_404_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_916_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1940_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n355);
   U14883 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_308_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_820_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1844_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n569);
   U14884 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_372_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_884_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1908_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n427);
   U14885 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_213_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_725_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1749_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n779);
   U14886 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_117_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_629_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1653_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n993);
   U14887 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_53_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_565_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1589_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n111);
   U14888 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_181_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_693_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1717_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n851);
   U14889 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_85_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_597_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1621_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n41);
   U14890 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_21_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_533_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1557_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n765);
   U14891 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_149_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_661_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1685_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n923);
   U14892 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_245_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_757_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1781_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n709);
   U14893 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_437_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_949_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1973_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n283);
   U14894 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_341_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_853_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1877_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n495);
   U14895 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_277_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_789_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1813_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n639);
   U14896 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_405_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_917_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1941_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n353);
   U14897 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_309_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_821_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1845_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n567);
   U14898 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_373_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_885_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1909_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n425);
   U14899 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_214_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_726_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1750_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n777);
   U14900 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_118_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_630_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1654_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n991);
   U14901 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_54_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_566_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1590_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n109);
   U14902 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_182_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_694_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1718_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n849);
   U14903 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_86_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_598_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1622_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n39);
   U14904 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_22_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_534_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1558_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n743);
   U14905 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_150_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_662_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1686_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n919);
   U14906 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_246_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_758_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1782_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n707);
   U14907 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_438_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_950_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1974_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n281);
   U14908 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_342_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_854_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1878_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n493);
   U14909 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_278_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_790_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1814_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n637);
   U14910 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_406_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_918_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1942_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n351);
   U14911 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_310_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_822_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1846_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n563);
   U14912 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_374_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_886_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1910_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n423);
   U14913 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_215_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_727_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1751_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n775);
   U14914 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_119_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_631_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1655_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n989);
   U14915 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_55_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_567_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1591_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n107);
   U14916 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_183_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_695_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1719_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n847);
   U14917 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_87_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_599_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1623_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n37);
   U14918 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_23_port, A2 
                           => n3060, B1 => DataPath_RF_bus_reg_dataout_535_port
                           , B2 => n3115, C1 => 
                           DataPath_RF_bus_reg_dataout_1559_port, C2 => n3161, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n721);
   U14919 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_151_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_663_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1687_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n917);
   U14920 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_247_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_759_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1783_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n705);
   U14921 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_439_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_951_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1975_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n279);
   U14922 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_343_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_855_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1879_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n491);
   U14923 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_279_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_791_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1815_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n635);
   U14924 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_407_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_919_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1943_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n349);
   U14925 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_311_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_823_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1847_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n561);
   U14926 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_375_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_887_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1911_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n421);
   U14927 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_216_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_728_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1752_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n773);
   U14928 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_120_port, A2 
                           => n3049, B1 => DataPath_RF_bus_reg_dataout_632_port
                           , B2 => n3104, C1 => 
                           DataPath_RF_bus_reg_dataout_1656_port, C2 => n3150, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n985);
   U14929 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_56_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_568_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1592_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n105);
   U14930 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_184_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_696_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1720_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n845);
   U14931 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_88_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_600_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1624_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n35);
   U14932 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_24_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_536_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1560_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n699);
   U14933 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_152_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_664_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1688_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n915);
   U14934 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_248_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_760_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1784_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n703);
   U14935 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_440_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_952_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1976_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n275);
   U14936 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_344_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_856_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1880_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n489);
   U14937 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_280_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_792_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1816_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n631);
   U14938 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_408_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_920_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1944_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n347);
   U14939 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_312_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_824_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1848_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n559);
   U14940 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_376_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_888_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1912_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n419);
   U14941 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_217_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_729_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1753_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n771);
   U14942 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_121_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_633_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1657_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n983);
   U14943 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_57_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_569_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1593_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n103);
   U14944 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_185_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_697_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1721_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n843);
   U14945 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_89_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_601_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1625_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n33);
   U14946 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_25_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_537_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1561_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n677);
   U14947 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_153_port, A2 
                           => n3052, B1 => DataPath_RF_bus_reg_dataout_665_port
                           , B2 => n3107, C1 => 
                           DataPath_RF_bus_reg_dataout_1689_port, C2 => n3153, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n913);
   U14948 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_249_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_761_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1785_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n701);
   U14949 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_441_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_953_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1977_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n273);
   U14950 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_345_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_857_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1881_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n487);
   U14951 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_281_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_793_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1817_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n629);
   U14952 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_409_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_921_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1945_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n345);
   U14953 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_313_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_825_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1849_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n557);
   U14954 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_377_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_889_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1913_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n417);
   U14955 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_218_port, A2 
                           => n3058, B1 => DataPath_RF_bus_reg_dataout_730_port
                           , B2 => n3113, C1 => 
                           DataPath_RF_bus_reg_dataout_1754_port, C2 => n3159, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n769);
   U14956 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_122_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_634_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1658_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n981);
   U14957 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_58_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_570_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1594_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n101);
   U14958 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_186_port, A2 
                           => n3055, B1 => DataPath_RF_bus_reg_dataout_698_port
                           , B2 => n3110, C1 => 
                           DataPath_RF_bus_reg_dataout_1722_port, C2 => n3156, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n841);
   U14959 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_90_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_602_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1626_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n29);
   U14960 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_26_port, A2 
                           => n3063, B1 => DataPath_RF_bus_reg_dataout_538_port
                           , B2 => n3118, C1 => 
                           DataPath_RF_bus_reg_dataout_1562_port, C2 => n3164, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n655);
   U14961 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_154_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_666_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1690_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n911);
   U14962 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_250_port, A2 
                           => n3061, B1 => DataPath_RF_bus_reg_dataout_762_port
                           , B2 => n3116, C1 => 
                           DataPath_RF_bus_reg_dataout_1786_port, C2 => n3162, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n697);
   U14963 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_442_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_954_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1978_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n271);
   U14964 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_346_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_858_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1882_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n485);
   U14965 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_282_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_794_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1818_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n627);
   U14966 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_410_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_922_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1946_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n341);
   U14967 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_314_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_826_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1850_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n555);
   U14968 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_378_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_890_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1914_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n415);
   U14969 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_219_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_731_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1755_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n767);
   U14970 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_123_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_635_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1659_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n979);
   U14971 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_59_port, A2 
                           => n3086, B1 => DataPath_RF_bus_reg_dataout_571_port
                           , B2 => n3141, C1 => 
                           DataPath_RF_bus_reg_dataout_1595_port, C2 => n3187, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n99);
   U14972 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_187_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_699_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1723_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n839);
   U14973 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_91_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_603_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1627_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n27);
   U14974 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_27_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_539_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1563_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n633);
   U14975 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_155_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_667_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1691_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n909);
   U14976 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_251_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_763_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1787_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n695);
   U14977 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_443_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_955_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1979_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n269);
   U14978 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_347_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_859_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1883_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n483);
   U14979 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_283_port, A2 
                           => n3064, B1 => DataPath_RF_bus_reg_dataout_795_port
                           , B2 => n3119, C1 => 
                           DataPath_RF_bus_reg_dataout_1819_port, C2 => n3165, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n625);
   U14980 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_411_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_923_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1947_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n339);
   U14981 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_315_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_827_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1851_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n553);
   U14982 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_379_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_891_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1915_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n413);
   U14983 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_220_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_732_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1756_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n763);
   U14984 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_124_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_636_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1660_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n977);
   U14985 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_60_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_572_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1596_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n95);
   U14986 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_188_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_700_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1724_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n837);
   U14987 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_92_port, A2 
                           => n3089, B1 => DataPath_RF_bus_reg_dataout_604_port
                           , B2 => n3144, C1 => 
                           DataPath_RF_bus_reg_dataout_1628_port, C2 => n3190, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n25);
   U14988 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_28_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_540_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1564_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n611);
   U14989 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_156_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_668_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1692_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n907);
   U14990 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_252_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_764_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1788_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n693);
   U14991 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_444_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_956_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1980_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n267);
   U14992 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_348_port, A2 
                           => n3070, B1 => DataPath_RF_bus_reg_dataout_860_port
                           , B2 => n3125, C1 => 
                           DataPath_RF_bus_reg_dataout_1884_port, C2 => n3171, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n481);
   U14993 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_284_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_796_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1820_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n623);
   U14994 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_412_port, A2 
                           => n3076, B1 => DataPath_RF_bus_reg_dataout_924_port
                           , B2 => n3131, C1 => 
                           DataPath_RF_bus_reg_dataout_1948_port, C2 => n3177, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n337);
   U14995 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_316_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_828_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1852_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n551);
   U14996 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_380_port, A2 
                           => n3073, B1 => DataPath_RF_bus_reg_dataout_892_port
                           , B2 => n3128, C1 => 
                           DataPath_RF_bus_reg_dataout_1916_port, C2 => n3174, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n409);
   U14997 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_221_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_733_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1757_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n761);
   U14998 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_125_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_637_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1661_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n975);
   U14999 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_61_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_573_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1597_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n93);
   U15000 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_189_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_701_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1725_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n835);
   U15001 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_29_port, A2 
                           => n3066, B1 => DataPath_RF_bus_reg_dataout_541_port
                           , B2 => n3121, C1 => 
                           DataPath_RF_bus_reg_dataout_1565_port, C2 => n3167, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n589);
   U15002 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_157_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_669_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1693_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n905);
   U15003 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_253_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_765_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1789_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n691);
   U15004 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_445_port, A2 
                           => n3079, B1 => DataPath_RF_bus_reg_dataout_957_port
                           , B2 => n3134, C1 => 
                           DataPath_RF_bus_reg_dataout_1981_port, C2 => n3180, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n265);
   U15005 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_349_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_861_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1885_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n479);
   U15006 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_285_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_797_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1821_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n621);
   U15007 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_413_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_925_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1949_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n335);
   U15008 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_317_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_829_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1853_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n549);
   U15009 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_381_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_893_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1917_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n407);
   U15010 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_222_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_734_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1758_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n759);
   U15011 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_126_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_638_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1662_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n973);
   U15012 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_62_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_574_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1598_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n91);
   U15013 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_190_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_702_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1726_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n831);
   U15014 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_30_port, A2 
                           => n3067, B1 => DataPath_RF_bus_reg_dataout_542_port
                           , B2 => n3122, C1 => 
                           DataPath_RF_bus_reg_dataout_1566_port, C2 => n3168, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n565);
   U15015 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_158_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_670_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1694_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n903);
   U15016 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_254_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_766_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1790_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n689);
   U15017 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_446_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_958_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1982_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n263);
   U15018 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_350_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_862_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1886_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n475);
   U15019 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_286_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_798_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1822_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n619);
   U15020 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_414_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_926_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1950_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n333);
   U15021 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_318_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_830_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1854_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n547);
   U15022 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_382_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_894_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1918_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n405);
   U15023 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_223_port, A2 
                           => n3059, B1 => DataPath_RF_bus_reg_dataout_735_port
                           , B2 => n3114, C1 => 
                           DataPath_RF_bus_reg_dataout_1759_port, C2 => n3160, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n757);
   U15024 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_127_port, A2 
                           => n3050, B1 => DataPath_RF_bus_reg_dataout_639_port
                           , B2 => n3105, C1 => 
                           DataPath_RF_bus_reg_dataout_1663_port, C2 => n3151, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n971);
   U15025 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_63_port, A2 
                           => n3087, B1 => DataPath_RF_bus_reg_dataout_575_port
                           , B2 => n3142, C1 => 
                           DataPath_RF_bus_reg_dataout_1599_port, C2 => n3188, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n89);
   U15026 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_191_port, A2 
                           => n3056, B1 => DataPath_RF_bus_reg_dataout_703_port
                           , B2 => n3111, C1 => 
                           DataPath_RF_bus_reg_dataout_1727_port, C2 => n3157, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n829);
   U15027 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_31_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_543_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1567_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n543);
   U15028 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_159_port, A2 
                           => n3053, B1 => DataPath_RF_bus_reg_dataout_671_port
                           , B2 => n3108, C1 => 
                           DataPath_RF_bus_reg_dataout_1695_port, C2 => n3154, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n901);
   U15029 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_255_port, A2 
                           => n3062, B1 => DataPath_RF_bus_reg_dataout_767_port
                           , B2 => n3117, C1 => 
                           DataPath_RF_bus_reg_dataout_1791_port, C2 => n3163, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n687);
   U15030 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_447_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_959_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1983_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n261);
   U15031 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_351_port, A2 
                           => n3071, B1 => DataPath_RF_bus_reg_dataout_863_port
                           , B2 => n3126, C1 => 
                           DataPath_RF_bus_reg_dataout_1887_port, C2 => n3172, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n473);
   U15032 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_287_port, A2 
                           => n3065, B1 => DataPath_RF_bus_reg_dataout_799_port
                           , B2 => n3120, C1 => 
                           DataPath_RF_bus_reg_dataout_1823_port, C2 => n3166, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n617);
   U15033 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_415_port, A2 
                           => n3077, B1 => DataPath_RF_bus_reg_dataout_927_port
                           , B2 => n3132, C1 => 
                           DataPath_RF_bus_reg_dataout_1951_port, C2 => n3178, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n331);
   U15034 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_319_port, A2 
                           => n3068, B1 => DataPath_RF_bus_reg_dataout_831_port
                           , B2 => n3123, C1 => 
                           DataPath_RF_bus_reg_dataout_1855_port, C2 => n3169, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n545);
   U15035 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_383_port, A2 
                           => n3074, B1 => DataPath_RF_bus_reg_dataout_895_port
                           , B2 => n3129, C1 => 
                           DataPath_RF_bus_reg_dataout_1919_port, C2 => n3175, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n403);
   U15036 : OAI22_X1 port map( A1 => n3904, A2 => DataPath_RF_PUSH_ADDRGEN_n12,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n39, B2 => 
                           DataPath_RF_n10, ZN => 
                           DataPath_RF_spill_address_ext_6_port);
   U15037 : OAI22_X1 port map( A1 => n3904, A2 => DataPath_RF_PUSH_ADDRGEN_n11,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n38, B2 => 
                           DataPath_RF_n10, ZN => 
                           DataPath_RF_spill_address_ext_7_port);
   U15038 : OAI22_X1 port map( A1 => n3902, A2 => DataPath_RF_PUSH_ADDRGEN_n5, 
                           B1 => DataPath_RF_PUSH_ADDRGEN_n47, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_13_port);
   U15039 : OAI22_X1 port map( A1 => n3902, A2 => DataPath_RF_PUSH_ADDRGEN_n8, 
                           B1 => DataPath_RF_PUSH_ADDRGEN_n50, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_10_port);
   U15040 : OAI22_X1 port map( A1 => n3902, A2 => DataPath_RF_PUSH_ADDRGEN_n6, 
                           B1 => DataPath_RF_PUSH_ADDRGEN_n48, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_12_port);
   U15041 : OAI22_X1 port map( A1 => n3905, A2 => DataPath_RF_PUSH_ADDRGEN_n9, 
                           B1 => DataPath_RF_PUSH_ADDRGEN_n36, B2 => 
                           DataPath_RF_n10, ZN => 
                           DataPath_RF_spill_address_ext_9_port);
   U15042 : OAI22_X1 port map( A1 => n3905, A2 => DataPath_RF_PUSH_ADDRGEN_n10,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n37, B2 => 
                           DataPath_RF_n10, ZN => 
                           DataPath_RF_spill_address_ext_8_port);
   U15043 : OAI22_X1 port map( A1 => n3901, A2 => DataPath_RF_PUSH_ADDRGEN_n18,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n51, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_0_port);
   U15044 : OAI22_X1 port map( A1 => n3903, A2 => DataPath_RF_PUSH_ADDRGEN_n16,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n43, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_2_port);
   U15045 : OAI22_X1 port map( A1 => n3903, A2 => DataPath_RF_PUSH_ADDRGEN_n17,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n44, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_1_port);
   U15046 : OAI22_X1 port map( A1 => n3903, A2 => DataPath_RF_PUSH_ADDRGEN_n15,
                           B1 => DataPath_RF_PUSH_ADDRGEN_n42, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_3_port);
   U15047 : OAI22_X1 port map( A1 => n3902, A2 => DataPath_RF_PUSH_ADDRGEN_n7, 
                           B1 => DataPath_RF_PUSH_ADDRGEN_n49, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_11_port);
   U15048 : OAI22_X1 port map( A1 => n3903, A2 => DataPath_RF_PUSH_ADDRGEN_n4, 
                           B1 => DataPath_RF_PUSH_ADDRGEN_n46, B2 => 
                           DataPath_RF_n10, ZN => 
                           DataPath_RF_spill_address_ext_14_port);
   U15049 : OAI22_X1 port map( A1 => n3905, A2 => DataPath_RF_PUSH_ADDRGEN_n1, 
                           B1 => DataPath_RF_PUSH_ADDRGEN_n45, B2 => n3900, ZN 
                           => DataPath_RF_spill_address_ext_15_port);
   U15050 : NOR3_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n3889, A3 
                           => n11604, ZN => DataPath_RF_SELBLOCK_INLOC_n9);
   U15051 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1120_port, A2 
                           => n3246, B1 => 
                           DataPath_RF_bus_reg_dataout_2144_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n16);
   U15052 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1121_port, A2 
                           => n3246, B1 => 
                           DataPath_RF_bus_reg_dataout_2145_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n14);
   U15053 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1122_port, A2 
                           => n3246, B1 => 
                           DataPath_RF_bus_reg_dataout_2146_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n12);
   U15054 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1123_port, A2 
                           => n3246, B1 => 
                           DataPath_RF_bus_reg_dataout_2147_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n10);
   U15055 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1033_port, A2 
                           => n3246, B1 => n3890, B2 => 
                           DataPath_RF_bus_reg_dataout_2057_port, ZN => 
                           DataPath_RF_SELBLOCK_INLOC_n4);
   U15056 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1117_port, A2 
                           => n3246, B1 => 
                           DataPath_RF_bus_reg_dataout_2141_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n22);
   U15057 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1118_port, A2 
                           => n3246, B1 => 
                           DataPath_RF_bus_reg_dataout_2142_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n20);
   U15058 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1119_port, A2 
                           => n3246, B1 => 
                           DataPath_RF_bus_reg_dataout_2143_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n18);
   U15059 : NOR3_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n3889, A3 
                           => DataPath_RF_c_swin_2_port, ZN => 
                           DataPath_RF_SELBLOCK_INLOC_n1032);
   U15060 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_195_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_99_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n89);
   U15061 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n820, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n821, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_195_port);
   U15062 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n10, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n11, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_99_port);
   U15063 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1219_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2243_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n820);
   U15064 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_419_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_323_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n85);
   U15065 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n534, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n535, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_323_port);
   U15066 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n322, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n323, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_419_port);
   U15067 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1347_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2371_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n534);
   U15068 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_196_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_100_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n79);
   U15069 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1028, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1029, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_100_port);
   U15070 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n818, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n819, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_196_port);
   U15071 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1124_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2148_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1028);
   U15072 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_420_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_324_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n75);
   U15073 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n532, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n533, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_324_port);
   U15074 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n318, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n319, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_420_port);
   U15075 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1348_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2372_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n532);
   U15076 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_197_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_101_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n69);
   U15077 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1026, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1027, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_101_port);
   U15078 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n816, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n817, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_197_port);
   U15079 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1125_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2149_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1026);
   U15080 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_421_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_325_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n65);
   U15081 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n530, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n531, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_325_port);
   U15082 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n316, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n317, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_421_port);
   U15083 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1349_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2373_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n530);
   U15084 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_198_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_102_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n59);
   U15085 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1024, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1025, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_102_port);
   U15086 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n814, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n815, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_198_port);
   U15087 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1126_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2150_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1024);
   U15088 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_422_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_326_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n55);
   U15089 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n528, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n529, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_326_port);
   U15090 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n314, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n315, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_422_port);
   U15091 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1350_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2374_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n528);
   U15092 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_199_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_103_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n49);
   U15093 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1022, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1023, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_103_port);
   U15094 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n812, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n813, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_199_port);
   U15095 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1127_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2151_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1022);
   U15096 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_423_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_327_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n45);
   U15097 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n526, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n527, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_327_port);
   U15098 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n312, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n313, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_423_port);
   U15099 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1351_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2375_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n526);
   U15100 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_200_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_104_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n39);
   U15101 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1020, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1021, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_104_port);
   U15102 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n806, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n807, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_200_port);
   U15103 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1128_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2152_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1020);
   U15104 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_424_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_328_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n35);
   U15105 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n524, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n525, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_328_port);
   U15106 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n310, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n311, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_424_port);
   U15107 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1352_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2376_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n524);
   U15108 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_201_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_105_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n21);
   U15109 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1018, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1019, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_105_port);
   U15110 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n804, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n805, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_201_port);
   U15111 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1129_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2153_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1018);
   U15112 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_425_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_329_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n9);
   U15113 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n522, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n523, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_329_port);
   U15114 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n308, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n309, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_425_port);
   U15115 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1353_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2377_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n522);
   U15116 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_223_port
                           , A2 => n3014, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_127_port, B2 => 
                           n3017, ZN => DataPath_RF_RDPORT_SPILL_n99);
   U15117 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n970, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n971, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_127_port);
   U15118 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n756, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n757, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_223_port);
   U15119 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1151_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2175_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n970);
   U15120 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_447_port
                           , A2 => n2990, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_351_port, B2 => 
                           n2993, ZN => DataPath_RF_RDPORT_SPILL_n95);
   U15121 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n472, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n473, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_351_port);
   U15122 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n260, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n261, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_447_port);
   U15123 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1375_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2399_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n472);
   U15124 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_192_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_96_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n345);
   U15125 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n826, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n827, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_192_port);
   U15126 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n16, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n17, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_96_port);
   U15127 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1216_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2240_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n826);
   U15128 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_416_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_320_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n335);
   U15129 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n540, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n541, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_320_port);
   U15130 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n328, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n329, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_416_port);
   U15131 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1344_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2368_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n540);
   U15132 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_193_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_97_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n229);
   U15133 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n824, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n825, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_193_port);
   U15134 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n14, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n15, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_97_port);
   U15135 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1217_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2241_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n824);
   U15136 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_417_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_321_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n225);
   U15137 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n538, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n539, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_321_port);
   U15138 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n326, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n327, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_417_port);
   U15139 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1345_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2369_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n538);
   U15140 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_194_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_98_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n119);
   U15141 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n822, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n823, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_194_port);
   U15142 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n12, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n13, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_98_port);
   U15143 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1218_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2242_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n822);
   U15144 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_418_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_322_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n115);
   U15145 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n536, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n537, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_322_port);
   U15146 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n324, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n325, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_418_port);
   U15147 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1346_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2370_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n536);
   U15148 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_202_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_106_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n329);
   U15149 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1016, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1017, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_106_port);
   U15150 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n802, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n803, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_202_port);
   U15151 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1130_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2154_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1016);
   U15152 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_426_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_330_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n325);
   U15153 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n518, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n519, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_330_port);
   U15154 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n306, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n307, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_426_port);
   U15155 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1354_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2378_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n518);
   U15156 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_203_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_107_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n319);
   U15157 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1014, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1015, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_107_port);
   U15158 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n800, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n801, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_203_port);
   U15159 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1131_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2155_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1014);
   U15160 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_427_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_331_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n315);
   U15161 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n516, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n517, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_331_port);
   U15162 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n304, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n305, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_427_port);
   U15163 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1355_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2379_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n516);
   U15164 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_204_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_108_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n309);
   U15165 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1012, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1013, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_108_port);
   U15166 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n798, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n799, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_204_port);
   U15167 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1132_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2156_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1012);
   U15168 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_428_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_332_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n305);
   U15169 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n514, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n515, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_332_port);
   U15170 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n302, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n303, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_428_port);
   U15171 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1356_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2380_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n514);
   U15172 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_205_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_109_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n299);
   U15173 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1010, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1011, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_109_port);
   U15174 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n796, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n797, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_205_port);
   U15175 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1133_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2157_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1010);
   U15176 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_429_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_333_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n295);
   U15177 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n512, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n513, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_333_port);
   U15178 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n300, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n301, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_429_port);
   U15179 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1357_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2381_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n512);
   U15180 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_206_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_110_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n289);
   U15181 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1006, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1007, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_110_port);
   U15182 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n794, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n795, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_206_port);
   U15183 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1134_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2158_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1006);
   U15184 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_430_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_334_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n285);
   U15185 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n510, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n511, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_334_port);
   U15186 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n296, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n297, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_430_port);
   U15187 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1358_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2382_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n510);
   U15188 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_207_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_111_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n279);
   U15189 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1004, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1005, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_111_port);
   U15190 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n792, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n793, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_207_port);
   U15191 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1135_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2159_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1004);
   U15192 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_431_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_335_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n275);
   U15193 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n508, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n509, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_335_port);
   U15194 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n294, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n295, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_431_port);
   U15195 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1359_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2383_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n508);
   U15196 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_208_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_112_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n269);
   U15197 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1002, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1003, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_112_port);
   U15198 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n790, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n791, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_208_port);
   U15199 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1136_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2160_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1002);
   U15200 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_432_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_336_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n265);
   U15201 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n506, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n507, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_336_port);
   U15202 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n292, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n293, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_432_port);
   U15203 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1360_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2384_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n506);
   U15204 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_209_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_113_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n259);
   U15205 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1000, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1001, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_113_port);
   U15206 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n788, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n789, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_209_port);
   U15207 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1137_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2161_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1000);
   U15208 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_433_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_337_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n255);
   U15209 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n504, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n505, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_337_port);
   U15210 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n290, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n291, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_433_port);
   U15211 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1361_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2385_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n504);
   U15212 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_210_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_114_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n249);
   U15213 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n998, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n999, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_114_port);
   U15214 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n784, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n785, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_210_port);
   U15215 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1138_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2162_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n998);
   U15216 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_434_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_338_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n245);
   U15217 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n502, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n503, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_338_port);
   U15218 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n288, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n289, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_434_port);
   U15219 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1362_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2386_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n502);
   U15220 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_211_port
                           , A2 => n3012, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_115_port, B2 => 
                           n3015, ZN => DataPath_RF_RDPORT_SPILL_n239);
   U15221 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n996, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n997, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_115_port);
   U15222 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n782, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n783, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_211_port);
   U15223 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1139_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2163_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n996);
   U15224 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_435_port
                           , A2 => n2988, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_339_port, B2 => 
                           n2991, ZN => DataPath_RF_RDPORT_SPILL_n235);
   U15225 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n500, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n501, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_339_port);
   U15226 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n286, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n287, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_435_port);
   U15227 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1363_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2387_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n500);
   U15228 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_212_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_116_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n219);
   U15229 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n994, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n995, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_116_port);
   U15230 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n780, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n781, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_212_port);
   U15231 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1140_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2164_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n994);
   U15232 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_436_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_340_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n215);
   U15233 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n496, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n497, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_340_port);
   U15234 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n284, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n285, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_436_port);
   U15235 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1364_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2388_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n496);
   U15236 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_213_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_117_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n209);
   U15237 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n992, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n993, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_117_port);
   U15238 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n778, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n779, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_213_port);
   U15239 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1141_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2165_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n992);
   U15240 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_437_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_341_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n205);
   U15241 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n494, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n495, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_341_port);
   U15242 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n282, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n283, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_437_port);
   U15243 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1365_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2389_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n494);
   U15244 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_214_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_118_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n199);
   U15245 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n990, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n991, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_118_port);
   U15246 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n776, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n777, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_214_port);
   U15247 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1142_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2166_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n990);
   U15248 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_438_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_342_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n195);
   U15249 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n492, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n493, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_342_port);
   U15250 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n280, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n281, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_438_port);
   U15251 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1366_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2390_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n492);
   U15252 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_215_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_119_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n189);
   U15253 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n988, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n989, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_119_port);
   U15254 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n774, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n775, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_215_port);
   U15255 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1143_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2167_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n988);
   U15256 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_439_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_343_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n185);
   U15257 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n490, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n491, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_343_port);
   U15258 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n278, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n279, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_439_port);
   U15259 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1367_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2391_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n490);
   U15260 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_216_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_120_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n179);
   U15261 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n984, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n985, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_120_port);
   U15262 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n772, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n773, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_216_port);
   U15263 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1144_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2168_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n984);
   U15264 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_440_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_344_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n175);
   U15265 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n488, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n489, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_344_port);
   U15266 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n274, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n275, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_440_port);
   U15267 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1368_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2392_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n488);
   U15268 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_217_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_121_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n169);
   U15269 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n982, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n983, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_121_port);
   U15270 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n770, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n771, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_217_port);
   U15271 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1145_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2169_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n982);
   U15272 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_441_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_345_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n165);
   U15273 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n486, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n487, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_345_port);
   U15274 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n272, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n273, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_441_port);
   U15275 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1369_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2393_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n486);
   U15276 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_218_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_122_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n159);
   U15277 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n980, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n981, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_122_port);
   U15278 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n768, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n769, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_218_port);
   U15279 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1146_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2170_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n980);
   U15280 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_442_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_346_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n155);
   U15281 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n484, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n485, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_346_port);
   U15282 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n270, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n271, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_442_port);
   U15283 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1370_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2394_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n484);
   U15284 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_219_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_123_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n149);
   U15285 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n978, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n979, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_123_port);
   U15286 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n766, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n767, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_219_port);
   U15287 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1147_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2171_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n978);
   U15288 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_443_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_347_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n145);
   U15289 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n482, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n483, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_347_port);
   U15290 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n268, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n269, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_443_port);
   U15291 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1371_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2395_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n482);
   U15292 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_220_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_124_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n139);
   U15293 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n976, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n977, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_124_port);
   U15294 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n762, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n763, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_220_port);
   U15295 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1148_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2172_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n976);
   U15296 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_444_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_348_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n135);
   U15297 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n480, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n481, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_348_port);
   U15298 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n266, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n267, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_444_port);
   U15299 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1372_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2396_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n480);
   U15300 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_221_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_125_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n129);
   U15301 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n974, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n975, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_125_port);
   U15302 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n760, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n761, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_221_port);
   U15303 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1149_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2173_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n974);
   U15304 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_445_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_349_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n125);
   U15305 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n478, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n479, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_349_port);
   U15306 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n264, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n265, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_445_port);
   U15307 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1373_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2397_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n478);
   U15308 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_222_port
                           , A2 => n3013, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_126_port, B2 => 
                           n3016, ZN => DataPath_RF_RDPORT_SPILL_n109);
   U15309 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n972, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n973, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_126_port);
   U15310 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n758, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n759, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_222_port);
   U15311 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1150_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2174_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n972);
   U15312 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_446_port
                           , A2 => n2989, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_350_port, B2 => 
                           n2992, ZN => DataPath_RF_RDPORT_SPILL_n105);
   U15313 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n474, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n475, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_350_port);
   U15314 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n262, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n263, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_446_port);
   U15315 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1374_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2398_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n474);
   U15316 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_35_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_163_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n88);
   U15317 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n890, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n891, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_163_port);
   U15318 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n454, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n455, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_35_port);
   U15319 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1187_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2211_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n890);
   U15320 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_259_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_387_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n84);
   U15321 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n394, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n395, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_387_port);
   U15322 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n678, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n679, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_259_port);
   U15323 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1411_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2435_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n394);
   U15324 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_36_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_164_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n78);
   U15325 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n888, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n889, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_164_port);
   U15326 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n432, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n433, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_36_port);
   U15327 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1188_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2212_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n888);
   U15328 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_260_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_388_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n74);
   U15329 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n392, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n393, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_388_port);
   U15330 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n674, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n675, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_260_port);
   U15331 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1412_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2436_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n392);
   U15332 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_37_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_165_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n68);
   U15333 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n886, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n887, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_165_port);
   U15334 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n410, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n411, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_37_port);
   U15335 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1189_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2213_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n886);
   U15336 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_261_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_389_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n64);
   U15337 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n390, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n391, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_389_port);
   U15338 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n672, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n673, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_261_port);
   U15339 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1413_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2437_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n390);
   U15340 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_38_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_166_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n58);
   U15341 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n884, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n885, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_166_port);
   U15342 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n388, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n389, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_38_port);
   U15343 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1190_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2214_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n884);
   U15344 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_262_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_390_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n54);
   U15345 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n386, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n387, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_390_port);
   U15346 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n670, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n671, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_262_port);
   U15347 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1414_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2438_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n386);
   U15348 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_39_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_167_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n48);
   U15349 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n882, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n883, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_167_port);
   U15350 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n366, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n367, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_39_port);
   U15351 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1191_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2215_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n882);
   U15352 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_263_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_391_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n44);
   U15353 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n384, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n385, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_391_port);
   U15354 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n668, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n669, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_263_port);
   U15355 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1415_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2439_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n384);
   U15356 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_40_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_168_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n38);
   U15357 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n880, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n881, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_168_port);
   U15358 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n342, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n343, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_40_port);
   U15359 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1192_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2216_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n880);
   U15360 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_264_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_392_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n34);
   U15361 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n382, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n383, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_392_port);
   U15362 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n666, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n667, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_264_port);
   U15363 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1416_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2440_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n382);
   U15364 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_41_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_169_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n20);
   U15365 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n878, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n879, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_169_port);
   U15366 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n320, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n321, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_41_port);
   U15367 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1193_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2217_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n878);
   U15368 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_265_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_393_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n8);
   U15369 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n380, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n381, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_393_port);
   U15370 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n664, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n665, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_265_port);
   U15371 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1417_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2441_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n380);
   U15372 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_63_port,
                           A2 => n3020, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_191_port, B2 => 
                           n3023, ZN => DataPath_RF_RDPORT_SPILL_n98);
   U15373 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n828, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n829, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_191_port);
   U15374 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n88, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n89, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_63_port);
   U15375 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1215_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2239_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n828);
   U15376 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_287_port
                           , A2 => n2996, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_415_port, B2 => 
                           n2999, ZN => DataPath_RF_RDPORT_SPILL_n94);
   U15377 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n330, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n331, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_415_port);
   U15378 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n616, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n617, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_287_port);
   U15379 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1439_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2463_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n330);
   U15380 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_67_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_3_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n87);
   U15381 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n364, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n365, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_3_port);
   U15382 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n80, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n81, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_67_port);
   U15383 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1027_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2051_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n364);
   U15384 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_291_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_355_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n83);
   U15385 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n464, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n465, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_355_port);
   U15386 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n606, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n607, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_291_port);
   U15387 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1379_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2403_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n464);
   U15388 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_68_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_4_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n77);
   U15389 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n142, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n143, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_4_port);
   U15390 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n78, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n79, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_68_port);
   U15391 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1028_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2052_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n142);
   U15392 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_292_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_356_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n73);
   U15393 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n462, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n463, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_356_port);
   U15394 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n604, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n605, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_292_port);
   U15395 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1380_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2404_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n462);
   U15396 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_69_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_5_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n67);
   U15397 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n96, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n97, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_5_port);
   U15398 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n76, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n77, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_69_port);
   U15399 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1029_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2053_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n96);
   U15400 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_293_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_357_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n63);
   U15401 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n460, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n461, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_357_port);
   U15402 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n602, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n603, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_293_port);
   U15403 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1381_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2405_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n460);
   U15404 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_70_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_6_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n57);
   U15405 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n74, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n75, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_6_port);
   U15406 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n72, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n73, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_70_port);
   U15407 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1030_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2054_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n74);
   U15408 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_294_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_358_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n53);
   U15409 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n458, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n459, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_358_port);
   U15410 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n600, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n601, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_294_port);
   U15411 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1382_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2406_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n458);
   U15412 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_71_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_7_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n47);
   U15413 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n52, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n53, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_7_port);
   U15414 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n70, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n71, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_71_port);
   U15415 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1031_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2055_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n52);
   U15416 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_295_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_359_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n43);
   U15417 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n456, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n457, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_359_port);
   U15418 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n598, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n599, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_295_port);
   U15419 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1383_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2407_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n456);
   U15420 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_72_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_8_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n37);
   U15421 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n30, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n31, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_8_port);
   U15422 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n68, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n69, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_72_port);
   U15423 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1032_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2056_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n30);
   U15424 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_296_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_360_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n33);
   U15425 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n452, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n453, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_360_port);
   U15426 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n596, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n597, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_296_port);
   U15427 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1384_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2408_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n452);
   U15428 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_73_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_9_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n19);
   U15429 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n66, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n67, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_73_port);
   U15430 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n4, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n5, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_9_port);
   U15431 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1097_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2121_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n66);
   U15432 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_297_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_361_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n7);
   U15433 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n450, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n451, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_361_port);
   U15434 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n594, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n595, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_297_port);
   U15435 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1385_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2409_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n450);
   U15436 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_95_port,
                           A2 => n3026, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_31_port, B2 => 
                           n3029, ZN => DataPath_RF_RDPORT_SPILL_n97);
   U15437 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n542, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n543, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_31_port);
   U15438 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n18, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n19, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_95_port);
   U15439 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1055_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2079_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n542);
   U15440 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_319_port
                           , A2 => n3002, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_383_port, B2 => 
                           n3005, ZN => DataPath_RF_RDPORT_SPILL_n93);
   U15441 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n402, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n403, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_383_port);
   U15442 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n544, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n545, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_319_port);
   U15443 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1407_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2431_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n402);
   U15444 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_32_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_160_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n344);
   U15445 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n896, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n897, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_160_port);
   U15446 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n520, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n521, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_32_port);
   U15447 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1184_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2208_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n896);
   U15448 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_256_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_384_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n334);
   U15449 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n400, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n401, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_384_port);
   U15450 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n684, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n685, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_256_port);
   U15451 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1408_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2432_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n400);
   U15452 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_33_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_161_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n228);
   U15453 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n894, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n895, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_161_port);
   U15454 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n498, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n499, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_33_port);
   U15455 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1185_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2209_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n894);
   U15456 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_257_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_385_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n224);
   U15457 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n398, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n399, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_385_port);
   U15458 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n682, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n683, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_257_port);
   U15459 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1409_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2433_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n398);
   U15460 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_34_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_162_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n118);
   U15461 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n892, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n893, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_162_port);
   U15462 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n476, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n477, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_34_port);
   U15463 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1186_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2210_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n892);
   U15464 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_258_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_386_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n114);
   U15465 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n396, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n397, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_386_port);
   U15466 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n680, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n681, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_258_port);
   U15467 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1410_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2434_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n396);
   U15468 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_42_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_170_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n328);
   U15469 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n874, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n875, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_170_port);
   U15470 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n298, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n299, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_42_port);
   U15471 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1194_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2218_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n874);
   U15472 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_266_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_394_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n324);
   U15473 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n378, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n379, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_394_port);
   U15474 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n662, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n663, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_266_port);
   U15475 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1418_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2442_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n378);
   U15476 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_43_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_171_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n318);
   U15477 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n872, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n873, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_171_port);
   U15478 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n276, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n277, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_43_port);
   U15479 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1195_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2219_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n872);
   U15480 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_267_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_395_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n314);
   U15481 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n376, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n377, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_395_port);
   U15482 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n660, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n661, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_267_port);
   U15483 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1419_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2443_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n376);
   U15484 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_44_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_172_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n308);
   U15485 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n870, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n871, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_172_port);
   U15486 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n254, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n255, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_44_port);
   U15487 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1196_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2220_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n870);
   U15488 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_268_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_396_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n304);
   U15489 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n374, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n375, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_396_port);
   U15490 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n658, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n659, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_268_port);
   U15491 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1420_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2444_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n374);
   U15492 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_45_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_173_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n298);
   U15493 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n868, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n869, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_173_port);
   U15494 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n232, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n233, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_45_port);
   U15495 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1197_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2221_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n868);
   U15496 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_269_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_397_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n294);
   U15497 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n372, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n373, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_397_port);
   U15498 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n656, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n657, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_269_port);
   U15499 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1421_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2445_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n372);
   U15500 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_46_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_174_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n288);
   U15501 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n866, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n867, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_174_port);
   U15502 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n210, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n211, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_46_port);
   U15503 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1198_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2222_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n866);
   U15504 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_270_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_398_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n284);
   U15505 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n370, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n371, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_398_port);
   U15506 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n652, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n653, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_270_port);
   U15507 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1422_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2446_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n370);
   U15508 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_47_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_175_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n278);
   U15509 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n864, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n865, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_175_port);
   U15510 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n188, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n189, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_47_port);
   U15511 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1199_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2223_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n864);
   U15512 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_271_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_399_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n274);
   U15513 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n368, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n369, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_399_port);
   U15514 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n650, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n651, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_271_port);
   U15515 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1423_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2447_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n368);
   U15516 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_48_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_176_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n268);
   U15517 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n862, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n863, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_176_port);
   U15518 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n166, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n167, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_48_port);
   U15519 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1200_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2224_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n862);
   U15520 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_272_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_400_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n264);
   U15521 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n362, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n363, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_400_port);
   U15522 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n648, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n649, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_272_port);
   U15523 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1424_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2448_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n362);
   U15524 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_49_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_177_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n258);
   U15525 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n860, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n861, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_177_port);
   U15526 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n144, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n145, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_49_port);
   U15527 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1201_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2225_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n860);
   U15528 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_273_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_401_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n254);
   U15529 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n360, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n361, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_401_port);
   U15530 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n646, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n647, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_273_port);
   U15531 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1425_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2449_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n360);
   U15532 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_50_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_178_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n248);
   U15533 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n858, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n859, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_178_port);
   U15534 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n120, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n121, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_50_port);
   U15535 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1202_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2226_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n858);
   U15536 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_274_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_402_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n244);
   U15537 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n358, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n359, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_402_port);
   U15538 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n644, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n645, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_274_port);
   U15539 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1426_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2450_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n358);
   U15540 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_51_port,
                           A2 => n3018, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_179_port, B2 => 
                           n3021, ZN => DataPath_RF_RDPORT_SPILL_n238);
   U15541 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n856, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n857, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_179_port);
   U15542 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n114, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n115, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_51_port);
   U15543 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1203_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2227_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n856);
   U15544 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_275_port
                           , A2 => n2994, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_403_port, B2 => 
                           n2997, ZN => DataPath_RF_RDPORT_SPILL_n234);
   U15545 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n356, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n357, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_403_port);
   U15546 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n642, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n643, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_275_port);
   U15547 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1427_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2451_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n356);
   U15548 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_52_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_180_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n218);
   U15549 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n852, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n853, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_180_port);
   U15550 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n112, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n113, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_52_port);
   U15551 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1204_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2228_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n852);
   U15552 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_276_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_404_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n214);
   U15553 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n354, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n355, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_404_port);
   U15554 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n640, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n641, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_276_port);
   U15555 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1428_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2452_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n354);
   U15556 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_53_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_181_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n208);
   U15557 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n850, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n851, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_181_port);
   U15558 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n110, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n111, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_53_port);
   U15559 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1205_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2229_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n850);
   U15560 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_277_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_405_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n204);
   U15561 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n352, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n353, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_405_port);
   U15562 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n638, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n639, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_277_port);
   U15563 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1429_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2453_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n352);
   U15564 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_54_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_182_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n198);
   U15565 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n848, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n849, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_182_port);
   U15566 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n108, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n109, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_54_port);
   U15567 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1206_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2230_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n848);
   U15568 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_278_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_406_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n194);
   U15569 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n350, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n351, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_406_port);
   U15570 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n636, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n637, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_278_port);
   U15571 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1430_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2454_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n350);
   U15572 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_55_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_183_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n188);
   U15573 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n846, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n847, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_183_port);
   U15574 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n106, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n107, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_55_port);
   U15575 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1207_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2231_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n846);
   U15576 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_279_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_407_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n184);
   U15577 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n348, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n349, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_407_port);
   U15578 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n634, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n635, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_279_port);
   U15579 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1431_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2455_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n348);
   U15580 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_56_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_184_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n178);
   U15581 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n844, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n845, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_184_port);
   U15582 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n104, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n105, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_56_port);
   U15583 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1208_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2232_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n844);
   U15584 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_280_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_408_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n174);
   U15585 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n346, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n347, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_408_port);
   U15586 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n630, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n631, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_280_port);
   U15587 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1432_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2456_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n346);
   U15588 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_57_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_185_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n168);
   U15589 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n842, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n843, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_185_port);
   U15590 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n102, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n103, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_57_port);
   U15591 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1209_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2233_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n842);
   U15592 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_281_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_409_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n164);
   U15593 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n344, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n345, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_409_port);
   U15594 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n628, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n629, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_281_port);
   U15595 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1433_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2457_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n344);
   U15596 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_58_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_186_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n158);
   U15597 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n840, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n841, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_186_port);
   U15598 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n100, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n101, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_58_port);
   U15599 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1210_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2234_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n840);
   U15600 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_282_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_410_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n154);
   U15601 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n340, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n341, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_410_port);
   U15602 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n626, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n627, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_282_port);
   U15603 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1434_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2458_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n340);
   U15604 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_59_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_187_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n148);
   U15605 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n838, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n839, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_187_port);
   U15606 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n98, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n99, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_59_port);
   U15607 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1211_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2235_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n838);
   U15608 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_283_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_411_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n144);
   U15609 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n338, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n339, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_411_port);
   U15610 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n624, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n625, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_283_port);
   U15611 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1435_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2459_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n338);
   U15612 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_60_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_188_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n138);
   U15613 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n836, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n837, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_188_port);
   U15614 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n94, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n95, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_60_port);
   U15615 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1212_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2236_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n836);
   U15616 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_284_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_412_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n134);
   U15617 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n336, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n337, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_412_port);
   U15618 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n622, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n623, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_284_port);
   U15619 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1436_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2460_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n336);
   U15620 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_61_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_189_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n128);
   U15621 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n834, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n835, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_189_port);
   U15622 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n92, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n93, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_61_port);
   U15623 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1213_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2237_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n834);
   U15624 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_285_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_413_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n124);
   U15625 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n334, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n335, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_413_port);
   U15626 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n620, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n621, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_285_port);
   U15627 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1437_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2461_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n334);
   U15628 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_62_port,
                           A2 => n3019, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_190_port, B2 => 
                           n3022, ZN => DataPath_RF_RDPORT_SPILL_n108);
   U15629 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n830, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n831, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_190_port);
   U15630 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n90, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n91, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_62_port);
   U15631 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1214_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2238_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n830);
   U15632 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_286_port
                           , A2 => n2995, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_414_port, B2 => 
                           n2998, ZN => DataPath_RF_RDPORT_SPILL_n104);
   U15633 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n332, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n333, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_414_port);
   U15634 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n618, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n619, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_286_port);
   U15635 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1438_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2462_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n332);
   U15636 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_64_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_0_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n343);
   U15637 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1030, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1031, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_0_port);
   U15638 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n86, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n87, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_64_port);
   U15639 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1024_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2048_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1030);
   U15640 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_288_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_352_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n333);
   U15641 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n470, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n471, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_352_port);
   U15642 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n614, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n615, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_288_port);
   U15643 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1376_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2400_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n470);
   U15644 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_65_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_1_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n227);
   U15645 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n808, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n809, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_1_port);
   U15646 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n84, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n85, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_65_port);
   U15647 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1025_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2049_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n808);
   U15648 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_289_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_353_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n223);
   U15649 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n468, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n469, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_353_port);
   U15650 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n612, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n613, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_289_port);
   U15651 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1377_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2401_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n468);
   U15652 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_66_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_2_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n117);
   U15653 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n586, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n587, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_2_port);
   U15654 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n82, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n83, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_66_port);
   U15655 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1026_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2050_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n586);
   U15656 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_290_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_354_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n113);
   U15657 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n466, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n467, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_354_port);
   U15658 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n608, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n609, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_290_port);
   U15659 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1378_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2402_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n466);
   U15660 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_74_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_10_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n327);
   U15661 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1008, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1009, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_10_port);
   U15662 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n64, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n65, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_74_port);
   U15663 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1034_port, A2 
                           => n3204, B1 => 
                           DataPath_RF_bus_reg_dataout_2058_port, B2 => n3858, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n1008);
   U15664 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_298_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_362_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n323);
   U15665 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n448, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n449, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_362_port);
   U15666 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n592, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n593, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_298_port);
   U15667 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1386_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2410_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n448);
   U15668 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_75_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_11_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n317);
   U15669 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n986, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n987, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_11_port);
   U15670 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n62, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n63, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_75_port);
   U15671 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1035_port, A2 
                           => n3205, B1 => 
                           DataPath_RF_bus_reg_dataout_2059_port, B2 => n3859, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n986);
   U15672 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_299_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_363_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n313);
   U15673 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n446, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n447, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_363_port);
   U15674 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n590, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n591, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_299_port);
   U15675 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1387_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2411_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n446);
   U15676 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_76_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_12_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n307);
   U15677 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n964, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n965, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_12_port);
   U15678 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n60, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n61, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_76_port);
   U15679 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1036_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2060_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n964);
   U15680 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_300_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_364_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n303);
   U15681 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n444, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n445, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_364_port);
   U15682 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n584, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n585, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_300_port);
   U15683 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1388_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2412_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n444);
   U15684 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_77_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_13_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n297);
   U15685 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n942, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n943, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_13_port);
   U15686 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n58, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n59, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_77_port);
   U15687 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1037_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2061_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n942);
   U15688 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_301_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_365_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n293);
   U15689 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n442, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n443, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_365_port);
   U15690 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n582, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n583, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_301_port);
   U15691 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1389_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2413_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n442);
   U15692 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_78_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_14_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n287);
   U15693 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n920, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n921, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_14_port);
   U15694 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n56, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n57, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_78_port);
   U15695 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1038_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2062_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n920);
   U15696 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_302_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_366_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n283);
   U15697 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n440, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n441, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_366_port);
   U15698 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n580, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n581, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_302_port);
   U15699 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1390_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2414_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n440);
   U15700 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_79_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_15_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n277);
   U15701 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n898, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n899, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_15_port);
   U15702 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n54, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n55, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_79_port);
   U15703 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1039_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2063_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n898);
   U15704 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_303_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_367_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n273);
   U15705 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n438, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n439, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_367_port);
   U15706 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n578, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n579, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_303_port);
   U15707 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1391_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2415_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n438);
   U15708 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_80_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_16_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n267);
   U15709 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n876, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n877, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_16_port);
   U15710 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n50, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n51, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_80_port);
   U15711 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1040_port, A2 
                           => n3210, B1 => 
                           DataPath_RF_bus_reg_dataout_2064_port, B2 => n3864, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n876);
   U15712 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_304_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_368_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n263);
   U15713 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n436, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n437, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_368_port);
   U15714 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n576, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n577, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_304_port);
   U15715 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1392_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2416_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n436);
   U15716 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_81_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_17_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n257);
   U15717 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n854, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n855, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_17_port);
   U15718 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n48, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n49, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_81_port);
   U15719 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1041_port, A2 
                           => n3211, B1 => 
                           DataPath_RF_bus_reg_dataout_2065_port, B2 => n3865, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n854);
   U15720 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_305_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_369_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n253);
   U15721 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n434, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n435, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_369_port);
   U15722 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n574, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n575, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_305_port);
   U15723 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1393_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2417_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n434);
   U15724 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_82_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_18_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n247);
   U15725 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n832, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n833, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_18_port);
   U15726 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n46, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n47, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_82_port);
   U15727 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1042_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2066_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n832);
   U15728 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_306_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_370_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n243);
   U15729 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n430, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n431, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_370_port);
   U15730 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n572, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n573, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_306_port);
   U15731 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1394_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2418_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n430);
   U15732 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_83_port,
                           A2 => n3024, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_19_port, B2 => 
                           n3027, ZN => DataPath_RF_RDPORT_SPILL_n237);
   U15733 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n810, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n811, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_19_port);
   U15734 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n44, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n45, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_83_port);
   U15735 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1043_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2067_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n810);
   U15736 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_307_port
                           , A2 => n3000, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_371_port, B2 => 
                           n3003, ZN => DataPath_RF_RDPORT_SPILL_n233);
   U15737 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n428, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n429, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_371_port);
   U15738 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n570, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n571, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_307_port);
   U15739 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1395_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2419_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n428);
   U15740 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_84_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_20_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n217);
   U15741 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n786, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n787, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_20_port);
   U15742 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n42, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n43, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_84_port);
   U15743 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1044_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2068_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n786);
   U15744 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_308_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_372_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n213);
   U15745 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n426, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n427, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_372_port);
   U15746 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n568, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n569, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_308_port);
   U15747 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1396_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2420_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n426);
   U15748 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_85_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_21_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n207);
   U15749 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n764, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n765, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_21_port);
   U15750 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n40, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n41, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_85_port);
   U15751 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1045_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2069_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n764);
   U15752 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_309_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_373_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n203);
   U15753 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n424, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n425, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_373_port);
   U15754 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n566, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n567, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_309_port);
   U15755 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1397_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2421_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n424);
   U15756 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_86_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_22_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n197);
   U15757 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n742, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n743, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_22_port);
   U15758 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n38, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n39, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_86_port);
   U15759 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1046_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2070_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n742);
   U15760 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_310_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_374_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n193);
   U15761 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n422, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n423, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_374_port);
   U15762 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n562, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n563, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_310_port);
   U15763 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1398_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2422_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n422);
   U15764 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_87_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_23_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n187);
   U15765 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n720, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n721, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_23_port);
   U15766 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n36, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n37, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_87_port);
   U15767 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1047_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2071_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n720);
   U15768 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_311_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_375_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n183);
   U15769 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n420, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n421, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_375_port);
   U15770 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n560, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n561, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_311_port);
   U15771 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1399_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2423_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n420);
   U15772 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_88_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_24_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n177);
   U15773 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n698, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n699, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_24_port);
   U15774 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n34, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n35, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_88_port);
   U15775 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1048_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2072_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n698);
   U15776 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_312_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_376_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n173);
   U15777 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n418, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n419, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_376_port);
   U15778 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n558, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n559, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_312_port);
   U15779 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1400_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2424_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n418);
   U15780 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_89_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_25_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n167);
   U15781 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n676, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n677, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_25_port);
   U15782 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n32, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n33, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_89_port);
   U15783 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1049_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2073_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n676);
   U15784 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_313_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_377_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n163);
   U15785 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n416, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n417, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_377_port);
   U15786 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n556, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n557, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_313_port);
   U15787 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1401_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2425_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n416);
   U15788 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_90_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_26_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n157);
   U15789 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n654, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n655, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_26_port);
   U15790 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n28, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n29, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_90_port);
   U15791 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1050_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2074_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n654);
   U15792 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_314_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_378_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n153);
   U15793 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n414, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n415, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_378_port);
   U15794 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n554, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n555, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_314_port);
   U15795 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1402_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2426_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n414);
   U15796 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_91_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_27_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n147);
   U15797 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n632, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n633, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_27_port);
   U15798 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n26, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n27, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_91_port);
   U15799 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1051_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2075_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n632);
   U15800 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_315_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_379_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n143);
   U15801 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n412, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n413, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_379_port);
   U15802 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n552, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n553, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_315_port);
   U15803 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1403_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2427_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n412);
   U15804 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_92_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_28_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n137);
   U15805 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n610, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n611, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_28_port);
   U15806 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n24, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n25, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_92_port);
   U15807 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1052_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2076_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n610);
   U15808 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_316_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_380_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n133);
   U15809 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n408, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n409, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_380_port);
   U15810 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n550, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n551, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_316_port);
   U15811 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1404_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2428_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n408);
   U15812 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_93_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_29_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n127);
   U15813 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n588, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n589, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_29_port);
   U15814 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n22, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n23, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_93_port);
   U15815 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1053_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2077_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n588);
   U15816 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_317_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_381_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n123);
   U15817 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n406, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n407, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_381_port);
   U15818 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n548, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n549, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_317_port);
   U15819 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1405_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2429_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n406);
   U15820 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_94_port,
                           A2 => n3025, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_30_port, B2 => 
                           n3028, ZN => DataPath_RF_RDPORT_SPILL_n107);
   U15821 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n564, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n565, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_30_port);
   U15822 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n20, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n21, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_94_port);
   U15823 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1054_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2078_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n564);
   U15824 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_318_port
                           , A2 => n3001, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_382_port, B2 => 
                           n3004, ZN => DataPath_RF_RDPORT_SPILL_n103);
   U15825 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n404, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n405, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_382_port);
   U15826 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n546, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n547, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_318_port);
   U15827 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1406_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2430_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n404);
   U15828 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_131_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_227_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n86);
   U15829 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n748, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n749, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_227_port);
   U15830 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n960, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n961, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_131_port);
   U15831 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1251_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2275_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n748);
   U15832 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_132_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_228_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n76);
   U15833 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n746, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n747, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_228_port);
   U15834 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n958, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n959, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_132_port);
   U15835 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1252_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2276_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n746);
   U15836 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_133_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_229_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n66);
   U15837 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n744, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n745, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_229_port);
   U15838 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n956, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n957, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_133_port);
   U15839 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1253_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2277_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n744);
   U15840 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_134_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_230_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n56);
   U15841 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n740, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n741, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_230_port);
   U15842 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n954, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n955, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_134_port);
   U15843 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1254_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2278_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n740);
   U15844 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_135_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_231_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n46);
   U15845 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n738, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n739, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_231_port);
   U15846 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n952, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n953, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_135_port);
   U15847 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1255_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2279_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n738);
   U15848 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_136_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_232_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n36);
   U15849 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n736, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n737, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_232_port);
   U15850 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n950, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n951, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_136_port);
   U15851 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1256_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2280_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n736);
   U15852 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_137_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_233_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n18);
   U15853 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n734, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n735, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_233_port);
   U15854 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n948, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n949, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_137_port);
   U15855 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1257_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2281_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n734);
   U15856 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_159_port
                           , A2 => n3032, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_255_port, B2 => 
                           n3035, ZN => DataPath_RF_RDPORT_SPILL_n96);
   U15857 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n686, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n687, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_255_port);
   U15858 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n900, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n901, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_159_port);
   U15859 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1279_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2303_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n686);
   U15860 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1056_port, A2 
                           => n3225, B1 => 
                           DataPath_RF_bus_reg_dataout_2080_port, B2 => n3857, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n520);
   U15861 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1088_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2112_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n86);
   U15862 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1152_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2176_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n968);
   U15863 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1440_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2464_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n328);
   U15864 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1280_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2304_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n684);
   U15865 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1312_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2336_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n614);
   U15866 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1057_port, A2 
                           => n3226, B1 => 
                           DataPath_RF_bus_reg_dataout_2081_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n498);
   U15867 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1089_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2113_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n84);
   U15868 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1153_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2177_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n966);
   U15869 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1441_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2465_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n326);
   U15870 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1281_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2305_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n682);
   U15871 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1313_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2337_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n612);
   U15872 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1058_port, A2 
                           => n3227, B1 => 
                           DataPath_RF_bus_reg_dataout_2082_port, B2 => n3880, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n476);
   U15873 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1090_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2114_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n82);
   U15874 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1154_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2178_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n962);
   U15875 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1442_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2466_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n324);
   U15876 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1282_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2306_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n680);
   U15877 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1314_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2338_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n608);
   U15878 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1059_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2083_port, B2 => n3881, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n454);
   U15879 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1091_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2115_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n80);
   U15880 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1155_port, A2 
                           => n3206, B1 => 
                           DataPath_RF_bus_reg_dataout_2179_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n960);
   U15881 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1443_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2467_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n322);
   U15882 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1283_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2307_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n678);
   U15883 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1315_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2339_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n606);
   U15884 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1220_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2244_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n818);
   U15885 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1060_port, A2 
                           => n3228, B1 => 
                           DataPath_RF_bus_reg_dataout_2084_port, B2 => n3882, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n432);
   U15886 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1092_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2116_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n78);
   U15887 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1156_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2180_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n958);
   U15888 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1444_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2468_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n318);
   U15889 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1284_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2308_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n674);
   U15890 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1316_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2340_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n604);
   U15891 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1221_port, A2 
                           => n3212, B1 => 
                           DataPath_RF_bus_reg_dataout_2245_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n816);
   U15892 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1061_port, A2 
                           => n3229, B1 => 
                           DataPath_RF_bus_reg_dataout_2085_port, B2 => n3883, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n410);
   U15893 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1093_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2117_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n76);
   U15894 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1157_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2181_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n956);
   U15895 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1445_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2469_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n316);
   U15896 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1285_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2309_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n672);
   U15897 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1317_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2341_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n602);
   U15898 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1222_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2246_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n814);
   U15899 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1062_port, A2 
                           => n3230, B1 => 
                           DataPath_RF_bus_reg_dataout_2086_port, B2 => n3884, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n388);
   U15900 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1094_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2118_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n72);
   U15901 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1158_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2182_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n954);
   U15902 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1446_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2470_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n314);
   U15903 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1286_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2310_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n670);
   U15904 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1318_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2342_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n600);
   U15905 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1223_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2247_port, B2 => n3866, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n812);
   U15906 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1063_port, A2 
                           => n3231, B1 => 
                           DataPath_RF_bus_reg_dataout_2087_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n366);
   U15907 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1095_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2119_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n70);
   U15908 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1159_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2183_port, B2 => n3860, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n952);
   U15909 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1447_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2471_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n312);
   U15910 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1287_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2311_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n668);
   U15911 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1319_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2343_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n598);
   U15912 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1224_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2248_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n806);
   U15913 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1064_port, A2 
                           => n3232, B1 => 
                           DataPath_RF_bus_reg_dataout_2088_port, B2 => n3886, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n342);
   U15914 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1096_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2120_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n68);
   U15915 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1160_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2184_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n950);
   U15916 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1448_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2472_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n310);
   U15917 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1288_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2312_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n666);
   U15918 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1320_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2344_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n596);
   U15919 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1225_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2249_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n804);
   U15920 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1065_port, A2 
                           => n3233, B1 => 
                           DataPath_RF_bus_reg_dataout_2089_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n320);
   U15921 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1161_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2185_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n948);
   U15922 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1449_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2473_port, B2 => n3885, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n308);
   U15923 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1289_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2313_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n664);
   U15924 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1321_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2345_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n594);
   U15925 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1226_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2250_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n802);
   U15926 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1066_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2090_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n298);
   U15927 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1098_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2122_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n64);
   U15928 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1162_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2186_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n946);
   U15929 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1450_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2474_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n306);
   U15930 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1290_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2314_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n662);
   U15931 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1322_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2346_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n592);
   U15932 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1227_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2251_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n800);
   U15933 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1067_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2091_port, B2 => n3889, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n276);
   U15934 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1099_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2123_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n62);
   U15935 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1163_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2187_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n944);
   U15936 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1451_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2475_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n304);
   U15937 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1291_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2315_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n660);
   U15938 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1323_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2347_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n590);
   U15939 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1228_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2252_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n798);
   U15940 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1068_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2092_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n254);
   U15941 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1100_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2124_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n60);
   U15942 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1164_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2188_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n940);
   U15943 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1452_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2476_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n302);
   U15944 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1292_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2316_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n658);
   U15945 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1324_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2348_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n584);
   U15946 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1229_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2253_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n796);
   U15947 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1069_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2093_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n232);
   U15948 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1101_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2125_port, B2 => n3876, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n58);
   U15949 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1165_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2189_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n938);
   U15950 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1453_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2477_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n300);
   U15951 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1293_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2317_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n656);
   U15952 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1325_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2349_port, B2 => n3854, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n582);
   U15953 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1230_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2254_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n794);
   U15954 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1070_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2094_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n210);
   U15955 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1102_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2126_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n56);
   U15956 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1166_port, A2 
                           => n3207, B1 => 
                           DataPath_RF_bus_reg_dataout_2190_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n936);
   U15957 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1454_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2478_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n296);
   U15958 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1294_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2318_port, B2 => n3851, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n652);
   U15959 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1326_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2350_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n580);
   U15960 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1231_port, A2 
                           => n3213, B1 => 
                           DataPath_RF_bus_reg_dataout_2255_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n792);
   U15961 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1071_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2095_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n188);
   U15962 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1103_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2127_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n54);
   U15963 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1167_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2191_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n934);
   U15964 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1455_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2479_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n294);
   U15965 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1295_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2319_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n650);
   U15966 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1327_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2351_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n578);
   U15967 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1232_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2256_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n790);
   U15968 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1072_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2096_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n166);
   U15969 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1104_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2128_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n50);
   U15970 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1168_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2192_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n932);
   U15971 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1456_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2480_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n292);
   U15972 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1296_port, A2 
                           => n3219, B1 => 
                           DataPath_RF_bus_reg_dataout_2320_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n648);
   U15973 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1328_port, A2 
                           => n3222, B1 => 
                           DataPath_RF_bus_reg_dataout_2352_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n576);
   U15974 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1233_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2257_port, B2 => n3867, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n788);
   U15975 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1073_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2097_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n144);
   U15976 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1105_port, A2 
                           => n3244, B1 => 
                           DataPath_RF_bus_reg_dataout_2129_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n48);
   U15977 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1169_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2193_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n930);
   U15978 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1457_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2481_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n290);
   U15979 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1297_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2321_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n646);
   U15980 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1329_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2353_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n574);
   U15981 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1234_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2258_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n784);
   U15982 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1074_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2098_port, B2 => n3879, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n120);
   U15983 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1106_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2130_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n46);
   U15984 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1170_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2194_port, B2 => n3861, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n928);
   U15985 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1458_port, A2 
                           => n3234, B1 => 
                           DataPath_RF_bus_reg_dataout_2482_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n288);
   U15986 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1298_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2322_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n644);
   U15987 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1330_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2354_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n572);
   U15988 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1235_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2259_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n782);
   U15989 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1075_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2099_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n114);
   U15990 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1107_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2131_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n44);
   U15991 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1171_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2195_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n926);
   U15992 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1459_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2483_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n286);
   U15993 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1299_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2323_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n642);
   U15994 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1331_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2355_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n570);
   U15995 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1236_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2260_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n780);
   U15996 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1076_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2100_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n112);
   U15997 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1108_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2132_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n42);
   U15998 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1172_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2196_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n924);
   U15999 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1460_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2484_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n284);
   U16000 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1300_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2324_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n640);
   U16001 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1332_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2356_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n568);
   U16002 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1237_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2261_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n778);
   U16003 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1077_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2101_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n110);
   U16004 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1109_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2133_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n40);
   U16005 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1173_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2197_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n922);
   U16006 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1461_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2485_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n282);
   U16007 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1301_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2325_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n638);
   U16008 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1333_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2357_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n566);
   U16009 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1238_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2262_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n776);
   U16010 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1078_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2102_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n108);
   U16011 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1110_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2134_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n38);
   U16012 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1174_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2198_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n918);
   U16013 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1462_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2486_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n280);
   U16014 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1302_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2326_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n636);
   U16015 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1334_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2358_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n562);
   U16016 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1239_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2263_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n774);
   U16017 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1079_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2103_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n106);
   U16018 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1111_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2135_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n36);
   U16019 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1175_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2199_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n916);
   U16020 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1463_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2487_port, B2 => n3888, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n278);
   U16021 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1303_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2327_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n634);
   U16022 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1335_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2359_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n560);
   U16023 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1240_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2264_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n772);
   U16024 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1080_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2104_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n104);
   U16025 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1112_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2136_port, B2 => n3877, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n34);
   U16026 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1176_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2200_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n914);
   U16027 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1464_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2488_port, B2 => n3889, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n274);
   U16028 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1304_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2328_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n630);
   U16029 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1336_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2360_port, B2 => n3855, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n558);
   U16030 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1241_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2265_port, B2 => n3852, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n770);
   U16031 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1081_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2105_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n102);
   U16032 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1113_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2137_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n32);
   U16033 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1177_port, A2 
                           => n3208, B1 => 
                           DataPath_RF_bus_reg_dataout_2201_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n912);
   U16034 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1465_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2489_port, B2 => n3889, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n272);
   U16035 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1305_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2329_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n628);
   U16036 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1337_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2361_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n556);
   U16037 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1242_port, A2 
                           => n3214, B1 => 
                           DataPath_RF_bus_reg_dataout_2266_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n768);
   U16038 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1082_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2106_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n100);
   U16039 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1114_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2138_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n28);
   U16040 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1178_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2202_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n910);
   U16041 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1466_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2490_port, B2 => n3889, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n270);
   U16042 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1306_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2330_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n626);
   U16043 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1338_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2362_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n554);
   U16044 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1243_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2267_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n766);
   U16045 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1083_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2107_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n98);
   U16046 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1115_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2139_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n26);
   U16047 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1179_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2203_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n908);
   U16048 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1467_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2491_port, B2 => n3889, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n268);
   U16049 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1307_port, A2 
                           => n3220, B1 => 
                           DataPath_RF_bus_reg_dataout_2331_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n624);
   U16050 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1339_port, A2 
                           => n3223, B1 => 
                           DataPath_RF_bus_reg_dataout_2363_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n552);
   U16051 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1244_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2268_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n762);
   U16052 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1084_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2108_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n94);
   U16053 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1116_port, A2 
                           => n3245, B1 => 
                           DataPath_RF_bus_reg_dataout_2140_port, B2 => n3878, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n24);
   U16054 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1180_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2204_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n906);
   U16055 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1468_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2492_port, B2 => n3889, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n266);
   U16056 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1308_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2332_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n622);
   U16057 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1340_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2364_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n550);
   U16058 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1245_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2269_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n760);
   U16059 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1085_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2109_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n92);
   U16060 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1181_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2205_port, B2 => n3862, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n904);
   U16061 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1469_port, A2 
                           => n3235, B1 => 
                           DataPath_RF_bus_reg_dataout_2493_port, B2 => n3889, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n264);
   U16062 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1309_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2333_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n620);
   U16063 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1341_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2365_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n548);
   U16064 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1246_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2270_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n758);
   U16065 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1086_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2110_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n90);
   U16066 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1182_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2206_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n902);
   U16067 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1470_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2494_port, B2 => n3887, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n262);
   U16068 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1310_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2334_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n618);
   U16069 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1342_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2366_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n546);
   U16070 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1247_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2271_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n756);
   U16071 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1087_port, A2 
                           => n3243, B1 => 
                           DataPath_RF_bus_reg_dataout_2111_port, B2 => n3875, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n88);
   U16072 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1183_port, A2 
                           => n3209, B1 => 
                           DataPath_RF_bus_reg_dataout_2207_port, B2 => n3863, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n900);
   U16073 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1471_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2495_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n260);
   U16074 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1311_port, A2 
                           => n3221, B1 => 
                           DataPath_RF_bus_reg_dataout_2335_port, B2 => n3853, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n616);
   U16075 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1343_port, A2 
                           => n3224, B1 => 
                           DataPath_RF_bus_reg_dataout_2367_port, B2 => n3856, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n544);
   U16076 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_128_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_224_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n342);
   U16077 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n754, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n755, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_224_port);
   U16078 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n968, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n969, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_128_port);
   U16079 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1248_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2272_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n754);
   U16080 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_129_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_225_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n226);
   U16081 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n752, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n753, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_225_port);
   U16082 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n966, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n967, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_129_port);
   U16083 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1249_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2273_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n752);
   U16084 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_130_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_226_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n116);
   U16085 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n750, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n751, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_226_port);
   U16086 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n962, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n963, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_130_port);
   U16087 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1250_port, A2 
                           => n3215, B1 => 
                           DataPath_RF_bus_reg_dataout_2274_port, B2 => n3847, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n750);
   U16088 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_138_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_234_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n326);
   U16089 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n732, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n733, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_234_port);
   U16090 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n946, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n947, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_138_port);
   U16091 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1258_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2282_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n732);
   U16092 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_139_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_235_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n316);
   U16093 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n730, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n731, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_235_port);
   U16094 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n944, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n945, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_139_port);
   U16095 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1259_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2283_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n730);
   U16096 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_140_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_236_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n306);
   U16097 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n728, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n729, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_236_port);
   U16098 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n940, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n941, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_140_port);
   U16099 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1260_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2284_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n728);
   U16100 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_141_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_237_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n296);
   U16101 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n726, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n727, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_237_port);
   U16102 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n938, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n939, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_141_port);
   U16103 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1261_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2285_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n726);
   U16104 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_142_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_238_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n286);
   U16105 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n724, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n725, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_238_port);
   U16106 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n936, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n937, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_142_port);
   U16107 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1262_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2286_port, B2 => n3848, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n724);
   U16108 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_143_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_239_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n276);
   U16109 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n722, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n723, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_239_port);
   U16110 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n934, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n935, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_143_port);
   U16111 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1263_port, A2 
                           => n3216, B1 => 
                           DataPath_RF_bus_reg_dataout_2287_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n722);
   U16112 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_144_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_240_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n266);
   U16113 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n718, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n719, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_240_port);
   U16114 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n932, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n933, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_144_port);
   U16115 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1264_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2288_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n718);
   U16116 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_145_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_241_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n256);
   U16117 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n716, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n717, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_241_port);
   U16118 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n930, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n931, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_145_port);
   U16119 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1265_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2289_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n716);
   U16120 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_146_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_242_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n246);
   U16121 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n714, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n715, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_242_port);
   U16122 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n928, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n929, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_146_port);
   U16123 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1266_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2290_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n714);
   U16124 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_147_port
                           , A2 => n3030, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_243_port, B2 => 
                           n3033, ZN => DataPath_RF_RDPORT_SPILL_n236);
   U16125 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n712, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n713, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_243_port);
   U16126 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n926, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n927, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_147_port);
   U16127 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1267_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2291_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n712);
   U16128 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_148_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_244_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n216);
   U16129 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n710, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n711, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_244_port);
   U16130 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n924, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n925, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_148_port);
   U16131 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1268_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2292_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n710);
   U16132 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_149_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_245_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n206);
   U16133 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n708, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n709, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_245_port);
   U16134 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n922, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n923, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_149_port);
   U16135 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1269_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2293_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n708);
   U16136 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_150_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_246_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n196);
   U16137 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n706, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n707, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_246_port);
   U16138 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n918, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n919, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_150_port);
   U16139 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1270_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2294_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n706);
   U16140 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_151_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_247_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n186);
   U16141 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n704, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n705, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_247_port);
   U16142 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n916, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n917, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_151_port);
   U16143 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1271_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2295_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n704);
   U16144 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_152_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_248_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n176);
   U16145 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n702, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n703, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_248_port);
   U16146 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n914, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n915, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_152_port);
   U16147 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1272_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2296_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n702);
   U16148 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_153_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_249_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n166);
   U16149 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n700, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n701, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_249_port);
   U16150 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n912, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n913, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_153_port);
   U16151 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1273_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2297_port, B2 => n3849, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n700);
   U16152 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_154_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_250_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n156);
   U16153 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n696, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n697, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_250_port);
   U16154 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n910, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n911, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_154_port);
   U16155 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1274_port, A2 
                           => n3217, B1 => 
                           DataPath_RF_bus_reg_dataout_2298_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n696);
   U16156 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_155_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_251_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n146);
   U16157 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n694, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n695, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_251_port);
   U16158 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n908, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n909, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_155_port);
   U16159 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1275_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2299_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n694);
   U16160 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_156_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_252_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n136);
   U16161 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n692, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n693, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_252_port);
   U16162 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n906, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n907, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_156_port);
   U16163 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1276_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2300_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n692);
   U16164 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_157_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_253_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n126);
   U16165 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n690, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n691, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_253_port);
   U16166 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n904, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n905, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_157_port);
   U16167 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1277_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2301_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n690);
   U16168 : AOI22_X1 port map( A1 => DataPath_RF_bus_sel_savedwin_data_158_port
                           , A2 => n3031, B1 => 
                           DataPath_RF_bus_sel_savedwin_data_254_port, B2 => 
                           n3034, ZN => DataPath_RF_RDPORT_SPILL_n106);
   U16169 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n688, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n689, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_254_port);
   U16170 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n902, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n903, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_158_port);
   U16171 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1278_port, A2 
                           => n3218, B1 => 
                           DataPath_RF_bus_reg_dataout_2302_port, B2 => n3850, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n688);
   U16172 : NOR2_X1 port map( A1 => n11605, A2 => n3889, ZN => 
                           DataPath_RF_SELBLOCK_INLOC_n8);
   U16173 : AND3_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n1032, A2 => 
                           n11603, A3 => DataPath_RF_c_swin_0_port, ZN => 
                           DataPath_RF_SELBLOCK_INLOC_n6);
   U16174 : AND2_X1 port map( A1 => DataPath_RF_c_swin_1_port, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n1032, ZN => 
                           DataPath_RF_SELBLOCK_INLOC_n7);
   U16175 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n258, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n259, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_448_port);
   U16176 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1472_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2496_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n258);
   U16177 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_448_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_960_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1984_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n259);
   U16178 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n256, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n257, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_449_port);
   U16179 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1473_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2497_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n256);
   U16180 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_449_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_961_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1985_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n257);
   U16181 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n252, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n253, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_450_port);
   U16182 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1474_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2498_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n252);
   U16183 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_450_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_962_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1986_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n253);
   U16184 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n250, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n251, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_451_port);
   U16185 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1475_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2499_port, B2 => n3868, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n250);
   U16186 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_451_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_963_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1987_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n251);
   U16187 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n248, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n249, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_452_port);
   U16188 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1476_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2500_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n248);
   U16189 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_452_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_964_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1988_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n249);
   U16190 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n246, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n247, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_453_port);
   U16191 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1477_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2501_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n246);
   U16192 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_453_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_965_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1989_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n247);
   U16193 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n244, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n245, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_454_port);
   U16194 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1478_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2502_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n244);
   U16195 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_454_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_966_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1990_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n245);
   U16196 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n242, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n243, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_455_port);
   U16197 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1479_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2503_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n242);
   U16198 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_455_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_967_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1991_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n243);
   U16199 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n240, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n241, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_456_port);
   U16200 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1480_port, A2 
                           => n3236, B1 => 
                           DataPath_RF_bus_reg_dataout_2504_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n240);
   U16201 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_456_port, A2 
                           => n3080, B1 => DataPath_RF_bus_reg_dataout_968_port
                           , B2 => n3135, C1 => 
                           DataPath_RF_bus_reg_dataout_1992_port, C2 => n3181, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n241);
   U16202 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n238, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n239, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_457_port);
   U16203 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1481_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2505_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n238);
   U16204 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_457_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_969_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1993_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n239);
   U16205 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n236, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n237, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_458_port);
   U16206 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1482_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2506_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n236);
   U16207 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_458_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_970_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1994_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n237);
   U16208 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n234, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n235, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_459_port);
   U16209 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1483_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2507_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n234);
   U16210 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_459_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_971_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1995_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n235);
   U16211 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n230, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n231, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_460_port);
   U16212 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1484_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2508_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n230);
   U16213 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_460_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_972_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1996_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n231);
   U16214 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n228, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n229, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_461_port);
   U16215 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1485_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2509_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n228);
   U16216 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_461_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_973_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1997_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n229);
   U16217 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n226, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n227, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_462_port);
   U16218 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1486_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2510_port, B2 => n3869, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n226);
   U16219 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_462_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_974_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1998_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n227);
   U16220 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n224, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n225, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_463_port);
   U16221 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1487_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2511_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n224);
   U16222 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_463_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_975_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_1999_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n225);
   U16223 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n222, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n223, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_464_port);
   U16224 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1488_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2512_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n222);
   U16225 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_464_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_976_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_2000_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n223);
   U16226 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n220, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n221, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_465_port);
   U16227 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1489_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2513_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n220);
   U16228 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_465_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_977_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_2001_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n221);
   U16229 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n218, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n219, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_466_port);
   U16230 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1490_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2514_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n218);
   U16231 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_466_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_978_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_2002_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n219);
   U16232 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n216, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n217, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_467_port);
   U16233 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1491_port, A2 
                           => n3237, B1 => 
                           DataPath_RF_bus_reg_dataout_2515_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n216);
   U16234 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_467_port, A2 
                           => n3081, B1 => DataPath_RF_bus_reg_dataout_979_port
                           , B2 => n3136, C1 => 
                           DataPath_RF_bus_reg_dataout_2003_port, C2 => n3182, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n217);
   U16235 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n214, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n215, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_468_port);
   U16236 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1492_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2516_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n214);
   U16237 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_468_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_980_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2004_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n215);
   U16238 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n212, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n213, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_469_port);
   U16239 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1493_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2517_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n212);
   U16240 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_469_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_981_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2005_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n213);
   U16241 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n208, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n209, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_470_port);
   U16242 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1494_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2518_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n208);
   U16243 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_470_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_982_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2006_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n209);
   U16244 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n206, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n207, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_471_port);
   U16245 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1495_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2519_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n206);
   U16246 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_471_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_983_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2007_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n207);
   U16247 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n204, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n205, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_472_port);
   U16248 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1496_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2520_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n204);
   U16249 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_472_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_984_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2008_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n205);
   U16250 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n202, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n203, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_473_port);
   U16251 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1497_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2521_port, B2 => n3870, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n202);
   U16252 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_473_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_985_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2009_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n203);
   U16253 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n200, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n201, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_474_port);
   U16254 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1498_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2522_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n200);
   U16255 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_474_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_986_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2010_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n201);
   U16256 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n196, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n197, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_476_port);
   U16257 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1500_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2524_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n196);
   U16258 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_476_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_988_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2012_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n197);
   U16259 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n194, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n195, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_477_port);
   U16260 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1501_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2525_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n194);
   U16261 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_477_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_989_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2013_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n195);
   U16262 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n192, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n193, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_478_port);
   U16263 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1502_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2526_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n192);
   U16264 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_478_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_990_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2014_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n193);
   U16265 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n190, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n191, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_479_port);
   U16266 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1503_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2527_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n190);
   U16267 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_479_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_991_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2015_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n191);
   U16268 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n198, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n199, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_475_port);
   U16269 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1499_port, A2 
                           => n3238, B1 => 
                           DataPath_RF_bus_reg_dataout_2523_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n198);
   U16270 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_475_port, A2 
                           => n3082, B1 => DataPath_RF_bus_reg_dataout_987_port
                           , B2 => n3137, C1 => 
                           DataPath_RF_bus_reg_dataout_2011_port, C2 => n3183, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n199);
   U16271 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n186, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n187, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_480_port);
   U16272 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1504_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2528_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n186);
   U16273 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_480_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_992_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2016_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n187);
   U16274 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n184, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n185, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_481_port);
   U16275 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1505_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2529_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n184);
   U16276 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_481_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_993_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2017_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n185);
   U16277 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n182, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n183, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_482_port);
   U16278 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1506_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2530_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n182);
   U16279 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_482_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_994_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2018_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n183);
   U16280 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n180, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n181, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_483_port);
   U16281 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1507_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2531_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n180);
   U16282 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_483_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_995_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2019_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n181);
   U16283 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n178, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n179, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_484_port);
   U16284 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1508_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2532_port, B2 => n3871, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n178);
   U16285 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_484_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_996_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2020_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n179);
   U16286 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n176, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n177, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_485_port);
   U16287 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1509_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2533_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n176);
   U16288 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_485_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_997_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2021_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n177);
   U16289 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n174, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n175, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_486_port);
   U16290 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1510_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2534_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n174);
   U16291 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_486_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_998_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2022_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n175);
   U16292 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n172, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n173, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_487_port);
   U16293 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1511_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2535_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n172);
   U16294 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_487_port, A2 
                           => n3083, B1 => DataPath_RF_bus_reg_dataout_999_port
                           , B2 => n3138, C1 => 
                           DataPath_RF_bus_reg_dataout_2023_port, C2 => n3184, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n173);
   U16295 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n170, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n171, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_488_port);
   U16296 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1512_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2536_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n170);
   U16297 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_488_port, A2 
                           => n3083, B1 => 
                           DataPath_RF_bus_reg_dataout_1000_port, B2 => n3138, 
                           C1 => DataPath_RF_bus_reg_dataout_2024_port, C2 => 
                           n3184, ZN => DataPath_RF_SELBLOCK_INLOC_n171);
   U16298 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n168, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n169, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_489_port);
   U16299 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1513_port, A2 
                           => n3239, B1 => 
                           DataPath_RF_bus_reg_dataout_2537_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n168);
   U16300 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_489_port, A2 
                           => n3083, B1 => 
                           DataPath_RF_bus_reg_dataout_1001_port, B2 => n3138, 
                           C1 => DataPath_RF_bus_reg_dataout_2025_port, C2 => 
                           n3184, ZN => DataPath_RF_SELBLOCK_INLOC_n169);
   U16301 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n164, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n165, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_490_port);
   U16302 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1514_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2538_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n164);
   U16303 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_490_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1002_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2026_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n165);
   U16304 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n162, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n163, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_491_port);
   U16305 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1515_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2539_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n162);
   U16306 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_491_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1003_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2027_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n163);
   U16307 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n160, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n161, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_492_port);
   U16308 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1516_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2540_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n160);
   U16309 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_492_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1004_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2028_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n161);
   U16310 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n158, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n159, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_493_port);
   U16311 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1517_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2541_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n158);
   U16312 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_493_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1005_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2029_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n159);
   U16313 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n156, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n157, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_494_port);
   U16314 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1518_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2542_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n156);
   U16315 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_494_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1006_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2030_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n157);
   U16316 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n154, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n155, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_495_port);
   U16317 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1519_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2543_port, B2 => n3872, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n154);
   U16318 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_495_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1007_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2031_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n155);
   U16319 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n152, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n153, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_496_port);
   U16320 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1520_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2544_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n152);
   U16321 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_496_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1008_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2032_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n153);
   U16322 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n150, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n151, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_497_port);
   U16323 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1521_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2545_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n150);
   U16324 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_497_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1009_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2033_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n151);
   U16325 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n148, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n149, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_498_port);
   U16326 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1522_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2546_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n148);
   U16327 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_498_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1010_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2034_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n149);
   U16328 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n146, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n147, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_499_port);
   U16329 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1523_port, A2 
                           => n3240, B1 => 
                           DataPath_RF_bus_reg_dataout_2547_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n146);
   U16330 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_499_port, A2 
                           => n3084, B1 => 
                           DataPath_RF_bus_reg_dataout_1011_port, B2 => n3139, 
                           C1 => DataPath_RF_bus_reg_dataout_2035_port, C2 => 
                           n3185, ZN => DataPath_RF_SELBLOCK_INLOC_n147);
   U16331 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n140, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n141, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_500_port);
   U16332 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1524_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2548_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n140);
   U16333 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_500_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1012_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2036_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n141);
   U16334 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n138, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n139, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_501_port);
   U16335 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1525_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2549_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n138);
   U16336 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_501_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1013_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2037_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n139);
   U16337 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n136, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n137, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_502_port);
   U16338 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1526_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2550_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n136);
   U16339 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_502_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1014_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2038_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n137);
   U16340 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n134, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n135, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_503_port);
   U16341 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1527_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2551_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n134);
   U16342 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_503_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1015_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2039_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n135);
   U16343 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n132, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n133, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_504_port);
   U16344 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1528_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2552_port, B2 => n3873, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n132);
   U16345 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_504_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1016_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2040_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n133);
   U16346 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n130, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n131, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_505_port);
   U16347 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1529_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2553_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n130);
   U16348 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_505_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1017_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2041_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n131);
   U16349 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n128, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n129, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_506_port);
   U16350 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1530_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2554_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n128);
   U16351 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_506_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1018_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2042_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n129);
   U16352 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n126, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n127, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_507_port);
   U16353 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1531_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2555_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n126);
   U16354 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_507_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1019_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2043_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n127);
   U16355 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n124, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n125, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_508_port);
   U16356 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1532_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2556_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n124);
   U16357 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_508_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1020_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2044_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n125);
   U16358 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n122, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n123, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_509_port);
   U16359 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1533_port, A2 
                           => n3241, B1 => 
                           DataPath_RF_bus_reg_dataout_2557_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n122);
   U16360 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_509_port, A2 
                           => n3085, B1 => 
                           DataPath_RF_bus_reg_dataout_1021_port, B2 => n3140, 
                           C1 => DataPath_RF_bus_reg_dataout_2045_port, C2 => 
                           n3186, ZN => DataPath_RF_SELBLOCK_INLOC_n123);
   U16361 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n118, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n119, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_510_port);
   U16362 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1534_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2558_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n118);
   U16363 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_510_port, A2 
                           => n3086, B1 => 
                           DataPath_RF_bus_reg_dataout_1022_port, B2 => n3141, 
                           C1 => DataPath_RF_bus_reg_dataout_2046_port, C2 => 
                           n3187, ZN => DataPath_RF_SELBLOCK_INLOC_n119);
   U16364 : NAND2_X1 port map( A1 => DataPath_RF_SELBLOCK_INLOC_n116, A2 => 
                           DataPath_RF_SELBLOCK_INLOC_n117, ZN => 
                           DataPath_RF_bus_sel_savedwin_data_511_port);
   U16365 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1535_port, A2 
                           => n3242, B1 => 
                           DataPath_RF_bus_reg_dataout_2559_port, B2 => n3874, 
                           ZN => DataPath_RF_SELBLOCK_INLOC_n116);
   U16366 : AOI222_X1 port map( A1 => DataPath_RF_bus_reg_dataout_511_port, A2 
                           => n3086, B1 => 
                           DataPath_RF_bus_reg_dataout_1023_port, B2 => n3141, 
                           C1 => DataPath_RF_bus_reg_dataout_2047_port, C2 => 
                           n3187, ZN => DataPath_RF_SELBLOCK_INLOC_n117);
   U16367 : INV_X1 port map( A => DRAMRF_DATA_IN(31), ZN => n11447);
   U16368 : INV_X1 port map( A => DRAMRF_DATA_IN(30), ZN => n11448);
   U16369 : INV_X1 port map( A => DRAMRF_DATA_IN(29), ZN => n11449);
   U16370 : INV_X1 port map( A => DRAMRF_DATA_IN(28), ZN => n11450);
   U16371 : INV_X1 port map( A => DRAMRF_DATA_IN(27), ZN => n11451);
   U16372 : INV_X1 port map( A => DRAMRF_DATA_IN(26), ZN => n11452);
   U16373 : INV_X1 port map( A => DRAMRF_DATA_IN(25), ZN => n11453);
   U16374 : INV_X1 port map( A => DRAMRF_DATA_IN(24), ZN => n11454);
   U16375 : INV_X1 port map( A => DRAMRF_DATA_IN(23), ZN => n11455);
   U16376 : INV_X1 port map( A => DRAMRF_DATA_IN(22), ZN => n11456);
   U16377 : INV_X1 port map( A => DRAMRF_DATA_IN(21), ZN => n11457);
   U16378 : INV_X1 port map( A => DRAMRF_DATA_IN(20), ZN => n11458);
   U16379 : INV_X1 port map( A => DRAMRF_DATA_IN(19), ZN => n11459);
   U16380 : INV_X1 port map( A => DRAMRF_DATA_IN(18), ZN => n11460);
   U16381 : INV_X1 port map( A => DRAMRF_DATA_IN(17), ZN => n11461);
   U16382 : INV_X1 port map( A => DRAMRF_DATA_IN(16), ZN => n11462);
   U16383 : INV_X1 port map( A => DRAMRF_DATA_IN(15), ZN => n11463);
   U16384 : INV_X1 port map( A => DRAMRF_DATA_IN(14), ZN => n11464);
   U16385 : INV_X1 port map( A => DRAMRF_DATA_IN(13), ZN => n11465);
   U16386 : INV_X1 port map( A => DRAMRF_DATA_IN(12), ZN => n11466);
   U16387 : INV_X1 port map( A => DRAMRF_DATA_IN(11), ZN => n11467);
   U16388 : INV_X1 port map( A => DRAMRF_DATA_IN(10), ZN => n11468);
   U16389 : INV_X1 port map( A => DRAMRF_DATA_IN(9), ZN => n11469);
   U16390 : INV_X1 port map( A => DRAMRF_DATA_IN(8), ZN => n11470);
   U16391 : INV_X1 port map( A => DRAMRF_DATA_IN(7), ZN => n11471);
   U16392 : INV_X1 port map( A => DRAMRF_DATA_IN(6), ZN => n11472);
   U16393 : INV_X1 port map( A => DRAMRF_DATA_IN(5), ZN => n11473);
   U16394 : INV_X1 port map( A => DRAMRF_DATA_IN(4), ZN => n11474);
   U16395 : INV_X1 port map( A => DRAMRF_DATA_IN(3), ZN => n11475);
   U16396 : INV_X1 port map( A => DRAMRF_DATA_IN(2), ZN => n11476);
   U16397 : INV_X1 port map( A => DRAMRF_DATA_IN(1), ZN => n11477);
   U16398 : INV_X1 port map( A => DRAMRF_DATA_IN(0), ZN => n11478);
   U16399 : BUF_X1 port map( A => DataPath_RF_c_swin_4_port, Z => n3845);
   U16400 : BUF_X1 port map( A => DRAMRF_READY, Z => n4153);
   U16401 : BUF_X1 port map( A => DRAMRF_READY, Z => n4154);
   U16402 : BUF_X1 port map( A => DRAMRF_READY, Z => n4152);
   U16403 : BUF_X1 port map( A => RST, Z => n4254);
   U16404 : BUF_X1 port map( A => RST, Z => n4255);
   U16405 : BUF_X1 port map( A => DataPath_RF_c_swin_4_port, Z => n3846);
   U16406 : BUF_X1 port map( A => RST, Z => n4256);
   U16407 : AND2_X1 port map( A1 => 
                           DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_0_port, A2 =>
                           DATA_SIZE_1_port, ZN => DRAM_ADDRESS_0_port);
   U16408 : INV_X1 port map( A => DataPath_MEM_ADDR_MASK_n2, ZN => 
                           DRAM_ADDRESS_1_port);
   U16409 : OAI21_X1 port map( B1 => DATA_SIZE_1_port, B2 => DATA_SIZE_0_port, 
                           A => DataPath_i_REG_ALU_OUT_ADDRESS_DATAMEM_1_port, 
                           ZN => DataPath_MEM_ADDR_MASK_n2);
   U16410 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_3_port, A2 => n2488, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_3_port, B2 => 
                           n2489, ZN => n14264);
   OPCODE_5_port <= '0';
   OPCODE_3_port <= '0';
   OPCODE_1_port <= '0';
   RS1(4) <= '0';
   IRO_25_port <= '0';
   RS1(3) <= '0';
   IRO_24_port <= '0';
   RS1(2) <= '0';
   IRO_23_port <= '0';
   RS1(1) <= '0';
   IRO_22_port <= '0';
   RS1(0) <= '0';
   IRO_21_port <= '0';
   IRO_20_port <= '0';
   IRO_19_port <= '0';
   IRO_18_port <= '0';
   IRO_17_port <= '0';
   IRO_16_port <= '0';
   IRO_15_port <= '0';
   IRO_14_port <= '0';
   IRO_13_port <= '0';
   IRO_12_port <= '0';
   IRO_11_port <= '0';
   IRO_10_port <= '0';
   IRO_9_port <= '0';
   IRO_8_port <= '0';
   IRO_7_port <= '0';
   IRO_6_port <= '0';
   IRO_5_port <= '0';
   IRO_4_port <= '0';
   IRO_3_port <= '0';
   IRO_2_port <= '0';
   IRO_1_port <= '0';
   IRO_0_port <= '0';
   OPCODE_4_port <= '1';
   OPCODE_2_port <= '1';
   OPCODE_0_port <= '1';
   U16448 : AOI22_X1 port map( A1 => n4830, A2 => n4952, B1 => n4912, B2 => 
                           n1427, ZN => n4915);
   U16449 : XNOR2_X1 port map( A => n5152, B => n1197, ZN => n5161);
   U16450 : INV_X1 port map( A => n5187, ZN => n4830);
   U16451 : MUX2_X2 port map( A => n5591, B => n5590, S => n2244, Z => n5987);
   U16452 : XNOR2_X1 port map( A => n5128, B => n448, ZN => n5133);
   U16453 : XNOR2_X1 port map( A => n4711, B => n4712, ZN => n4713);
   U16454 : INV_X1 port map( A => n7688, ZN => n2235);
   U16455 : XNOR2_X1 port map( A => n5158, B => n5159, ZN => n5160);
   U16456 : CLKBUF_X1 port map( A => n17194, Z => n2132);
   U16457 : NAND2_X1 port map( A1 => i_S2, A2 => n1745, ZN => n4449);
   U16458 : INV_X1 port map( A => n2144, ZN => n2133);
   U16459 : BUF_X1 port map( A => n2150, Z => n2143);
   U16460 : CLKBUF_X1 port map( A => n6858, Z => n2135);
   U16461 : BUF_X1 port map( A => n2136, Z => n2137);
   U16462 : CLKBUF_X1 port map( A => n8023, Z => n2134);
   U16463 : AOI21_X1 port map( B1 => n848, B2 => n5123, A => n5121, ZN => n5126
                           );
   U16464 : AOI22_X1 port map( A1 => n1266, A2 => n2488, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_0_port, B2 => n2489, 
                           ZN => n14259);
   U16465 : NAND2_X1 port map( A1 => n5147, A2 => n5148, ZN => n5150);
   U16466 : INV_X2 port map( A => n2146, ZN => n2147);
   U16467 : XNOR2_X1 port map( A => n998, B => n5376, ZN => n5378);
   U16468 : NAND2_X1 port map( A1 => n4893, A2 => n4894, ZN => n4895);
   U16469 : NAND2_X1 port map( A1 => n17174, A2 => n5484, ZN => n5487);
   U16470 : NAND2_X1 port map( A1 => n1189, A2 => n5146, ZN => n5151);
   U16471 : XNOR2_X1 port map( A => n5256, B => n5756, ZN => n5258);
   U16472 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_1_port, A2 => n2488, 
                           B1 => DataPath_i_REG_ME_DATA_DATAMEM_1_port, B2 => 
                           n2489, ZN => n14262);
   U16473 : OAI221_X1 port map( B1 => DataPath_i_PIPLIN_B_0_port, B2 => i_S2, 
                           C1 => n4450, C2 => n4451, A => n4449, ZN => n4547);
   U16474 : NAND2_X1 port map( A1 => n7747, A2 => n1208, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n192);
   U16475 : NAND2_X1 port map( A1 => n5660, A2 => n5659, ZN => n5661);
   U16476 : OAI22_X1 port map( A1 => n1716, A2 => i_S2, B1 => n1745, B2 => 
                           CU_I_n107, ZN => n7318);
   U16477 : INV_X1 port map( A => n4142, ZN => n2150);
   U16478 : INV_X1 port map( A => n4142, ZN => n2151);
   U16479 : OAI33_X1 port map( A1 => n4594, A2 => n4882, A3 => n804, B1 => 
                           n4881, B2 => n4879, B3 => n4880, ZN => n2153);
   U16480 : MUX2_X1 port map( A => DataPath_i_PIPLIN_B_3_port, B => 
                           DataPath_i_PIPLIN_IN2_3_port, S => i_S2, Z => n2155)
                           ;
   U16481 : INV_X1 port map( A => n669, ZN => n2157);
   U16482 : XNOR2_X1 port map( A => n1262, B => n662, ZN => n5961);
   U16483 : XOR2_X1 port map( A => n740, B => n6312, Z => n2158);
   U16484 : XNOR2_X1 port map( A => n6172, B => n2160, ZN => n6173);
   U16485 : XNOR2_X1 port map( A => n1236, B => n5345, ZN => n5347);
   U16486 : NAND2_X1 port map( A1 => n6128, A2 => n6127, ZN => n6017);
   U16487 : OR2_X1 port map( A1 => n2162, A2 => n5948, ZN => n5940);
   U16488 : XNOR2_X1 port map( A => n5684, B => n728, ZN => n2164);
   U16489 : NOR2_X1 port map( A1 => n1577, A2 => n6183, ZN => n2166);
   U16490 : INV_X1 port map( A => n2167, ZN => n2191);
   U16491 : XNOR2_X1 port map( A => n5248, B => n5226, ZN => n5228);
   U16492 : XNOR2_X1 port map( A => n4691, B => n5218, ZN => n4693);
   U16493 : XNOR2_X1 port map( A => n17173, B => n4780, ZN => n4782);
   U16494 : XNOR2_X1 port map( A => n4787, B => n4785, ZN => n4789);
   U16495 : AOI21_X1 port map( B1 => n5488, B2 => n5487, A => n5486, ZN => 
                           n5492);
   U16496 : NOR2_X1 port map( A1 => n1785, A2 => n1011, ZN => n5488);
   U16497 : NAND2_X1 port map( A1 => n5183, A2 => n5184, ZN => n4913);
   U16498 : OAI22_X1 port map( A1 => n1213, A2 => n6352, B1 => n6440, B2 => 
                           n950, ZN => n6435);
   U16499 : NOR2_X1 port map( A1 => n6439, A2 => n6346, ZN => n6352);
   U16500 : XNOR2_X1 port map( A => n801, B => n5382, ZN => n5384);
   U16501 : MUX2_X2 port map( A => n5636, B => n5635, S => n2244, Z => n5908);
   U16502 : INV_X1 port map( A => n2169, ZN => n6002);
   U16503 : MUX2_X2 port map( A => n5104, B => n5103, S => n2248, Z => n5436);
   U16504 : XNOR2_X1 port map( A => n5131, B => n1356, ZN => n5132);
   U16505 : NAND2_X1 port map( A1 => n1253, A2 => n5130, ZN => n5131);
   U16506 : XNOR2_X1 port map( A => n5952, B => n5951, ZN => n2170);
   U16507 : XNOR2_X1 port map( A => n5492, B => n5491, ZN => n5493);
   U16508 : NAND2_X1 port map( A1 => n5481, A2 => n5480, ZN => n5482);
   U16509 : NOR2_X1 port map( A1 => n6205, A2 => n6204, ZN => n6210);
   U16510 : NAND2_X1 port map( A1 => n6165, A2 => n6152, ZN => n6156);
   U16511 : XNOR2_X1 port map( A => n5937, B => n5938, ZN => n5947);
   U16512 : OAI211_X1 port map( C1 => n1485, C2 => n1848, A => n6125, B => 
                           n6124, ZN => n6014);
   U16513 : NAND2_X1 port map( A1 => n1116, A2 => n5949, ZN => n5935);
   U16514 : XNOR2_X1 port map( A => n6434, B => n994, ZN => n2173);
   U16515 : XNOR2_X1 port map( A => n6437, B => n994, ZN => n2174);
   U16516 : XNOR2_X1 port map( A => n842, B => n2157, ZN => n6205);
   U16517 : INV_X1 port map( A => n215, ZN => n6194);
   U16518 : XNOR2_X1 port map( A => n6781, B => n6033, ZN => n6035);
   U16519 : XNOR2_X1 port map( A => n5767, B => n1282, ZN => n5268);
   U16520 : XNOR2_X1 port map( A => n4698, B => n4696, ZN => n4700);
   U16521 : XNOR2_X1 port map( A => n4703, B => n4705, ZN => n4707);
   U16522 : XNOR2_X1 port map( A => n4718, B => n4716, ZN => n4720);
   U16523 : XNOR2_X1 port map( A => n4725, B => n4723, ZN => n4727);
   U16524 : XNOR2_X1 port map( A => n4773, B => n4772, ZN => n4775);
   U16525 : XNOR2_X1 port map( A => n4792, B => n4794, ZN => n4796);
   U16526 : XNOR2_X1 port map( A => n708, B => n6555, ZN => n6554);
   U16527 : NAND2_X1 port map( A1 => n5301, A2 => n5300, ZN => n5343);
   U16528 : XNOR2_X1 port map( A => n5067, B => n5069, ZN => n5071);
   U16529 : OAI22_X1 port map( A1 => n1117, A2 => n602, B1 => n747, B2 => n6221
                           , ZN => n6245);
   U16530 : OAI211_X1 port map( C1 => n1608, C2 => n1794, A => n5913, B => 
                           n5969, ZN => n5741);
   U16532 : OAI22_X1 port map( A1 => n6692, A2 => n993, B1 => n7010, B2 => 
                           n7012, ZN => n7028);
   U16533 : INV_X1 port map( A => n6329, ZN => n6209);
   U16534 : XNOR2_X1 port map( A => n5655, B => n5656, ZN => n5663);
   U16535 : XNOR2_X1 port map( A => n5047, B => n5049, ZN => n5051);
   U16536 : OAI22_X1 port map( A1 => n5298, A2 => n5299, B1 => n5350, B2 => 
                           n1837, ZN => n5301);
   U16537 : OAI22_X1 port map( A1 => n6225, A2 => n6224, B1 => n6222, B2 => 
                           n6223, ZN => n6238);
   U16538 : INV_X1 port map( A => n6245, ZN => n6224);
   U16539 : NAND2_X1 port map( A1 => n939, A2 => n7576, ZN => n7072);
   U16540 : OAI211_X1 port map( C1 => n1433, C2 => n5808, A => n5972, B => 
                           n5741, ZN => n5903);
   U16541 : NAND2_X1 port map( A1 => n7070, A2 => n7578, ZN => n7071);
   U16542 : XNOR2_X1 port map( A => n551, B => n5943, ZN => n5944);
   U16543 : XNOR2_X1 port map( A => n1753, B => n5936, ZN => n5937);
   U16544 : NAND2_X1 port map( A1 => n7496, A2 => n7547, ZN => n7501);
   U16545 : OAI22_X1 port map( A1 => n7042, A2 => n1305, B1 => n7041, B2 => 
                           n7641, ZN => n7058);
   U16546 : NOR2_X1 port map( A1 => n1660, A2 => n7032, ZN => n6692);
   U16547 : INV_X1 port map( A => n840, ZN => n6351);
   U16548 : AOI21_X1 port map( B1 => n5126, B2 => n5125, A => n5124, ZN => 
                           n5128);
   U16549 : AOI22_X1 port map( A1 => n7494, A2 => n1292, B1 => n7493, B2 => 
                           n7492, ZN => n7513);
   U16550 : NOR2_X1 port map( A1 => n7492, A2 => n7498, ZN => n7494);
   U16551 : NOR2_X1 port map( A1 => n756, A2 => n7039, ZN => n7042);
   U16552 : XNOR2_X1 port map( A => n6687, B => n582, ZN => n6689);
   U16553 : XNOR2_X1 port map( A => n17213, B => n1385, ZN => n6639);
   U16554 : XNOR2_X1 port map( A => n6443, B => n1490, ZN => n6445);
   U16555 : XNOR2_X1 port map( A => n6179, B => n911, ZN => n6181);
   U16556 : INV_X2 port map( A => n2203, ZN => n2200);
   U16557 : INV_X2 port map( A => n2228, ZN => n2227);
   U16558 : INV_X2 port map( A => n2241, ZN => n2240);
   U16559 : BUF_X4 port map( A => n7295, Z => n2182);
   U16560 : XOR2_X2 port map( A => n8232, B => n2265, Z => n7284);
   U16561 : OAI221_X4 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n600, B2 => 
                           n7987, C1 => n7986, C2 => n8089, A => n7985, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n146);
   U16562 : INV_X1 port map( A => n1873, ZN => n2190);
   U16563 : INV_X1 port map( A => n548, ZN => n2192);
   U16565 : INV_X1 port map( A => n1208, ZN => n2194);
   U16566 : INV_X1 port map( A => n703, ZN => n2195);
   U16567 : INV_X1 port map( A => n1374, ZN => n2198);
   U16568 : INV_X1 port map( A => n2203, ZN => n2201);
   U16569 : INV_X1 port map( A => n7249, ZN => n2202);
   U16570 : INV_X1 port map( A => n7249, ZN => n2203);
   U16571 : INV_X1 port map( A => n252, ZN => n2206);
   U16572 : INV_X1 port map( A => n2212, ZN => n2210);
   U16573 : INV_X1 port map( A => n7259, ZN => n2211);
   U16574 : INV_X1 port map( A => n7259, ZN => n2212);
   U16575 : CLKBUF_X1 port map( A => n7312, Z => n2223);
   U16576 : INV_X1 port map( A => n2229, ZN => n2231);
   U16577 : INV_X1 port map( A => n7658, ZN => n2232);
   U16578 : INV_X1 port map( A => n7658, ZN => n2233);
   U16580 : INV_X1 port map( A => n1542, ZN => n2241);
   U16581 : CLKBUF_X1 port map( A => n3044, Z => n3090);
   U16582 : CLKBUF_X1 port map( A => n3099, Z => n3145);
   U16583 : CLKBUF_X1 port map( A => n3192, Z => n3191);
   U16584 : CLKBUF_X1 port map( A => n3247, Z => n3246);
   U16585 : INV_X1 port map( A => n3278, ZN => n3270);
   U16586 : INV_X1 port map( A => n3370, ZN => n3295);
   U16587 : INV_X1 port map( A => n3371, ZN => n3299);
   U16588 : INV_X1 port map( A => n3482, ZN => n3409);
   U16589 : INV_X1 port map( A => n3483, ZN => n3411);
   U16590 : INV_X1 port map( A => n3594, ZN => n3521);
   U16591 : INV_X1 port map( A => n3595, ZN => n3523);
   U16592 : INV_X1 port map( A => n3706, ZN => n3632);
   U16593 : INV_X1 port map( A => n3707, ZN => n3635);
   U16594 : INV_X1 port map( A => n3819, ZN => n3746);
   U16595 : CLKBUF_X1 port map( A => n3891, Z => n3890);
   U16596 : INV_X1 port map( A => n2148, ZN => n4142);
   U16597 : INV_X1 port map( A => n4220, ZN => n4257);
   U16598 : NAND2_X1 port map( A1 => n1302, A2 => DataPath_i_PIPLIN_B_1_port, 
                           ZN => n4444);
   U16599 : NAND2_X1 port map( A1 => i_S2, A2 => DataPath_i_PIPLIN_IN2_1_port, 
                           ZN => n4443);
   U16600 : XOR2_X1 port map( A => n2259, B => n4129, Z => n4271);
   U16601 : XOR2_X1 port map( A => n17175, B => n4130, Z => n4270);
   U16602 : MUX2_X1 port map( A => n4269, B => n4268, S => i_S1, Z => n8091);
   U16603 : INV_X1 port map( A => n8091, ZN => n8277);
   U16604 : NAND2_X1 port map( A1 => n4270, A2 => n2154, ZN => n4284);
   U16605 : NAND2_X1 port map( A1 => n4271, A2 => n2146, ZN => n4285);
   U16606 : OAI21_X1 port map( B1 => n1797, B2 => n370, A => n4285, ZN => n4279
                           );
   U16607 : NAND2_X1 port map( A1 => n259, A2 => n7196, ZN => n4428);
   U16608 : OAI21_X1 port map( B1 => n259, B2 => n7196, A => n4428, ZN => n4274
                           );
   U16609 : MUX2_X1 port map( A => n4273, B => n4272, S => i_S1, Z => n7658);
   U16610 : XOR2_X1 port map( A => n4274, B => n2231, Z => n4276);
   U16611 : NAND2_X1 port map( A1 => n4279, A2 => n4276, ZN => n4283);
   U16612 : NAND2_X1 port map( A1 => n4274, A2 => n2231, ZN => n4290);
   U16613 : NAND2_X1 port map( A1 => n4283, A2 => n4290, ZN => n4275);
   U16614 : XOR2_X1 port map( A => n818, B => n4130, Z => n4292);
   U16615 : XOR2_X1 port map( A => n4292, B => n2228, Z => n4291);
   U16616 : INV_X1 port map( A => n4291, ZN => n4287);
   U16617 : XOR2_X1 port map( A => n4275, B => n4287, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_3_port
                           );
   U16618 : INV_X1 port map( A => n4276, ZN => n4282);
   U16619 : OAI21_X1 port map( B1 => n1797, B2 => n4284, A => n4285, ZN => 
                           n4277);
   U16620 : INV_X1 port map( A => n4277, ZN => n4281);
   U16621 : OAI21_X1 port map( B1 => n4282, B2 => n4281, A => n4290, ZN => 
                           n4278);
   U16622 : XOR2_X1 port map( A => n4278, B => n4287, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_3_port
                           );
   U16623 : INV_X1 port map( A => n4279, ZN => n4280);
   U16624 : XOR2_X1 port map( A => n4282, B => n4280, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_2_port
                           );
   U16625 : XOR2_X1 port map( A => n4282, B => n4281, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_2_port
                           );
   U16626 : XOR2_X1 port map( A => n1797, B => n370, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_1_1_port
                           );
   U16627 : XOR2_X1 port map( A => n4284, B => n1797, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_0_sum_mux21_0_1_port
                           );
   U16628 : INV_X1 port map( A => n4283, ZN => n4288);
   U16629 : NAND3_X1 port map( A1 => n4285, A2 => n4135, A3 => n4284, ZN => 
                           n4286);
   U16630 : NAND3_X1 port map( A1 => n4288, A2 => n4287, A3 => n4286, ZN => 
                           n4289);
   U16631 : OAI221_X1 port map( B1 => n2227, B2 => n4292, C1 => n4291, C2 => 
                           n4290, A => n4289, ZN => n11516);
   U16632 : MUX2_X1 port map( A => n263, B => n323, S => n527, Z => n4985);
   U16633 : XOR2_X1 port map( A => n4985, B => n4129, Z => n4299);
   U16634 : XOR2_X1 port map( A => n4299, B => n1933, Z => n4308);
   U16635 : XOR2_X1 port map( A => n6890, B => n4129, Z => n4296);
   U16636 : XOR2_X1 port map( A => n4296, B => n788, Z => n4376);
   U16637 : MUX2_X1 port map( A => n4293, B => n324, S => n2152, Z => n7109);
   U16638 : XOR2_X1 port map( A => n7109, B => n4130, Z => n4294);
   U16639 : XOR2_X1 port map( A => n4294, B => n2241, Z => n8186);
   U16640 : INV_X1 port map( A => n4294, ZN => n4295);
   U16641 : NAND2_X1 port map( A1 => n4295, A2 => n2241, ZN => n4311);
   U16642 : NAND2_X1 port map( A1 => n8186, A2 => n4311, ZN => n4310);
   U16643 : INV_X1 port map( A => n4310, ZN => n4298);
   U16644 : INV_X1 port map( A => n4296, ZN => n4297);
   U16645 : NAND2_X1 port map( A1 => n4297, A2 => n788, ZN => n4305);
   U16646 : OAI21_X1 port map( B1 => n4376, B2 => n4298, A => n4305, ZN => 
                           n4309);
   U16647 : INV_X1 port map( A => n4309, ZN => n4301);
   U16648 : INV_X1 port map( A => n4299, ZN => n4300);
   U16649 : NAND2_X1 port map( A1 => n4300, A2 => n1933, ZN => n4378);
   U16650 : OAI21_X1 port map( B1 => n4308, B2 => n4301, A => n4378, ZN => 
                           n4304);
   U16651 : MUX2_X1 port map( A => n4302, B => n254, S => n2152, Z => n6920);
   U16652 : XOR2_X1 port map( A => n6920, B => n4129, Z => n4377);
   U16653 : XOR2_X1 port map( A => n4377, B => n1520, Z => n4379);
   U16654 : INV_X1 port map( A => n4379, ZN => n4374);
   U16655 : XOR2_X1 port map( A => n4304, B => n4374, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_3_port
                           );
   U16656 : OAI21_X1 port map( B1 => n4376, B2 => n4311, A => n4305, ZN => 
                           n11535);
   U16657 : INV_X1 port map( A => n11535, ZN => n4306);
   U16658 : OAI21_X1 port map( B1 => n4308, B2 => n4306, A => n4378, ZN => 
                           n4307);
   U16659 : XOR2_X1 port map( A => n4307, B => n4374, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_3_port
                           );
   U16660 : INV_X1 port map( A => n11516, ZN => n12926);
   U16661 : INV_X1 port map( A => n4308, ZN => n4375);
   U16662 : XOR2_X1 port map( A => n4309, B => n4375, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_2_port
                           );
   U16663 : XOR2_X1 port map( A => n11535, B => n4375, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_2_port
                           );
   U16664 : INV_X1 port map( A => n4376, ZN => n4313);
   U16665 : XOR2_X1 port map( A => n4310, B => n4313, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_1_1_port
                           );
   U16666 : INV_X1 port map( A => n4311, ZN => n4312);
   U16667 : XOR2_X1 port map( A => n4313, B => n4312, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_1_sum_mux21_0_1_port
                           );
   U16668 : INV_X1 port map( A => n12927, ZN => n11511);
   U16669 : MUX2_X1 port map( A => n272, B => n325, S => n525, Z => n8270);
   U16670 : XOR2_X1 port map( A => n8270, B => n4129, Z => n4321);
   U16671 : MUX2_X1 port map( A => n4314, B => n326, S => n2148, Z => n7259);
   U16672 : XOR2_X1 port map( A => n4321, B => n2211, Z => n4328);
   U16673 : MUX2_X1 port map( A => n257, B => n261, S => n524, Z => n6912);
   U16674 : XOR2_X1 port map( A => n6912, B => n4130, Z => n4318);
   U16675 : XOR2_X1 port map( A => n4318, B => n797, Z => n4382);
   U16676 : MUX2_X1 port map( A => n264, B => n327, S => n526, Z => n8143);
   U16677 : XOR2_X1 port map( A => n8143, B => n4129, Z => n4316);
   U16678 : MUX2_X1 port map( A => n4315, B => n328, S => i_S1, Z => n7249);
   U16679 : XOR2_X1 port map( A => n4316, B => n2202, Z => n8149);
   U16680 : INV_X1 port map( A => n4316, ZN => n4317);
   U16681 : NAND2_X1 port map( A1 => n4317, A2 => n2202, ZN => n4331);
   U16682 : NAND2_X1 port map( A1 => n8149, A2 => n4331, ZN => n4330);
   U16683 : INV_X1 port map( A => n4330, ZN => n4320);
   U16684 : INV_X1 port map( A => n4318, ZN => n4319);
   U16685 : NAND2_X1 port map( A1 => n4319, A2 => n797, ZN => n4325);
   U16686 : OAI21_X1 port map( B1 => n4382, B2 => n4320, A => n4325, ZN => 
                           n4329);
   U16687 : INV_X1 port map( A => n4329, ZN => n4323);
   U16688 : INV_X1 port map( A => n4321, ZN => n4322);
   U16689 : NAND2_X1 port map( A1 => n4322, A2 => n2212, ZN => n4384);
   U16690 : OAI21_X1 port map( B1 => n4328, B2 => n4323, A => n4384, ZN => 
                           n4324);
   U16691 : XOR2_X1 port map( A => n6776, B => n4130, Z => n4383);
   U16692 : XOR2_X1 port map( A => n4383, B => n2207, Z => n4385);
   U16693 : INV_X1 port map( A => n4385, ZN => n4380);
   U16694 : XOR2_X1 port map( A => n4324, B => n4380, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_3_port
                           );
   U16695 : OAI21_X1 port map( B1 => n4382, B2 => n4331, A => n4325, ZN => 
                           n11537);
   U16696 : INV_X1 port map( A => n11537, ZN => n4326);
   U16697 : OAI21_X1 port map( B1 => n4328, B2 => n4326, A => n4384, ZN => 
                           n4327);
   U16698 : XOR2_X1 port map( A => n4327, B => n4380, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_3_port
                           );
   U16699 : INV_X1 port map( A => n4328, ZN => n4381);
   U16700 : XOR2_X1 port map( A => n4329, B => n4381, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_2_port
                           );
   U16701 : XOR2_X1 port map( A => n11537, B => n4381, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_2_port
                           );
   U16702 : INV_X1 port map( A => n4382, ZN => n4333);
   U16703 : XOR2_X1 port map( A => n4330, B => n4333, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_1_1_port
                           );
   U16704 : INV_X1 port map( A => n4331, ZN => n4332);
   U16705 : XOR2_X1 port map( A => n4333, B => n4332, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_2_sum_mux21_0_1_port
                           );
   U16706 : INV_X1 port map( A => n12928, ZN => n11506);
   U16707 : MUX2_X1 port map( A => n273, B => n351, S => n525, Z => n8232);
   U16708 : XOR2_X1 port map( A => n8232, B => n4130, Z => n4340);
   U16709 : MUX2_X1 port map( A => n4334, B => n329, S => n2150, Z => n7275);
   U16710 : INV_X1 port map( A => n7275, ZN => n8234);
   U16711 : XOR2_X1 port map( A => n4340, B => n8234, Z => n4348);
   U16712 : XOR2_X1 port map( A => n6967, B => n4130, Z => n4337);
   U16713 : XOR2_X1 port map( A => n4337, B => n1935, Z => n4388);
   U16714 : MUX2_X1 port map( A => n274, B => n352, S => n527, Z => n8250);
   U16715 : XOR2_X1 port map( A => n8250, B => n4130, Z => n4335);
   U16716 : XOR2_X1 port map( A => n4335, B => n1934, Z => n8256);
   U16717 : INV_X1 port map( A => n4335, ZN => n4336);
   U16718 : NAND2_X1 port map( A1 => n4336, A2 => n1934, ZN => n4351);
   U16719 : NAND2_X1 port map( A1 => n8256, A2 => n4351, ZN => n4350);
   U16720 : INV_X1 port map( A => n4350, ZN => n4339);
   U16721 : INV_X1 port map( A => n4337, ZN => n4338);
   U16722 : NAND2_X1 port map( A1 => n4338, A2 => n1935, ZN => n4345);
   U16723 : OAI21_X1 port map( B1 => n4388, B2 => n4339, A => n4345, ZN => 
                           n4349);
   U16724 : INV_X1 port map( A => n4349, ZN => n4342);
   U16725 : INV_X1 port map( A => n4340, ZN => n4341);
   U16726 : NAND2_X1 port map( A1 => n4341, A2 => n8234, ZN => n4390);
   U16727 : OAI21_X1 port map( B1 => n4348, B2 => n4342, A => n4390, ZN => 
                           n4344);
   U16728 : MUX2_X1 port map( A => n275, B => n353, S => n526, Z => n6839);
   U16729 : XOR2_X1 port map( A => n6839, B => n4130, Z => n4389);
   U16730 : MUX2_X1 port map( A => n4343, B => n330, S => n2143, Z => n7273);
   U16731 : INV_X1 port map( A => n7273, ZN => n8223);
   U16732 : XOR2_X1 port map( A => n4389, B => n8223, Z => n4391);
   U16733 : INV_X1 port map( A => n4391, ZN => n4386);
   U16734 : XOR2_X1 port map( A => n4344, B => n4386, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_3_port
                           );
   U16735 : OAI21_X1 port map( B1 => n4388, B2 => n4351, A => n4345, ZN => 
                           n11521);
   U16736 : INV_X1 port map( A => n11521, ZN => n4346);
   U16737 : OAI21_X1 port map( B1 => n4348, B2 => n4346, A => n4390, ZN => 
                           n4347);
   U16738 : XOR2_X1 port map( A => n4347, B => n4386, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_3_port
                           );
   U16739 : INV_X1 port map( A => n4348, ZN => n4387);
   U16740 : XOR2_X1 port map( A => n4349, B => n4387, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_2_port
                           );
   U16741 : XOR2_X1 port map( A => n11521, B => n4387, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_2_port
                           );
   U16742 : INV_X1 port map( A => n4388, ZN => n4353);
   U16743 : XOR2_X1 port map( A => n4350, B => n4353, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_1_1_port
                           );
   U16744 : INV_X1 port map( A => n4351, ZN => n4352);
   U16745 : XOR2_X1 port map( A => n4353, B => n4352, Z => 
                           DataPath_ALUhw_ADDER_SUMGEM_csb_3_sum_mux21_0_1_port
                           );
   U16746 : MUX2_X1 port map( A => n4355, B => n4354, S => n527, Z => n4436);
   U16747 : XOR2_X1 port map( A => n4436, B => n4130, Z => n4362);
   U16748 : MUX2_X1 port map( A => n4356, B => n354, S => n2145, Z => n7311);
   U16749 : INV_X1 port map( A => n7311, ZN => n7709);
   U16750 : XOR2_X1 port map( A => n4362, B => n7709, Z => n7637);
   U16751 : INV_X1 port map( A => n7637, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_26_port);
   U16752 : MUX2_X1 port map( A => n4358, B => n4357, S => n525, Z => n7737);
   U16753 : XOR2_X1 port map( A => n7737, B => n4130, Z => n4360);
   U16754 : MUX2_X1 port map( A => n4359, B => n355, S => n2144, Z => n8094);
   U16755 : INV_X1 port map( A => n8094, ZN => n7736);
   U16756 : XOR2_X1 port map( A => n4360, B => n7736, Z => n7618);
   U16757 : INV_X1 port map( A => n7618, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_25_port);
   U16758 : INV_X1 port map( A => n4360, ZN => n4361);
   U16759 : NAND2_X1 port map( A1 => n4361, A2 => n7736, ZN => n7702);
   U16760 : INV_X1 port map( A => n7702, ZN => n8324);
   U16761 : INV_X1 port map( A => n4362, ZN => n4363);
   U16762 : NAND2_X1 port map( A1 => n4363, A2 => n7709, ZN => n7636);
   U16763 : INV_X1 port map( A => n7636, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_26_port);
   U16764 : XOR2_X1 port map( A => n7471, B => n4130, Z => n4373);
   U16765 : MUX2_X1 port map( A => n4367, B => n4366, S => n2145, Z => n7315);
   U16766 : INV_X1 port map( A => n7315, ZN => n7644);
   U16767 : MUX2_X1 port map( A => n4369, B => n4368, S => n525, Z => n7678);
   U16768 : XOR2_X1 port map( A => n7678, B => n4130, Z => n4371);
   U16769 : MUX2_X1 port map( A => n4370, B => n356, S => n2145, Z => n7670);
   U16770 : INV_X1 port map( A => n7670, ZN => n7677);
   U16771 : XOR2_X1 port map( A => n4371, B => n7677, Z => n7622);
   U16772 : INV_X1 port map( A => n7622, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_27_port);
   U16773 : INV_X1 port map( A => n4371, ZN => n4372);
   U16774 : NAND2_X1 port map( A1 => n4372, A2 => n7677, ZN => n7620);
   U16775 : INV_X1 port map( A => n7620, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_27_port);
   U16776 : NOR2_X1 port map( A1 => n7315, A2 => n4373, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_28_port);
   U16777 : NOR2_X1 port map( A1 => n8186, A2 => n4376, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_6_port);
   U16778 : OAI22_X1 port map( A1 => n4379, A2 => n4378, B1 => n17239, B2 => 
                           n4377, ZN => n11536);
   U16779 : NOR2_X1 port map( A1 => n8149, A2 => n4382, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_10_port);
   U16780 : OAI22_X1 port map( A1 => n4385, A2 => n4384, B1 => n2205, B2 => 
                           n4383, ZN => n11519);
   U16781 : NOR2_X1 port map( A1 => n8256, A2 => n4388, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_14_port);
   U16782 : OAI22_X1 port map( A1 => n4391, A2 => n4390, B1 => n2178, B2 => 
                           n4389, ZN => n11522);
   U16783 : XOR2_X1 port map( A => n6369, B => n4130, Z => n4404);
   U16784 : MUX2_X1 port map( A => n4392, B => n331, S => n2144, Z => n7289);
   U16785 : INV_X1 port map( A => n7289, ZN => n7899);
   U16786 : XOR2_X1 port map( A => n4404, B => n7899, Z => n4405);
   U16787 : INV_X1 port map( A => n4405, ZN => n7892);
   U16788 : MUX2_X1 port map( A => n4394, B => n4393, S => n525, Z => n7933);
   U16789 : XOR2_X1 port map( A => n7933, B => n259, Z => n4402);
   U16790 : MUX2_X1 port map( A => n4395, B => n332, S => n2144, Z => n7923);
   U16791 : INV_X1 port map( A => n7923, ZN => n7932);
   U16792 : XOR2_X1 port map( A => n4402, B => n7932, Z => n7883);
   U16793 : INV_X1 port map( A => n7883, ZN => n7918);
   U16794 : MUX2_X1 port map( A => n277, B => n358, S => n525, Z => n8215);
   U16795 : XOR2_X1 port map( A => n8215, B => n4130, Z => n4398);
   U16796 : MUX2_X1 port map( A => n4396, B => n333, S => n2143, Z => n7286);
   U16797 : INV_X1 port map( A => n7286, ZN => n8217);
   U16798 : XOR2_X1 port map( A => n4398, B => n8217, Z => n8222);
   U16799 : XOR2_X1 port map( A => n529, B => n4130, Z => n4400);
   U16800 : MUX2_X1 port map( A => n4397, B => n334, S => n2145, Z => n7283);
   U16801 : INV_X1 port map( A => n7283, ZN => n7968);
   U16802 : XOR2_X1 port map( A => n4400, B => n7968, Z => n7951);
   U16803 : NOR2_X1 port map( A1 => n8222, A2 => n7951, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_18_port);
   U16804 : INV_X1 port map( A => n4398, ZN => n4399);
   U16805 : NAND2_X1 port map( A1 => n4399, A2 => n8217, ZN => n7960);
   U16806 : INV_X1 port map( A => n4400, ZN => n4401);
   U16807 : NAND2_X1 port map( A1 => n4401, A2 => n7968, ZN => n7880);
   U16808 : OAI21_X1 port map( B1 => n7951, B2 => n7960, A => n7880, ZN => 
                           n11526);
   U16809 : INV_X1 port map( A => n4402, ZN => n4403);
   U16810 : NAND2_X1 port map( A1 => n4403, A2 => n7932, ZN => n7889);
   U16811 : OAI22_X1 port map( A1 => n4405, A2 => n7889, B1 => n7289, B2 => 
                           n4404, ZN => n11527);
   U16812 : XOR2_X1 port map( A => n6594, B => n259, Z => n4424);
   U16813 : MUX2_X1 port map( A => n4408, B => n359, S => n2144, Z => n7302);
   U16814 : INV_X1 port map( A => n7302, ZN => n7768);
   U16815 : XOR2_X1 port map( A => n4424, B => n7768, Z => n4425);
   U16816 : INV_X1 port map( A => n4425, ZN => n7761);
   U16817 : MUX2_X1 port map( A => n4410, B => n4409, S => n525, Z => n7800);
   U16818 : XOR2_X1 port map( A => n7800, B => n259, Z => n4422);
   U16819 : MUX2_X1 port map( A => n4411, B => n335, S => n2144, Z => n7792);
   U16820 : INV_X1 port map( A => n7792, ZN => n7799);
   U16821 : XOR2_X1 port map( A => n4422, B => n7799, Z => n7752);
   U16822 : INV_X1 port map( A => n7752, ZN => n7787);
   U16823 : MUX2_X1 port map( A => n4413, B => n4412, S => n527, Z => n7865);
   U16824 : XOR2_X1 port map( A => n7865, B => n259, Z => n4418);
   U16825 : MUX2_X1 port map( A => n4414, B => n336, S => n2144, Z => n7864);
   U16826 : INV_X1 port map( A => n7864, ZN => n7863);
   U16827 : XOR2_X1 port map( A => n4418, B => n7863, Z => n7860);
   U16828 : XOR2_X1 port map( A => n6495, B => n259, Z => n4420);
   U16829 : MUX2_X1 port map( A => n4417, B => n337, S => n2144, Z => n7294);
   U16830 : INV_X1 port map( A => n7294, ZN => n7832);
   U16831 : XOR2_X1 port map( A => n4420, B => n7832, Z => n7817);
   U16832 : NOR2_X1 port map( A1 => n7860, A2 => n7817, ZN => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_1_22_port);
   U16833 : INV_X1 port map( A => n4418, ZN => n4419);
   U16834 : NAND2_X1 port map( A1 => n4419, A2 => n7863, ZN => n7825);
   U16835 : INV_X1 port map( A => n4420, ZN => n4421);
   U16836 : NAND2_X1 port map( A1 => n4421, A2 => n7832, ZN => n7749);
   U16837 : OAI21_X1 port map( B1 => n7817, B2 => n7825, A => n7749, ZN => 
                           n11529);
   U16838 : INV_X1 port map( A => n4422, ZN => n4423);
   U16839 : NAND2_X1 port map( A1 => n4423, A2 => n7799, ZN => n7758);
   U16840 : OAI22_X1 port map( A1 => n4425, A2 => n7758, B1 => n7302, B2 => 
                           n4424, ZN => n11530);
   U16841 : INV_X1 port map( A => n12918, ZN => n11518);
   U16842 : INV_X1 port map( A => n12920, ZN => n11525);
   U16843 : INV_X1 port map( A => n12917, ZN => n11534);
   U16844 : INV_X1 port map( A => n12929, ZN => n8326);
   U16845 : INV_X1 port map( A => CU_I_n71, ZN => n4427);
   U16846 : NAND2_X1 port map( A1 => n4427, A2 => n4426, ZN => n7077);
   U16847 : INV_X1 port map( A => n7077, ZN => i_EN2);
   U16848 : NAND3_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n549, A2 => 
                           n8181, A3 => n2250, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n600);
   U16849 : INV_X1 port map( A => n4428, ZN => n7747);
   U16850 : OAI21_X1 port map( B1 => DataPath_i_PIPLIN_B_0_port, B2 => n2140, A
                           => CU_I_n107, ZN => n4430);
   U16851 : OAI21_X1 port map( B1 => DataPath_i_PIPLIN_IN2_0_port, B2 => n2139,
                           A => i_S2, ZN => n4429);
   U16852 : NAND2_X1 port map( A1 => n1907, A2 => n1208, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n155);
   U16853 : MUX2_X1 port map( A => n4432, B => n4431, S => n527, Z => n7579);
   U16854 : INV_X1 port map( A => n7579, ZN => n7581);
   U16855 : XOR2_X1 port map( A => n7647, B => n7581, Z => n4435);
   U16856 : MUX2_X1 port map( A => n4434, B => n4433, S => n525, Z => n7608);
   U16857 : XOR2_X1 port map( A => n7608, B => n7647, Z => n7230);
   U16858 : NAND2_X1 port map( A1 => n4435, A2 => n7230, ZN => n7231);
   U16859 : OAI22_X1 port map( A1 => n2147, A2 => n7231, B1 => n2230, B2 => 
                           n7230, ZN => n7487);
   U16860 : INV_X1 port map( A => n7487, ZN => n7229);
   U16861 : XOR2_X1 port map( A => n7712, B => n7647, Z => n4437);
   U16862 : XOR2_X1 port map( A => n7678, B => n7712, Z => n7236);
   U16863 : NAND2_X1 port map( A1 => n4437, A2 => n7236, ZN => n7237);
   U16864 : OAI22_X1 port map( A1 => n2227, A2 => n7237, B1 => n2240, B2 => 
                           n7236, ZN => n7478);
   U16865 : NAND2_X1 port map( A1 => n7110, A2 => n8181, ZN => n8023);
   U16866 : NAND2_X1 port map( A1 => n8089, A2 => n8023, ZN => n4899);
   U16867 : XOR2_X1 port map( A => n2247, B => n609, Z => n4438);
   U16868 : NAND2_X1 port map( A1 => n1242, A2 => n4438, ZN => n7316);
   U16869 : OAI22_X1 port map( A1 => n7864, A2 => n2226, B1 => n2224, B2 => 
                           n7294, ZN => n5236);
   U16870 : NAND2_X1 port map( A1 => n4444, A2 => n4443, ZN => n4570);
   U16871 : OAI22_X1 port map( A1 => n731, A2 => n4442, B1 => n4441, B2 => n838
                           , ZN => n4552);
   U16872 : OAI22_X1 port map( A1 => n7792, A2 => n2141, B1 => n2188, B2 => 
                           n7302, ZN => n5225);
   U16873 : NAND2_X1 port map( A1 => n703, A2 => n1619, ZN => n4575);
   U16874 : NAND2_X1 port map( A1 => n2149, A2 => n834, ZN => n4574);
   U16875 : NAND2_X1 port map( A1 => n4575, A2 => n4574, ZN => n4583);
   U16876 : OAI22_X1 port map( A1 => n1716, A2 => i_S2, B1 => n1302, B2 => 
                           n1745, ZN => n4448);
   U16877 : AOI22_X1 port map( A1 => n2148, A2 => DataPath_i_PIPLIN_IN1_2_port,
                           B1 => n544, B2 => DataPath_i_PIPLIN_A_2_port, ZN => 
                           n4447);
   U16878 : OAI21_X1 port map( B1 => DataPath_i_PIPLIN_IN1_0_port, B2 => 
                           DataPath_i_PIPLIN_IN1_1_port, A => n2148, ZN => 
                           n4446);
   U16879 : OAI21_X1 port map( B1 => DataPath_i_PIPLIN_A_0_port, B2 => 
                           DataPath_i_PIPLIN_A_1_port, A => n547, ZN => n4445);
   U16881 : OAI21_X1 port map( B1 => n1155, B2 => n703, A => n4576, ZN => n4556
                           );
   U16882 : NAND2_X1 port map( A1 => n703, A2 => n812, ZN => n4549);
   U16883 : NAND2_X1 port map( A1 => n2149, A2 => n1619, ZN => n4548);
   U16884 : OAI21_X1 port map( B1 => n7658, B2 => n841, A => n4547, ZN => n4555
                           );
   U16885 : INV_X1 port map( A => n4555, ZN => n4452);
   U16886 : NAND3_X1 port map( A1 => n4557, A2 => n4548, A3 => n4549, ZN => 
                           n4579);
   U16887 : OAI22_X1 port map( A1 => n8045, A2 => n6858, B1 => n2270, B2 => 
                           n2201, ZN => n4598);
   U16888 : INV_X1 port map( A => n4598, ZN => n4538);
   U16889 : INV_X1 port map( A => n4453, ZN => n4599);
   U16890 : OAI22_X1 port map( A1 => n1146, A2 => n6858, B1 => n2270, B2 => 
                           n809, ZN => n4528);
   U16891 : OAI22_X1 port map( A1 => n2196, A2 => n2195, B1 => n830, B2 => 
                           n2210, ZN => n4629);
   U16892 : INV_X1 port map( A => n4629, ZN => n4630);
   U16893 : OAI22_X1 port map( A1 => n2208, A2 => n2194, B1 => n2269, B2 => 
                           n2206, ZN => n4455);
   U16894 : INV_X1 port map( A => n4455, ZN => n4532);
   U16895 : NAND2_X1 port map( A1 => n680, A2 => n4532, ZN => n4534);
   U16896 : OAI22_X1 port map( A1 => n2204, A2 => n2194, B1 => n2269, B2 => 
                           n2216, ZN => n4456);
   U16897 : INV_X1 port map( A => n4456, ZN => n4524);
   U16898 : OAI22_X1 port map( A1 => n2216, A2 => n2136, B1 => n2269, B2 => 
                           n2214, ZN => n4457);
   U16899 : INV_X1 port map( A => n4457, ZN => n4520);
   U16900 : OAI22_X1 port map( A1 => n2213, A2 => n2135, B1 => n2269, B2 => 
                           n2175, ZN => n4458);
   U16901 : INV_X1 port map( A => n4458, ZN => n4516);
   U16902 : OAI22_X1 port map( A1 => n2175, A2 => n2137, B1 => n2269, B2 => 
                           n2177, ZN => n4459);
   U16903 : INV_X1 port map( A => n4459, ZN => n4510);
   U16904 : OAI22_X1 port map( A1 => n2177, A2 => n2136, B1 => n2269, B2 => 
                           n2179, ZN => n4460);
   U16905 : INV_X1 port map( A => n4460, ZN => n4506);
   U16906 : OAI22_X1 port map( A1 => n2179, A2 => n2136, B1 => n2269, B2 => 
                           n7283, ZN => n4461);
   U16907 : INV_X1 port map( A => n4461, ZN => n4501);
   U16908 : OAI22_X1 port map( A1 => n7283, A2 => n2136, B1 => n2269, B2 => 
                           n7923, ZN => n4462);
   U16909 : OAI22_X1 port map( A1 => n7923, A2 => n2136, B1 => n2269, B2 => 
                           n7289, ZN => n4463);
   U16910 : OAI22_X1 port map( A1 => n7289, A2 => n2136, B1 => n2269, B2 => 
                           n7864, ZN => n4464);
   U16911 : INV_X1 port map( A => n4464, ZN => n4491);
   U16912 : OAI22_X1 port map( A1 => n7864, A2 => n2136, B1 => n2269, B2 => 
                           n7294, ZN => n4465);
   U16913 : INV_X1 port map( A => n4465, ZN => n4487);
   U16914 : OAI22_X1 port map( A1 => n7294, A2 => n2136, B1 => n2269, B2 => 
                           n7792, ZN => n4466);
   U16915 : INV_X1 port map( A => n4466, ZN => n4483);
   U16916 : OAI22_X1 port map( A1 => n7792, A2 => n2136, B1 => n2269, B2 => 
                           n7302, ZN => n4467);
   U16917 : INV_X1 port map( A => n4467, ZN => n4479);
   U16919 : OAI22_X1 port map( A1 => n7302, A2 => n2136, B1 => n2269, B2 => 
                           n8094, ZN => n4468);
   U16920 : INV_X1 port map( A => n4468, ZN => n4475);
   U16922 : NAND2_X1 port map( A1 => n4477, A2 => n2259, ZN => n4471);
   U16923 : OAI22_X1 port map( A1 => n8094, A2 => n2136, B1 => n2269, B2 => 
                           n7311, ZN => n4470);
   U16924 : INV_X1 port map( A => n4470, ZN => n4472);
   U16925 : MUX2_X1 port map( A => n4471, B => n2261, S => n4472, Z => n4474);
   U16928 : NAND2_X1 port map( A1 => n4474, A2 => n5214, ZN => n5224);
   U16929 : INV_X1 port map( A => n5224, ZN => n5222);
   U16931 : OAI22_X1 port map( A1 => n7294, A2 => n2141, B1 => n2190, B2 => 
                           n7792, ZN => n4695);
   U16932 : INV_X1 port map( A => n4695, ZN => n4688);
   U16933 : NAND2_X1 port map( A1 => n4481, A2 => n2259, ZN => n4476);
   U16934 : MUX2_X1 port map( A => n4476, B => n2259, S => n4475, Z => n4478);
   U16935 : NAND2_X1 port map( A1 => n4478, A2 => n4477, ZN => n4690);
   U16936 : INV_X1 port map( A => n4690, ZN => n4694);
   U16937 : OAI22_X1 port map( A1 => n7864, A2 => n2141, B1 => n2188, B2 => 
                           n7294, ZN => n4702);
   U16938 : INV_X1 port map( A => n4702, ZN => n4685);
   U16939 : NAND2_X1 port map( A1 => n4485, A2 => n2259, ZN => n4480);
   U16940 : MUX2_X1 port map( A => n4480, B => n2259, S => n4479, Z => n4482);
   U16941 : NAND2_X1 port map( A1 => n4482, A2 => n4481, ZN => n4687);
   U16942 : INV_X1 port map( A => n4687, ZN => n4701);
   U16943 : OAI22_X1 port map( A1 => n7289, A2 => n2142, B1 => n2190, B2 => 
                           n7864, ZN => n4709);
   U16944 : INV_X1 port map( A => n4709, ZN => n4682);
   U16945 : NAND2_X1 port map( A1 => n4489, A2 => n2259, ZN => n4484);
   U16946 : MUX2_X1 port map( A => n4484, B => n2259, S => n4483, Z => n4486);
   U16947 : NAND2_X1 port map( A1 => n4486, A2 => n4485, ZN => n4684);
   U16948 : INV_X1 port map( A => n4684, ZN => n4708);
   U16949 : OAI22_X1 port map( A1 => n7923, A2 => n2142, B1 => n2188, B2 => 
                           n7289, ZN => n4715);
   U16950 : INV_X1 port map( A => n4715, ZN => n4679);
   U16951 : NAND2_X1 port map( A1 => n4493, A2 => n2259, ZN => n4488);
   U16952 : MUX2_X1 port map( A => n4488, B => n2259, S => n4487, Z => n4490);
   U16953 : OAI22_X1 port map( A1 => n7283, A2 => n2141, B1 => n2190, B2 => 
                           n7923, ZN => n4722);
   U16954 : INV_X1 port map( A => n4722, ZN => n4676);
   U16955 : NAND2_X1 port map( A1 => n4496, A2 => n2259, ZN => n4492);
   U16956 : MUX2_X1 port map( A => n4492, B => n2259, S => n4491, Z => n4494);
   U16957 : NAND2_X1 port map( A1 => n4494, A2 => n4493, ZN => n4678);
   U16958 : INV_X1 port map( A => n4678, ZN => n4721);
   U16959 : INV_X1 port map( A => n4729, ZN => n4673);
   U16960 : NAND2_X1 port map( A1 => n4499, A2 => n2259, ZN => n4495);
   U16961 : NAND2_X1 port map( A1 => n4497, A2 => n4496, ZN => n4675);
   U16962 : INV_X1 port map( A => n4675, ZN => n4728);
   U16963 : NAND2_X1 port map( A1 => n4503, A2 => n2259, ZN => n4498);
   U16964 : NAND2_X1 port map( A1 => n4500, A2 => n4499, ZN => n4624);
   U16965 : OAI22_X1 port map( A1 => n2178, A2 => n2141, B1 => n2190, B2 => 
                           n2179, ZN => n4733);
   U16966 : NAND2_X1 port map( A1 => n682, A2 => n4733, ZN => n4610);
   U16967 : INV_X1 port map( A => n4610, ZN => n4613);
   U16968 : INV_X1 port map( A => n4733, ZN => n4621);
   U16969 : OAI22_X1 port map( A1 => n2175, A2 => n2142, B1 => n2190, B2 => 
                           n2178, ZN => n4750);
   U16970 : INV_X1 port map( A => n4750, ZN => n4627);
   U16971 : NAND2_X1 port map( A1 => n4508, A2 => n2260, ZN => n4502);
   U16972 : MUX2_X1 port map( A => n4502, B => n2261, S => n4501, Z => n4504);
   U16973 : NAND2_X1 port map( A1 => n4504, A2 => n4503, ZN => n4622);
   U16974 : NAND2_X1 port map( A1 => n4627, A2 => n4622, ZN => n4738);
   U16975 : INV_X1 port map( A => n4738, ZN => n4505);
   U16976 : AOI21_X1 port map( B1 => n4624, B2 => n4621, A => n4505, ZN => 
                           n4612);
   U16977 : OAI22_X1 port map( A1 => n2213, A2 => n2142, B1 => n2190, B2 => 
                           n2176, ZN => n4757);
   U16978 : INV_X1 port map( A => n4757, ZN => n4514);
   U16979 : NAND2_X1 port map( A1 => n4512, A2 => n2260, ZN => n4507);
   U16980 : MUX2_X1 port map( A => n4507, B => n2261, S => n4506, Z => n4509);
   U16981 : NAND2_X1 port map( A1 => n4509, A2 => n4508, ZN => n4756);
   U16982 : NAND2_X1 port map( A1 => n4518, A2 => n2260, ZN => n4511);
   U16983 : MUX2_X1 port map( A => n4511, B => n2261, S => n4510, Z => n4513);
   U16984 : NAND2_X1 port map( A1 => n4513, A2 => n4512, ZN => n4628);
   U16985 : INV_X1 port map( A => n4628, ZN => n4770);
   U16986 : OAI22_X1 port map( A1 => n2215, A2 => n2141, B1 => n2188, B2 => 
                           n2213, ZN => n4771);
   U16987 : NAND2_X1 port map( A1 => n4770, A2 => n4771, ZN => n4758);
   U16988 : OAI22_X1 port map( A1 => n4514, A2 => n4756, B1 => n1060, B2 => 
                           n4758, ZN => n4515);
   U16989 : INV_X1 port map( A => n4515, ZN => n4735);
   U16990 : INV_X1 port map( A => n4622, ZN => n4749);
   U16991 : NAND2_X1 port map( A1 => n4749, A2 => n4750, ZN => n4736);
   U16992 : INV_X1 port map( A => n4771, ZN => n4625);
   U16993 : NAND2_X1 port map( A1 => n4625, A2 => n4628, ZN => n4760);
   U16994 : OAI22_X1 port map( A1 => n2204, A2 => n2141, B1 => n2190, B2 => 
                           n2215, ZN => n4777);
   U16995 : INV_X1 port map( A => n4777, ZN => n4666);
   U16996 : NAND2_X1 port map( A1 => n4522, A2 => n2260, ZN => n4517);
   U16997 : MUX2_X1 port map( A => n4517, B => n2261, S => n4516, Z => n4519);
   U16998 : NAND2_X1 port map( A1 => n4519, A2 => n4518, ZN => n4668);
   U16999 : INV_X1 port map( A => n4668, ZN => n4776);
   U17000 : OAI22_X1 port map( A1 => n2208, A2 => n2142, B1 => n2190, B2 => 
                           n2206, ZN => n4784);
   U17001 : INV_X1 port map( A => n4784, ZN => n4663);
   U17002 : NAND2_X1 port map( A1 => n4526, A2 => n2260, ZN => n4521);
   U17003 : MUX2_X1 port map( A => n4521, B => n2261, S => n4520, Z => n4523);
   U17004 : NAND2_X1 port map( A1 => n4523, A2 => n4522, ZN => n4665);
   U17005 : INV_X1 port map( A => n4665, ZN => n4783);
   U17006 : OAI22_X1 port map( A1 => n2196, A2 => n2141, B1 => n2188, B2 => 
                           n2210, ZN => n4791);
   U17007 : INV_X1 port map( A => n4791, ZN => n4660);
   U17008 : NAND2_X1 port map( A1 => n4534, A2 => n2260, ZN => n4525);
   U17009 : MUX2_X1 port map( A => n4525, B => n2261, S => n4524, Z => n4527);
   U17010 : NAND2_X1 port map( A1 => n4527, A2 => n4526, ZN => n4662);
   U17011 : INV_X1 port map( A => n4662, ZN => n4790);
   U17012 : OAI22_X1 port map( A1 => n2200, A2 => n2142, B1 => n2188, B2 => 
                           n2198, ZN => n4798);
   U17013 : INV_X1 port map( A => n4798, ZN => n4606);
   U17014 : INV_X1 port map( A => n596, ZN => n4580);
   U17015 : NAND3_X1 port map( A1 => n1891, A2 => n4580, A3 => n831, ZN => 
                           n4854);
   U17016 : INV_X1 port map( A => n4854, ZN => n4541);
   U17017 : INV_X1 port map( A => n4857, ZN => n4543);
   U17018 : INV_X1 port map( A => n4529, ZN => n4530);
   U17019 : NAND4_X1 port map( A1 => n4541, A2 => n4543, A3 => n4630, A4 => 
                           n4530, ZN => n4531);
   U17020 : NAND2_X1 port map( A1 => n4531, A2 => n2260, ZN => n4533);
   U17021 : MUX2_X1 port map( A => n4533, B => n2261, S => n4532, Z => n4535);
   U17022 : NAND4_X1 port map( A1 => n1730, A2 => n831, A3 => n4580, A4 => 
                           n4543, ZN => n4536);
   U17023 : NAND2_X1 port map( A1 => n4536, A2 => n2260, ZN => n4537);
   U17024 : MUX2_X1 port map( A => n4537, B => n2261, S => n4538, Z => n4540);
   U17025 : NAND3_X1 port map( A1 => n4541, A2 => n4538, A3 => n4543, ZN => 
                           n4539);
   U17026 : NAND2_X1 port map( A1 => n4540, A2 => n4539, ZN => n4654);
   U17027 : INV_X1 port map( A => n4654, ZN => n4849);
   U17028 : OAI22_X1 port map( A1 => n2138, A2 => n2141, B1 => n2190, B2 => 
                           n2238, ZN => n4850);
   U17029 : NAND2_X1 port map( A1 => n4849, A2 => n4850, ZN => n4831);
   U17030 : NAND2_X1 port map( A1 => n4541, A2 => n4543, ZN => n4855);
   U17031 : INV_X1 port map( A => n4855, ZN => n4546);
   U17032 : NAND2_X1 port map( A1 => n1891, A2 => n831, ZN => n4587);
   U17033 : INV_X1 port map( A => n4587, ZN => n4542);
   U17035 : INV_X1 port map( A => n17247, ZN => n4635);
   U17036 : OAI22_X1 port map( A1 => n2240, A2 => n2142, B1 => n2239, B2 => 
                           n2188, ZN => n4651);
   U17037 : NAND2_X1 port map( A1 => n4635, A2 => n4651, ZN => n4844);
   U17038 : INV_X1 port map( A => n4651, ZN => n4858);
   U17039 : NAND2_X1 port map( A1 => n4858, A2 => n17247, ZN => n4843);
   U17040 : OAI21_X1 port map( B1 => n6858, B2 => n7658, A => n761, ZN => n4585
                           );
   U17041 : INV_X1 port map( A => n4555, ZN => n4557);
   U17042 : NAND2_X1 port map( A1 => n573, A2 => n1833, ZN => n4586);
   U17043 : INV_X1 port map( A => n4586, ZN => n4550);
   U17044 : NAND2_X1 port map( A1 => n835, A2 => n4550, ZN => n4571);
   U17045 : OAI22_X1 port map( A1 => n2262, A2 => n4557, B1 => n573, B2 => 
                           n17165, ZN => n4551);
   U17046 : XOR2_X1 port map( A => n4552, B => n1906, Z => n4558);
   U17047 : NAND2_X1 port map( A1 => n555, A2 => n1315, ZN => n4871);
   U17048 : NAND4_X1 port map( A1 => n4561, A2 => n7196, A3 => n609, A4 => 
                           n8277, ZN => n4554);
   U17049 : NAND4_X1 port map( A1 => n8277, A2 => n8208, A3 => n7110, A4 => 
                           n2130, ZN => n4553);
   U17050 : OAI211_X1 port map( C1 => n17195, C2 => n4558, A => n4554, B => 
                           n4553, ZN => n4643);
   U17051 : INV_X1 port map( A => n546, ZN => n8187);
   U17052 : NAND2_X1 port map( A1 => n4641, A2 => n1870, ZN => n4642);
   U17053 : INV_X1 port map( A => n216, ZN => n4559);
   U17054 : OAI22_X1 port map( A1 => n2131, A2 => n6858, B1 => n519, B2 => 
                           n7688, ZN => n8204);
   U17055 : NAND2_X1 port map( A1 => n8277, A2 => n2149, ZN => n8206);
   U17056 : INV_X1 port map( A => n8206, ZN => n8280);
   U17057 : NOR3_X1 port map( A1 => n8204, A2 => n8280, A3 => n4561, ZN => 
                           n4566);
   U17058 : AOI22_X1 port map( A1 => n2233, A2 => n2149, B1 => n703, B2 => 
                           n2235, ZN => n4560);
   U17059 : OAI22_X1 port map( A1 => n8276, A2 => n7688, B1 => n841, B2 => 
                           n8091, ZN => n4562);
   U17060 : INV_X1 port map( A => n4562, ZN => n4568);
   U17061 : OAI22_X1 port map( A1 => n841, A2 => n7688, B1 => n8276, B2 => 
                           n7658, ZN => n4563);
   U17062 : INV_X1 port map( A => n4563, ZN => n4569);
   U17063 : NAND3_X1 port map( A1 => n4568, A2 => n8206, A3 => n4569, ZN => 
                           n4564);
   U17064 : INV_X1 port map( A => n1549, ZN => n4567);
   U17065 : NAND2_X1 port map( A1 => n4567, A2 => n1878, ZN => n8189);
   U17066 : INV_X1 port map( A => n8188, ZN => n4645);
   U17067 : NAND2_X1 port map( A1 => n4645, A2 => n691, ZN => n4889);
   U17068 : OAI21_X1 port map( B1 => n8189, B2 => n1825, A => n4889, ZN => 
                           n4573);
   U17069 : INV_X1 port map( A => n493, ZN => n4891);
   U17070 : OAI21_X1 port map( B1 => n4647, B2 => n1199, A => n4891, ZN => 
                           n4572);
   U17071 : NAND2_X1 port map( A1 => n4573, A2 => n4572, ZN => n4870);
   U17072 : NAND2_X1 port map( A1 => n4870, A2 => n4871, ZN => n4861);
   U17073 : INV_X1 port map( A => n4861, ZN => n4594);
   U17074 : INV_X1 port map( A => n4884, ZN => n4592);
   U17075 : INV_X1 port map( A => n4574, ZN => n4578);
   U17076 : INV_X1 port map( A => n4575, ZN => n4577);
   U17077 : NOR4_X1 port map( A1 => n4579, A2 => n4578, A3 => n4577, A4 => 
                           n1552, ZN => n4582);
   U17078 : NAND2_X1 port map( A1 => n597, A2 => n2232, ZN => n4591);
   U17079 : NAND2_X1 port map( A1 => n1873, A2 => n2228, ZN => n4590);
   U17080 : NAND2_X1 port map( A1 => n17243, A2 => n4590, ZN => n4885);
   U17081 : XOR2_X1 port map( A => n4583, B => n2262, Z => n4584);
   U17082 : OAI21_X1 port map( B1 => n4586, B2 => n819, A => n4584, ZN => n4588
                           );
   U17083 : NAND2_X1 port map( A1 => n4588, A2 => n4587, ZN => n4639);
   U17084 : NAND2_X1 port map( A1 => n4637, A2 => n17228, ZN => n4872);
   U17085 : NAND2_X1 port map( A1 => n4589, A2 => n4872, ZN => n4860);
   U17086 : NAND2_X1 port map( A1 => n4591, A2 => n4590, ZN => n4636);
   U17087 : NAND2_X1 port map( A1 => n1564, A2 => n4636, ZN => n4877);
   U17088 : OAI22_X1 port map( A1 => n827, A2 => n4877, B1 => n753, B2 => n4592
                           , ZN => n4593);
   U17089 : INV_X1 port map( A => n4593, ZN => n4865);
   U17090 : NAND2_X1 port map( A1 => n475, A2 => n4843, ZN => n4834);
   U17091 : NAND3_X1 port map( A1 => n4834, A2 => n4844, A3 => n4831, ZN => 
                           n4820);
   U17092 : OAI22_X1 port map( A1 => n17238, A2 => n2141, B1 => n2189, B2 => 
                           n2200, ZN => n4829);
   U17093 : INV_X1 port map( A => n4829, ZN => n4631);
   U17094 : NAND2_X1 port map( A1 => n4600, A2 => n2260, ZN => n4595);
   U17095 : MUX2_X1 port map( A => n4595, B => n2261, S => n4630, Z => n4597);
   U17096 : NAND2_X1 port map( A1 => n4597, A2 => n4596, ZN => n4633);
   U17097 : NAND2_X1 port map( A1 => n4631, A2 => n4633, ZN => n4809);
   U17098 : INV_X1 port map( A => n4850, ZN => n4634);
   U17099 : NAND2_X1 port map( A1 => n4634, A2 => n4654, ZN => n4835);
   U17100 : NAND2_X1 port map( A1 => n4606, A2 => n4797, ZN => n4603);
   U17101 : OAI22_X1 port map( A1 => n2238, A2 => n2141, B1 => n2188, B2 => 
                           n17239, ZN => n4842);
   U17102 : INV_X1 port map( A => n4842, ZN => n4632);
   U17103 : XOR2_X1 port map( A => n2262, B => n4599, Z => n4601);
   U17104 : OAI21_X1 port map( B1 => n4602, B2 => n4601, A => n4600, ZN => 
                           n4655);
   U17105 : NAND2_X1 port map( A1 => n17217, A2 => n4632, ZN => n4819);
   U17106 : NAND4_X1 port map( A1 => n4809, A2 => n4835, A3 => n4603, A4 => 
                           n4819, ZN => n4605);
   U17107 : INV_X1 port map( A => n4655, ZN => n4841);
   U17108 : INV_X1 port map( A => n4633, ZN => n4828);
   U17109 : OAI21_X1 port map( B1 => n1602, B2 => n941, A => n4603, ZN => n4604
                           );
   U17110 : OAI221_X1 port map( B1 => n4606, B2 => n4797, C1 => n474, C2 => 
                           n4605, A => n4604, ZN => n4792);
   U17111 : NAND3_X1 port map( A1 => n4760, A2 => n4772, A3 => n4609, ZN => 
                           n4734);
   U17112 : OAI21_X1 port map( B1 => n4613, B2 => n4612, A => n4611, ZN => 
                           n4614);
   U17113 : OAI21_X1 port map( B1 => n4708, B2 => n4709, A => n4710, ZN => 
                           n4618);
   U17114 : NAND2_X1 port map( A1 => n4750, A2 => n4622, ZN => n4745);
   U17115 : INV_X1 port map( A => n4745, ZN => n4623);
   U17116 : AOI21_X1 port map( B1 => n4733, B2 => n4624, A => n4623, ZN => 
                           n4671);
   U17117 : NAND2_X1 port map( A1 => n4757, A2 => n4756, ZN => n4669);
   U17118 : NAND2_X1 port map( A1 => n4770, A2 => n4625, ZN => n4763);
   U17119 : OAI22_X1 port map( A1 => n4757, A2 => n4756, B1 => n463, B2 => 
                           n4763, ZN => n4626);
   U17120 : INV_X1 port map( A => n4626, ZN => n4742);
   U17121 : NAND2_X1 port map( A1 => n4749, A2 => n4627, ZN => n4743);
   U17122 : NAND2_X1 port map( A1 => n4771, A2 => n4628, ZN => n4765);
   U17123 : OAI33_X1 port map( A1 => n4631, A2 => n2264, A3 => n4630, B1 => 
                           n4631, B2 => n2261, B3 => n450, ZN => n4653);
   U17124 : INV_X1 port map( A => n4806, ZN => n4659);
   U17125 : NAND2_X1 port map( A1 => n4798, A2 => n4797, ZN => n4656);
   U17126 : INV_X1 port map( A => n4656, ZN => n4658);
   U17127 : NAND2_X1 port map( A1 => n1270, A2 => n4858, ZN => n4848);
   U17128 : NAND2_X1 port map( A1 => n4883, A2 => n608, ZN => n4640);
   U17129 : INV_X1 port map( A => n4640, ZN => n4638);
   U17130 : INV_X1 port map( A => n4636, ZN => n4637);
   U17131 : NAND2_X1 port map( A1 => n17212, A2 => n1564, ZN => n4876);
   U17132 : OAI22_X1 port map( A1 => n4638, A2 => n4876, B1 => n753, B2 => 
                           n1141, ZN => n4864);
   U17133 : INV_X1 port map( A => n4864, ZN => n4650);
   U17134 : NAND2_X1 port map( A1 => n4639, A2 => n4885, ZN => n4875);
   U17135 : NAND2_X1 port map( A1 => n555, A2 => n772, ZN => n4874);
   U17136 : NAND2_X1 port map( A1 => n8199, A2 => n1878, ZN => n8198);
   U17137 : INV_X1 port map( A => n4641, ZN => n4644);
   U17138 : OAI211_X1 port map( C1 => n4644, C2 => n792, A => n4642, B => n4643
                           , ZN => n4892);
   U17139 : INV_X1 port map( A => n4892, ZN => n4646);
   U17140 : OAI21_X1 port map( B1 => n4646, B2 => n1636, A => n4894, ZN => 
                           n4649);
   U17141 : OAI21_X1 port map( B1 => n4647, B2 => n1199, A => n4896, ZN => 
                           n4648);
   U17142 : NAND2_X1 port map( A1 => n4649, A2 => n4648, ZN => n4873);
   U17143 : NAND2_X1 port map( A1 => n452, A2 => n4873, ZN => n4863);
   U17144 : NAND2_X1 port map( A1 => n17262, A2 => n1851, ZN => n4845);
   U17145 : NAND2_X1 port map( A1 => n4650, A2 => n4845, ZN => n4799);
   U17146 : NAND2_X1 port map( A1 => n4652, A2 => n4651, ZN => n4846);
   U17147 : NAND2_X1 port map( A1 => n4799, A2 => n4846, ZN => n4836);
   U17148 : NAND2_X1 port map( A1 => n4836, A2 => n1274, ZN => n4821);
   U17149 : INV_X1 port map( A => n17226, ZN => n4802);
   U17150 : NAND2_X1 port map( A1 => n4850, A2 => n4654, ZN => n4823);
   U17151 : NAND2_X1 port map( A1 => n17217, A2 => n4842, ZN => n4822);
   U17152 : NAND4_X1 port map( A1 => n4802, A2 => n4823, A3 => n4656, A4 => 
                           n4822, ZN => n4657);
   U17153 : OAI222_X1 port map( A1 => n4798, A2 => n4797, B1 => n4659, B2 => 
                           n4658, C1 => n1144, C2 => n4657, ZN => n4793);
   U17154 : INV_X1 port map( A => n4730, ZN => n4672);
   U17155 : XOR2_X1 port map( A => n4691, B => n5220, Z => n4692);
   U17156 : INV_X1 port map( A => n5235, ZN => n5233);
   U17157 : OAI22_X1 port map( A1 => n7289, A2 => n2226, B1 => n2224, B2 => 
                           n7864, ZN => n4988);
   U17158 : INV_X1 port map( A => n4988, ZN => n4979);
   U17160 : XOR2_X1 port map( A => n4698, B => n4697, Z => n4699);
   U17161 : INV_X1 port map( A => n4981, ZN => n4987);
   U17162 : OAI22_X1 port map( A1 => n7923, A2 => n2225, B1 => n2224, B2 => 
                           n7289, ZN => n5006);
   U17163 : INV_X1 port map( A => n5006, ZN => n4931);
   U17164 : XOR2_X1 port map( A => n4701, B => n4702, Z => n4705);
   U17165 : XOR2_X1 port map( A => n4705, B => n4704, Z => n4706);
   U17166 : MUX2_X1 port map( A => n4707, B => n4706, S => n804, Z => n4930);
   U17167 : NAND2_X1 port map( A1 => n4931, A2 => n4930, ZN => n4993);
   U17168 : INV_X1 port map( A => n4930, ZN => n5005);
   U17169 : NAND2_X1 port map( A1 => n5005, A2 => n5006, ZN => n4991);
   U17170 : XOR2_X1 port map( A => n4709, B => n4708, Z => n4712);
   U17171 : XOR2_X1 port map( A => n4712, B => n4710, Z => n4714);
   U17172 : OAI22_X1 port map( A1 => n7283, A2 => n2226, B1 => n2224, B2 => 
                           n7923, ZN => n5013);
   U17173 : NAND2_X1 port map( A1 => n5012, A2 => n5013, ZN => n4990);
   U17174 : OAI22_X1 port map( A1 => n2179, A2 => n2225, B1 => n2224, B2 => 
                           n7283, ZN => n5020);
   U17175 : INV_X1 port map( A => n5020, ZN => n4974);
   U17176 : XOR2_X1 port map( A => n4715, B => n251, Z => n4718);
   U17177 : XOR2_X1 port map( A => n4718, B => n17235, Z => n4719);
   U17178 : INV_X1 port map( A => n4976, ZN => n5019);
   U17179 : OAI22_X1 port map( A1 => n2177, A2 => n2226, B1 => n2224, B2 => 
                           n2179, ZN => n4972);
   U17180 : INV_X1 port map( A => n4972, ZN => n5038);
   U17181 : XOR2_X1 port map( A => n4725, B => n786, Z => n4726);
   U17182 : NAND2_X1 port map( A1 => n5038, A2 => n5037, ZN => n4924);
   U17183 : INV_X1 port map( A => n4924, ZN => n4926);
   U17184 : XOR2_X1 port map( A => n1742, B => n311, Z => n4732);
   U17185 : XOR2_X1 port map( A => n4730, B => n311, Z => n4731);
   U17186 : OAI22_X1 port map( A1 => n2176, A2 => n2225, B1 => n2224, B2 => 
                           n2177, ZN => n5041);
   U17187 : NAND2_X1 port map( A1 => n779, A2 => n5041, ZN => n5031);
   U17188 : INV_X1 port map( A => n5041, ZN => n4932);
   U17189 : NAND2_X1 port map( A1 => n4932, A2 => n4933, ZN => n5027);
   U17190 : OAI22_X1 port map( A1 => n2213, A2 => n2226, B1 => n2224, B2 => 
                           n2176, ZN => n5046);
   U17191 : INV_X1 port map( A => n5046, ZN => n4967);
   U17192 : XOR2_X1 port map( A => n4733, B => n682, Z => n4740);
   U17193 : NAND2_X1 port map( A1 => n4735, A2 => n4734, ZN => n4751);
   U17194 : INV_X1 port map( A => n4736, ZN => n4737);
   U17195 : AOI21_X1 port map( B1 => n4738, B2 => n4751, A => n4737, ZN => 
                           n4739);
   U17196 : XOR2_X1 port map( A => n4739, B => n4740, Z => n4748);
   U17197 : NAND2_X1 port map( A1 => n4741, A2 => n4742, ZN => n4752);
   U17198 : INV_X1 port map( A => n4743, ZN => n4744);
   U17199 : AOI21_X1 port map( B1 => n4745, B2 => n4752, A => n4744, ZN => 
                           n4746);
   U17200 : INV_X1 port map( A => n4969, ZN => n5045);
   U17201 : OAI22_X1 port map( A1 => n2215, A2 => n2225, B1 => n2224, B2 => 
                           n2213, ZN => n5053);
   U17202 : INV_X1 port map( A => n5053, ZN => n4921);
   U17203 : XOR2_X1 port map( A => n4750, B => n4749, Z => n4753);
   U17204 : XOR2_X1 port map( A => n4753, B => n4752, Z => n4754);
   U17205 : NAND2_X1 port map( A1 => n4921, A2 => n5052, ZN => n4919);
   U17206 : INV_X1 port map( A => n4919, ZN => n4922);
   U17207 : INV_X1 port map( A => n4758, ZN => n4759);
   U17208 : AOI21_X1 port map( B1 => n4760, B2 => n4772, A => n4759, ZN => 
                           n4761);
   U17209 : XOR2_X1 port map( A => n4762, B => n4761, Z => n4769);
   U17210 : INV_X1 port map( A => n4762, ZN => n4767);
   U17211 : INV_X1 port map( A => n4763, ZN => n4764);
   U17212 : AOI21_X1 port map( B1 => n1057, B2 => n4765, A => n4764, ZN => 
                           n4766);
   U17213 : XOR2_X1 port map( A => n4767, B => n4766, Z => n4768);
   U17214 : INV_X1 port map( A => n4935, ZN => n5065);
   U17215 : OAI22_X1 port map( A1 => n2204, A2 => n2226, B1 => n2224, B2 => 
                           n2215, ZN => n5066);
   U17216 : NAND2_X1 port map( A1 => n5065, A2 => n5066, ZN => n5054);
   U17217 : INV_X1 port map( A => n5066, ZN => n4934);
   U17218 : NAND2_X1 port map( A1 => n4934, A2 => n4935, ZN => n5056);
   U17219 : OAI22_X1 port map( A1 => n2208, A2 => n2225, B1 => n2224, B2 => 
                           n2205, ZN => n5072);
   U17220 : INV_X1 port map( A => n5072, ZN => n4918);
   U17221 : XOR2_X1 port map( A => n4771, B => n4770, Z => n4773);
   U17222 : OAI22_X1 port map( A1 => n2196, A2 => n2226, B1 => n2224, B2 => 
                           n2209, ZN => n5084);
   U17223 : INV_X1 port map( A => n5084, ZN => n4936);
   U17224 : XOR2_X1 port map( A => n4777, B => n4776, Z => n4780);
   U17225 : XOR2_X1 port map( A => n4780, B => n4779, Z => n4781);
   U17226 : XOR2_X1 port map( A => n4784, B => n4783, Z => n4787);
   U17227 : XOR2_X1 port map( A => n621, B => n4787, Z => n4788);
   U17228 : INV_X1 port map( A => n4960, ZN => n5090);
   U17229 : OAI22_X1 port map( A1 => n2199, A2 => n2225, B1 => n2224, B2 => 
                           n2198, ZN => n5091);
   U17230 : NAND2_X1 port map( A1 => n5090, A2 => n5091, ZN => n5086);
   U17231 : OAI22_X1 port map( A1 => n17239, A2 => n2226, B1 => n2224, B2 => 
                           n2200, ZN => n5100);
   U17232 : INV_X1 port map( A => n5100, ZN => n4955);
   U17233 : XOR2_X1 port map( A => n4791, B => n4790, Z => n4794);
   U17234 : XOR2_X1 port map( A => n4793, B => n4794, Z => n4795);
   U17235 : INV_X1 port map( A => n4954, ZN => n5099);
   U17236 : INV_X1 port map( A => n4823, ZN => n4833);
   U17237 : NAND3_X1 port map( A1 => n4846, A2 => n4823, A3 => n4799, ZN => 
                           n4800);
   U17238 : OAI21_X1 port map( B1 => n1774, B2 => n4833, A => n4800, ZN => 
                           n4801);
   U17239 : INV_X1 port map( A => n4813, ZN => n4810);
   U17240 : OAI33_X1 port map( A1 => n449, A2 => n646, A3 => n472, B1 => n4810,
                           B2 => n4803, B3 => n818, ZN => n4818);
   U17241 : NAND3_X1 port map( A1 => n818, A2 => n4805, A3 => n4804, ZN => 
                           n4808);
   U17242 : NAND3_X1 port map( A1 => n449, A2 => n2250, A3 => n4806, ZN => 
                           n4807);
   U17243 : OAI211_X1 port map( C1 => n804, C2 => n449, A => n4808, B => n4807,
                           ZN => n4817);
   U17244 : INV_X1 port map( A => n4808, ZN => n4811);
   U17245 : NAND4_X1 port map( A1 => n4820, A2 => n4835, A3 => n4809, A4 => 
                           n4819, ZN => n4812);
   U17246 : NAND3_X1 port map( A1 => n4811, A2 => n4810, A3 => n4812, ZN => 
                           n4816);
   U17247 : INV_X1 port map( A => n4812, ZN => n4814);
   U17248 : NAND3_X1 port map( A1 => n4814, A2 => n1606, A3 => n449, ZN => 
                           n4815);
   U17249 : OAI211_X1 port map( C1 => n17185, C2 => n4817, A => n4816, B => 
                           n4815, ZN => n5187);
   U17250 : OAI22_X1 port map( A1 => n2238, A2 => n2225, B1 => n2224, B2 => 
                           n17240, ZN => n4952);
   U17251 : INV_X1 port map( A => n4952, ZN => n5186);
   U17252 : NAND2_X1 port map( A1 => n5186, A2 => n833, ZN => n4912);
   U17253 : NAND4_X1 port map( A1 => n4820, A2 => n4835, A3 => n818, A4 => 
                           n4819, ZN => n4827);
   U17254 : OAI211_X1 port map( C1 => n1839, C2 => n804, A => n4824, B => n4825
                           , ZN => n4826);
   U17255 : OAI22_X1 port map( A1 => n2138, A2 => n2226, B1 => n2224, B2 => 
                           n2238, ZN => n4949);
   U17256 : NAND2_X1 port map( A1 => n729, A2 => n4949, ZN => n5182);
   U17257 : INV_X1 port map( A => n4949, ZN => n5117);
   U17258 : NAND2_X1 port map( A1 => n5116, A2 => n5117, ZN => n5181);
   U17259 : NAND3_X1 port map( A1 => n4831, A2 => n4844, A3 => n818, ZN => 
                           n4832);
   U17260 : OAI211_X1 port map( C1 => n818, C2 => n4833, A => n4832, B => n4835
                           , ZN => n4840);
   U17261 : NAND4_X1 port map( A1 => n4836, A2 => n2250, A3 => n4837, A4 => 
                           n4848, ZN => n4838);
   U17262 : OAI22_X1 port map( A1 => n2240, A2 => n2225, B1 => n2224, B2 => 
                           n2239, ZN => n4944);
   U17263 : OAI22_X1 port map( A1 => n2227, A2 => n2226, B1 => n2224, B2 => 
                           n2240, ZN => n4947);
   U17264 : INV_X1 port map( A => n4947, ZN => n5127);
   U17265 : NAND3_X1 port map( A1 => n1569, A2 => n4843, A3 => n818, ZN => 
                           n4853);
   U17266 : OAI211_X1 port map( C1 => n1705, C2 => n1093, A => n2129, B => 
                           n4846, ZN => n4847);
   U17267 : OAI211_X1 port map( C1 => n1257, C2 => n2250, A => n4847, B => 
                           n4848, ZN => n4852);
   U17268 : NAND2_X1 port map( A1 => n4948, A2 => n5127, ZN => n5165);
   U17269 : OAI21_X1 port map( B1 => n1166, B2 => n4944, A => n5165, ZN => 
                           n4851);
   U17270 : INV_X1 port map( A => n17257, ZN => n5108);
   U17271 : NAND2_X1 port map( A1 => n4945, A2 => n4947, ZN => n5163);
   U17272 : NAND3_X1 port map( A1 => n637, A2 => n2260, A3 => n1566, ZN => 
                           n4856);
   U17273 : OAI211_X1 port map( C1 => n637, C2 => n2261, A => n4856, B => n4855
                           , ZN => n4859);
   U17274 : NOR2_X1 port map( A1 => n4904, A2 => n5145, ZN => n4869);
   U17275 : INV_X1 port map( A => n4860, ZN => n4862);
   U17276 : NAND3_X1 port map( A1 => n4862, A2 => n17181, A3 => n1606, ZN => 
                           n4908);
   U17278 : NAND3_X1 port map( A1 => n17262, A2 => n804, A3 => n1851, ZN => 
                           n4907);
   U17279 : NAND2_X1 port map( A1 => n4864, A2 => n2129, ZN => n4906);
   U17280 : NAND3_X1 port map( A1 => n4906, A2 => n4907, A3 => n4905, ZN => 
                           n4903);
   U17281 : INV_X1 port map( A => n4909, ZN => n4866);
   U17282 : NOR3_X1 port map( A1 => n5145, A2 => n17252, A3 => n4866, ZN => 
                           n4868);
   U17283 : XOR2_X1 port map( A => n4869, B => n4868, Z => n4902);
   U17284 : OAI22_X1 port map( A1 => n2147, A2 => n7316, B1 => n2229, B2 => 
                           n1242, ZN => n4941);
   U17285 : INV_X1 port map( A => n4941, ZN => n5134);
   U17286 : INV_X1 port map( A => n4872, ZN => n4882);
   U17287 : INV_X1 port map( A => n4876, ZN => n4880);
   U17288 : INV_X1 port map( A => n4877, ZN => n4878);
   U17289 : NOR2_X1 port map( A1 => n4878, A2 => n2250, ZN => n4879);
   U17290 : OAI33_X1 port map( A1 => n2251, A2 => n4882, A3 => n17241, B1 => 
                           n4881, B2 => n4880, B3 => n4879, ZN => n4910);
   U17291 : INV_X1 port map( A => n5135, ZN => n4938);
   U17292 : NAND2_X1 port map( A1 => n4911, A2 => n5134, ZN => n5149);
   U17293 : XOR2_X1 port map( A => n1564, B => n4885, Z => n4886);
   U17294 : XOR2_X1 port map( A => n1795, B => n4886, Z => n4888);
   U17295 : OAI22_X1 port map( A1 => n17194, A2 => n7316, B1 => n2147, B2 => 
                           n1242, ZN => n4943);
   U17296 : NAND2_X1 port map( A1 => n5140, A2 => n4943, ZN => n5146);
   U17297 : FA_X1 port map( A => n772, B => n1467, CI => n4890, CO => n_3778, S
                           => n4898);
   U17298 : FA_X1 port map( A => n1315, B => n1467, CI => n4895, CO => n_3779, 
                           S => n4897);
   U17302 : NAND3_X1 port map( A1 => n5147, A2 => n5146, A3 => n5148, ZN => 
                           n4901);
   U17303 : OAI211_X1 port map( C1 => n4902, C2 => n5145, A => n5149, B => 
                           n4901, ZN => n5166);
   U17305 : NAND3_X1 port map( A1 => n4906, A2 => n4905, A3 => n4907, ZN => 
                           n4909);
   U17306 : INV_X1 port map( A => n1222, ZN => n5136);
   U17307 : NAND2_X1 port map( A1 => n5164, A2 => n1288, ZN => n5124);
   U17308 : NAND3_X1 port map( A1 => n5166, A2 => n5163, A3 => n1621, ZN => 
                           n5107);
   U17309 : NAND2_X1 port map( A1 => n5107, A2 => n1269, ZN => n5183);
   U17310 : NAND2_X1 port map( A1 => n1166, A2 => n4944, ZN => n5184);
   U17311 : NAND3_X1 port map( A1 => n4913, A2 => n969, A3 => n4912, ZN => 
                           n4914);
   U17312 : OAI211_X1 port map( C1 => n4936, C2 => n4937, A => n5085, B => 
                           n5086, ZN => n5074);
   U17313 : NAND2_X1 port map( A1 => n4936, A2 => n4937, ZN => n5073);
   U17314 : NAND3_X1 port map( A1 => n5067, A2 => n5056, A3 => n4919, ZN => 
                           n4920);
   U17315 : NAND3_X1 port map( A1 => n5027, A2 => n5026, A3 => n4924, ZN => 
                           n4925);
   U17318 : NAND3_X1 port map( A1 => n4991, A2 => n4990, A3 => n4989, ZN => 
                           n4928);
   U17319 : OAI211_X1 port map( C1 => n4987, C2 => n4988, A => n4993, B => 
                           n4928, ZN => n4929);
   U17320 : NAND2_X1 port map( A1 => n5006, A2 => n4930, ZN => n5000);
   U17321 : INV_X1 port map( A => n5013, ZN => n4977);
   U17322 : NAND2_X1 port map( A1 => n5012, A2 => n4977, ZN => n4997);
   U17323 : NAND2_X1 port map( A1 => n4972, A2 => n5037, ZN => n4970);
   U17324 : INV_X1 port map( A => n4970, ZN => n4973);
   U17325 : NAND2_X1 port map( A1 => n779, A2 => n4932, ZN => n5030);
   U17326 : NAND2_X1 port map( A1 => n5041, A2 => n4933, ZN => n5029);
   U17327 : INV_X1 port map( A => n4964, ZN => n4966);
   U17328 : NAND2_X1 port map( A1 => n5065, A2 => n4934, ZN => n5059);
   U17329 : NAND2_X1 port map( A1 => n5066, A2 => n4935, ZN => n5061);
   U17330 : NAND2_X1 port map( A1 => n5072, A2 => n4963, ZN => n4961);
   U17331 : INV_X1 port map( A => n4937, ZN => n5083);
   U17332 : NAND2_X1 port map( A1 => n5083, A2 => n4936, ZN => n5077);
   U17333 : NAND2_X1 port map( A1 => n5084, A2 => n4937, ZN => n5076);
   U17334 : INV_X1 port map( A => n5091, ZN => n4958);
   U17335 : NAND2_X1 port map( A1 => n5187, A2 => n4952, ZN => n4950);
   U17336 : INV_X1 port map( A => n4950, ZN => n4953);
   U17337 : INV_X1 port map( A => n5145, ZN => n5123);
   U17338 : NAND2_X1 port map( A1 => n4939, A2 => n5134, ZN => n5153);
   U17339 : OAI21_X1 port map( B1 => n5123, B2 => n1567, A => n926, ZN => n4940
                           );
   U17340 : NAND2_X1 port map( A1 => n4911, A2 => n1322, ZN => n5156);
   U17341 : NAND2_X1 port map( A1 => n4942, A2 => n5145, ZN => n5129);
   U17342 : NAND2_X1 port map( A1 => n1875, A2 => n8180, ZN => n8179);
   U17343 : INV_X1 port map( A => n4943, ZN => n8171);
   U17344 : NAND2_X1 port map( A1 => n802, A2 => n1059, ZN => n5111);
   U17345 : INV_X1 port map( A => n4944, ZN => n5168);
   U17346 : NAND2_X1 port map( A1 => n1813, A2 => n5168, ZN => n5112);
   U17347 : NAND2_X1 port map( A1 => n4945, A2 => n5127, ZN => n5171);
   U17348 : NAND4_X1 port map( A1 => n1253, A2 => n5111, A3 => n5112, A4 => 
                           n5171, ZN => n5192);
   U17349 : NAND2_X1 port map( A1 => n4948, A2 => n4947, ZN => n5174);
   U17350 : OAI21_X1 port map( B1 => n5168, B2 => n1813, A => n5174, ZN => 
                           n5110);
   U17351 : NAND2_X1 port map( A1 => n5110, A2 => n5112, ZN => n5190);
   U17352 : NAND2_X1 port map( A1 => n5105, A2 => n4949, ZN => n5189);
   U17353 : NAND4_X1 port map( A1 => n4950, A2 => n5192, A3 => n5190, A4 => 
                           n5189, ZN => n4951);
   U17354 : OAI221_X1 port map( B1 => n4953, B2 => n5191, C1 => n1579, C2 => 
                           n4952, A => n4951, ZN => n5096);
   U17355 : INV_X1 port map( A => n5096, ZN => n5102);
   U17356 : NAND2_X1 port map( A1 => n5100, A2 => n4954, ZN => n5097);
   U17357 : INV_X1 port map( A => n5097, ZN => n4956);
   U17358 : NAND2_X1 port map( A1 => n5099, A2 => n4955, ZN => n5094);
   U17359 : OAI21_X1 port map( B1 => n5102, B2 => n4956, A => n5094, ZN => 
                           n4957);
   U17360 : NAND3_X1 port map( A1 => n4961, A2 => n5075, A3 => n5076, ZN => 
                           n4962);
   U17361 : NAND3_X1 port map( A1 => n4964, A2 => n5068, A3 => n5061, ZN => 
                           n4965);
   U17362 : NAND3_X1 port map( A1 => n5029, A2 => n5028, A3 => n4970, ZN => 
                           n4971);
   U17363 : OAI21_X1 port map( B1 => n5020, B2 => n4976, A => n4975, ZN => 
                           n5015);
   U17364 : OAI21_X1 port map( B1 => n5012, B2 => n4977, A => n5015, ZN => 
                           n4996);
   U17365 : NAND3_X1 port map( A1 => n4998, A2 => n4997, A3 => n4996, ZN => 
                           n4978);
   U17366 : OAI211_X1 port map( C1 => n4987, C2 => n4979, A => n5000, B => 
                           n4978, ZN => n4980);
   U17367 : OAI21_X1 port map( B1 => n4988, B2 => n4981, A => n4980, ZN => 
                           n5231);
   U17368 : XOR2_X1 port map( A => n4982, B => n5231, Z => n4983);
   U17369 : INV_X1 port map( A => n6920, ZN => n8158);
   U17370 : XOR2_X1 port map( A => n8158, B => n2247, Z => n4986);
   U17371 : INV_X1 port map( A => n4985, ZN => n8166);
   U17372 : NAND2_X1 port map( A1 => n4986, A2 => n2220, ZN => n7312);
   U17373 : OAI22_X1 port map( A1 => n7923, A2 => n2223, B1 => n2220, B2 => 
                           n7289, ZN => n5304);
   U17374 : OAI22_X1 port map( A1 => n7283, A2 => n2222, B1 => n2220, B2 => 
                           n7923, ZN => n5302);
   U17375 : INV_X1 port map( A => n5302, ZN => n5341);
   U17376 : NAND2_X1 port map( A1 => n4990, A2 => n4989, ZN => n5007);
   U17377 : INV_X1 port map( A => n4991, ZN => n4992);
   U17378 : AOI21_X1 port map( B1 => n4993, B2 => n5007, A => n4992, ZN => 
                           n4994);
   U17379 : XOR2_X1 port map( A => n4995, B => n4994, Z => n5004);
   U17380 : INV_X1 port map( A => n4995, ZN => n5002);
   U17381 : NAND2_X1 port map( A1 => n4997, A2 => n4996, ZN => n5008);
   U17382 : INV_X1 port map( A => n4998, ZN => n4999);
   U17383 : AOI21_X1 port map( B1 => n5000, B2 => n5008, A => n4999, ZN => 
                           n5001);
   U17384 : XOR2_X1 port map( A => n5002, B => n5001, Z => n5003);
   U17385 : MUX2_X1 port map( A => n5004, B => n5003, S => n2249, Z => n5342);
   U17386 : INV_X1 port map( A => n5342, ZN => n5303);
   U17387 : NAND2_X1 port map( A1 => n5341, A2 => n5303, ZN => n5338);
   U17388 : XOR2_X1 port map( A => n5009, B => n5008, Z => n5010);
   U17389 : OAI22_X1 port map( A1 => n2179, A2 => n2222, B1 => n2220, B2 => 
                           n7283, ZN => n5299);
   U17390 : INV_X1 port map( A => n5349, ZN => n5298);
   U17391 : XOR2_X1 port map( A => n5016, B => n5015, Z => n5017);
   U17392 : OAI22_X1 port map( A1 => n2178, A2 => n2222, B1 => n2220, B2 => 
                           n2179, ZN => n5296);
   U17393 : INV_X1 port map( A => n5296, ZN => n5356);
   U17394 : INV_X1 port map( A => n5357, ZN => n5297);
   U17395 : XOR2_X1 port map( A => n5023, B => n635, Z => n5024);
   U17396 : OAI22_X1 port map( A1 => n2176, A2 => n2222, B1 => n2220, B2 => 
                           n2178, ZN => n5364);
   U17397 : NAND2_X1 port map( A1 => n5365, A2 => n5364, ZN => n5206);
   U17398 : INV_X1 port map( A => n5206, ZN => n5208);
   U17399 : OAI22_X1 port map( A1 => n2213, A2 => n2222, B1 => n2220, B2 => 
                           n2175, ZN => n5292);
   U17400 : INV_X1 port map( A => n5292, ZN => n5373);
   U17401 : INV_X1 port map( A => n5027, ZN => n5036);
   U17402 : INV_X1 port map( A => n5030, ZN => n5034);
   U17403 : INV_X1 port map( A => n5031, ZN => n5032);
   U17404 : NOR2_X1 port map( A1 => n5032, A2 => n2249, ZN => n5033);
   U17405 : OAI33_X1 port map( A1 => n622, A2 => n5036, A3 => n2249, B1 => 
                           n5035, B2 => n5034, B3 => n5033, ZN => n5040);
   U17406 : INV_X1 port map( A => n5037, ZN => n5039);
   U17407 : NAND2_X1 port map( A1 => n1370, A2 => n5373, ZN => n5367);
   U17408 : NAND2_X1 port map( A1 => n5374, A2 => n5292, ZN => n5369);
   U17409 : OAI22_X1 port map( A1 => n2215, A2 => n2222, B1 => n2220, B2 => 
                           n2213, ZN => n5289);
   U17410 : INV_X1 port map( A => n5289, ZN => n5379);
   U17411 : INV_X1 port map( A => n778, ZN => n5290);
   U17412 : XOR2_X1 port map( A => n5048, B => n5049, Z => n5050);
   U17413 : OAI22_X1 port map( A1 => n2204, A2 => n2222, B1 => n2220, B2 => 
                           n2215, ZN => n5269);
   U17414 : NAND2_X1 port map( A1 => n5386, A2 => n5269, ZN => n5202);
   U17415 : INV_X1 port map( A => n5202, ZN => n5204);
   U17416 : OAI22_X1 port map( A1 => n2208, A2 => n2222, B1 => n2220, B2 => 
                           n2205, ZN => n5270);
   U17417 : INV_X1 port map( A => n5270, ZN => n5401);
   U17418 : INV_X1 port map( A => n5054, ZN => n5055);
   U17419 : AOI21_X1 port map( B1 => n485, B2 => n5056, A => n5055, ZN => n5057
                           );
   U17420 : XOR2_X1 port map( A => n5057, B => n5058, Z => n5064);
   U17421 : INV_X1 port map( A => n5059, ZN => n5060);
   U17422 : AOI21_X1 port map( B1 => n5061, B2 => n847, A => n5060, ZN => n5062
                           );
   U17423 : INV_X1 port map( A => n5397, ZN => n5400);
   U17424 : NAND2_X1 port map( A1 => n5401, A2 => n5400, ZN => n5391);
   U17425 : NAND2_X1 port map( A1 => n17214, A2 => n5270, ZN => n5393);
   U17427 : OAI22_X1 port map( A1 => n2196, A2 => n2222, B1 => n2220, B2 => 
                           n2209, ZN => n5284);
   U17428 : INV_X1 port map( A => n5284, ZN => n5498);
   U17429 : INV_X1 port map( A => n5499, ZN => n5285);
   U17430 : INV_X1 port map( A => n5076, ZN => n5078);
   U17431 : OAI21_X1 port map( B1 => n1337, B2 => n5078, A => n5077, ZN => 
                           n5080);
   U17432 : INV_X1 port map( A => n5405, ZN => n5417);
   U17433 : OAI22_X1 port map( A1 => n2200, A2 => n2222, B1 => n2220, B2 => 
                           n2197, ZN => n5282);
   U17434 : NAND2_X1 port map( A1 => n5417, A2 => n5282, ZN => n5513);
   U17435 : INV_X1 port map( A => n5282, ZN => n5418);
   U17436 : NAND2_X1 port map( A1 => n5418, A2 => n5405, ZN => n5510);
   U17437 : OAI22_X1 port map( A1 => n17240, A2 => n2222, B1 => n2219, B2 => 
                           n2200, ZN => n5281);
   U17438 : INV_X1 port map( A => n5422, ZN => n5425);
   U17439 : NAND2_X1 port map( A1 => n5426, A2 => n5425, ZN => n5508);
   U17440 : NAND2_X1 port map( A1 => n5422, A2 => n5281, ZN => n5414);
   U17441 : INV_X1 port map( A => n5094, ZN => n5095);
   U17442 : AOI21_X1 port map( B1 => n5097, B2 => n1379, A => n5095, ZN => 
                           n5098);
   U17443 : OAI22_X1 port map( A1 => n2238, A2 => n2222, B1 => n2219, B2 => 
                           n17240, ZN => n5431);
   U17444 : INV_X1 port map( A => n5431, ZN => n5199);
   U17445 : NAND2_X1 port map( A1 => n1822, A2 => n5199, ZN => n5413);
   U17446 : OAI22_X1 port map( A1 => n2138, A2 => n2221, B1 => n2219, B2 => 
                           n2238, ZN => n5437);
   U17447 : NAND2_X1 port map( A1 => n5437, A2 => n5436, ZN => n5433);
   U17448 : INV_X1 port map( A => n5184, ZN => n5106);
   U17449 : AOI21_X1 port map( B1 => n821, B2 => n5108, A => n5106, ZN => n5109
                           );
   U17450 : INV_X1 port map( A => n5110, ZN => n5115);
   U17451 : NAND3_X1 port map( A1 => n1350, A2 => n5171, A3 => n5111, ZN => 
                           n5114);
   U17452 : INV_X1 port map( A => n5112, ZN => n5113);
   U17453 : AOI21_X1 port map( B1 => n5115, B2 => n5114, A => n5113, ZN => 
                           n5118);
   U17454 : INV_X1 port map( A => n552, ZN => n5489);
   U17455 : OAI22_X1 port map( A1 => n2227, A2 => n2221, B1 => n2219, B2 => 
                           n2240, ZN => n5490);
   U17456 : INV_X1 port map( A => n5490, ZN => n5279);
   U17457 : NAND2_X1 port map( A1 => n5489, A2 => n5279, ZN => n5442);
   U17458 : INV_X1 port map( A => n5149, ZN => n5121);
   U17459 : NAND3_X1 port map( A1 => n5147, A2 => n828, A3 => n5146, ZN => 
                           n5125);
   U17460 : NAND3_X1 port map( A1 => n5129, A2 => n5156, A3 => n802, ZN => 
                           n5130);
   U17461 : OAI22_X1 port map( A1 => n2147, A2 => n2221, B1 => n2229, B2 => 
                           n2219, ZN => n5274);
   U17462 : NAND2_X1 port map( A1 => n5458, A2 => n5274, ZN => n5472);
   U17463 : INV_X1 port map( A => n5472, ZN => n5179);
   U17464 : OAI22_X1 port map( A1 => n2132, A2 => n2221, B1 => n2147, B2 => 
                           n2219, ZN => n5460);
   U17465 : INV_X1 port map( A => n5460, ZN => n8150);
   U17466 : NAND2_X1 port map( A1 => n1899, A2 => n2154, ZN => n8152);
   U17467 : INV_X1 port map( A => n8152, ZN => n8165);
   U17468 : NAND2_X1 port map( A1 => n8171, A2 => n1358, ZN => n5137);
   U17469 : AOI21_X1 port map( B1 => n1237, B2 => n5137, A => n1539, ZN => 
                           n5138);
   U17470 : XOR2_X1 port map( A => n5138, B => n5139, Z => n5143);
   U17471 : OAI21_X1 port map( B1 => n8171, B2 => n832, A => n8179, ZN => n5154
                           );
   U17472 : NAND2_X1 port map( A1 => n8164, A2 => n8165, ZN => n8163);
   U17473 : NAND3_X1 port map( A1 => n5154, A2 => n5155, A3 => n5153, ZN => 
                           n5157);
   U17474 : INV_X1 port map( A => n8151, ZN => n5273);
   U17475 : AOI21_X1 port map( B1 => n5167, B2 => n5166, A => n894, ZN => n5170
                           );
   U17476 : INV_X1 port map( A => n802, ZN => n5172);
   U17477 : OAI211_X1 port map( C1 => n5172, C2 => n1162, A => n1350, B => 
                           n5171, ZN => n5173);
   U17478 : NAND2_X1 port map( A1 => n5173, A2 => n1042, ZN => n5175);
   U17479 : OAI22_X1 port map( A1 => n2229, A2 => n2221, B1 => n2219, B2 => 
                           n2227, ZN => n5465);
   U17480 : INV_X1 port map( A => n5458, ZN => n5275);
   U17481 : INV_X1 port map( A => n5274, ZN => n5457);
   U17482 : NAND2_X1 port map( A1 => n1530, A2 => n5457, ZN => n5471);
   U17483 : OAI221_X1 port map( B1 => n5179, B2 => n5178, C1 => n678, C2 => 
                           n5465, A => n5471, ZN => n5180);
   U17484 : NAND2_X1 port map( A1 => n5276, A2 => n5465, ZN => n5485);
   U17485 : OAI211_X1 port map( C1 => n5489, C2 => n5279, A => n5485, B => 
                           n5180, ZN => n5441);
   U17486 : OAI22_X1 port map( A1 => n2240, A2 => n2221, B1 => n2219, B2 => 
                           n2239, ZN => n5453);
   U17487 : INV_X1 port map( A => n5181, ZN => n5185);
   U17488 : OAI221_X1 port map( B1 => n5185, B2 => n5184, C1 => n1227, C2 => 
                           n5185, A => n5182, ZN => n5188);
   U17489 : XOR2_X1 port map( A => n5188, B => n1821, Z => n5196);
   U17490 : AOI21_X1 port map( B1 => n5193, B2 => n5192, A => n17225, ZN => 
                           n5194);
   U17491 : XOR2_X1 port map( A => n5194, B => n1821, Z => n5195);
   U17492 : NAND2_X1 port map( A1 => n17259, A2 => n5453, ZN => n5443);
   U17493 : INV_X1 port map( A => n5443, ZN => n5198);
   U17495 : OAI221_X1 port map( B1 => n5437, B2 => n5436, C1 => n1773, C2 => 
                           n5198, A => n5440, ZN => n5432);
   U17496 : OAI211_X1 port map( C1 => n5199, C2 => n1822, A => n5433, B => 
                           n5432, ZN => n5412);
   U17497 : NAND2_X1 port map( A1 => n5412, A2 => n5413, ZN => n5424);
   U17498 : NAND2_X1 port map( A1 => n5424, A2 => n5414, ZN => n5509);
   U17499 : NAND3_X1 port map( A1 => n5509, A2 => n5508, A3 => n5510, ZN => 
                           n5200);
   U17500 : OAI211_X1 port map( C1 => n5498, C2 => n5285, A => n5200, B => 
                           n5513, ZN => n5201);
   U17501 : NAND3_X1 port map( A1 => n5399, A2 => n5202, A3 => n5393, ZN => 
                           n5203);
   U17502 : OAI21_X1 port map( B1 => n5379, B2 => n5290, A => n5381, ZN => 
                           n5205);
   U17503 : NAND3_X1 port map( A1 => n707, A2 => n5206, A3 => n5369, ZN => 
                           n5207);
   U17504 : OAI21_X1 port map( B1 => n5356, B2 => n5297, A => n5360, ZN => 
                           n5209);
   U17505 : INV_X1 port map( A => n5304, ZN => n5333);
   U17506 : INV_X1 port map( A => n5334, ZN => n5305);
   U17507 : NAND2_X1 port map( A1 => n5333, A2 => n5305, ZN => n5784);
   U17508 : OAI221_X1 port map( B1 => n1883, B2 => n5338, C1 => n1883, C2 => 
                           n5337, A => n5784, ZN => n5211);
   U17509 : INV_X1 port map( A => n5211, ZN => n5327);
   U17510 : OAI22_X1 port map( A1 => n7294, A2 => n2225, B1 => n2224, B2 => 
                           n7792, ZN => n5266);
   U17511 : OAI22_X1 port map( A1 => n7302, A2 => n2142, B1 => n2190, B2 => 
                           n8094, ZN => n5255);
   U17512 : NAND2_X1 port map( A1 => n5214, A2 => n2260, ZN => n5213);
   U17513 : OAI22_X1 port map( A1 => n7311, A2 => n2136, B1 => n2269, B2 => 
                           n7670, ZN => n5212);
   U17514 : INV_X1 port map( A => n5212, ZN => n5215);
   U17515 : MUX2_X1 port map( A => n5213, B => n2261, S => n5215, Z => n5217);
   U17516 : INV_X1 port map( A => n5214, ZN => n5216);
   U17517 : NAND2_X1 port map( A1 => n5216, A2 => n5215, ZN => n5244);
   U17518 : NAND2_X1 port map( A1 => n5217, A2 => n5244, ZN => n5254);
   U17519 : INV_X1 port map( A => n5254, ZN => n5252);
   U17521 : INV_X1 port map( A => n5225, ZN => n5221);
   U17522 : OAI21_X1 port map( B1 => n5222, B2 => n5221, A => n5220, ZN => 
                           n5223);
   U17523 : XOR2_X1 port map( A => n5250, B => n5226, Z => n5227);
   U17524 : INV_X1 port map( A => n5265, ZN => n5263);
   U17525 : INV_X1 port map( A => n5236, ZN => n5232);
   U17526 : OAI21_X1 port map( B1 => n5232, B2 => n5235, A => n5230, ZN => 
                           n5259);
   U17527 : OAI21_X1 port map( B1 => n5233, B2 => n5232, A => n5231, ZN => 
                           n5234);
   U17528 : OAI21_X1 port map( B1 => n5236, B2 => n5235, A => n5234, ZN => 
                           n5261);
   U17529 : XOR2_X1 port map( A => n5237, B => n5261, Z => n5238);
   U17530 : OAI22_X1 port map( A1 => n7289, A2 => n2221, B1 => n2219, B2 => 
                           n7864, ZN => n5306);
   U17531 : NAND2_X1 port map( A1 => n5326, A2 => n5306, ZN => n5786);
   U17532 : INV_X1 port map( A => n5786, ZN => n5240);
   U17533 : INV_X1 port map( A => n5326, ZN => n5330);
   U17534 : INV_X1 port map( A => n5306, ZN => n5328);
   U17535 : NAND2_X1 port map( A1 => n906, A2 => n5328, ZN => n5783);
   U17536 : OAI21_X1 port map( B1 => n5327, B2 => n5240, A => n5783, ZN => 
                           n5241);
   U17537 : OAI22_X1 port map( A1 => n7864, A2 => n2221, B1 => n2219, B2 => 
                           n7294, ZN => n5791);
   U17538 : INV_X1 port map( A => n5791, ZN => n5787);
   U17539 : OAI22_X1 port map( A1 => n7792, A2 => n2226, B1 => n2224, B2 => 
                           n7302, ZN => n5774);
   U17540 : OAI22_X1 port map( A1 => n8094, A2 => n2142, B1 => n2188, B2 => 
                           n7311, ZN => n5763);
   U17541 : NAND2_X1 port map( A1 => n5244, A2 => n2260, ZN => n5243);
   U17542 : OAI22_X1 port map( A1 => n7670, A2 => n2136, B1 => n2269, B2 => 
                           n7315, ZN => n5242);
   U17543 : INV_X1 port map( A => n5242, ZN => n5245);
   U17544 : MUX2_X1 port map( A => n5243, B => n2261, S => n5245, Z => n5247);
   U17545 : INV_X1 port map( A => n5244, ZN => n5246);
   U17546 : NAND2_X1 port map( A1 => n5246, A2 => n5245, ZN => n5752);
   U17547 : NAND2_X1 port map( A1 => n5247, A2 => n5752, ZN => n5762);
   U17548 : INV_X1 port map( A => n5762, ZN => n5760);
   U17549 : XOR2_X1 port map( A => n5763, B => n5760, Z => n5256);
   U17550 : INV_X1 port map( A => n5255, ZN => n5251);
   U17551 : XOR2_X1 port map( A => n5256, B => n5758, Z => n5257);
   U17552 : INV_X1 port map( A => n5773, ZN => n5771);
   U17553 : INV_X1 port map( A => n5266, ZN => n5262);
   U17554 : OAI21_X1 port map( B1 => n5263, B2 => n5262, A => n5261, ZN => 
                           n5264);
   U17555 : INV_X1 port map( A => n5790, ZN => n5788);
   U17556 : INV_X1 port map( A => n584, ZN => n5314);
   U17557 : NAND2_X1 port map( A1 => n5328, A2 => n5326, ZN => n5313);
   U17558 : NAND2_X1 port map( A1 => n5341, A2 => n5342, ZN => n5319);
   U17559 : INV_X1 port map( A => n5365, ZN => n5294);
   U17560 : INV_X1 port map( A => n5269, ZN => n5385);
   U17561 : NAND2_X1 port map( A1 => n5386, A2 => n5385, ZN => n5287);
   U17562 : NAND2_X1 port map( A1 => n5400, A2 => n5270, ZN => n5387);
   U17563 : NAND2_X1 port map( A1 => n5401, A2 => n17214, ZN => n5388);
   U17564 : NAND2_X1 port map( A1 => n5418, A2 => n5417, ZN => n5505);
   U17565 : NAND2_X1 port map( A1 => n5422, A2 => n5426, ZN => n5408);
   U17566 : NAND2_X1 port map( A1 => n1822, A2 => n5431, ZN => n5407);
   U17567 : INV_X1 port map( A => n5437, ZN => n5280);
   U17568 : NAND2_X1 port map( A1 => n1276, A2 => n5453, ZN => n5439);
   U17569 : NAND2_X1 port map( A1 => n1040, A2 => n5457, ZN => n5479);
   U17570 : INV_X1 port map( A => n8164, ZN => n5272);
   U17571 : NAND2_X1 port map( A1 => n943, A2 => n1790, ZN => n5468);
   U17572 : NAND2_X1 port map( A1 => n5273, A2 => n5460, ZN => n5466);
   U17573 : NAND4_X1 port map( A1 => n762, A2 => n5467, A3 => n5468, A4 => 
                           n5466, ZN => n5477);
   U17574 : INV_X1 port map( A => n5465, ZN => n5484);
   U17575 : NAND2_X1 port map( A1 => n5276, A2 => n5484, ZN => n5478);
   U17576 : NAND3_X1 port map( A1 => n5477, A2 => n5478, A3 => n5479, ZN => 
                           n5277);
   U17578 : NAND2_X1 port map( A1 => n17174, A2 => n5465, ZN => n5481);
   U17579 : NAND3_X1 port map( A1 => n5277, A2 => n5278, A3 => n5481, ZN => 
                           n5450);
   U17580 : NAND2_X1 port map( A1 => n657, A2 => n5279, ZN => n5449);
   U17581 : OAI211_X1 port map( C1 => n1276, C2 => n5453, A => n5450, B => 
                           n5449, ZN => n5438);
   U17582 : OAI211_X1 port map( C1 => n5280, C2 => n5436, A => n5438, B => 
                           n5439, ZN => n5430);
   U17583 : NAND2_X1 port map( A1 => n5280, A2 => n5436, ZN => n5429);
   U17584 : NAND2_X1 port map( A1 => n5406, A2 => n5407, ZN => n5423);
   U17585 : NAND2_X1 port map( A1 => n5423, A2 => n5408, ZN => n5501);
   U17586 : NAND2_X1 port map( A1 => n5425, A2 => n5281, ZN => n5500);
   U17587 : NAND2_X1 port map( A1 => n5405, A2 => n5282, ZN => n5502);
   U17588 : NAND3_X1 port map( A1 => n5501, A2 => n5500, A3 => n5502, ZN => 
                           n5283);
   U17589 : OAI211_X1 port map( C1 => n5285, C2 => n5284, A => n5283, B => 
                           n5505, ZN => n5286);
   U17590 : NAND3_X1 port map( A1 => n5398, A2 => n5287, A3 => n5388, ZN => 
                           n5288);
   U17592 : OAI21_X1 port map( B1 => n5290, B2 => n5289, A => n5380, ZN => 
                           n5291);
   U17593 : OAI22_X1 port map( A1 => n5294, A2 => n5364, B1 => n694, B2 => 
                           n1836, ZN => n5293);
   U17594 : INV_X1 port map( A => n5293, ZN => n5358);
   U17595 : OAI22_X1 port map( A1 => n5297, A2 => n5296, B1 => n5358, B2 => 
                           n1835, ZN => n5295);
   U17596 : INV_X1 port map( A => n5295, ZN => n5350);
   U17597 : NAND2_X1 port map( A1 => n5303, A2 => n5302, ZN => n5322);
   U17598 : INV_X1 port map( A => n5322, ZN => n5335);
   U17599 : NAND2_X1 port map( A1 => n5333, A2 => n5334, ZN => n5318);
   U17600 : OAI21_X1 port map( B1 => n1390, B2 => n5335, A => n5318, ZN => 
                           n5307);
   U17601 : NAND2_X1 port map( A1 => n5305, A2 => n5304, ZN => n5321);
   U17602 : NAND2_X1 port map( A1 => n5330, A2 => n5306, ZN => n5778);
   U17603 : NAND3_X1 port map( A1 => n5307, A2 => n5321, A3 => n5778, ZN => 
                           n5308);
   U17604 : INV_X1 port map( A => n5308, ZN => n5311);
   U17605 : INV_X1 port map( A => n5313, ZN => n5779);
   U17606 : NOR2_X1 port map( A1 => n5310, A2 => n5779, ZN => n5309);
   U17607 : AOI22_X1 port map( A1 => n5311, A2 => n5310, B1 => n5309, B2 => 
                           n5308, ZN => n5312);
   U17608 : OAI211_X1 port map( C1 => n5314, C2 => n5313, A => n6920, B => 
                           n5312, ZN => n5315);
   U17609 : INV_X1 port map( A => n6912, ZN => n8135);
   U17610 : XOR2_X1 port map( A => n2243, B => n2246, Z => n5317);
   U17611 : NAND2_X1 port map( A1 => n5317, A2 => n2218, ZN => n7303);
   U17612 : OAI22_X1 port map( A1 => n7923, A2 => n2180, B1 => n2218, B2 => 
                           n7289, ZN => n5796);
   U17613 : INV_X1 port map( A => n5796, ZN => n5800);
   U17614 : OAI22_X1 port map( A1 => n7283, A2 => n2180, B1 => n2218, B2 => 
                           n7923, ZN => n5526);
   U17615 : INV_X1 port map( A => n5318, ZN => n5323);
   U17616 : NAND3_X1 port map( A1 => n5343, A2 => n5319, A3 => n5318, ZN => 
                           n5320);
   U17617 : OAI211_X1 port map( C1 => n5323, C2 => n5322, A => n5321, B => 
                           n5320, ZN => n5324);
   U17618 : INV_X1 port map( A => n5324, ZN => n5780);
   U17619 : XOR2_X1 port map( A => n5325, B => n5326, Z => n5332);
   U17620 : XOR2_X1 port map( A => n5330, B => n5329, Z => n5331);
   U17621 : OAI22_X1 port map( A1 => n2179, A2 => n2181, B1 => n2218, B2 => 
                           n7283, ZN => n5567);
   U17622 : INV_X1 port map( A => n5567, ZN => n5569);
   U17623 : XOR2_X1 port map( A => n5334, B => n5333, Z => n5336);
   U17624 : INV_X1 port map( A => n5570, ZN => n5572);
   U17625 : OAI22_X1 port map( A1 => n2177, A2 => n2181, B1 => n2218, B2 => 
                           n2179, ZN => n5523);
   U17626 : XOR2_X1 port map( A => n5342, B => n5341, Z => n5345);
   U17627 : XOR2_X1 port map( A => n5345, B => n5344, Z => n5346);
   U17628 : INV_X1 port map( A => n5579, ZN => n5587);
   U17629 : OAI22_X1 port map( A1 => n2175, A2 => n2180, B1 => n2218, B2 => 
                           n2177, ZN => n5521);
   U17630 : INV_X1 port map( A => n5521, ZN => n5592);
   U17631 : NOR2_X1 port map( A1 => n5350, A2 => n1837, ZN => n5351);
   U17632 : XOR2_X1 port map( A => n5351, B => n5352, Z => n5355);
   U17633 : NAND2_X1 port map( A1 => n5592, A2 => n5593, ZN => n5584);
   U17634 : XOR2_X1 port map( A => n5357, B => n5356, Z => n5359);
   U17636 : INV_X1 port map( A => n5600, ZN => n5551);
   U17637 : OAI22_X1 port map( A1 => n2213, A2 => n2180, B1 => n2218, B2 => 
                           n2175, ZN => n5553);
   U17638 : NAND2_X1 port map( A1 => n5551, A2 => n5553, ZN => n5581);
   U17639 : INV_X1 port map( A => n5549, ZN => n5608);
   U17640 : INV_X1 port map( A => n5367, ZN => n5368);
   U17641 : AOI21_X1 port map( B1 => n5369, B2 => n707, A => n5368, ZN => n5370
                           );
   U17642 : INV_X1 port map( A => n5609, ZN => n5528);
   U17643 : OAI22_X1 port map( A1 => n2204, A2 => n2181, B1 => n2218, B2 => 
                           n2215, ZN => n5529);
   U17644 : INV_X1 port map( A => n5529, ZN => n5624);
   U17645 : XOR2_X1 port map( A => n5374, B => n5373, Z => n5376);
   U17646 : XOR2_X1 port map( A => n5376, B => n5375, Z => n5377);
   U17647 : INV_X1 port map( A => n5617, ZN => n5623);
   U17648 : OAI22_X1 port map( A1 => n2208, A2 => n2180, B1 => n2218, B2 => 
                           n2205, ZN => n5548);
   U17649 : INV_X1 port map( A => n5548, ZN => n5633);
   U17650 : XOR2_X1 port map( A => n5382, B => n505, Z => n5383);
   U17651 : NAND2_X1 port map( A1 => n5633, A2 => n664, ZN => n5621);
   U17652 : XOR2_X1 port map( A => n5386, B => n5385, Z => n5390);
   U17653 : XOR2_X1 port map( A => n5389, B => n5390, Z => n5396);
   U17654 : INV_X1 port map( A => n5391, ZN => n5392);
   U17655 : AOI21_X1 port map( B1 => n5393, B2 => n5399, A => n5392, ZN => 
                           n5394);
   U17656 : INV_X1 port map( A => n706, ZN => n5544);
   U17657 : OAI22_X1 port map( A1 => n2196, A2 => n2180, B1 => n2218, B2 => 
                           n2209, ZN => n5546);
   U17658 : NAND2_X1 port map( A1 => n5544, A2 => n5546, ZN => n5630);
   U17659 : OAI22_X1 port map( A1 => n2199, A2 => n2181, B1 => n2217, B2 => 
                           n2197, ZN => n5530);
   U17660 : INV_X1 port map( A => n5530, ZN => n5734);
   U17661 : NAND2_X1 port map( A1 => n5734, A2 => n929, ZN => n5641);
   U17662 : INV_X1 port map( A => n5408, ZN => n5409);
   U17663 : AOI21_X1 port map( B1 => n5410, B2 => n5500, A => n5409, ZN => 
                           n5411);
   U17664 : INV_X1 port map( A => n5414, ZN => n5415);
   U17665 : AOI21_X1 port map( B1 => n5508, B2 => n5416, A => n5415, ZN => 
                           n5419);
   U17666 : INV_X1 port map( A => n726, ZN => n5652);
   U17667 : OAI22_X1 port map( A1 => n2238, A2 => n2181, B1 => n2217, B2 => 
                           n17240, ZN => n5658);
   U17668 : OAI22_X1 port map( A1 => n2138, A2 => n2180, B1 => n2217, B2 => 
                           n2238, ZN => n5664);
   U17669 : INV_X1 port map( A => n5664, ZN => n5671);
   U17670 : OAI22_X1 port map( A1 => n2240, A2 => n2180, B1 => n2217, B2 => 
                           n2239, ZN => n5673);
   U17671 : NAND2_X1 port map( A1 => n689, A2 => n5673, ZN => n5666);
   U17672 : OAI22_X1 port map( A1 => n2227, A2 => n2181, B1 => n2217, B2 => 
                           n2240, ZN => n5537);
   U17673 : NAND3_X1 port map( A1 => n5441, A2 => n5442, A3 => n5440, ZN => 
                           n5444);
   U17674 : NAND2_X1 port map( A1 => n5444, A2 => n5443, ZN => n5446);
   U17675 : INV_X1 port map( A => n1157, ZN => n5535);
   U17676 : OAI22_X1 port map( A1 => n2229, A2 => n2181, B1 => n2217, B2 => 
                           n2227, ZN => n5683);
   U17677 : INV_X1 port map( A => n5683, ZN => n5696);
   U17678 : OAI22_X1 port map( A1 => n771, A2 => n2180, B1 => n2147, B2 => 
                           n2218, ZN => n5456);
   U17679 : INV_X1 port map( A => n5456, ZN => n8128);
   U17680 : NAND3_X1 port map( A1 => n5467, A2 => n5468, A3 => n5466, ZN => 
                           n5459);
   U17682 : OAI21_X1 port map( B1 => n8154, B2 => n5460, A => n503, ZN => n5473
                           );
   U17683 : XOR2_X1 port map( A => n5461, B => n1139, Z => n5462);
   U17684 : INV_X1 port map( A => n17169, ZN => n5464);
   U17685 : NAND3_X1 port map( A1 => n5467, A2 => n898, A3 => n5466, ZN => 
                           n5469);
   U17686 : AOI21_X1 port map( B1 => n5479, B2 => n5469, A => n1221, ZN => 
                           n5470);
   U17687 : OAI22_X1 port map( A1 => n2147, A2 => n2180, B1 => n2217, B2 => 
                           n2230, ZN => n5707);
   U17688 : INV_X1 port map( A => n5707, ZN => n5533);
   U17689 : NAND3_X1 port map( A1 => n1048, A2 => n5478, A3 => n5479, ZN => 
                           n5480);
   U17690 : NAND2_X1 port map( A1 => n942, A2 => n5533, ZN => n5693);
   U17691 : INV_X1 port map( A => n5693, ZN => n5680);
   U17692 : INV_X1 port map( A => n5698, ZN => n5706);
   U17693 : NAND2_X1 port map( A1 => n5706, A2 => n5707, ZN => n5691);
   U17694 : OAI221_X1 port map( B1 => n5694, B2 => n5696, C1 => n1216, C2 => 
                           n5680, A => n5691, ZN => n5495);
   U17695 : OAI211_X1 port map( C1 => n5671, C2 => n790, A => n5665, B => n5666
                           , ZN => n5653);
   U17696 : NAND2_X1 port map( A1 => n790, A2 => n5671, ZN => n5654);
   U17697 : OAI211_X1 port map( C1 => n5652, C2 => n5658, A => n5653, B => 
                           n5654, ZN => n5497);
   U17698 : INV_X1 port map( A => n5497, ZN => n5728);
   U17699 : OAI22_X1 port map( A1 => n17240, A2 => n2181, B1 => n2217, B2 => 
                           n2200, ZN => n5540);
   U17700 : INV_X1 port map( A => n5540, ZN => n5722);
   U17701 : XOR2_X1 port map( A => n5499, B => n5498, Z => n5507);
   U17702 : NAND2_X1 port map( A1 => n1318, A2 => n5500, ZN => n5504);
   U17703 : INV_X1 port map( A => n5502, ZN => n5503);
   U17704 : AOI21_X1 port map( B1 => n5504, B2 => n5505, A => n5503, ZN => 
                           n5506);
   U17705 : XOR2_X1 port map( A => n5506, B => n5507, Z => n5516);
   U17706 : NAND2_X1 port map( A1 => n5509, A2 => n5508, ZN => n5512);
   U17707 : INV_X1 port map( A => n5510, ZN => n5511);
   U17708 : AOI21_X1 port map( B1 => n5513, B2 => n5512, A => n5511, ZN => 
                           n5514);
   U17709 : NAND2_X1 port map( A1 => n5723, A2 => n5722, ZN => n5729);
   U17710 : OAI21_X1 port map( B1 => n1807, B2 => n5728, A => n5729, ZN => 
                           n5639);
   U17711 : INV_X1 port map( A => n601, ZN => n5541);
   U17712 : NAND2_X1 port map( A1 => n476, A2 => n5540, ZN => n5731);
   U17713 : NAND3_X1 port map( A1 => n5639, A2 => n5731, A3 => n5640, ZN => 
                           n5517);
   U17714 : OAI211_X1 port map( C1 => n5544, C2 => n5546, A => n5641, B => 
                           n5517, ZN => n5629);
   U17715 : INV_X1 port map( A => n5628, ZN => n5632);
   U17716 : NAND2_X1 port map( A1 => n5632, A2 => n5548, ZN => n5618);
   U17717 : NAND3_X1 port map( A1 => n17227, A2 => n5630, A3 => n5618, ZN => 
                           n5518);
   U17718 : OAI211_X1 port map( C1 => n5623, C2 => n5529, A => n5621, B => 
                           n5518, ZN => n5519);
   U17719 : NAND2_X1 port map( A1 => n1647, A2 => n5521, ZN => n5582);
   U17720 : NAND3_X1 port map( A1 => n5581, A2 => n5580, A3 => n5582, ZN => 
                           n5522);
   U17721 : OAI211_X1 port map( C1 => n5587, C2 => n5523, A => n5584, B => 
                           n5522, ZN => n5524);
   U17722 : OAI21_X1 port map( B1 => n5567, B2 => n5572, A => n5566, ZN => 
                           n5525);
   U17723 : OAI21_X1 port map( B1 => n683, B2 => n5526, A => n5560, ZN => n5527
                           );
   U17724 : INV_X1 port map( A => n5553, ZN => n5599);
   U17725 : NAND2_X1 port map( A1 => n5617, A2 => n5529, ZN => n5611);
   U17726 : INV_X1 port map( A => n5546, ZN => n5637);
   U17727 : NAND2_X1 port map( A1 => n929, A2 => n5530, ZN => n5647);
   U17728 : INV_X1 port map( A => n5658, ZN => n5538);
   U17729 : NAND2_X1 port map( A1 => n5664, A2 => n790, ZN => n5659);
   U17730 : INV_X1 port map( A => n5673, ZN => n5675);
   U17731 : NAND2_X1 port map( A1 => n689, A2 => n5675, ZN => n5670);
   U17732 : NAND2_X1 port map( A1 => n1214, A2 => n5683, ZN => n5688);
   U17733 : INV_X1 port map( A => n663, ZN => n5531);
   U17734 : NAND2_X1 port map( A1 => n8142, A2 => n1872, ZN => n5532);
   U17735 : NAND2_X1 port map( A1 => n1428, A2 => n5532, ZN => n5710);
   U17736 : NAND2_X1 port map( A1 => n8128, A2 => n5532, ZN => n5711);
   U17737 : NAND2_X1 port map( A1 => n5706, A2 => n5533, ZN => n5699);
   U17738 : NAND2_X1 port map( A1 => n5697, A2 => n5696, ZN => n5686);
   U17739 : NAND3_X1 port map( A1 => n5685, A2 => n5686, A3 => n5699, ZN => 
                           n5534);
   U17740 : OAI211_X1 port map( C1 => n5664, C2 => n790, A => n5669, B => n5670
                           , ZN => n5660);
   U17741 : OAI211_X1 port map( C1 => n5652, C2 => n5538, A => n5660, B => 
                           n5659, ZN => n5539);
   U17742 : NAND2_X1 port map( A1 => n601, A2 => n5540, ZN => n5645);
   U17743 : INV_X1 port map( A => n5645, ZN => n5542);
   U17744 : NAND2_X1 port map( A1 => n5722, A2 => n5541, ZN => n5737);
   U17745 : OAI211_X1 port map( C1 => n5725, C2 => n5542, A => n5737, B => 
                           n5646, ZN => n5543);
   U17746 : OAI211_X1 port map( C1 => n5637, C2 => n5544, A => n5543, B => 
                           n5647, ZN => n5545);
   U17747 : NAND2_X1 port map( A1 => n1012, A2 => n5611, ZN => n5602);
   U17748 : AOI21_X1 port map( B1 => n5602, B2 => n5612, A => n1840, ZN => 
                           n5550);
   U17750 : OAI21_X1 port map( B1 => n5592, B2 => n1647, A => n5594, ZN => 
                           n5554);
   U17751 : INV_X1 port map( A => n5554, ZN => n5586);
   U17752 : OAI22_X1 port map( A1 => n5562, A2 => n683, B1 => n813, B2 => n1845
                           , ZN => n5798);
   U17753 : NAND2_X1 port map( A1 => n683, A2 => n5562, ZN => n5799);
   U17754 : INV_X1 port map( A => n6041, ZN => n5834);
   U17755 : INV_X1 port map( A => n6776, ZN => n8263);
   U17756 : XOR2_X1 port map( A => n2243, B => n2267, Z => n5558);
   U17757 : XOR2_X1 port map( A => n8270, B => n2243, Z => n7295);
   U17758 : NAND2_X1 port map( A1 => n5558, A2 => n2182, ZN => n7296);
   U17759 : OAI22_X1 port map( A1 => n2179, A2 => n2183, B1 => n2182, B2 => 
                           n7283, ZN => n5836);
   U17760 : NAND2_X1 port map( A1 => n5834, A2 => n5836, ZN => n6700);
   U17761 : INV_X1 port map( A => n6700, ZN => n5749);
   U17762 : INV_X1 port map( A => n5836, ZN => n6038);
   U17763 : NAND2_X1 port map( A1 => n6038, A2 => n6041, ZN => n5837);
   U17764 : INV_X1 port map( A => n5837, ZN => n5559);
   U17765 : NOR2_X1 port map( A1 => n5559, A2 => n2268, ZN => n5748);
   U17766 : INV_X1 port map( A => n5845, ZN => n5848);
   U17767 : NOR2_X1 port map( A1 => n1845, A2 => n17157, ZN => n5563);
   U17768 : NAND3_X1 port map( A1 => n5576, A2 => n233, A3 => n1809, ZN => 
                           n5575);
   U17769 : NOR2_X1 port map( A1 => n5567, A2 => n5568, ZN => n5573);
   U17770 : NOR2_X1 port map( A1 => n5569, A2 => n5568, ZN => n5571);
   U17771 : AOI221_X1 port map( B1 => n5572, B2 => n5573, C1 => n5571, C2 => 
                           n471, A => n6912, ZN => n5574);
   U17772 : INV_X1 port map( A => n5856, ZN => n5859);
   U17773 : OAI22_X1 port map( A1 => n2175, A2 => n2184, B1 => n2182, B2 => 
                           n2178, ZN => n5805);
   U17774 : OAI22_X1 port map( A1 => n2213, A2 => n2184, B1 => n2182, B2 => 
                           n2176, ZN => n5831);
   U17775 : INV_X1 port map( A => n5831, ZN => n5990);
   U17776 : INV_X1 port map( A => n5582, ZN => n5583);
   U17777 : AOI21_X1 port map( B1 => n5584, B2 => n1088, A => n5583, ZN => 
                           n5585);
   U17778 : NOR2_X1 port map( A1 => n5586, A2 => n1787, ZN => n5589);
   U17779 : INV_X1 port map( A => n5987, ZN => n5989);
   U17780 : OAI22_X1 port map( A1 => n2215, A2 => n2183, B1 => n2182, B2 => 
                           n2213, ZN => n5829);
   U17781 : INV_X1 port map( A => n951, ZN => n5867);
   U17782 : OAI22_X1 port map( A1 => n2204, A2 => n2183, B1 => n2182, B2 => 
                           n2215, ZN => n5827);
   U17783 : INV_X1 port map( A => n5827, ZN => n5878);
   U17784 : INV_X1 port map( A => n5612, ZN => n5601);
   U17785 : NOR2_X1 port map( A1 => n5601, A2 => n1791, ZN => n5603);
   U17786 : AOI21_X1 port map( B1 => n5603, B2 => n5602, A => n1840, ZN => 
                           n5604);
   U17787 : XOR2_X1 port map( A => n5605, B => n5604, Z => n5606);
   U17788 : INV_X1 port map( A => n1058, ZN => n5875);
   U17789 : INV_X1 port map( A => n5611, ZN => n5613);
   U17790 : OAI21_X1 port map( B1 => n1062, B2 => n5613, A => n5612, ZN => 
                           n5614);
   U17791 : XOR2_X1 port map( A => n1778, B => n5614, Z => n5615);
   U17792 : INV_X1 port map( A => n867, ZN => n5806);
   U17793 : OAI22_X1 port map( A1 => n2208, A2 => n2184, B1 => n2182, B2 => 
                           n2205, ZN => n5824);
   U17794 : NAND2_X1 port map( A1 => n5806, A2 => n5824, ZN => n5873);
   U17795 : INV_X1 port map( A => n5873, ZN => n5743);
   U17796 : NAND2_X1 port map( A1 => n17227, A2 => n5630, ZN => n5620);
   U17797 : INV_X1 port map( A => n5618, ZN => n5619);
   U17798 : AOI21_X1 port map( B1 => n5621, B2 => n5620, A => n5619, ZN => 
                           n5622);
   U17799 : INV_X1 port map( A => n5897, ZN => n5894);
   U17800 : OAI22_X1 port map( A1 => n2196, A2 => n2184, B1 => n2209, B2 => 
                           n2182, ZN => n5807);
   U17801 : NAND2_X1 port map( A1 => n1514, A2 => n5807, ZN => n5872);
   U17802 : OAI22_X1 port map( A1 => n2199, A2 => n2183, B1 => n2197, B2 => 
                           n2182, ZN => n5823);
   U17803 : INV_X1 port map( A => n5823, ZN => n5909);
   U17804 : NAND2_X1 port map( A1 => n5639, A2 => n5731, ZN => n5642);
   U17805 : AOI21_X1 port map( B1 => n5642, B2 => n5641, A => n460, ZN => n5643
                           );
   U17806 : NAND2_X1 port map( A1 => n5645, A2 => n5644, ZN => n5736);
   U17807 : NAND3_X1 port map( A1 => n5736, A2 => n5737, A3 => n957, ZN => 
                           n5648);
   U17808 : NAND2_X1 port map( A1 => n5648, A2 => n5647, ZN => n5649);
   U17809 : OAI22_X1 port map( A1 => n17239, A2 => n2183, B1 => n2200, B2 => 
                           n2182, ZN => n5808);
   U17810 : NAND2_X1 port map( A1 => n1433, A2 => n5808, ZN => n5904);
   U17811 : OAI22_X1 port map( A1 => n2240, A2 => n2184, B1 => n2239, B2 => 
                           n2182, ZN => n5925);
   U17812 : INV_X1 port map( A => n5925, ZN => n5927);
   U17813 : INV_X1 port map( A => n660, ZN => n5928);
   U17814 : OAI22_X1 port map( A1 => n2227, A2 => n2184, B1 => n2240, B2 => 
                           n2182, ZN => n5936);
   U17815 : INV_X1 port map( A => n5936, ZN => n5943);
   U17816 : OAI22_X1 port map( A1 => n2229, A2 => n2183, B1 => n2227, B2 => 
                           n2182, ZN => n5811);
   U17817 : NAND2_X1 port map( A1 => n5955, A2 => n1352, ZN => n5934);
   U17818 : OAI21_X1 port map( B1 => n5680, B2 => n1216, A => n5691, ZN => 
                           n5682);
   U17819 : AOI22_X1 port map( A1 => n5697, A2 => n5683, B1 => n5681, B2 => 
                           n5682, ZN => n5684);
   U17820 : NAND2_X1 port map( A1 => n5685, A2 => n5699, ZN => n5689);
   U17821 : INV_X1 port map( A => n5686, ZN => n5687);
   U17822 : OAI22_X1 port map( A1 => n2147, A2 => n2183, B1 => n2230, B2 => 
                           n2182, ZN => n5957);
   U17823 : INV_X1 port map( A => n5957, ZN => n5812);
   U17824 : NAND2_X1 port map( A1 => n5812, A2 => n972, ZN => n5950);
   U17825 : OAI22_X1 port map( A1 => n2132, A2 => n2184, B1 => n2147, B2 => 
                           n2182, ZN => n8258);
   U17826 : INV_X1 port map( A => n8258, ZN => n5813);
   U17827 : AOI21_X1 port map( B1 => n5693, B2 => n5692, A => n495, ZN => n5695
                           );
   U17828 : NAND2_X1 port map( A1 => n5707, A2 => n942, ZN => n5702);
   U17829 : NAND3_X1 port map( A1 => n5709, A2 => n5710, A3 => n5711, ZN => 
                           n5701);
   U17830 : INV_X1 port map( A => n5699, ZN => n5700);
   U17831 : INV_X1 port map( A => n5711, ZN => n5712);
   U17832 : NOR3_X1 port map( A1 => n1010, A2 => n775, A3 => n5712, ZN => n5713
                           );
   U17833 : INV_X1 port map( A => n8269, ZN => n5717);
   U17834 : INV_X1 port map( A => n7295, ZN => n5716);
   U17835 : OAI21_X1 port map( B1 => n8257, B2 => n8258, A => n1826, ZN => 
                           n5718);
   U17836 : NAND2_X1 port map( A1 => n5958, A2 => n5950, ZN => n5932);
   U17837 : NAND3_X1 port map( A1 => n5932, A2 => n5949, A3 => n5933, ZN => 
                           n5719);
   U17838 : OAI211_X1 port map( C1 => n5936, C2 => n456, A => n5719, B => n5934
                           , ZN => n5720);
   U17839 : INV_X1 port map( A => n5919, ZN => n5920);
   U17841 : NOR2_X1 port map( A1 => n5728, A2 => n1807, ZN => n5732);
   U17842 : INV_X1 port map( A => n5729, ZN => n5730);
   U17843 : AOI21_X1 port map( B1 => n5732, B2 => n5731, A => n5730, ZN => 
                           n5733);
   U17844 : OAI22_X1 port map( A1 => n2238, A2 => n2183, B1 => n17239, B2 => 
                           n2182, ZN => n5809);
   U17845 : NAND2_X1 port map( A1 => n5915, A2 => n5809, ZN => n5969);
   U17846 : INV_X1 port map( A => n5809, ZN => n5914);
   U17847 : INV_X1 port map( A => n17183, ZN => n5810);
   U17848 : NAND2_X1 port map( A1 => n5914, A2 => n5810, ZN => n5972);
   U17849 : OAI211_X1 port map( C1 => n5909, C2 => n5908, A => n5903, B => 
                           n5904, ZN => n5893);
   U17850 : NAND2_X1 port map( A1 => n5909, A2 => n5908, ZN => n5892);
   U17851 : INV_X1 port map( A => n5824, ZN => n5887);
   U17852 : AOI21_X1 port map( B1 => n5871, B2 => n5872, A => n1886, ZN => 
                           n5742);
   U17853 : OAI22_X1 port map( A1 => n5827, A2 => n5875, B1 => n5742, B2 => 
                           n5743, ZN => n5744);
   U17854 : OAI21_X1 port map( B1 => n1445, B2 => n5831, A => n5988, ZN => 
                           n5745);
   U17855 : OAI21_X1 port map( B1 => n5990, B2 => n1744, A => n5745, ZN => 
                           n5857);
   U17856 : INV_X1 port map( A => n5852, ZN => n5746);
   U17857 : INV_X1 port map( A => n5833, ZN => n5854);
   U17858 : OAI22_X1 port map( A1 => n5746, A2 => n1812, B1 => n5854, B2 => 
                           n5845, ZN => n5747);
   U17859 : AOI22_X1 port map( A1 => n5749, A2 => n6776, B1 => n5748, B2 => 
                           n6045, ZN => n5841);
   U17860 : OAI22_X1 port map( A1 => n7302, A2 => n2225, B1 => n2224, B2 => 
                           n8094, ZN => n6733);
   U17861 : OAI22_X1 port map( A1 => n7311, A2 => n2142, B1 => n2190, B2 => 
                           n7670, ZN => n6726);
   U17862 : NAND2_X1 port map( A1 => n5752, A2 => n2259, ZN => n5751);
   U17863 : MUX2_X1 port map( A => n278, B => n360, S => n2145, Z => n7607);
   U17864 : OAI22_X1 port map( A1 => n7315, A2 => n2137, B1 => n2269, B2 => 
                           n7607, ZN => n5750);
   U17865 : INV_X1 port map( A => n5750, ZN => n5753);
   U17866 : MUX2_X1 port map( A => n5751, B => n2261, S => n5753, Z => n5755);
   U17867 : INV_X1 port map( A => n5752, ZN => n5754);
   U17868 : NAND2_X1 port map( A1 => n5754, A2 => n5753, ZN => n6715);
   U17869 : NAND2_X1 port map( A1 => n5755, A2 => n6715, ZN => n6725);
   U17870 : INV_X1 port map( A => n6725, ZN => n6723);
   U17871 : XOR2_X1 port map( A => n6726, B => n6723, Z => n5764);
   U17872 : INV_X1 port map( A => n5763, ZN => n5759);
   U17873 : OAI21_X1 port map( B1 => n5759, B2 => n5762, A => n5757, ZN => 
                           n6719);
   U17874 : OAI21_X1 port map( B1 => n5763, B2 => n5762, A => n5761, ZN => 
                           n6721);
   U17875 : XOR2_X1 port map( A => n5764, B => n6721, Z => n5765);
   U17876 : INV_X1 port map( A => n6736, ZN => n6734);
   U17877 : INV_X1 port map( A => n5774, ZN => n5770);
   U17878 : OAI21_X1 port map( B1 => n5771, B2 => n5774, A => n5767, ZN => 
                           n5768);
   U17880 : OAI21_X1 port map( B1 => n5771, B2 => n5770, A => n5769, ZN => 
                           n5772);
   U17881 : XOR2_X1 port map( A => n5775, B => n6711, Z => n5776);
   U17882 : OAI21_X1 port map( B1 => n5780, B2 => n5779, A => n5778, ZN => 
                           n5781);
   U17883 : INV_X1 port map( A => n5781, ZN => n6708);
   U17884 : AOI21_X1 port map( B1 => n6708, B2 => n6707, A => n1842, ZN => 
                           n5782);
   U17885 : OAI22_X1 port map( A1 => n7294, A2 => n2221, B1 => n2219, B2 => 
                           n7792, ZN => n6710);
   U17886 : INV_X1 port map( A => n6710, ZN => n6747);
   U17887 : OAI211_X1 port map( C1 => n1780, C2 => n1883, A => n5784, B => 
                           n5783, ZN => n5785);
   U17888 : OAI211_X1 port map( C1 => n5788, C2 => n5787, A => n5786, B => 
                           n5785, ZN => n5789);
   U17889 : OAI21_X1 port map( B1 => n5791, B2 => n1109, A => n5789, ZN => 
                           n6745);
   U17890 : INV_X1 port map( A => n6706, ZN => n6746);
   U17891 : XOR2_X1 port map( A => n5792, B => n796, Z => n5793);
   U17892 : OAI22_X1 port map( A1 => n7289, A2 => n2181, B1 => n2217, B2 => 
                           n7864, ZN => n6705);
   U17893 : INV_X1 port map( A => n6705, ZN => n6755);
   U17894 : INV_X1 port map( A => n6704, ZN => n5803);
   U17895 : NAND2_X1 port map( A1 => n869, A2 => n5796, ZN => n6703);
   U17896 : NOR2_X1 port map( A1 => n6912, A2 => n1887, ZN => n5801);
   U17897 : NAND2_X1 port map( A1 => n5798, A2 => n5799, ZN => n6751);
   U17898 : AOI221_X1 port map( B1 => n6912, B2 => n6703, C1 => n6751, C2 => 
                           n5801, A => n1377, ZN => n5802);
   U17899 : AOI21_X1 port map( B1 => n5803, B2 => n6912, A => n5802, ZN => 
                           n5804);
   U17900 : OAI22_X1 port map( A1 => n7283, A2 => n2183, B1 => n2182, B2 => 
                           n7923, ZN => n6765);
   U17901 : NAND2_X1 port map( A1 => n5887, A2 => n5806, ZN => n5882);
   U17902 : INV_X1 port map( A => n5808, ZN => n5979);
   U17903 : NAND2_X1 port map( A1 => n5979, A2 => n5978, ZN => n5907);
   U17904 : NAND2_X1 port map( A1 => n5810, A2 => n5809, ZN => n5977);
   U17905 : NAND2_X1 port map( A1 => n1352, A2 => n5811, ZN => n5941);
   U17906 : NAND2_X1 port map( A1 => n1290, A2 => n5812, ZN => n5953);
   U17907 : NAND2_X1 port map( A1 => n5957, A2 => n784, ZN => n5954);
   U17908 : NAND2_X1 port map( A1 => n1893, A2 => n8269, ZN => n8268);
   U17909 : OAI21_X1 port map( B1 => n1431, B2 => n5813, A => n8268, ZN => 
                           n5814);
   U17910 : NAND2_X1 port map( A1 => n5959, A2 => n5954, ZN => n5939);
   U17911 : NAND3_X1 port map( A1 => n5939, A2 => n5953, A3 => n5940, ZN => 
                           n5816);
   U17912 : OAI211_X1 port map( C1 => n5943, C2 => n456, A => n5816, B => n5941
                           , ZN => n5817);
   U17913 : NAND2_X1 port map( A1 => n5915, A2 => n5914, ZN => n5974);
   U17914 : OAI211_X1 port map( C1 => n648, C2 => n1834, A => n690, B => n5974,
                           ZN => n5822);
   U17915 : OAI211_X1 port map( C1 => n5979, C2 => n5978, A => n5977, B => 
                           n5822, ZN => n5906);
   U17916 : OAI211_X1 port map( C1 => n620, C2 => n5823, A => n5906, B => n5907
                           , ZN => n5899);
   U17917 : NAND2_X1 port map( A1 => n620, A2 => n5823, ZN => n5898);
   U17918 : OAI211_X1 port map( C1 => n5896, C2 => n5894, A => n5899, B => 
                           n5898, ZN => n5880);
   U17919 : AOI21_X1 port map( B1 => n5880, B2 => n5881, A => n1885, ZN => 
                           n5825);
   U17920 : OAI22_X1 port map( A1 => n17158, A2 => n5878, B1 => n5825, B2 => 
                           n865, ZN => n5826);
   U17921 : OAI22_X1 port map( A1 => n1816, A2 => n895, B1 => n5854, B2 => 
                           n5848, ZN => n5832);
   U17922 : OAI21_X1 port map( B1 => n6038, B2 => n5834, A => n5843, ZN => 
                           n5835);
   U17923 : NAND2_X1 port map( A1 => n5837, A2 => n6045, ZN => n6701);
   U17924 : NAND4_X1 port map( A1 => n6776, A2 => n6700, A3 => n6701, A4 => 
                           n5840, ZN => n5838);
   U17926 : INV_X1 port map( A => n6967, ZN => n8245);
   U17927 : XOR2_X1 port map( A => n2267, B => n2265, Z => n5842);
   U17928 : XOR2_X1 port map( A => n8250, B => n2267, Z => n7290);
   U17929 : NAND2_X1 port map( A1 => n5842, A2 => n2185, ZN => n7291);
   U17930 : OAI22_X1 port map( A1 => n2177, A2 => n7291, B1 => n2185, B2 => 
                           n2179, ZN => n6784);
   U17931 : INV_X1 port map( A => n6784, ZN => n6783);
   U17932 : OAI22_X1 port map( A1 => n2176, A2 => n7291, B1 => n2185, B2 => 
                           n2177, ZN => n6031);
   U17933 : INV_X1 port map( A => n6031, ZN => n6039);
   U17934 : INV_X1 port map( A => n1081, ZN => n6044);
   U17935 : INV_X1 port map( A => n5843, ZN => n6042);
   U17936 : OAI22_X1 port map( A1 => n2213, A2 => n7291, B1 => n2185, B2 => 
                           n2176, ZN => n6057);
   U17937 : INV_X1 port map( A => n6057, ZN => n6060);
   U17938 : NAND2_X1 port map( A1 => n5848, A2 => n6776, ZN => n5853);
   U17939 : INV_X1 port map( A => n5853, ZN => n5847);
   U17940 : NOR3_X1 port map( A1 => n1812, A2 => n5848, A3 => n2268, ZN => 
                           n5849);
   U17941 : AOI22_X1 port map( A1 => n895, A2 => n1858, B1 => n5849, B2 => 
                           n5852, ZN => n5850);
   U17942 : OAI211_X1 port map( C1 => n5853, C2 => n5852, A => n5851, B => 
                           n5850, ZN => n5855);
   U17943 : INV_X1 port map( A => n930, ZN => n5861);
   U17944 : OAI22_X1 port map( A1 => n2215, A2 => n7291, B1 => n2185, B2 => 
                           n2213, ZN => n6079);
   U17945 : OAI22_X1 port map( A1 => n2208, A2 => n7291, B1 => n2205, B2 => 
                           n2185, ZN => n5997);
   U17946 : INV_X1 port map( A => n5997, ZN => n6100);
   U17947 : INV_X1 port map( A => n5864, ZN => n5865);
   U17948 : NAND2_X1 port map( A1 => n1112, A2 => n6100, ZN => n6073);
   U17949 : OAI22_X1 port map( A1 => n2196, A2 => n7291, B1 => n2209, B2 => 
                           n2185, ZN => n6022);
   U17950 : INV_X1 port map( A => n6022, ZN => n6108);
   U17951 : AOI21_X1 port map( B1 => n5874, B2 => n5873, A => n1886, ZN => 
                           n5877);
   U17953 : INV_X1 port map( A => n6103, ZN => n6107);
   U17954 : OAI22_X1 port map( A1 => n2199, A2 => n7291, B1 => n2197, B2 => 
                           n2185, ZN => n6019);
   U17955 : INV_X1 port map( A => n6019, ZN => n6115);
   U17956 : INV_X1 port map( A => n6112, ZN => n6114);
   U17957 : OAI22_X1 port map( A1 => n17239, A2 => n7291, B1 => n2200, B2 => 
                           n2185, ZN => n6016);
   U17958 : INV_X1 port map( A => n6016, ZN => n6128);
   U17959 : INV_X1 port map( A => n6118, ZN => n6127);
   U17960 : OAI22_X1 port map( A1 => n2238, A2 => n7291, B1 => n17239, B2 => 
                           n2185, ZN => n6013);
   U17961 : INV_X1 port map( A => n6013, ZN => n6136);
   U17962 : NAND2_X1 port map( A1 => n6136, A2 => n461, ZN => n6122);
   U17963 : INV_X1 port map( A => n6142, ZN => n6145);
   U17964 : OAI21_X1 port map( B1 => n1608, B2 => n1794, A => n5913, ZN => 
                           n5971);
   U17965 : OAI21_X1 port map( B1 => n1834, B2 => n705, A => n690, ZN => n5976)
                           ;
   U17966 : INV_X1 port map( A => n17163, ZN => n6146);
   U17967 : OAI22_X1 port map( A1 => n2227, A2 => n7291, B1 => n2240, B2 => 
                           n2185, ZN => n6160);
   U17968 : INV_X1 port map( A => n6160, ZN => n6151);
   U17969 : INV_X1 port map( A => n6008, ZN => n6168);
   U17970 : OAI22_X1 port map( A1 => n2230, A2 => n7291, B1 => n2227, B2 => 
                           n2185, ZN => n6169);
   U17971 : INV_X1 port map( A => n6169, ZN => n6171);
   U17972 : NAND2_X1 port map( A1 => n2159, A2 => n6171, ZN => n6158);
   U17973 : INV_X1 port map( A => n6158, ZN => n5965);
   U17974 : OAI22_X1 port map( A1 => n2147, A2 => n7291, B1 => n2229, B2 => 
                           n2185, ZN => n6176);
   U17975 : INV_X1 port map( A => n6176, ZN => n6003);
   U17976 : NAND2_X1 port map( A1 => n776, A2 => n6003, ZN => n6157);
   U17977 : OAI22_X1 port map( A1 => n771, A2 => n7291, B1 => n2147, B2 => 
                           n2185, ZN => n8240);
   U17978 : INV_X1 port map( A => n8240, ZN => n6000);
   U17979 : AOI21_X1 port map( B1 => n662, B2 => n1095, A => n744, ZN => n5951)
                           ;
   U17980 : INV_X1 port map( A => n7290, ZN => n5962);
   U17981 : OAI21_X1 port map( B1 => n1711, B2 => n8240, A => n1827, ZN => 
                           n5963);
   U17982 : OAI21_X1 port map( B1 => n6002, B2 => n6000, A => n5963, ZN => 
                           n6177);
   U17983 : INV_X1 port map( A => n5999, ZN => n6175);
   U17984 : AOI21_X1 port map( B1 => n508, B2 => n911, A => n17170, ZN => n5964
                           );
   U17985 : NAND2_X1 port map( A1 => n1196, A2 => n6169, ZN => n6159);
   U17986 : OAI21_X1 port map( B1 => n5964, B2 => n5965, A => n6159, ZN => 
                           n5966);
   U17987 : OAI21_X1 port map( B1 => n6168, B2 => n6160, A => n5966, ZN => 
                           n5967);
   U17988 : OAI21_X1 port map( B1 => n6146, B2 => n6142, A => n6143, ZN => 
                           n5968);
   U17989 : OAI22_X1 port map( A1 => n2138, A2 => n7291, B1 => n2238, B2 => 
                           n2185, ZN => n6012);
   U17990 : INV_X1 port map( A => n6012, ZN => n6141);
   U17991 : INV_X1 port map( A => n656, ZN => n5970);
   U17992 : AOI21_X1 port map( B1 => n5971, B2 => n5972, A => n5970, ZN => 
                           n5973);
   U17993 : INV_X1 port map( A => n5974, ZN => n5975);
   U17994 : AOI21_X1 port map( B1 => n5976, B2 => n5977, A => n5975, ZN => 
                           n5980);
   U17995 : INV_X1 port map( A => n1134, ZN => n6140);
   U17996 : NAND2_X1 port map( A1 => n6140, A2 => n6012, ZN => n6119);
   U17997 : OAI211_X1 port map( C1 => n1607, C2 => n1793, A => n6120, B => 
                           n6119, ZN => n5983);
   U17998 : OAI211_X1 port map( C1 => n6127, C2 => n6016, A => n5983, B => 
                           n6122, ZN => n5984);
   U17999 : NAND2_X1 port map( A1 => n6096, A2 => n6073, ZN => n6094);
   U18000 : INV_X1 port map( A => n6095, ZN => n6099);
   U18001 : OAI22_X1 port map( A1 => n2204, A2 => n7291, B1 => n2215, B2 => 
                           n2185, ZN => n6085);
   U18002 : NAND2_X1 port map( A1 => n6198, A2 => n6085, ZN => n6078);
   U18003 : NAND3_X1 port map( A1 => n6094, A2 => n6074, A3 => n6078, ZN => 
                           n6053);
   U18004 : INV_X1 port map( A => n6085, ZN => n6089);
   U18005 : NAND2_X1 port map( A1 => n6089, A2 => n6023, ZN => n6075);
   U18006 : INV_X1 port map( A => n6079, ZN => n6070);
   U18007 : NAND2_X1 port map( A1 => n6070, A2 => n1297, ZN => n6054);
   U18008 : OAI22_X1 port map( A1 => n1219, A2 => n5994, B1 => n6027, B2 => 
                           n6057, ZN => n5995);
   U18009 : OAI21_X1 port map( B1 => n1106, B2 => n6031, A => n6037, ZN => 
                           n5996);
   U18010 : OAI21_X1 port map( B1 => n6039, B2 => n6032, A => n5996, ZN => 
                           n6781);
   U18011 : NAND2_X1 port map( A1 => n1112, A2 => n5997, ZN => n6084);
   U18012 : NAND2_X1 port map( A1 => n2159, A2 => n6169, ZN => n6150);
   U18013 : INV_X1 port map( A => n6150, ZN => n6005);
   U18014 : NAND2_X1 port map( A1 => n5999, A2 => n6176, ZN => n6149);
   U18015 : NAND2_X1 port map( A1 => n1892, A2 => n8255, ZN => n8254);
   U18016 : OAI21_X1 port map( B1 => n2169, B2 => n6000, A => n8254, ZN => 
                           n6001);
   U18017 : OAI21_X1 port map( B1 => n6002, B2 => n8240, A => n6001, ZN => 
                           n6178);
   U18018 : AOI21_X1 port map( B1 => n6149, B2 => n1481, A => n1772, ZN => 
                           n6004);
   U18019 : NAND2_X1 port map( A1 => n1196, A2 => n6171, ZN => n6152);
   U18020 : OAI21_X1 port map( B1 => n6004, B2 => n6005, A => n6152, ZN => 
                           n6006);
   U18021 : OAI21_X1 port map( B1 => n6146, B2 => n6145, A => n6144, ZN => 
                           n6009);
   U18022 : NAND2_X1 port map( A1 => n6141, A2 => n6140, ZN => n6124);
   U18023 : NAND2_X1 port map( A1 => n512, A2 => n6013, ZN => n6126);
   U18024 : NAND3_X1 port map( A1 => n6014, A2 => n6015, A3 => n6126, ZN => 
                           n6018);
   U18025 : OAI21_X1 port map( B1 => n6108, B2 => n6107, A => n858, ZN => n6021
                           );
   U18026 : NAND2_X1 port map( A1 => n571, A2 => n6084, ZN => n6067);
   U18027 : NAND2_X1 port map( A1 => n6099, A2 => n6100, ZN => n6066);
   U18028 : NAND2_X1 port map( A1 => n1220, A2 => n6089, ZN => n6072);
   U18029 : NAND3_X1 port map( A1 => n6072, A2 => n439, A3 => n6067, ZN => 
                           n6055);
   U18030 : INV_X1 port map( A => n6055, ZN => n6026);
   U18031 : NAND2_X1 port map( A1 => n6085, A2 => n6023, ZN => n6068);
   U18032 : INV_X1 port map( A => n6068, ZN => n6025);
   U18033 : NAND2_X1 port map( A1 => n1297, A2 => n6079, ZN => n6056);
   U18034 : NOR3_X1 port map( A1 => n6026, A2 => n6025, A3 => n1223, ZN => 
                           n6028);
   U18035 : OAI22_X1 port map( A1 => n6028, A2 => n1226, B1 => n6027, B2 => 
                           n6060, ZN => n6029);
   U18036 : OAI21_X1 port map( B1 => n6039, B2 => n1684, A => n6050, ZN => 
                           n6030);
   U18037 : OAI21_X1 port map( B1 => n6032, B2 => n6031, A => n6030, ZN => 
                           n6956);
   U18038 : XOR2_X1 port map( A => n6033, B => n6956, Z => n6034);
   U18039 : XOR2_X1 port map( A => n2265, B => n8229, Z => n6036);
   U18040 : NAND2_X1 port map( A1 => n6036, A2 => n7284, ZN => n7285);
   U18041 : OAI22_X1 port map( A1 => n2213, A2 => n7285, B1 => n2175, B2 => 
                           n7284, ZN => n6696);
   U18042 : INV_X1 port map( A => n6696, ZN => n6695);
   U18043 : OAI22_X1 port map( A1 => n2215, A2 => n7285, B1 => n2213, B2 => 
                           n7284, ZN => n6233);
   U18044 : INV_X1 port map( A => n6233, ZN => n6237);
   U18045 : XOR2_X1 port map( A => n6039, B => n6038, Z => n6040);
   U18046 : XOR2_X1 port map( A => n1500, B => n6042, Z => n6048);
   U18047 : NAND3_X1 port map( A1 => n6044, A2 => n6043, A3 => n6776, ZN => 
                           n6047);
   U18048 : NAND3_X1 port map( A1 => n1500, A2 => n1081, A3 => n6776, ZN => 
                           n6046);
   U18049 : OAI211_X1 port map( C1 => n6776, C2 => n6048, A => n6047, B => 
                           n6046, ZN => n6049);
   U18050 : INV_X1 port map( A => n6234, ZN => n6236);
   U18051 : NAND2_X1 port map( A1 => n6060, A2 => n6967, ZN => n6065);
   U18052 : NAND3_X1 port map( A1 => n6053, A2 => n6075, A3 => n6054, ZN => 
                           n6064);
   U18053 : INV_X1 port map( A => n6065, ZN => n6059);
   U18054 : AOI22_X1 port map( A1 => n339, A2 => n1009, B1 => n6061, B2 => 
                           n6064, ZN => n6062);
   U18055 : OAI211_X1 port map( C1 => n6065, C2 => n6064, A => n6062, B => 
                           n6063, ZN => n6242);
   U18056 : XOR2_X1 port map( A => n6242, B => n1681, Z => n6223);
   U18057 : OAI22_X1 port map( A1 => n2205, A2 => n7285, B1 => n2215, B2 => 
                           n7284, ZN => n6222);
   U18058 : INV_X1 port map( A => n6221, ZN => n6252);
   U18059 : NAND2_X1 port map( A1 => n6079, A2 => n2266, ZN => n6081);
   U18060 : NAND2_X1 port map( A1 => n6070, A2 => n6967, ZN => n6076);
   U18061 : INV_X1 port map( A => n6066, ZN => n6088);
   U18062 : INV_X1 port map( A => n6067, ZN => n6069);
   U18063 : OAI21_X1 port map( B1 => n6088, B2 => n1601, A => n6068, ZN => 
                           n6082);
   U18064 : NAND4_X1 port map( A1 => n6082, A2 => n2266, A3 => n6072, A4 => 
                           n6070, ZN => n6071);
   U18065 : NAND3_X1 port map( A1 => n557, A2 => n6250, A3 => n973, ZN => n6083
                           );
   U18066 : OAI22_X1 port map( A1 => n2197, A2 => n7285, B1 => n2209, B2 => 
                           n7284, ZN => n6220);
   U18067 : INV_X1 port map( A => n6220, ZN => n6258);
   U18068 : NAND2_X1 port map( A1 => n6089, A2 => n6967, ZN => n6093);
   U18069 : INV_X1 port map( A => n6093, ZN => n6087);
   U18070 : AOI22_X1 port map( A1 => n338, A2 => n6069, B1 => n6094, B2 => 
                           n6090, ZN => n6091);
   U18071 : OAI211_X1 port map( C1 => n1087, C2 => n6093, A => n6091, B => 
                           n1151, ZN => n6199);
   U18072 : INV_X1 port map( A => n6218, ZN => n6192);
   U18073 : INV_X1 port map( A => n6217, ZN => n6267);
   U18074 : INV_X1 port map( A => n6262, ZN => n6266);
   U18075 : OAI22_X1 port map( A1 => n17239, A2 => n7285, B1 => n2200, B2 => 
                           n7284, ZN => n6215);
   U18076 : INV_X1 port map( A => n6215, ZN => n6271);
   U18077 : OAI22_X1 port map( A1 => n2238, A2 => n7285, B1 => n17240, B2 => 
                           n7284, ZN => n6200);
   U18078 : NAND2_X1 port map( A1 => n6292, A2 => n1178, ZN => n6276);
   U18079 : OAI21_X1 port map( B1 => n1793, B2 => n1607, A => n6119, ZN => 
                           n6133);
   U18080 : INV_X1 port map( A => n6120, ZN => n6121);
   U18081 : AOI21_X1 port map( B1 => n985, B2 => n6122, A => n6121, ZN => n6123
                           );
   U18082 : OAI21_X1 port map( B1 => n1485, B2 => n1848, A => n6124, ZN => 
                           n6135);
   U18083 : AOI21_X1 port map( B1 => n6135, B2 => n6126, A => n671, ZN => n6129
                           );
   U18084 : INV_X1 port map( A => n6296, ZN => n6201);
   U18085 : OAI22_X1 port map( A1 => n2138, A2 => n7285, B1 => n2238, B2 => 
                           n7284, ZN => n6202);
   U18086 : NAND2_X1 port map( A1 => n6201, A2 => n6202, ZN => n6289);
   U18087 : INV_X1 port map( A => n6202, ZN => n6295);
   U18088 : NAND2_X1 port map( A1 => n6296, A2 => n6295, ZN => n6274);
   U18089 : OAI22_X1 port map( A1 => n2240, A2 => n7285, B1 => n2239, B2 => 
                           n7284, ZN => n6309);
   U18090 : INV_X1 port map( A => n6309, ZN => n6312);
   U18091 : XOR2_X1 port map( A => n512, B => n6136, Z => n6134);
   U18092 : NAND2_X1 port map( A1 => n6312, A2 => n739, ZN => n6301);
   U18093 : OAI22_X1 port map( A1 => n2227, A2 => n7285, B1 => n2240, B2 => 
                           n7284, ZN => n6316);
   U18094 : NAND2_X1 port map( A1 => n1718, A2 => n6316, ZN => n6298);
   U18095 : OAI22_X1 port map( A1 => n2229, A2 => n7285, B1 => n2227, B2 => 
                           n7284, ZN => n6323);
   U18096 : INV_X1 port map( A => n6323, ZN => n6325);
   U18097 : OAI22_X1 port map( A1 => n2147, A2 => n7285, B1 => n2229, B2 => 
                           n7284, ZN => n6328);
   U18098 : INV_X1 port map( A => n6328, ZN => n6204);
   U18099 : NAND2_X1 port map( A1 => n6151, A2 => n6967, ZN => n6163);
   U18100 : NAND2_X1 port map( A1 => n6160, A2 => n2266, ZN => n6164);
   U18101 : OAI21_X1 port map( B1 => n1161, B2 => n17170, A => n6158, ZN => 
                           n6162);
   U18102 : INV_X1 port map( A => n8227, ZN => n6206);
   U18103 : NOR2_X1 port map( A1 => n1788, A2 => n1775, ZN => n6170);
   U18104 : NOR2_X1 port map( A1 => n1789, A2 => n17208, ZN => n6172);
   U18105 : INV_X1 port map( A => n6208, ZN => n8226);
   U18106 : XOR2_X1 port map( A => n1481, B => n6179, Z => n6180);
   U18107 : INV_X1 port map( A => n7284, ZN => n6182);
   U18108 : NAND2_X1 port map( A1 => n6182, A2 => n2154, ZN => n6183);
   U18109 : INV_X1 port map( A => n6183, ZN => n8239);
   U18110 : INV_X1 port map( A => n6203, ZN => n6313);
   U18111 : NAND3_X1 port map( A1 => n6299, A2 => n6297, A3 => n6298, ZN => 
                           n6273);
   U18112 : NAND3_X1 port map( A1 => n6273, A2 => n6301, A3 => n6274, ZN => 
                           n6187);
   U18113 : NAND3_X1 port map( A1 => n208, A2 => n6275, A3 => n6289, ZN => 
                           n6188);
   U18114 : OAI211_X1 port map( C1 => n1442, C2 => n6215, A => n6188, B => 
                           n6276, ZN => n6189);
   U18115 : OAI21_X1 port map( B1 => n6266, B2 => n6217, A => n6263, ZN => 
                           n6190);
   U18116 : OAI21_X1 port map( B1 => n6218, B2 => n6220, A => n1013, ZN => 
                           n6191);
   U18117 : OAI21_X1 port map( B1 => n6192, B2 => n6258, A => n6191, ZN => 
                           n6249);
   U18119 : NAND2_X1 port map( A1 => n1178, A2 => n6200, ZN => n6283);
   U18120 : NAND2_X1 port map( A1 => n1150, A2 => n6292, ZN => n6281);
   U18121 : NAND2_X1 port map( A1 => n6295, A2 => n6201, ZN => n6291);
   U18122 : NAND2_X1 port map( A1 => n6296, A2 => n6202, ZN => n6280);
   U18123 : NAND2_X1 port map( A1 => n6309, A2 => n740, ZN => n6307);
   U18124 : NAND2_X1 port map( A1 => n17164, A2 => n6319, ZN => n6304);
   U18125 : NAND2_X1 port map( A1 => n8238, A2 => n8239, ZN => n8237);
   U18126 : OAI21_X1 port map( B1 => n8226, B2 => n6206, A => n8237, ZN => 
                           n6207);
   U18128 : OAI21_X1 port map( B1 => n743, B2 => n6325, A => n642, ZN => n6211)
                           ;
   U18129 : NAND2_X1 port map( A1 => n6313, A2 => n6312, ZN => n6305);
   U18130 : NAND3_X1 port map( A1 => n6305, A2 => n6303, A3 => n6304, ZN => 
                           n6279);
   U18131 : NAND3_X1 port map( A1 => n6279, A2 => n6307, A3 => n6280, ZN => 
                           n6212);
   U18132 : NAND3_X1 port map( A1 => n6281, A2 => n6291, A3 => n6212, ZN => 
                           n6213);
   U18133 : OAI211_X1 port map( C1 => n6271, C2 => n1442, A => n6213, B => 
                           n6283, ZN => n6214);
   U18134 : OAI21_X1 port map( B1 => n732, B2 => n6267, A => n6265, ZN => n6216
                           );
   U18135 : OAI21_X1 port map( B1 => n6258, B2 => n6218, A => n6259, ZN => 
                           n6219);
   U18136 : XOR2_X1 port map( A => n8229, B => n7973, Z => n6232);
   U18137 : OAI22_X1 port map( A1 => n2204, A2 => n7274, B1 => n2215, B2 => 
                           n7272, ZN => n6793);
   U18138 : OAI22_X1 port map( A1 => n2208, A2 => n7274, B1 => n2205, B2 => 
                           n7272, ZN => n6365);
   U18139 : INV_X1 port map( A => n6365, ZN => n6374);
   U18140 : INV_X1 port map( A => n897, ZN => n6373);
   U18141 : OAI22_X1 port map( A1 => n2196, A2 => n7274, B1 => n2209, B2 => 
                           n7272, ZN => n6363);
   U18142 : INV_X1 port map( A => n6363, ZN => n6392);
   U18143 : INV_X1 port map( A => n6244, ZN => n6246);
   U18144 : OAI22_X1 port map( A1 => n2199, A2 => n7274, B1 => n2197, B2 => 
                           n7272, ZN => n6343);
   U18145 : NAND3_X1 port map( A1 => n506, A2 => n6250, A3 => n557, ZN => n6253
                           );
   U18146 : NAND2_X1 port map( A1 => n1007, A2 => n6396, ZN => n6384);
   U18147 : INV_X1 port map( A => n6459, ZN => n6460);
   U18148 : OAI22_X1 port map( A1 => n17239, A2 => n7274, B1 => n2200, B2 => 
                           n7272, ZN => n6344);
   U18149 : INV_X1 port map( A => n6344, ZN => n6461);
   U18150 : NAND2_X1 port map( A1 => n6459, A2 => n6461, ZN => n6380);
   U18151 : OAI22_X1 port map( A1 => n2238, A2 => n7274, B1 => n17240, B2 => 
                           n7272, ZN => n6360);
   U18152 : INV_X1 port map( A => n6360, ZN => n6406);
   U18153 : XOR2_X1 port map( A => n1003, B => n6267, Z => n6264);
   U18154 : XOR2_X1 port map( A => n6268, B => n1252, Z => n6269);
   U18155 : INV_X1 port map( A => n6403, ZN => n6405);
   U18156 : OAI22_X1 port map( A1 => n2138, A2 => n7274, B1 => n2238, B2 => 
                           n7272, ZN => n6358);
   U18157 : INV_X1 port map( A => n6358, ZN => n6421);
   U18158 : AOI21_X1 port map( B1 => n1727, B2 => n6276, A => n946, ZN => n6277
                           );
   U18159 : XOR2_X1 port map( A => n6278, B => n6277, Z => n6287);
   U18160 : NAND3_X1 port map( A1 => n6279, A2 => n6307, A3 => n6280, ZN => 
                           n6290);
   U18161 : NAND2_X1 port map( A1 => n6291, A2 => n6212, ZN => n6284);
   U18162 : INV_X1 port map( A => n6281, ZN => n6282);
   U18163 : AOI21_X1 port map( B1 => n6284, B2 => n6283, A => n6282, ZN => 
                           n6285);
   U18164 : OAI22_X1 port map( A1 => n2240, A2 => n7274, B1 => n2239, B2 => 
                           n7272, ZN => n6345);
   U18165 : INV_X1 port map( A => n6345, ZN => n6430);
   U18166 : NAND2_X1 port map( A1 => n6430, A2 => n1032, ZN => n6413);
   U18167 : NAND2_X1 port map( A1 => n242, A2 => n6298, ZN => n6310);
   U18168 : INV_X1 port map( A => n6299, ZN => n6300);
   U18169 : AOI21_X1 port map( B1 => n6301, B2 => n6310, A => n6300, ZN => 
                           n6302);
   U18170 : NAND2_X1 port map( A1 => n6304, A2 => n6303, ZN => n6311);
   U18171 : INV_X1 port map( A => n6305, ZN => n6306);
   U18172 : AOI21_X1 port map( B1 => n6307, B2 => n6311, A => n6306, ZN => 
                           n6308);
   U18173 : OAI22_X1 port map( A1 => n2227, A2 => n7274, B1 => n2240, B2 => 
                           n7272, ZN => n6448);
   U18174 : NAND2_X1 port map( A1 => n1888, A2 => n6448, ZN => n6426);
   U18175 : OAI22_X1 port map( A1 => n2230, A2 => n7274, B1 => n2227, B2 => 
                           n7272, ZN => n6355);
   U18176 : INV_X1 port map( A => n6354, ZN => n6438);
   U18177 : OAI22_X1 port map( A1 => n2147, A2 => n7274, B1 => n2229, B2 => 
                           n7272, ZN => n6440);
   U18178 : INV_X1 port map( A => n6440, ZN => n6346);
   U18179 : INV_X1 port map( A => n6350, ZN => n6439);
   U18180 : OAI22_X1 port map( A1 => n2132, A2 => n7274, B1 => n2147, B2 => 
                           n7272, ZN => n7964);
   U18181 : INV_X1 port map( A => n7964, ZN => n6347);
   U18182 : XOR2_X1 port map( A => n2161, B => n822, Z => n6330);
   U18183 : INV_X1 port map( A => n7272, ZN => n6332);
   U18184 : OAI21_X1 port map( B1 => n953, B2 => n7964, A => n1830, ZN => n6333
                           );
   U18185 : OAI21_X1 port map( B1 => n6347, B2 => n6349, A => n6333, ZN => 
                           n6441);
   U18186 : OAI21_X1 port map( B1 => n1028, B2 => n6440, A => n6441, ZN => 
                           n6334);
   U18187 : OAI21_X1 port map( B1 => n6438, B2 => n6355, A => n6433, ZN => 
                           n6335);
   U18188 : INV_X1 port map( A => n1031, ZN => n6429);
   U18189 : NAND2_X1 port map( A1 => n6429, A2 => n6345, ZN => n6411);
   U18190 : NAND3_X1 port map( A1 => n655, A2 => n6426, A3 => n6411, ZN => 
                           n6336);
   U18191 : OAI211_X1 port map( C1 => n6420, C2 => n6358, A => n6413, B => 
                           n6336, ZN => n6337);
   U18192 : NAND3_X1 port map( A1 => n652, A2 => n606, A3 => n6382, ZN => n6339
                           );
   U18193 : OAI211_X1 port map( C1 => n220, C2 => n6363, A => n6339, B => n6384
                           , ZN => n6340);
   U18195 : OAI21_X1 port map( B1 => n647, B2 => n6365, A => n6372, ZN => n6341
                           );
   U18196 : NAND2_X1 port map( A1 => n1007, A2 => n6343, ZN => n6390);
   U18197 : NAND2_X1 port map( A1 => n6459, A2 => n6344, ZN => n6388);
   U18198 : NAND2_X1 port map( A1 => n1032, A2 => n6345, ZN => n6418);
   U18199 : INV_X1 port map( A => n6448, ZN => n6451);
   U18200 : NAND2_X1 port map( A1 => n909, A2 => n6451, ZN => n6428);
   U18201 : NAND2_X1 port map( A1 => n1894, A2 => n8221, ZN => n8220);
   U18202 : OAI21_X1 port map( B1 => n1050, B2 => n6347, A => n8220, ZN => 
                           n6348);
   U18203 : OAI21_X1 port map( B1 => n6349, B2 => n7964, A => n6348, ZN => 
                           n6442);
   U18204 : OAI21_X1 port map( B1 => n6438, B2 => n6436, A => n6435, ZN => 
                           n6353);
   U18205 : NAND3_X1 port map( A1 => n1396, A2 => n6428, A3 => n6416, ZN => 
                           n6356);
   U18206 : OAI211_X1 port map( C1 => n6421, C2 => n6420, A => n6356, B => 
                           n6418, ZN => n6357);
   U18207 : OAI21_X1 port map( B1 => n6410, B2 => n6358, A => n6357, ZN => 
                           n6404);
   U18208 : NAND2_X1 port map( A1 => n6388, A2 => n6387, ZN => n6399);
   U18209 : NAND3_X1 port map( A1 => n6399, A2 => n919, A3 => n6400, ZN => 
                           n6361);
   U18210 : OAI211_X1 port map( C1 => n6392, C2 => n815, A => n6390, B => n6361
                           , ZN => n6362);
   U18211 : OAI21_X1 port map( B1 => n6374, B2 => n6373, A => n980, ZN => n6364
                           );
   U18212 : OAI21_X1 port map( B1 => n250, B2 => n6365, A => n6364, ZN => n6795
                           );
   U18213 : XOR2_X1 port map( A => n7973, B => n1702, Z => n6370);
   U18214 : OAI22_X1 port map( A1 => n2197, A2 => n7266, B1 => n2209, B2 => 
                           n7265, ZN => n6802);
   U18215 : OAI22_X1 port map( A1 => n2199, A2 => n7266, B1 => n2197, B2 => 
                           n7265, ZN => n6490);
   U18216 : INV_X1 port map( A => n6490, ZN => n6501);
   U18217 : INV_X1 port map( A => n1094, ZN => n6500);
   U18218 : OAI22_X1 port map( A1 => n17239, A2 => n7266, B1 => n2200, B2 => 
                           n7265, ZN => n6488);
   U18219 : INV_X1 port map( A => n6380, ZN => n6381);
   U18220 : OAI21_X1 port map( B1 => n653, B2 => n6381, A => n606, ZN => n6385)
                           ;
   U18222 : AOI21_X1 port map( B1 => n6385, B2 => n6384, A => n17171, ZN => 
                           n6386);
   U18223 : OAI21_X1 port map( B1 => n610, B2 => n997, A => n6400, ZN => n6391)
                           ;
   U18224 : INV_X1 port map( A => n919, ZN => n6389);
   U18225 : AOI21_X1 port map( B1 => n6391, B2 => n6390, A => n6389, ZN => 
                           n6393);
   U18226 : INV_X1 port map( A => n850, ZN => n6514);
   U18227 : OAI22_X1 port map( A1 => n2238, A2 => n7266, B1 => n17240, B2 => 
                           n7265, ZN => n6468);
   U18228 : NAND2_X1 port map( A1 => n1124, A2 => n6522, ZN => n6508);
   U18229 : OAI22_X1 port map( A1 => n2240, A2 => n7266, B1 => n2239, B2 => 
                           n7265, ZN => n6482);
   U18230 : INV_X1 port map( A => n6482, ZN => n6530);
   U18231 : INV_X1 port map( A => n6404, ZN => n6407);
   U18232 : INV_X1 port map( A => n1120, ZN => n6529);
   U18233 : OAI22_X1 port map( A1 => n2227, A2 => n7266, B1 => n2240, B2 => 
                           n7265, ZN => n6480);
   U18234 : INV_X1 port map( A => n6480, ZN => n6548);
   U18235 : NAND2_X1 port map( A1 => n6426, A2 => n655, ZN => n6414);
   U18236 : INV_X1 port map( A => n6411, ZN => n6412);
   U18237 : AOI21_X1 port map( B1 => n6414, B2 => n6413, A => n6412, ZN => 
                           n6415);
   U18238 : NAND2_X1 port map( A1 => n6428, A2 => n1396, ZN => n6419);
   U18239 : INV_X1 port map( A => n6416, ZN => n6417);
   U18240 : AOI21_X1 port map( B1 => n6419, B2 => n6418, A => n6417, ZN => 
                           n6422);
   U18241 : INV_X1 port map( A => n6534, ZN => n6547);
   U18242 : OAI22_X1 port map( A1 => n2229, A2 => n7266, B1 => n2227, B2 => 
                           n7265, ZN => n6555);
   U18243 : INV_X1 port map( A => n6555, ZN => n6476);
   U18244 : NAND2_X1 port map( A1 => n1540, A2 => n6476, ZN => n6539);
   U18245 : OAI22_X1 port map( A1 => n771, A2 => n7266, B1 => n2147, B2 => 
                           n7265, ZN => n7895);
   U18246 : INV_X1 port map( A => n7895, ZN => n6471);
   U18247 : INV_X1 port map( A => n6469, ZN => n7936);
   U18248 : INV_X1 port map( A => n7265, ZN => n6446);
   U18249 : NAND2_X1 port map( A1 => n6446, A2 => n2154, ZN => n7935);
   U18250 : INV_X1 port map( A => n7935, ZN => n6470);
   U18251 : OAI21_X1 port map( B1 => n1517, B2 => n7895, A => n1783, ZN => 
                           n6447);
   U18252 : INV_X1 port map( A => n1406, ZN => n6561);
   U18253 : OAI22_X1 port map( A1 => n2147, A2 => n7266, B1 => n2229, B2 => 
                           n7265, ZN => n6560);
   U18254 : INV_X1 port map( A => n6560, ZN => n6475);
   U18255 : XOR2_X1 port map( A => n1888, B => n6451, Z => n6452);
   U18256 : NAND2_X1 port map( A1 => n6475, A2 => n1713, ZN => n6536);
   U18257 : INV_X1 port map( A => n6536, ZN => n6455);
   U18258 : INV_X1 port map( A => n6474, ZN => n6559);
   U18259 : NAND2_X1 port map( A1 => n6559, A2 => n6560, ZN => n6552);
   U18260 : INV_X1 port map( A => n6551, ZN => n6556);
   U18261 : NAND2_X1 port map( A1 => n852, A2 => n6555, ZN => n6537);
   U18262 : OAI211_X1 port map( C1 => n6561, C2 => n6455, A => n6537, B => 
                           n6552, ZN => n6456);
   U18263 : OAI211_X1 port map( C1 => n6547, C2 => n6480, A => n6539, B => 
                           n6456, ZN => n6457);
   U18264 : OAI22_X1 port map( A1 => n2138, A2 => n7266, B1 => n2238, B2 => 
                           n7265, ZN => n6484);
   U18267 : OAI211_X1 port map( C1 => n1104, C2 => n1849, A => n6506, B => 
                           n6507, ZN => n6464);
   U18268 : OAI211_X1 port map( C1 => n6514, C2 => n6488, A => n6464, B => 
                           n6508, ZN => n6465);
   U18269 : OAI21_X1 port map( B1 => n6515, B2 => n1594, A => n6465, ZN => 
                           n6498);
   U18270 : OAI21_X1 port map( B1 => n6500, B2 => n6490, A => n6498, ZN => 
                           n6466);
   U18271 : NAND2_X1 port map( A1 => n1124, A2 => n6468, ZN => n6513);
   U18272 : NAND2_X1 port map( A1 => n6555, A2 => n1540, ZN => n6546);
   U18273 : NAND2_X1 port map( A1 => n6470, A2 => n6469, ZN => n7898);
   U18274 : OAI21_X1 port map( B1 => n1517, B2 => n6471, A => n7898, ZN => 
                           n6472);
   U18275 : OAI21_X1 port map( B1 => n6473, B2 => n7895, A => n6472, ZN => 
                           n6543);
   U18276 : INV_X1 port map( A => n6543, ZN => n6563);
   U18277 : NAND2_X1 port map( A1 => n6560, A2 => n1713, ZN => n6544);
   U18278 : INV_X1 port map( A => n6544, ZN => n6477);
   U18279 : NAND2_X1 port map( A1 => n6559, A2 => n6475, ZN => n6557);
   U18280 : NAND2_X1 port map( A1 => n6556, A2 => n6476, ZN => n6545);
   U18281 : OAI211_X1 port map( C1 => n6477, C2 => n6563, A => n6545, B => 
                           n6557, ZN => n6478);
   U18282 : OAI211_X1 port map( C1 => n6548, C2 => n6547, A => n6546, B => 
                           n6478, ZN => n6479);
   U18283 : OAI211_X1 port map( C1 => n1847, C2 => n764, A => n6510, B => n6511
                           , ZN => n6486);
   U18284 : OAI211_X1 port map( C1 => n631, C2 => n6515, A => n6513, B => n6486
                           , ZN => n6487);
   U18285 : INV_X1 port map( A => n6491, ZN => n6805);
   U18286 : XOR2_X1 port map( A => n1702, B => n7835, Z => n6496);
   U18287 : NAND2_X1 port map( A1 => n6496, A2 => n7256, ZN => n7258);
   U18288 : OAI22_X1 port map( A1 => n17239, A2 => n7258, B1 => n2200, B2 => 
                           n7256, ZN => n6809);
   U18289 : INV_X1 port map( A => n6809, ZN => n6812);
   U18290 : OAI22_X1 port map( A1 => n2238, A2 => n7258, B1 => n17240, B2 => 
                           n7256, ZN => n6590);
   U18291 : INV_X1 port map( A => n6590, ZN => n6599);
   U18292 : INV_X1 port map( A => n6596, ZN => n6598);
   U18293 : OAI22_X1 port map( A1 => n2239, A2 => n7258, B1 => n2238, B2 => 
                           n7256, ZN => n6589);
   U18294 : OAI21_X1 port map( B1 => n1849, B2 => n1104, A => n6506, ZN => 
                           n6520);
   U18295 : AOI21_X1 port map( B1 => n6508, B2 => n1650, A => n1172, ZN => 
                           n6509);
   U18296 : OAI21_X1 port map( B1 => n1097, B2 => n1847, A => n6510, ZN => 
                           n6521);
   U18297 : INV_X1 port map( A => n6511, ZN => n6512);
   U18298 : AOI21_X1 port map( B1 => n6513, B2 => n6521, A => n6512, ZN => 
                           n6516);
   U18299 : INV_X1 port map( A => n6604, ZN => n6587);
   U18300 : OAI22_X1 port map( A1 => n2240, A2 => n7258, B1 => n2239, B2 => 
                           n7256, ZN => n6574);
   U18301 : OAI22_X1 port map( A1 => n2227, A2 => n7258, B1 => n2240, B2 => 
                           n7256, ZN => n6575);
   U18302 : NAND2_X1 port map( A1 => n1651, A2 => n6575, ZN => n6605);
   U18303 : OAI22_X1 port map( A1 => n2229, A2 => n7258, B1 => n2227, B2 => 
                           n7256, ZN => n6629);
   U18304 : INV_X1 port map( A => n6629, ZN => n6632);
   U18305 : INV_X1 port map( A => n6585, ZN => n6633);
   U18306 : OAI22_X1 port map( A1 => n2147, A2 => n7258, B1 => n2230, B2 => 
                           n7256, ZN => n6634);
   U18307 : INV_X1 port map( A => n6634, ZN => n6581);
   U18308 : XOR2_X1 port map( A => n1070, B => n6548, Z => n6542);
   U18309 : NAND2_X1 port map( A1 => n6535, A2 => n6536, ZN => n6553);
   U18310 : NAND2_X1 port map( A1 => n6553, A2 => n6552, ZN => n6540);
   U18311 : INV_X1 port map( A => n6537, ZN => n6538);
   U18312 : AOI21_X1 port map( B1 => n6539, B2 => n6540, A => n6538, ZN => 
                           n6541);
   U18313 : NAND2_X1 port map( A1 => n6543, A2 => n6544, ZN => n6558);
   U18314 : AOI21_X1 port map( B1 => n6546, B2 => n1098, A => n1016, ZN => 
                           n6550);
   U18315 : OAI22_X1 port map( A1 => n2132, A2 => n7258, B1 => n2147, B2 => 
                           n7256, ZN => n7828);
   U18316 : INV_X1 port map( A => n7828, ZN => n6578);
   U18317 : INV_X1 port map( A => n7256, ZN => n6566);
   U18318 : NAND2_X1 port map( A1 => n6566, A2 => n2154, ZN => n7850);
   U18319 : INV_X1 port map( A => n7850, ZN => n6577);
   U18320 : OAI21_X1 port map( B1 => n1324, B2 => n7828, A => n1829, ZN => 
                           n6567);
   U18321 : OAI21_X1 port map( B1 => n6580, B2 => n6578, A => n6567, ZN => 
                           n6635);
   U18322 : OAI21_X1 port map( B1 => n1069, B2 => n6634, A => n6635, ZN => 
                           n6568);
   U18323 : OAI21_X1 port map( B1 => n982, B2 => n6629, A => n6630, ZN => n6569
                           );
   U18324 : NAND2_X1 port map( A1 => n1132, A2 => n6574, ZN => n6606);
   U18325 : NAND3_X1 port map( A1 => n6606, A2 => n6605, A3 => n970, ZN => 
                           n6570);
   U18326 : OAI211_X1 port map( C1 => n6587, C2 => n6589, A => n1254, B => 
                           n6570, ZN => n6571);
   U18327 : OAI21_X1 port map( B1 => n6598, B2 => n6590, A => n6597, ZN => 
                           n6572);
   U18328 : INV_X1 port map( A => n6575, ZN => n6625);
   U18329 : NAND2_X1 port map( A1 => n6625, A2 => n1651, ZN => n6610);
   U18330 : NAND2_X1 port map( A1 => n6576, A2 => n6577, ZN => n7831);
   U18331 : OAI21_X1 port map( B1 => n1324, B2 => n6578, A => n7831, ZN => 
                           n6579);
   U18332 : OAI21_X1 port map( B1 => n17167, B2 => n7828, A => n6579, ZN => 
                           n6636);
   U18333 : OAI21_X1 port map( B1 => n1069, B2 => n6581, A => n6636, ZN => 
                           n6582);
   U18334 : OAI21_X1 port map( B1 => n6633, B2 => n6632, A => n6631, ZN => 
                           n6584);
   U18335 : OAI21_X1 port map( B1 => n6625, B2 => n1651, A => n6624, ZN => 
                           n6609);
   U18336 : NAND2_X1 port map( A1 => n6619, A2 => n1132, ZN => n6611);
   U18337 : NAND3_X1 port map( A1 => n6609, A2 => n6611, A3 => n6610, ZN => 
                           n6586);
   U18338 : OAI211_X1 port map( C1 => n6603, C2 => n17224, A => n6612, B => 
                           n6586, ZN => n6588);
   U18339 : OAI21_X1 port map( B1 => n1586, B2 => n6590, A => n572, ZN => n6991
                           );
   U18340 : INV_X1 port map( A => n6810, ZN => n6811);
   U18341 : XOR2_X1 port map( A => n7835, B => n7771, Z => n6595);
   U18342 : OAI22_X1 port map( A1 => n2239, A2 => n7248, B1 => n2238, B2 => 
                           n7247, ZN => n6822);
   U18343 : INV_X1 port map( A => n6822, ZN => n6820);
   U18344 : OAI22_X1 port map( A1 => n2240, A2 => n7248, B1 => n2239, B2 => 
                           n7247, ZN => n6657);
   U18345 : INV_X1 port map( A => n6657, ZN => n6673);
   U18346 : INV_X1 port map( A => n6661, ZN => n6672);
   U18347 : OAI22_X1 port map( A1 => n2227, A2 => n7248, B1 => n2240, B2 => 
                           n7247, ZN => n6646);
   U18348 : NAND2_X1 port map( A1 => n970, A2 => n6605, ZN => n6617);
   U18349 : AOI21_X1 port map( B1 => n6617, B2 => n6607, A => n625, ZN => n6608
                           );
   U18350 : NAND2_X1 port map( A1 => n6609, A2 => n6610, ZN => n6618);
   U18351 : AOI21_X1 port map( B1 => n6612, B2 => n6618, A => n722, ZN => n6613
                           );
   U18352 : NAND2_X1 port map( A1 => n6681, A2 => n1175, ZN => n6665);
   U18353 : OAI22_X1 port map( A1 => n2229, A2 => n7248, B1 => n2227, B2 => 
                           n7247, ZN => n6682);
   U18354 : NAND2_X1 port map( A1 => n566, A2 => n6682, ZN => n6662);
   U18355 : OAI22_X1 port map( A1 => n2147, A2 => n7248, B1 => n2230, B2 => 
                           n7247, ZN => n6684);
   U18356 : INV_X1 port map( A => n6684, ZN => n6652);
   U18357 : OAI22_X1 port map( A1 => n2132, A2 => n7248, B1 => n2147, B2 => 
                           n7247, ZN => n7764);
   U18358 : INV_X1 port map( A => n7764, ZN => n6649);
   U18359 : XOR2_X1 port map( A => n1069, B => n6634, Z => n6637);
   U18360 : XOR2_X1 port map( A => n6637, B => n1615, Z => n6638);
   U18361 : INV_X1 port map( A => n6647, ZN => n7803);
   U18362 : INV_X1 port map( A => n7247, ZN => n6640);
   U18363 : NAND2_X1 port map( A1 => n6640, A2 => n2154, ZN => n7802);
   U18364 : INV_X1 port map( A => n7802, ZN => n6648);
   U18365 : OAI21_X1 port map( B1 => n1391, B2 => n7764, A => n1782, ZN => 
                           n6641);
   U18366 : OAI21_X1 port map( B1 => n6649, B2 => n6651, A => n6641, ZN => 
                           n6685);
   U18367 : OAI21_X1 port map( B1 => n1712, B2 => n6684, A => n6685, ZN => 
                           n6642);
   U18368 : INV_X1 port map( A => n6677, ZN => n6680);
   U18369 : NAND3_X1 port map( A1 => n634, A2 => n6663, A3 => n6662, ZN => 
                           n6643);
   U18370 : OAI211_X1 port map( C1 => n6672, C2 => n6657, A => n6643, B => 
                           n6665, ZN => n6644);
   U18371 : NAND2_X1 port map( A1 => n1175, A2 => n6646, ZN => n6671);
   U18372 : INV_X1 port map( A => n6682, ZN => n6683);
   U18373 : NAND2_X1 port map( A1 => n1867, A2 => n6683, ZN => n6668);
   U18374 : NAND2_X1 port map( A1 => n6648, A2 => n6647, ZN => n7767);
   U18375 : OAI21_X1 port map( B1 => n1391, B2 => n6649, A => n7767, ZN => 
                           n6650);
   U18376 : OAI21_X1 port map( B1 => n7764, B2 => n6651, A => n6650, ZN => 
                           n6686);
   U18377 : OAI21_X1 port map( B1 => n1712, B2 => n6652, A => n6686, ZN => 
                           n6653);
   U18378 : NAND3_X1 port map( A1 => n6669, A2 => n668, A3 => n6668, ZN => 
                           n6655);
   U18379 : OAI211_X1 port map( C1 => n6673, C2 => n6672, A => n6655, B => 
                           n6671, ZN => n6656);
   U18380 : INV_X1 port map( A => n6823, ZN => n6819);
   U18381 : INV_X1 port map( A => n7023, ZN => n7024);
   U18382 : XOR2_X1 port map( A => n7771, B => n7712, Z => n6660);
   U18383 : XOR2_X1 port map( A => n7737, B => n7771, Z => n7243);
   U18384 : NAND2_X1 port map( A1 => n6660, A2 => n7243, ZN => n7244);
   U18385 : INV_X1 port map( A => n7014, ZN => n7031);
   U18386 : NAND2_X1 port map( A1 => n634, A2 => n6662, ZN => n6678);
   U18387 : INV_X1 port map( A => n6663, ZN => n6664);
   U18388 : AOI21_X1 port map( B1 => n1039, B2 => n6665, A => n6664, ZN => 
                           n6666);
   U18389 : NAND2_X1 port map( A1 => n6667, A2 => n6668, ZN => n6679);
   U18390 : INV_X1 port map( A => n6669, ZN => n6670);
   U18391 : AOI21_X1 port map( B1 => n6679, B2 => n6671, A => n6670, ZN => 
                           n6674);
   U18392 : INV_X1 port map( A => n7027, ZN => n7030);
   U18393 : OAI22_X1 port map( A1 => n2147, A2 => n7244, B1 => n2230, B2 => 
                           n7243, ZN => n7032);
   U18394 : OAI22_X1 port map( A1 => n771, A2 => n7244, B1 => n2147, B2 => 
                           n7243, ZN => n7705);
   U18395 : XOR2_X1 port map( A => n6687, B => n615, Z => n6688);
   U18396 : INV_X1 port map( A => n7243, ZN => n6690);
   U18397 : NAND2_X1 port map( A1 => n6690, A2 => n2154, ZN => n7726);
   U18398 : INV_X1 port map( A => n7726, ZN => n7007);
   U18399 : INV_X1 port map( A => n7032, ZN => n7010);
   U18400 : NAND2_X1 port map( A1 => n1291, A2 => n7005, ZN => n7021);
   U18401 : INV_X1 port map( A => n7021, ZN => n7239);
   U18402 : NOR2_X1 port map( A1 => n1259, A2 => n7239, ZN => n6828);
   U18403 : OAI22_X1 port map( A1 => n2238, A2 => n7248, B1 => n17239, B2 => 
                           n7247, ZN => n7003);
   U18404 : OAI22_X1 port map( A1 => n2199, A2 => n7258, B1 => n2197, B2 => 
                           n7256, ZN => n6994);
   U18405 : OAI22_X1 port map( A1 => n2208, A2 => n7266, B1 => n2205, B2 => 
                           n7265, ZN => n6984);
   U18406 : OAI22_X1 port map( A1 => n2215, A2 => n7274, B1 => n2213, B2 => 
                           n7272, ZN => n6978);
   U18407 : NOR3_X1 port map( A1 => n570, A2 => n6839, A3 => n1844, ZN => n6699
                           );
   U18408 : NAND2_X1 port map( A1 => n1287, A2 => n6695, ZN => n6837);
   U18409 : INV_X1 port map( A => n6837, ZN => n6698);
   U18410 : NAND2_X1 port map( A1 => n1446, A2 => n6696, ZN => n6834);
   U18412 : OAI22_X1 port map( A1 => n2179, A2 => n7291, B1 => n2185, B2 => 
                           n7283, ZN => n6960);
   U18413 : NAND2_X1 port map( A1 => n6701, A2 => n6700, ZN => n6942);
   U18414 : NAND2_X1 port map( A1 => n6774, A2 => n1314, ZN => n6941);
   U18415 : AOI21_X1 port map( B1 => n6942, B2 => n6941, A => n1876, ZN => 
                           n6771);
   U18416 : INV_X1 port map( A => n6754, ZN => n6702);
   U18417 : NAND2_X1 port map( A1 => n6754, A2 => n6705, ZN => n6918);
   U18418 : OAI21_X1 port map( B1 => n1852, B2 => n1843, A => n6918, ZN => 
                           n6760);
   U18419 : INV_X1 port map( A => n6760, ZN => n6908);
   U18420 : NAND2_X1 port map( A1 => n6747, A2 => n6706, ZN => n6919);
   U18421 : INV_X1 port map( A => n6919, ZN => n6893);
   U18422 : OAI21_X1 port map( B1 => n6708, B2 => n1842, A => n6707, ZN => 
                           n6709);
   U18423 : INV_X1 port map( A => n6709, ZN => n6892);
   U18424 : NAND2_X1 port map( A1 => n6746, A2 => n6710, ZN => n6891);
   U18425 : NOR2_X1 port map( A1 => n6893, A2 => n749, ZN => n6744);
   U18426 : INV_X1 port map( A => n6733, ZN => n6737);
   U18427 : OAI21_X1 port map( B1 => n6734, B2 => n6737, A => n6711, ZN => 
                           n6712);
   U18428 : INV_X1 port map( A => n560, ZN => n6852);
   U18429 : OAI22_X1 port map( A1 => n7670, A2 => n2142, B1 => n2188, B2 => 
                           n7315, ZN => n6872);
   U18430 : NAND2_X1 port map( A1 => n6715, A2 => n2259, ZN => n6714);
   U18431 : MUX2_X1 port map( A => n279, B => n361, S => n2145, Z => n7166);
   U18432 : OAI22_X1 port map( A1 => n7607, A2 => n2137, B1 => n2269, B2 => 
                           n7166, ZN => n6713);
   U18433 : INV_X1 port map( A => n6713, ZN => n6716);
   U18434 : MUX2_X1 port map( A => n6714, B => n2261, S => n6716, Z => n6718);
   U18435 : INV_X1 port map( A => n6715, ZN => n6717);
   U18436 : NAND2_X1 port map( A1 => n6717, A2 => n6716, ZN => n6861);
   U18437 : NAND2_X1 port map( A1 => n6718, A2 => n6861, ZN => n6871);
   U18438 : INV_X1 port map( A => n6871, ZN => n6869);
   U18439 : XOR2_X1 port map( A => n6872, B => n6869, Z => n6727);
   U18440 : INV_X1 port map( A => n6726, ZN => n6722);
   U18441 : OAI21_X1 port map( B1 => n6723, B2 => n6726, A => n6719, ZN => 
                           n6720);
   U18442 : OAI21_X1 port map( B1 => n6722, B2 => n6725, A => n6720, ZN => 
                           n6865);
   U18443 : OAI21_X1 port map( B1 => n6723, B2 => n6722, A => n6721, ZN => 
                           n6724);
   U18444 : OAI21_X1 port map( B1 => n6726, B2 => n6725, A => n6724, ZN => 
                           n6867);
   U18445 : XOR2_X1 port map( A => n6727, B => n6867, Z => n6728);
   U18446 : OAI22_X1 port map( A1 => n8094, A2 => n2225, B1 => n2224, B2 => 
                           n7311, ZN => n6879);
   U18447 : OAI22_X1 port map( A1 => n7792, A2 => n2221, B1 => n2219, B2 => 
                           n7302, ZN => n6895);
   U18448 : INV_X1 port map( A => n6895, ZN => n6854);
   U18449 : XOR2_X1 port map( A => n6879, B => n6854, Z => n6738);
   U18450 : INV_X1 port map( A => n6738, ZN => n6730);
   U18452 : INV_X1 port map( A => n6878, ZN => n6849);
   U18453 : NAND3_X1 port map( A1 => n6849, A2 => n6739, A3 => n6890, ZN => 
                           n6742);
   U18454 : INV_X1 port map( A => n6739, ZN => n6740);
   U18455 : NAND3_X1 port map( A1 => n6740, A2 => n6878, A3 => n6890, ZN => 
                           n6741);
   U18456 : INV_X1 port map( A => n6922, ZN => n6748);
   U18457 : NAND2_X1 port map( A1 => n6747, A2 => n796, ZN => n6923);
   U18458 : OAI21_X1 port map( B1 => n6747, B2 => n6746, A => n6745, ZN => 
                           n6926);
   U18459 : NAND2_X1 port map( A1 => n6923, A2 => n6926, ZN => n6853);
   U18460 : OAI22_X1 port map( A1 => n7923, A2 => n2184, B1 => n2182, B2 => 
                           n7289, ZN => n6949);
   U18461 : INV_X1 port map( A => n6949, ZN => n6947);
   U18462 : OAI22_X1 port map( A1 => n7864, A2 => n2180, B1 => n2217, B2 => 
                           n7294, ZN => n6903);
   U18463 : INV_X1 port map( A => n6903, ZN => n6921);
   U18464 : NAND3_X1 port map( A1 => n6908, A2 => n1454, A3 => n6912, ZN => 
                           n6764);
   U18465 : NAND2_X1 port map( A1 => n6755, A2 => n6754, ZN => n6898);
   U18466 : OAI21_X1 port map( B1 => n5555, B2 => n1887, A => n6752, ZN => 
                           n6753);
   U18467 : INV_X1 port map( A => n1127, ZN => n6758);
   U18468 : INV_X1 port map( A => n6898, ZN => n6756);
   U18469 : NOR2_X1 port map( A1 => n6756, A2 => n6761, ZN => n6757);
   U18470 : AOI22_X1 port map( A1 => n6758, A2 => n1207, B1 => n6757, B2 => 
                           n1127, ZN => n6759);
   U18471 : OAI211_X1 port map( C1 => n1454, C2 => n6898, A => n2244, B => 
                           n6759, ZN => n6763);
   U18472 : NAND3_X1 port map( A1 => n1207, A2 => n976, A3 => n6912, ZN => 
                           n6762);
   U18473 : NAND3_X1 port map( A1 => n6763, A2 => n6764, A3 => n6762, ZN => 
                           n6775);
   U18474 : NOR2_X1 port map( A1 => n6766, A2 => n2268, ZN => n6770);
   U18475 : NAND2_X1 port map( A1 => n1314, A2 => n6765, ZN => n6944);
   U18476 : INV_X1 port map( A => n6942, ZN => n6768);
   U18477 : INV_X1 port map( A => n6941, ZN => n6767);
   U18478 : NAND2_X1 port map( A1 => n6766, A2 => n6776, ZN => n6772);
   U18479 : NOR3_X1 port map( A1 => n6768, A2 => n6767, A3 => n6772, ZN => 
                           n6769);
   U18480 : INV_X1 port map( A => n6772, ZN => n6778);
   U18481 : NAND2_X1 port map( A1 => n6779, A2 => n6780, ZN => n6959);
   U18482 : OAI22_X1 port map( A1 => n2176, A2 => n7285, B1 => n7284, B2 => 
                           n2178, ZN => n6842);
   U18483 : INV_X1 port map( A => n6842, ZN => n6841);
   U18484 : XOR2_X1 port map( A => n1879, B => n6841, Z => n6790);
   U18485 : INV_X1 port map( A => n17152, ZN => n6782);
   U18486 : OAI21_X1 port map( B1 => n6782, B2 => n6784, A => n17182, ZN => 
                           n6846);
   U18487 : NAND2_X1 port map( A1 => n6782, A2 => n6784, ZN => n6847);
   U18488 : INV_X1 port map( A => n6847, ZN => n6787);
   U18489 : NAND2_X1 port map( A1 => n6783, A2 => n6782, ZN => n6961);
   U18490 : NAND2_X1 port map( A1 => n17152, A2 => n6784, ZN => n6957);
   U18491 : OAI211_X1 port map( C1 => n6787, C2 => n2266, A => n6961, B => 
                           n6786, ZN => n6788);
   U18492 : INV_X1 port map( A => n6836, ZN => n6789);
   U18493 : OAI21_X1 port map( B1 => n6796, B2 => n6793, A => n1303, ZN => 
                           n6792);
   U18494 : INV_X1 port map( A => n6792, ZN => n7268);
   U18495 : OAI21_X1 port map( B1 => n6797, B2 => n440, A => n6795, ZN => n7414
                           );
   U18496 : INV_X1 port map( A => n7414, ZN => n6975);
   U18497 : NAND2_X1 port map( A1 => n440, A2 => n6797, ZN => n7415);
   U18498 : INV_X1 port map( A => n7415, ZN => n6974);
   U18499 : INV_X1 port map( A => n6978, ZN => n6976);
   U18502 : NAND2_X1 port map( A1 => n6806, A2 => n1083, ZN => n7427);
   U18503 : NAND2_X1 port map( A1 => n1159, A2 => n6812, ZN => n6830);
   U18504 : AOI21_X1 port map( B1 => n1066, B2 => n6830, A => n1811, ZN => 
                           n6807);
   U18505 : NAND2_X1 port map( A1 => n1159, A2 => n6809, ZN => n6992);
   U18506 : AOI21_X1 port map( B1 => n6992, B2 => n1345, A => n1035, ZN => 
                           n6814);
   U18507 : INV_X1 port map( A => n6994, ZN => n6990);
   U18508 : OAI21_X1 port map( B1 => n6822, B2 => n6819, A => n6815, ZN => 
                           n6816);
   U18509 : OAI21_X1 port map( B1 => n6819, B2 => n6820, A => n6818, ZN => 
                           n6821);
   U18510 : INV_X1 port map( A => n7003, ZN => n7000);
   U18511 : OAI22_X1 port map( A1 => n2240, A2 => n7244, B1 => n2239, B2 => 
                           n7243, ZN => n7022);
   U18512 : NAND2_X1 port map( A1 => n1672, A2 => n7022, ZN => n7240);
   U18513 : NAND2_X1 port map( A1 => n17189, A2 => n1630, ZN => n7238);
   U18514 : INV_X1 port map( A => n7238, ZN => n6827);
   U18515 : AOI21_X1 port map( B1 => n7240, B2 => n6828, A => n6827, ZN => 
                           n7004);
   U18516 : OAI22_X1 port map( A1 => n17240, A2 => n7248, B1 => n2200, B2 => 
                           n7247, ZN => n7453);
   U18517 : NOR2_X1 port map( A1 => n1422, A2 => n1811, ZN => n6831);
   U18518 : NAND2_X1 port map( A1 => n6830, A2 => n1066, ZN => n7250);
   U18519 : NAND2_X1 port map( A1 => n6990, A2 => n6993, ZN => n7251);
   U18520 : AOI21_X1 port map( B1 => n6831, B2 => n7250, A => n962, ZN => n6989
                           );
   U18521 : NOR2_X1 port map( A1 => n7261, A2 => n1815, ZN => n6833);
   U18522 : NAND2_X1 port map( A1 => n1599, A2 => n6984, ZN => n7262);
   U18523 : NAND2_X1 port map( A1 => n6982, A2 => n1415, ZN => n7260);
   U18524 : INV_X1 port map( A => n7260, ZN => n6832);
   U18525 : AOI21_X1 port map( B1 => n579, B2 => n7262, A => n6832, ZN => n6981
                           );
   U18526 : OAI22_X1 port map( A1 => n2213, A2 => n7274, B1 => n2175, B2 => 
                           n7272, ZN => n7420);
   U18527 : OAI21_X1 port map( B1 => n1154, B2 => n1846, A => n1565, ZN => 
                           n6835);
   U18528 : INV_X1 port map( A => n6835, ZN => n7280);
   U18529 : OAI21_X1 port map( B1 => n17192, B2 => n1844, A => n6837, ZN => 
                           n6838);
   U18530 : INV_X1 port map( A => n6838, ZN => n7401);
   U18531 : NOR3_X1 port map( A1 => n7401, A2 => n6839, A3 => n1838, ZN => 
                           n6845);
   U18532 : INV_X1 port map( A => n7400, ZN => n6844);
   U18533 : NOR2_X1 port map( A1 => n1513, A2 => n8229, ZN => n6843);
   U18534 : OAI33_X1 port map( A1 => n7280, A2 => n1792, A3 => n8229, B1 => 
                           n6845, B2 => n6843, B3 => n6844, ZN => n6970);
   U18535 : INV_X1 port map( A => n6960, ZN => n6848);
   U18536 : INV_X1 port map( A => n7287, ZN => n6954);
   U18537 : OAI22_X1 port map( A1 => n7289, A2 => n2184, B1 => n2182, B2 => 
                           n7864, ZN => n7382);
   U18538 : NAND2_X1 port map( A1 => n6921, A2 => n517, ZN => n6901);
   U18539 : INV_X1 port map( A => n6901, ZN => n6917);
   U18540 : INV_X1 port map( A => n6850, ZN => n6851);
   U18541 : NAND2_X1 port map( A1 => n1803, A2 => n6895, ZN => n7308);
   U18542 : OAI21_X1 port map( B1 => n6854, B2 => n1803, A => n6853, ZN => 
                           n7350);
   U18543 : NAND2_X1 port map( A1 => n6854, A2 => n1803, ZN => n7351);
   U18544 : NAND3_X1 port map( A1 => n7350, A2 => n2246, A3 => n7351, ZN => 
                           n6855);
   U18545 : INV_X1 port map( A => n6879, ZN => n6883);
   U18546 : OAI21_X1 port map( B1 => n6880, B2 => n6883, A => n6856, ZN => 
                           n6857);
   U18547 : OAI22_X1 port map( A1 => n7315, A2 => n2192, B1 => n2188, B2 => 
                           n7607, ZN => n7327);
   U18548 : NAND2_X1 port map( A1 => n6861, A2 => n2259, ZN => n6860);
   U18549 : MUX2_X1 port map( A => n280, B => n362, S => n2145, Z => n7515);
   U18550 : OAI22_X1 port map( A1 => n7166, A2 => n2136, B1 => n2269, B2 => 
                           n7515, ZN => n6859);
   U18551 : INV_X1 port map( A => n6859, ZN => n6862);
   U18552 : MUX2_X1 port map( A => n6860, B => n2261, S => n6862, Z => n6864);
   U18553 : INV_X1 port map( A => n6861, ZN => n6863);
   U18554 : NAND2_X1 port map( A1 => n6863, A2 => n6862, ZN => n7317);
   U18555 : NAND2_X1 port map( A1 => n6864, A2 => n7317, ZN => n7326);
   U18556 : INV_X1 port map( A => n7326, ZN => n7329);
   U18557 : XOR2_X1 port map( A => n7327, B => n7329, Z => n6873);
   U18558 : INV_X1 port map( A => n6872, ZN => n6868);
   U18559 : OAI21_X1 port map( B1 => n6869, B2 => n6872, A => n6865, ZN => 
                           n6866);
   U18560 : OAI21_X1 port map( B1 => n6869, B2 => n6868, A => n6867, ZN => 
                           n6870);
   U18561 : OAI21_X1 port map( B1 => n6872, B2 => n6871, A => n6870, ZN => 
                           n7330);
   U18562 : XOR2_X1 port map( A => n6873, B => n7330, Z => n6874);
   U18563 : INV_X1 port map( A => n7342, ZN => n7340);
   U18564 : OAI22_X1 port map( A1 => n7311, A2 => n2226, B1 => n2224, B2 => 
                           n7670, ZN => n7343);
   U18565 : OAI22_X1 port map( A1 => n7302, A2 => n2221, B1 => n2219, B2 => 
                           n8094, ZN => n7357);
   U18566 : INV_X1 port map( A => n7357, ZN => n7355);
   U18567 : XOR2_X1 port map( A => n7343, B => n7355, Z => n6884);
   U18568 : INV_X1 port map( A => n6884, ZN => n6876);
   U18569 : XOR2_X1 port map( A => n6877, B => n6876, Z => n6889);
   U18570 : OAI21_X1 port map( B1 => n6880, B2 => n6879, A => n6878, ZN => 
                           n6881);
   U18572 : INV_X1 port map( A => n7313, ZN => n7304);
   U18573 : XOR2_X1 port map( A => n6884, B => n7340, Z => n6885);
   U18574 : NAND3_X1 port map( A1 => n7304, A2 => n6885, A3 => n6890, ZN => 
                           n6888);
   U18575 : INV_X1 port map( A => n6885, ZN => n6886);
   U18576 : NAND3_X1 port map( A1 => n6886, A2 => n7313, A3 => n6890, ZN => 
                           n6887);
   U18577 : OAI211_X1 port map( C1 => n6890, C2 => n6889, A => n6888, B => 
                           n6887, ZN => n7298);
   U18578 : OAI22_X1 port map( A1 => n7294, A2 => n2180, B1 => n2217, B2 => 
                           n7792, ZN => n7369);
   U18579 : INV_X1 port map( A => n7369, ZN => n7367);
   U18580 : OAI21_X1 port map( B1 => n6893, B2 => n6892, A => n6891, ZN => 
                           n6894);
   U18581 : OAI21_X1 port map( B1 => n1803, B2 => n6895, A => n6894, ZN => 
                           n7309);
   U18582 : INV_X1 port map( A => n7309, ZN => n6896);
   U18583 : NAND2_X1 port map( A1 => n6896, A2 => n6920, ZN => n7297);
   U18584 : NAND3_X1 port map( A1 => n7297, A2 => n1863, A3 => n310, ZN => 
                           n6897);
   U18585 : NAND2_X1 port map( A1 => n6911, A2 => n2244, ZN => n6900);
   U18586 : INV_X1 port map( A => n6900, ZN => n6916);
   U18587 : NOR2_X1 port map( A1 => n1126, A2 => n6900, ZN => n6915);
   U18588 : INV_X1 port map( A => n6904, ZN => n6905);
   U18589 : NAND2_X1 port map( A1 => n6905, A2 => n6903, ZN => n6914);
   U18590 : INV_X1 port map( A => n6914, ZN => n6902);
   U18591 : OAI21_X1 port map( B1 => n1126, B2 => n6902, A => n6901, ZN => 
                           n7365);
   U18592 : INV_X1 port map( A => n6911, ZN => n6907);
   U18593 : NAND2_X1 port map( A1 => n518, A2 => n6903, ZN => n6906);
   U18594 : OAI21_X1 port map( B1 => n1108, B2 => n1850, A => n6906, ZN => 
                           n7300);
   U18595 : OAI22_X1 port map( A1 => n6907, A2 => n6906, B1 => n7300, B2 => 
                           n6911, ZN => n6910);
   U18596 : NOR3_X1 port map( A1 => n6907, A2 => n6908, A3 => n1850, ZN => 
                           n6909);
   U18597 : OAI33_X1 port map( A1 => n6912, A2 => n6911, A3 => n7365, B1 => 
                           n6910, B2 => n6909, B3 => n2244, ZN => n6913);
   U18598 : AOI21_X1 port map( B1 => n1843, B2 => n6918, A => n1852, ZN => 
                           n6938);
   U18599 : NAND2_X1 port map( A1 => n6920, A2 => n6919, ZN => n6929);
   U18600 : INV_X1 port map( A => n6934, ZN => n6924);
   U18601 : NOR3_X1 port map( A1 => n6929, A2 => n749, A3 => n17246, ZN => 
                           n6936);
   U18602 : NAND2_X1 port map( A1 => n6923, A2 => n2246, ZN => n6927);
   U18603 : INV_X1 port map( A => n6927, ZN => n6925);
   U18604 : OAI22_X1 port map( A1 => n6925, A2 => n6924, B1 => n6924, B2 => 
                           n6926, ZN => n6932);
   U18605 : INV_X1 port map( A => n6926, ZN => n6928);
   U18606 : NOR3_X1 port map( A1 => n6928, A2 => n6934, A3 => n6927, ZN => 
                           n6931);
   U18607 : INV_X1 port map( A => n6929, ZN => n6930);
   U18608 : OAI33_X1 port map( A1 => n2246, A2 => n6934, A3 => n6933, B1 => 
                           n6932, B2 => n6931, B3 => n6930, ZN => n6935);
   U18609 : INV_X1 port map( A => n6946, ZN => n6950);
   U18610 : OAI221_X1 port map( B1 => n6946, B2 => n6949, C1 => n1876, C2 => 
                           n6942, A => n6941, ZN => n6943);
   U18611 : OAI21_X1 port map( B1 => n6947, B2 => n6950, A => n6943, ZN => 
                           n7292);
   U18613 : XOR2_X1 port map( A => n6951, B => n17245, Z => n6952);
   U18614 : OAI22_X1 port map( A1 => n2178, A2 => n7285, B1 => n7284, B2 => 
                           n2179, ZN => n7406);
   U18615 : INV_X1 port map( A => n7406, ZN => n7404);
   U18616 : OAI22_X1 port map( A1 => n7283, A2 => n7291, B1 => n2185, B2 => 
                           n7923, ZN => n7393);
   U18617 : INV_X1 port map( A => n7393, ZN => n7391);
   U18618 : NOR2_X1 port map( A1 => n6954, A2 => n6963, ZN => n6968);
   U18619 : NAND2_X1 port map( A1 => n6960, A2 => n6959, ZN => n6955);
   U18620 : INV_X1 port map( A => n6955, ZN => n6962);
   U18621 : NAND3_X1 port map( A1 => n574, A2 => n6955, A3 => n6957, ZN => 
                           n6958);
   U18622 : OAI221_X1 port map( B1 => n6962, B2 => n6961, C1 => n6960, C2 => 
                           n1449, A => n6958, ZN => n7389);
   U18623 : INV_X1 port map( A => n6963, ZN => n6964);
   U18624 : XOR2_X1 port map( A => n1209, B => n6964, Z => n6966);
   U18625 : NOR3_X1 port map( A1 => n2266, A2 => n6964, A3 => n589, ZN => n6965
                           );
   U18626 : AOI221_X1 port map( B1 => n6968, B2 => n6967, C1 => n6966, C2 => 
                           n2266, A => n6965, ZN => n6969);
   U18627 : NOR2_X1 port map( A1 => n7268, A2 => n1814, ZN => n6972);
   U18628 : NAND2_X1 port map( A1 => n6977, A2 => n6976, ZN => n7267);
   U18629 : INV_X1 port map( A => n7267, ZN => n6971);
   U18630 : AOI21_X1 port map( B1 => n6972, B2 => n7269, A => n6971, ZN => 
                           n6973);
   U18631 : NOR2_X1 port map( A1 => n6974, A2 => n6975, ZN => n6979);
   U18632 : NAND2_X1 port map( A1 => n6976, A2 => n1447, ZN => n7413);
   U18633 : AOI21_X1 port map( B1 => n6979, B2 => n7413, A => n1831, ZN => 
                           n6980);
   U18634 : OAI22_X1 port map( A1 => n2204, A2 => n7266, B1 => n2215, B2 => 
                           n7265, ZN => n7433);
   U18635 : INV_X1 port map( A => n7433, ZN => n7430);
   U18636 : INV_X1 port map( A => n7445, ZN => n7443);
   U18637 : OAI22_X1 port map( A1 => n2196, A2 => n7258, B1 => n2209, B2 => 
                           n7256, ZN => n7446);
   U18638 : NOR2_X1 port map( A1 => n1786, A2 => n559, ZN => n6995);
   U18639 : NAND2_X1 port map( A1 => n6992, A2 => n1345, ZN => n7441);
   U18640 : AOI21_X1 port map( B1 => n6995, B2 => n7441, A => n1179, ZN => 
                           n6996);
   U18641 : OAI21_X1 port map( B1 => n1732, B2 => n7000, A => n599, ZN => n7001
                           );
   U18642 : OAI22_X1 port map( A1 => n2138, A2 => n7244, B1 => n2238, B2 => 
                           n7243, ZN => n7465);
   U18643 : INV_X1 port map( A => n7005, ZN => n7025);
   U18644 : NAND2_X1 port map( A1 => n7006, A2 => n7007, ZN => n7708);
   U18645 : OAI21_X1 port map( B1 => n1639, B2 => n1612, A => n7708, ZN => 
                           n7008);
   U18646 : OAI21_X1 port map( B1 => n7705, B2 => n7009, A => n7008, ZN => 
                           n7033);
   U18647 : OAI21_X1 port map( B1 => n1536, B2 => n7010, A => n7033, ZN => 
                           n7011);
   U18648 : OAI21_X1 port map( B1 => n7025, B2 => n1291, A => n595, ZN => n7459
                           );
   U18649 : NAND2_X1 port map( A1 => n7025, A2 => n457, ZN => n7460);
   U18650 : NAND2_X1 port map( A1 => n1174, A2 => n1630, ZN => n7458);
   U18651 : AOI21_X1 port map( B1 => n7015, B2 => n7458, A => n1828, ZN => 
                           n7016);
   U18652 : OAI22_X1 port map( A1 => n2229, A2 => n7237, B1 => n2227, B2 => 
                           n7236, ZN => n7051);
   U18653 : INV_X1 port map( A => n7051, ZN => n7054);
   U18654 : OAI22_X1 port map( A1 => n2147, A2 => n7237, B1 => n2230, B2 => 
                           n7236, ZN => n7045);
   U18655 : INV_X1 port map( A => n7045, ZN => n7059);
   U18656 : OAI22_X1 port map( A1 => n2132, A2 => n7237, B1 => n2147, B2 => 
                           n7236, ZN => n7641);
   U18657 : INV_X1 port map( A => n7641, ZN => n7039);
   U18658 : INV_X1 port map( A => n7236, ZN => n7035);
   U18659 : NAND2_X1 port map( A1 => n7035, A2 => n2154, ZN => n7679);
   U18660 : INV_X1 port map( A => n7679, ZN => n7040);
   U18661 : OAI21_X1 port map( B1 => n1347, B2 => n7641, A => n1796, ZN => 
                           n7036);
   U18662 : OAI21_X1 port map( B1 => n7039, B2 => n7041, A => n7036, ZN => 
                           n7057);
   U18663 : OAI21_X1 port map( B1 => n1723, B2 => n7045, A => n7057, ZN => 
                           n7037);
   U18664 : OAI21_X1 port map( B1 => n7059, B2 => n7044, A => n7037, ZN => 
                           n7052);
   U18665 : OAI21_X1 port map( B1 => n7051, B2 => n1192, A => n7052, ZN => 
                           n7038);
   U18666 : OAI21_X1 port map( B1 => n578, B2 => n7059, A => n7058, ZN => n7043
                           );
   U18667 : INV_X1 port map( A => n7478, ZN => n7474);
   U18668 : INV_X1 port map( A => n1507, ZN => n7073);
   U18669 : OAI22_X1 port map( A1 => n771, A2 => n7231, B1 => n2147, B2 => 
                           n7230, ZN => n7066);
   U18670 : NAND2_X1 port map( A1 => n7053, A2 => n7471, ZN => n7065);
   U18671 : NAND2_X1 port map( A1 => n7055, A2 => n7647, ZN => n7067);
   U18672 : NAND2_X1 port map( A1 => n7067, A2 => n1339, ZN => n7577);
   U18673 : INV_X1 port map( A => n7230, ZN => n7056);
   U18674 : NAND2_X1 port map( A1 => n7056, A2 => n2154, ZN => n7588);
   U18675 : INV_X1 port map( A => n7588, ZN => n7069);
   U18676 : INV_X1 port map( A => n7066, ZN => n7576);
   U18677 : AOI21_X1 port map( B1 => n7065, B2 => n7067, A => n7576, ZN => 
                           n7062);
   U18678 : OAI22_X1 port map( A1 => n7577, A2 => n7066, B1 => n7062, B2 => 
                           n1808, ZN => n7063);
   U18679 : INV_X1 port map( A => n877, ZN => n7488);
   U18680 : NAND2_X1 port map( A1 => n7064, A2 => n7581, ZN => n7508);
   U18681 : NAND3_X1 port map( A1 => n7065, A2 => n1336, A3 => n7066, ZN => 
                           n7070);
   U18682 : NAND2_X1 port map( A1 => n1235, A2 => n7508, ZN => n7496);
   U18683 : MUX2_X1 port map( A => n7076, B => n7075, S => n527, Z => n7516);
   U18684 : NAND2_X1 port map( A1 => n371, A2 => n2154, ZN => n7548);
   U18685 : INV_X1 port map( A => n7548, ZN => n7547);
   U18686 : NAND2_X1 port map( A1 => n1895, A2 => n8325, ZN => n7980);
   U18687 : INV_X1 port map( A => n7980, ZN => n7550);
   U18688 : MUX2_X1 port map( A => n7079, B => n7078, S => n526, Z => n7225);
   U18689 : INV_X1 port map( A => n7225, ZN => n7495);
   U18690 : NAND2_X1 port map( A1 => i_ALU_OP_0_port, A2 => n7080, ZN => n8205)
                           ;
   U18691 : NAND2_X1 port map( A1 => i_ALU_OP_1_port, A2 => n7081, ZN => n7083)
                           ;
   U18692 : NAND2_X1 port map( A1 => n2985, A2 => n8322, ZN => n7970);
   U18693 : NAND2_X1 port map( A1 => DataPath_ALUhw_BWISE_n72, A2 => n8322, ZN 
                           => n7969);
   U18694 : MUX2_X1 port map( A => n7082, B => n363, S => n2145, Z => n7193);
   U18695 : INV_X1 port map( A => n7193, ZN => n8049);
   U18696 : MUX2_X1 port map( A => n2187, B => n7969, S => n8049, Z => n7224);
   U18697 : NAND2_X1 port map( A1 => DataPath_ALUhw_BWISE_n71, A2 => n8322, ZN 
                           => n7965);
   U18698 : MUX2_X1 port map( A => n7965, B => n2187, S => n8049, Z => n7223);
   U18699 : NAND2_X1 port map( A1 => n12932, A2 => n2272, ZN => n7568);
   U18700 : INV_X1 port map( A => n7568, ZN => n7605);
   U18701 : XOR2_X1 port map( A => n7516, B => n259, Z => n7088);
   U18702 : INV_X1 port map( A => n7515, ZN => n8058);
   U18703 : XOR2_X1 port map( A => n7088, B => n8058, Z => n7096);
   U18704 : XOR2_X1 port map( A => n7579, B => n259, Z => n7085);
   U18705 : INV_X1 port map( A => n7166, ZN => n8067);
   U18706 : XOR2_X1 port map( A => n7085, B => n8067, Z => n7566);
   U18707 : XOR2_X1 port map( A => n7608, B => n259, Z => n7094);
   U18708 : INV_X1 port map( A => n7094, ZN => n7084);
   U18709 : INV_X1 port map( A => n7607, ZN => n8079);
   U18710 : NAND2_X1 port map( A1 => n7084, A2 => n8079, ZN => n7567);
   U18711 : INV_X1 port map( A => n7085, ZN => n7086);
   U18712 : NAND2_X1 port map( A1 => n7086, A2 => n8067, ZN => n7095);
   U18713 : OAI21_X1 port map( B1 => n7566, B2 => n7567, A => n7095, ZN => 
                           n7087);
   U18714 : INV_X1 port map( A => n7087, ZN => n7521);
   U18715 : INV_X1 port map( A => n7088, ZN => n7089);
   U18716 : NAND2_X1 port map( A1 => n7089, A2 => n8058, ZN => n7097);
   U18717 : OAI21_X1 port map( B1 => n7096, B2 => n7521, A => n7097, ZN => 
                           n7092);
   U18718 : XOR2_X1 port map( A => n7193, B => n259, Z => n7090);
   U18719 : XOR2_X1 port map( A => n7090, B => n7495, Z => n7100);
   U18720 : INV_X1 port map( A => n7100, ZN => n7091);
   U18721 : XOR2_X1 port map( A => n7092, B => n7091, Z => n7221);
   U18722 : INV_X1 port map( A => n12932, ZN => n7093);
   U18723 : NAND2_X1 port map( A1 => n2272, A2 => n7093, ZN => n7572);
   U18724 : INV_X1 port map( A => n7572, ZN => n7606);
   U18725 : XOR2_X1 port map( A => n7094, B => n8079, Z => n7603);
   U18726 : OAI21_X1 port map( B1 => n7566, B2 => n369, A => n7095, ZN => n7522
                           );
   U18727 : INV_X1 port map( A => n7096, ZN => n7524);
   U18728 : INV_X1 port map( A => n7097, ZN => n7098);
   U18729 : AOI21_X1 port map( B1 => n7522, B2 => n7524, A => n7098, ZN => 
                           n7099);
   U18730 : XOR2_X1 port map( A => n7100, B => n7099, Z => n7220);
   U18731 : NAND3_X1 port map( A1 => n259, A2 => n1208, A3 => n2130, ZN => 
                           n8032);
   U18732 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n155, A2 => 
                           n8032, ZN => n7697);
   U18733 : OAI22_X1 port map( A1 => n2196, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n7283, B2 => 
                           n7207, ZN => n7101);
   U18734 : INV_X1 port map( A => n7101, ZN => n7988);
   U18735 : OAI22_X1 port map( A1 => n7283, A2 => n4136, B1 => n7311, B2 => 
                           n4131, ZN => n7102);
   U18736 : INV_X1 port map( A => n7102, ZN => n7695);
   U18737 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n641, ZN => n7103);
   U18738 : NAND2_X1 port map( A1 => n8049, A2 => n7103, ZN => n7203);
   U18739 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n7311, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n2147, A => n7203, ZN => n8117);
   U18740 : NAND2_X1 port map( A1 => n8117, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n478, ZN => n7107);
   U18741 : OAI221_X1 port map( B1 => n11497, B2 => n7988, C1 => n2275, C2 => 
                           n7695, A => n7107, ZN => n7111);
   U18742 : INV_X1 port map( A => n7111, ZN => n7106);
   U18743 : OAI22_X1 port map( A1 => n2147, A2 => n4138, B1 => n2197, B2 => 
                           n4131, ZN => n7104);
   U18744 : INV_X1 port map( A => n7104, ZN => n8002);
   U18745 : OAI22_X1 port map( A1 => n2277, A2 => n7695, B1 => n2273, B2 => 
                           n8002, ZN => n7105);
   U18746 : INV_X1 port map( A => n7105, ZN => n7998);
   U18747 : OAI22_X1 port map( A1 => n2276, A2 => n7106, B1 => n2273, B2 => 
                           n7998, ZN => n7995);
   U18748 : INV_X1 port map( A => n7995, ZN => n7696);
   U18749 : NAND3_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n548, A2 => 
                           n8181, A3 => n804, ZN => n7997);
   U18750 : NAND3_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n349, A2 => 
                           n8181, A3 => n2250, ZN => n7144);
   U18751 : INV_X1 port map( A => n7144, ZN => n7210);
   U18752 : OAI22_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n597, A2 => 
                           n2147, B1 => DataPath_ALUhw_SHIFTER_HW_n576, B2 => 
                           n7311, ZN => n8119);
   U18753 : INV_X1 port map( A => n2134, ZN => n8043);
   U18754 : INV_X1 port map( A => n8117, ZN => n7690);
   U18755 : OAI22_X1 port map( A1 => n2196, A2 => n4139, B1 => n7283, B2 => 
                           n4131, ZN => n7993);
   U18756 : INV_X1 port map( A => n7993, ZN => n7689);
   U18757 : OAI22_X1 port map( A1 => n2276, A2 => n7690, B1 => n2273, B2 => 
                           n7689, ZN => n7693);
   U18758 : INV_X1 port map( A => n7693, ZN => n7691);
   U18759 : OAI22_X1 port map( A1 => n2196, A2 => n7207, B1 => n7283, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8126);
   U18760 : INV_X1 port map( A => n8126, ZN => n7108);
   U18761 : OAI211_X1 port map( C1 => n2274, C2 => n7691, A => n7108, B => 
                           n7107, ZN => n7692);
   U18762 : AOI22_X1 port map( A1 => n7210, A2 => n8119, B1 => n8043, B2 => 
                           n7692, ZN => n7113);
   U18763 : NAND2_X1 port map( A1 => n818, A2 => n7109, ZN => n8037);
   U18764 : INV_X1 port map( A => n8037, ZN => n7994);
   U18765 : NAND2_X1 port map( A1 => n7994, A2 => n259, ZN => n8082);
   U18766 : INV_X1 port map( A => n8082, ZN => n8118);
   U18767 : INV_X1 port map( A => n8089, ZN => n8116);
   U18768 : NAND2_X1 port map( A1 => n4136, A2 => n7994, ZN => n8102);
   U18769 : NAND2_X1 port map( A1 => n11499, A2 => n8102, ZN => n7211);
   U18770 : AOI222_X1 port map( A1 => n8118, A2 => n7709, B1 => n8116, B2 => 
                           n7111, C1 => n7211, C2 => n8117, ZN => n7112);
   U18771 : OAI211_X1 port map( C1 => n7696, C2 => n7997, A => n7113, B => 
                           n7112, ZN => n7563);
   U18772 : OAI22_X1 port map( A1 => n2208, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n7923, B2 => 
                           n7207, ZN => n7114);
   U18773 : INV_X1 port map( A => n7114, ZN => n7944);
   U18774 : OAI22_X1 port map( A1 => n7923, A2 => n4139, B1 => n7670, B2 => 
                           n4131, ZN => n7115);
   U18775 : INV_X1 port map( A => n7115, ZN => n7665);
   U18776 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n7670, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n2230, A => n7203, ZN => n8109);
   U18777 : NAND2_X1 port map( A1 => n8109, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n478, ZN => n7119);
   U18778 : OAI221_X1 port map( B1 => n11497, B2 => n7944, C1 => n2275, C2 => 
                           n7665, A => n7119, ZN => n7121);
   U18779 : INV_X1 port map( A => n7121, ZN => n7118);
   U18780 : OAI22_X1 port map( A1 => n2230, A2 => n4139, B1 => n2209, B2 => 
                           n4131, ZN => n7116);
   U18781 : INV_X1 port map( A => n7116, ZN => n8006);
   U18782 : OAI22_X1 port map( A1 => n2276, A2 => n7665, B1 => n2274, B2 => 
                           n8006, ZN => n7117);
   U18783 : INV_X1 port map( A => n7117, ZN => n7950);
   U18784 : OAI22_X1 port map( A1 => n2276, A2 => n7118, B1 => n2274, B2 => 
                           n7950, ZN => n7948);
   U18785 : INV_X1 port map( A => n7948, ZN => n7666);
   U18786 : OAI22_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n597, A2 => 
                           n2229, B1 => DataPath_ALUhw_SHIFTER_HW_n576, B2 => 
                           n7670, ZN => n8110);
   U18787 : INV_X1 port map( A => n8109, ZN => n7659);
   U18788 : OAI22_X1 port map( A1 => n2208, A2 => n4138, B1 => n7923, B2 => 
                           n4131, ZN => n7947);
   U18789 : INV_X1 port map( A => n7947, ZN => n7660);
   U18790 : OAI22_X1 port map( A1 => n7659, A2 => n7991, B1 => n7660, B2 => 
                           n7989, ZN => n7663);
   U18791 : INV_X1 port map( A => n7663, ZN => n7661);
   U18792 : OAI22_X1 port map( A1 => n2208, A2 => n7207, B1 => n7923, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8114);
   U18793 : INV_X1 port map( A => n8114, ZN => n7120);
   U18794 : OAI211_X1 port map( C1 => n2274, C2 => n7661, A => n7120, B => 
                           n7119, ZN => n7662);
   U18795 : AOI22_X1 port map( A1 => n7210, A2 => n8110, B1 => n8043, B2 => 
                           n7662, ZN => n7123);
   U18796 : AOI222_X1 port map( A1 => n8118, A2 => n7677, B1 => n8116, B2 => 
                           n7121, C1 => n7211, C2 => n8109, ZN => n7122);
   U18797 : OAI211_X1 port map( C1 => n7666, C2 => n7997, A => n7123, B => 
                           n7122, ZN => n7536);
   U18798 : INV_X1 port map( A => n1769, ZN => n8310);
   U18799 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n7515, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n2238, A => n7203, ZN => n7132);
   U18800 : INV_X1 port map( A => n7132, ZN => n8061);
   U18801 : OAI22_X1 port map( A1 => n2175, A2 => n4138, B1 => n7792, B2 => 
                           n259, ZN => n7813);
   U18802 : INV_X1 port map( A => n7813, ZN => n7526);
   U18803 : OAI22_X1 port map( A1 => n2276, A2 => n8061, B1 => n2274, B2 => 
                           n7526, ZN => n7530);
   U18804 : INV_X1 port map( A => n7530, ZN => n7528);
   U18805 : OAI22_X1 port map( A1 => n2175, A2 => n7207, B1 => n7792, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8057);
   U18806 : INV_X1 port map( A => n8057, ZN => n7124);
   U18807 : NAND2_X1 port map( A1 => n7132, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n478, ZN => n7127);
   U18808 : OAI211_X1 port map( C1 => n2274, C2 => n7528, A => n7124, B => 
                           n7127, ZN => n7529);
   U18809 : INV_X1 port map( A => n7529, ZN => n7135);
   U18810 : OAI21_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n576, B2 => 
                           n7144, A => n8082, ZN => n7164);
   U18811 : AOI22_X1 port map( A1 => n368, A2 => n1933, B1 => n7164, B2 => 
                           n8058, ZN => n7134);
   U18812 : INV_X1 port map( A => n7997, ZN => n8034);
   U18813 : OAI22_X1 port map( A1 => n2176, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n7792, B2 => 
                           n7207, ZN => n7125);
   U18814 : INV_X1 port map( A => n7125, ZN => n7811);
   U18815 : OAI22_X1 port map( A1 => n7792, A2 => n4138, B1 => n7515, B2 => 
                           n259, ZN => n7126);
   U18816 : INV_X1 port map( A => n7126, ZN => n7532);
   U18817 : OAI221_X1 port map( B1 => n11497, B2 => n7811, C1 => n2275, C2 => 
                           n7532, A => n7127, ZN => n7131);
   U18818 : INV_X1 port map( A => n7131, ZN => n7130);
   U18819 : OAI22_X1 port map( A1 => n2238, A2 => n4136, B1 => n2176, B2 => 
                           n259, ZN => n7128);
   U18820 : INV_X1 port map( A => n7128, ZN => n8014);
   U18821 : OAI22_X1 port map( A1 => n2276, A2 => n7532, B1 => n2274, B2 => 
                           n8014, ZN => n7129);
   U18822 : INV_X1 port map( A => n7129, ZN => n7815);
   U18823 : OAI22_X1 port map( A1 => n2276, A2 => n7130, B1 => n2274, B2 => 
                           n7815, ZN => n7525);
   U18824 : AOI222_X1 port map( A1 => n7211, A2 => n7132, B1 => n8034, B2 => 
                           n7525, C1 => n8116, C2 => n7131, ZN => n7133);
   U18825 : OAI211_X1 port map( C1 => n7135, C2 => n2134, A => n7134, B => 
                           n7133, ZN => n7215);
   U18826 : OAI22_X1 port map( A1 => n2199, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n2179, B2 => 
                           n7207, ZN => n7136);
   U18827 : INV_X1 port map( A => n7136, ZN => n7982);
   U18828 : OAI22_X1 port map( A1 => n2179, A2 => n4139, B1 => n8094, B2 => 
                           n4131, ZN => n7722);
   U18829 : INV_X1 port map( A => n7722, ZN => n7139);
   U18830 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n8094, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n2132, A => n7203, ZN => n7146);
   U18831 : NAND2_X1 port map( A1 => n7146, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n478, ZN => n7143);
   U18832 : OAI221_X1 port map( B1 => n11497, B2 => n7982, C1 => n2274, C2 => 
                           n7139, A => n7143, ZN => n7137);
   U18833 : INV_X1 port map( A => n7137, ZN => n7148);
   U18834 : OAI22_X1 port map( A1 => n771, A2 => n4138, B1 => n2200, B2 => 
                           n4131, ZN => n7138);
   U18835 : INV_X1 port map( A => n7138, ZN => n8038);
   U18836 : OAI22_X1 port map( A1 => n2276, A2 => n7139, B1 => n2274, B2 => 
                           n8038, ZN => n7140);
   U18837 : INV_X1 port map( A => n7140, ZN => n7986);
   U18838 : OAI22_X1 port map( A1 => n2276, A2 => n7148, B1 => n2274, B2 => 
                           n7986, ZN => n7141);
   U18839 : INV_X1 port map( A => n7141, ZN => n7987);
   U18840 : INV_X1 port map( A => n7146, ZN => n7721);
   U18841 : OAI22_X1 port map( A1 => n2199, A2 => n4138, B1 => n2179, B2 => 
                           n4131, ZN => n7984);
   U18842 : INV_X1 port map( A => n7984, ZN => n7720);
   U18843 : OAI22_X1 port map( A1 => n7721, A2 => n7991, B1 => n7720, B2 => 
                           n7989, ZN => n7142);
   U18844 : INV_X1 port map( A => n7142, ZN => n7725);
   U18845 : OAI22_X1 port map( A1 => n2199, A2 => n7207, B1 => n2179, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8033);
   U18846 : INV_X1 port map( A => n8033, ZN => n8093);
   U18847 : OAI211_X1 port map( C1 => n2274, C2 => n7725, A => n8093, B => 
                           n7143, ZN => n7723);
   U18848 : AOI21_X1 port map( B1 => n7144, B2 => n8082, A => n8094, ZN => 
                           n7145);
   U18849 : AOI221_X1 port map( B1 => n8043, B2 => n7723, C1 => n7211, C2 => 
                           n7146, A => n7145, ZN => n7147);
   U18850 : OAI221_X1 port map( B1 => n7987, B2 => n7997, C1 => n7148, C2 => 
                           n8089, A => n7147, ZN => n7561);
   U18851 : AOI22_X1 port map( A1 => n7215, A2 => n259, B1 => n7561, B2 => 
                           n4135, ZN => n7162);
   U18852 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n7607, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n2240, A => n7203, ZN => n7157);
   U18853 : INV_X1 port map( A => n7157, ZN => n8083);
   U18854 : OAI22_X1 port map( A1 => n2215, A2 => n4138, B1 => n7864, B2 => 
                           n4131, ZN => n7876);
   U18855 : INV_X1 port map( A => n7876, ZN => n7590);
   U18856 : OAI22_X1 port map( A1 => n8083, A2 => n7991, B1 => n7590, B2 => 
                           n7989, ZN => n7593);
   U18857 : INV_X1 port map( A => n7593, ZN => n7591);
   U18858 : OAI22_X1 port map( A1 => n2215, A2 => n7207, B1 => n7864, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8078);
   U18859 : INV_X1 port map( A => n8078, ZN => n7149);
   U18860 : NAND2_X1 port map( A1 => n7157, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n478, ZN => n7152);
   U18861 : OAI211_X1 port map( C1 => n2274, C2 => n7591, A => n7149, B => 
                           n7152, ZN => n7592);
   U18862 : INV_X1 port map( A => n7592, ZN => n7160);
   U18863 : AOI22_X1 port map( A1 => n368, A2 => n2241, B1 => n7164, B2 => 
                           n8079, ZN => n7159);
   U18864 : OAI22_X1 port map( A1 => n2215, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n7864, B2 => 
                           n7207, ZN => n7150);
   U18865 : INV_X1 port map( A => n7150, ZN => n7874);
   U18866 : OAI22_X1 port map( A1 => n7864, A2 => n4138, B1 => n7607, B2 => 
                           n4131, ZN => n7151);
   U18867 : INV_X1 port map( A => n7151, ZN => n7595);
   U18868 : OAI221_X1 port map( B1 => n11497, B2 => n7874, C1 => n2275, C2 => 
                           n7595, A => n7152, ZN => n7156);
   U18869 : INV_X1 port map( A => n7156, ZN => n7155);
   U18870 : OAI22_X1 port map( A1 => n2240, A2 => n4137, B1 => n2215, B2 => 
                           n4131, ZN => n7153);
   U18871 : INV_X1 port map( A => n7153, ZN => n8018);
   U18872 : OAI22_X1 port map( A1 => n2276, A2 => n7595, B1 => n2274, B2 => 
                           n8018, ZN => n7154);
   U18873 : INV_X1 port map( A => n7154, ZN => n7878);
   U18874 : OAI22_X1 port map( A1 => n2276, A2 => n7155, B1 => n2274, B2 => 
                           n7878, ZN => n7589);
   U18875 : AOI222_X1 port map( A1 => n7211, A2 => n7157, B1 => n8034, B2 => 
                           n7589, C1 => n8116, C2 => n7156, ZN => n7158);
   U18876 : OAI211_X1 port map( C1 => n7160, C2 => n2134, A => n7159, B => 
                           n7158, ZN => n7535);
   U18877 : AOI22_X1 port map( A1 => n7536, A2 => n259, B1 => n7535, B2 => 
                           n4135, ZN => n7161);
   U18878 : MUX2_X1 port map( A => n7162, B => n7161, S => n2130, Z => n7199);
   U18879 : NAND2_X1 port map( A1 => n2264, A2 => n17179, ZN => n7514);
   U18880 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n7166, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n2239, A => n7203, ZN => n7173);
   U18881 : INV_X1 port map( A => n7173, ZN => n8070);
   U18882 : OAI22_X1 port map( A1 => n2213, A2 => n4137, B1 => n7294, B2 => 
                           n4131, ZN => n7845);
   U18883 : INV_X1 port map( A => n7845, ZN => n7554);
   U18884 : OAI22_X1 port map( A1 => n2276, A2 => n8070, B1 => n2274, B2 => 
                           n7554, ZN => n7558);
   U18885 : INV_X1 port map( A => n7558, ZN => n7556);
   U18886 : OAI22_X1 port map( A1 => n2213, A2 => n7207, B1 => n7294, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8066);
   U18887 : INV_X1 port map( A => n8066, ZN => n7163);
   U18888 : NAND2_X1 port map( A1 => n7173, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n478, ZN => n7168);
   U18889 : OAI211_X1 port map( C1 => n2274, C2 => n7556, A => n7163, B => 
                           n7168, ZN => n7557);
   U18890 : INV_X1 port map( A => n7557, ZN => n7176);
   U18891 : AOI22_X1 port map( A1 => n368, A2 => n788, B1 => n7164, B2 => n8067
                           , ZN => n7175);
   U18892 : OAI22_X1 port map( A1 => n2213, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n7294, B2 => 
                           n7207, ZN => n7165);
   U18893 : INV_X1 port map( A => n7165, ZN => n7843);
   U18894 : OAI22_X1 port map( A1 => n7294, A2 => n4137, B1 => n7166, B2 => 
                           n4131, ZN => n7167);
   U18895 : INV_X1 port map( A => n7167, ZN => n7560);
   U18896 : OAI221_X1 port map( B1 => n11497, B2 => n7843, C1 => n2275, C2 => 
                           n7560, A => n7168, ZN => n7172);
   U18897 : INV_X1 port map( A => n7172, ZN => n7171);
   U18898 : OAI22_X1 port map( A1 => n2138, A2 => n4137, B1 => n2213, B2 => 
                           n4131, ZN => n7169);
   U18899 : INV_X1 port map( A => n7169, ZN => n8029);
   U18900 : OAI22_X1 port map( A1 => n2277, A2 => n7560, B1 => n2273, B2 => 
                           n8029, ZN => n7170);
   U18901 : INV_X1 port map( A => n7170, ZN => n7847);
   U18902 : OAI22_X1 port map( A1 => n2277, A2 => n7171, B1 => n2273, B2 => 
                           n7847, ZN => n7553);
   U18903 : AOI222_X1 port map( A1 => n7211, A2 => n7173, B1 => n8034, B2 => 
                           n7553, C1 => n8116, C2 => n7172, ZN => n7174);
   U18904 : OAI211_X1 port map( C1 => n7176, C2 => n2134, A => n7175, B => 
                           n7174, ZN => n7177);
   U18905 : INV_X1 port map( A => n7177, ZN => n8316);
   U18906 : NAND3_X1 port map( A1 => n4136, A2 => n1208, A3 => n2130, ZN => 
                           n8026);
   U18907 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n192, A2 => 
                           n8026, ZN => n7953);
   U18908 : INV_X1 port map( A => n7953, ZN => n7198);
   U18909 : OAI22_X1 port map( A1 => n7302, A2 => n4137, B1 => n7193, B2 => 
                           n4131, ZN => n7178);
   U18910 : INV_X1 port map( A => n7178, ZN => n7190);
   U18911 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n7193, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n17239, A => n7203, ZN => n7182);
   U18912 : INV_X1 port map( A => n7182, ZN => n8052);
   U18913 : OAI22_X1 port map( A1 => n2177, A2 => n4137, B1 => n7302, B2 => 
                           n4131, ZN => n7179);
   U18914 : INV_X1 port map( A => n7179, ZN => n7783);
   U18915 : OAI22_X1 port map( A1 => n8052, A2 => n7991, B1 => n7783, B2 => 
                           n7989, ZN => n7180);
   U18916 : INV_X1 port map( A => n7180, ZN => n7189);
   U18917 : OAI22_X1 port map( A1 => n2178, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n7302, B2 => 
                           n7207, ZN => n7181);
   U18918 : INV_X1 port map( A => n7181, ZN => n7779);
   U18919 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n478, A2 => 
                           n7182, ZN => n7186);
   U18920 : OAI211_X1 port map( C1 => n2274, C2 => n7190, A => n7779, B => 
                           n7186, ZN => n7192);
   U18921 : INV_X1 port map( A => n7192, ZN => n7185);
   U18922 : OAI22_X1 port map( A1 => n17240, A2 => n4137, B1 => n2177, B2 => 
                           n4131, ZN => n7183);
   U18923 : INV_X1 port map( A => n7183, ZN => n8010);
   U18924 : OAI22_X1 port map( A1 => n2277, A2 => n7190, B1 => n2273, B2 => 
                           n8010, ZN => n7184);
   U18925 : INV_X1 port map( A => n7184, ZN => n7784);
   U18926 : OAI22_X1 port map( A1 => n2277, A2 => n7185, B1 => n2273, B2 => 
                           n7784, ZN => n7781);
   U18927 : OAI222_X1 port map( A1 => n7783, A2 => n7991, B1 => n8052, B2 => 
                           n4135, C1 => n17240, C2 => n266, ZN => n8008);
   U18928 : INV_X1 port map( A => n8008, ZN => n8046);
   U18929 : OAI22_X1 port map( A1 => n2277, A2 => n7189, B1 => n2273, B2 => 
                           n8046, ZN => n8007);
   U18930 : OAI22_X1 port map( A1 => n2177, A2 => n7207, B1 => n7302, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8048);
   U18931 : INV_X1 port map( A => n8048, ZN => n7187);
   U18932 : OAI211_X1 port map( C1 => n2274, C2 => n7189, A => n7187, B => 
                           n7186, ZN => n7191);
   U18933 : AOI222_X1 port map( A1 => n8043, A2 => n7781, B1 => n8034, B2 => 
                           n8007, C1 => n7191, C2 => n8073, ZN => n7188);
   U18934 : OAI221_X1 port map( B1 => n7190, B2 => n8037, C1 => n7189, C2 => 
                           n8089, A => n7188, ZN => n7596);
   U18935 : INV_X1 port map( A => n7596, ZN => n8320);
   U18936 : AOI222_X1 port map( A1 => n8116, A2 => n7192, B1 => n8043, B2 => 
                           n7191, C1 => n8034, C2 => n7781, ZN => n7194);
   U18937 : OAI222_X1 port map( A1 => n259, A2 => n8320, B1 => n4135, B2 => 
                           n7194, C1 => n7193, C2 => n8082, ZN => n7195);
   U18938 : NAND3_X1 port map( A1 => n1861, A2 => n7196, A3 => n7195, ZN => 
                           n7197);
   U18939 : OAI221_X1 port map( B1 => n7199, B2 => n7514, C1 => n8316, C2 => 
                           n7198, A => n7197, ZN => n7200);
   U18940 : AOI221_X1 port map( B1 => n7697, B2 => n7563, C1 => n7536, C2 => 
                           n8310, A => n7200, ZN => n7218);
   U18941 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n191, ZN => n8309);
   U18942 : OAI22_X1 port map( A1 => n2204, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, B1 => n7289, B2 => 
                           n7207, ZN => n7201);
   U18943 : INV_X1 port map( A => n7201, ZN => n7909);
   U18944 : OAI22_X1 port map( A1 => n7289, A2 => n4137, B1 => n7315, B2 => 
                           n4131, ZN => n7202);
   U18945 : INV_X1 port map( A => n7202, ZN => n7631);
   U18946 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n7315, C1 => DataPath_ALUhw_SHIFTER_HW_n598, C2 => 
                           n2227, A => n7203, ZN => n8101);
   U18947 : NAND2_X1 port map( A1 => n8101, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n478, ZN => n7208);
   U18948 : OAI221_X1 port map( B1 => n11497, B2 => n7909, C1 => n2275, C2 => 
                           n7631, A => n7208, ZN => n7212);
   U18949 : INV_X1 port map( A => n7212, ZN => n7206);
   U18950 : OAI22_X1 port map( A1 => n2227, A2 => n4136, B1 => n2205, B2 => 
                           n4131, ZN => n7204);
   U18951 : INV_X1 port map( A => n7204, ZN => n8024);
   U18952 : OAI22_X1 port map( A1 => n2277, A2 => n7631, B1 => n2273, B2 => 
                           n8024, ZN => n7205);
   U18953 : INV_X1 port map( A => n7205, ZN => n7915);
   U18954 : OAI22_X1 port map( A1 => n2277, A2 => n7206, B1 => n2273, B2 => 
                           n7915, ZN => n7913);
   U18955 : INV_X1 port map( A => n7913, ZN => n7632);
   U18956 : OAI22_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n597, A2 => 
                           n2227, B1 => DataPath_ALUhw_SHIFTER_HW_n576, B2 => 
                           n7315, ZN => n8103);
   U18957 : INV_X1 port map( A => n8101, ZN => n7625);
   U18958 : OAI22_X1 port map( A1 => n2204, A2 => n4136, B1 => n7289, B2 => 
                           n4131, ZN => n7912);
   U18959 : INV_X1 port map( A => n7912, ZN => n7626);
   U18960 : OAI22_X1 port map( A1 => n7625, A2 => n7991, B1 => n7626, B2 => 
                           n7989, ZN => n7629);
   U18961 : INV_X1 port map( A => n7629, ZN => n7627);
   U18962 : OAI22_X1 port map( A1 => n2204, A2 => n7207, B1 => n7289, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n576, ZN => n8107);
   U18963 : INV_X1 port map( A => n8107, ZN => n7209);
   U18964 : OAI211_X1 port map( C1 => n2274, C2 => n7627, A => n7209, B => 
                           n7208, ZN => n7628);
   U18965 : AOI22_X1 port map( A1 => n7210, A2 => n8103, B1 => n8043, B2 => 
                           n7628, ZN => n7214);
   U18966 : AOI222_X1 port map( A1 => n8118, A2 => n7644, B1 => n8116, B2 => 
                           n7212, C1 => n7211, C2 => n8101, ZN => n7213);
   U18967 : OAI211_X1 port map( C1 => n7632, C2 => n7997, A => n7214, B => 
                           n7213, ZN => n7533);
   U18968 : INV_X1 port map( A => n7561, ZN => n8319);
   U18969 : NAND2_X1 port map( A1 => n1896, A2 => n259, ZN => n8030);
   U18970 : INV_X1 port map( A => n7215, ZN => n11492);
   U18971 : OAI22_X1 port map( A1 => n8319, A2 => n8030, B1 => n11492, B2 => 
                           n8031, ZN => n7216);
   U18972 : AOI221_X1 port map( B1 => n7535, B2 => n8309, C1 => n1859, C2 => 
                           n7533, A => n7216, ZN => n7217);
   U18973 : AOI21_X1 port map( B1 => n7218, B2 => n7217, A => n8140, ZN => 
                           n7219);
   U18974 : AOI221_X1 port map( B1 => n7605, B2 => n7221, C1 => n7606, C2 => 
                           n7220, A => n7219, ZN => n7222);
   U18975 : OAI221_X1 port map( B1 => n7225, B2 => n7224, C1 => n7495, C2 => 
                           n7223, A => n7222, ZN => n7226);
   U18976 : INV_X1 port map( A => n7226, ZN => n7499);
   U18977 : OAI21_X1 port map( B1 => n7495, B2 => n2255, A => n7499, ZN => 
                           n7227);
   U18978 : NAND2_X1 port map( A1 => n7550, A2 => n7227, ZN => n7498);
   U18979 : NAND2_X1 port map( A1 => n1507, A2 => n7229, ZN => n7483);
   U18980 : OAI21_X1 port map( B1 => n1507, B2 => n7229, A => n17223, ZN => 
                           n7482);
   U18981 : OAI22_X1 port map( A1 => n2229, A2 => n7231, B1 => n2227, B2 => 
                           n7230, ZN => n7235);
   U18982 : XOR2_X1 port map( A => n7581, B => n7495, Z => n7232);
   U18983 : NAND2_X1 port map( A1 => n7232, A2 => n2154, ZN => n7233);
   U18984 : MUX2_X1 port map( A => n7233, B => n2147, S => n371, Z => n7234);
   U18985 : XOR2_X1 port map( A => n7235, B => n7234, Z => n7489);
   U18986 : OAI22_X1 port map( A1 => n2240, A2 => n7237, B1 => n2239, B2 => 
                           n7236, ZN => n7470);
   U18987 : OAI21_X1 port map( B1 => n1259, B2 => n7239, A => n7238, ZN => 
                           n7241);
   U18988 : AOI22_X1 port map( A1 => n7241, A2 => n7240, B1 => n1726, B2 => 
                           n7464, ZN => n7242);
   U18989 : OAI22_X1 port map( A1 => n2238, A2 => n7244, B1 => n17239, B2 => 
                           n7243, ZN => n7457);
   U18990 : NAND2_X1 port map( A1 => n1717, A2 => n882, ZN => n7246);
   U18991 : AOI22_X1 port map( A1 => n7246, A2 => n7245, B1 => n1418, B2 => 
                           n7453, ZN => n7450);
   U18992 : INV_X1 port map( A => n7250, ZN => n7252);
   U18993 : OAI21_X1 port map( B1 => n1811, B2 => n7252, A => n7251, ZN => 
                           n7254);
   U18994 : AOI22_X1 port map( A1 => n7254, A2 => n7253, B1 => n763, B2 => 
                           n7445, ZN => n7255);
   U18995 : AOI21_X1 port map( B1 => n7443, B2 => n7446, A => n7255, ZN => 
                           n7439);
   U18996 : OAI22_X1 port map( A1 => n2209, A2 => n7258, B1 => n2205, B2 => 
                           n7256, ZN => n7438);
   U18997 : OAI21_X1 port map( B1 => n945, B2 => n1815, A => n7260, ZN => n7263
                           );
   U18998 : AOI22_X1 port map( A1 => n7263, A2 => n7262, B1 => n7430, B2 => 
                           n7432, ZN => n7264);
   U18999 : AOI21_X1 port map( B1 => n17221, B2 => n7433, A => n7264, ZN => 
                           n7425);
   U19000 : OAI22_X1 port map( A1 => n2215, A2 => n7266, B1 => n2213, B2 => 
                           n7265, ZN => n7424);
   U19001 : OAI21_X1 port map( B1 => n1814, B2 => n7268, A => n7267, ZN => 
                           n7270);
   U19002 : INV_X1 port map( A => n7420, ZN => n7417);
   U19003 : AOI22_X1 port map( A1 => n7270, A2 => n7269, B1 => n565, B2 => 
                           n7417, ZN => n7271);
   U19004 : AOI21_X1 port map( B1 => n7418, B2 => n7420, A => n7271, ZN => 
                           n7412);
   U19005 : OAI22_X1 port map( A1 => n2176, A2 => n7274, B1 => n2178, B2 => 
                           n7272, ZN => n7411);
   U19006 : XOR2_X1 port map( A => n7276, B => n7389, Z => n7277);
   U19007 : NAND2_X1 port map( A1 => n7404, A2 => n7407, ZN => n7282);
   U19008 : OAI21_X1 port map( B1 => n7280, B2 => n1792, A => n7279, ZN => 
                           n7281);
   U19009 : INV_X1 port map( A => n7407, ZN => n7403);
   U19010 : AOI22_X1 port map( A1 => n7282, A2 => n7281, B1 => n7403, B2 => 
                           n7406, ZN => n7399);
   U19011 : OAI22_X1 port map( A1 => n2179, A2 => n7285, B1 => n7284, B2 => 
                           n7283, ZN => n7398);
   U19012 : NAND2_X1 port map( A1 => n725, A2 => n7391, ZN => n7288);
   U19013 : INV_X1 port map( A => n725, ZN => n7390);
   U19014 : AOI22_X1 port map( A1 => n7288, A2 => n7287, B1 => n7390, B2 => 
                           n7393, ZN => n7388);
   U19015 : OAI22_X1 port map( A1 => n7923, A2 => n7291, B1 => n2185, B2 => 
                           n7289, ZN => n7387);
   U19016 : INV_X1 port map( A => n7382, ZN => n7378);
   U19018 : NAND2_X1 port map( A1 => n17219, A2 => n7378, ZN => n7293);
   U19019 : AOI22_X1 port map( A1 => n7293, A2 => n7292, B1 => n576, B2 => 
                           n7382, ZN => n7376);
   U19020 : OAI22_X1 port map( A1 => n7864, A2 => n2183, B1 => n2182, B2 => 
                           n7294, ZN => n7375);
   U19021 : NAND2_X1 port map( A1 => n310, A2 => n7297, ZN => n7299);
   U19022 : INV_X1 port map( A => n7366, ZN => n7370);
   U19023 : NAND2_X1 port map( A1 => n7367, A2 => n7370, ZN => n7301);
   U19024 : AOI22_X1 port map( A1 => n7301, A2 => n1334, B1 => n7366, B2 => 
                           n7369, ZN => n7364);
   U19025 : OAI22_X1 port map( A1 => n7792, A2 => n2181, B1 => n2217, B2 => 
                           n7302, ZN => n7363);
   U19026 : MUX2_X1 port map( A => n7307, B => n7306, S => n2247, Z => n7358);
   U19027 : INV_X1 port map( A => n7358, ZN => n7354);
   U19028 : AOI22_X1 port map( A1 => n7309, A2 => n7308, B1 => n7355, B2 => 
                           n7358, ZN => n7310);
   U19029 : AOI21_X1 port map( B1 => n7354, B2 => n7357, A => n7310, ZN => 
                           n7349);
   U19030 : OAI22_X1 port map( A1 => n8094, A2 => n2221, B1 => n2219, B2 => 
                           n7311, ZN => n7348);
   U19031 : INV_X1 port map( A => n7343, ZN => n7339);
   U19032 : NAND2_X1 port map( A1 => n7339, A2 => n7342, ZN => n7314);
   U19033 : AOI22_X1 port map( A1 => n7314, A2 => n7313, B1 => n7340, B2 => 
                           n7343, ZN => n7337);
   U19034 : OAI22_X1 port map( A1 => n7670, A2 => n2225, B1 => n2224, B2 => 
                           n7315, ZN => n7336);
   U19035 : NAND2_X1 port map( A1 => n7317, A2 => n2259, ZN => n7321);
   U19036 : AOI22_X1 port map( A1 => n8067, A2 => n924, B1 => n677, B2 => n8079
                           , ZN => n7320);
   U19037 : AOI22_X1 port map( A1 => n8049, A2 => n17175, B1 => n17193, B2 => 
                           n8058, ZN => n7319);
   U19038 : INV_X1 port map( A => n7327, ZN => n7328);
   U19039 : NAND2_X1 port map( A1 => n7328, A2 => n7326, ZN => n7323);
   U19040 : AOI22_X1 port map( A1 => n7323, A2 => n7322, B1 => n7329, B2 => 
                           n7327, ZN => n7324);
   U19041 : XOR2_X1 port map( A => n7325, B => n7324, Z => n7334);
   U19042 : NAND2_X1 port map( A1 => n7327, A2 => n7326, ZN => n7331);
   U19043 : AOI22_X1 port map( A1 => n7331, A2 => n7330, B1 => n7329, B2 => 
                           n7328, ZN => n7332);
   U19044 : XOR2_X1 port map( A => n7337, B => n1904, Z => n7346);
   U19045 : OAI21_X1 port map( B1 => n7340, B2 => n7339, A => n7338, ZN => 
                           n7341);
   U19046 : OAI21_X1 port map( B1 => n7343, B2 => n7342, A => n7341, ZN => 
                           n7344);
   U19047 : XOR2_X1 port map( A => n7344, B => n1904, Z => n7345);
   U19048 : MUX2_X1 port map( A => n7346, B => n7345, S => n2247, Z => n7347);
   U19049 : XOR2_X1 port map( A => n7349, B => n1903, Z => n7361);
   U19050 : INV_X1 port map( A => n7350, ZN => n7353);
   U19051 : INV_X1 port map( A => n7351, ZN => n7352);
   U19052 : OAI22_X1 port map( A1 => n7355, A2 => n7354, B1 => n7353, B2 => 
                           n7352, ZN => n7356);
   U19053 : OAI21_X1 port map( B1 => n7358, B2 => n7357, A => n7356, ZN => 
                           n7359);
   U19054 : XOR2_X1 port map( A => n7359, B => n1903, Z => n7360);
   U19055 : MUX2_X1 port map( A => n7361, B => n7360, S => n2245, Z => n7362);
   U19056 : XOR2_X1 port map( A => n1902, B => n7364, Z => n7373);
   U19057 : OAI21_X1 port map( B1 => n7367, B2 => n7366, A => n7365, ZN => 
                           n7368);
   U19059 : XOR2_X1 port map( A => n7371, B => n1902, Z => n7372);
   U19060 : XOR2_X1 port map( A => n17204, B => n7376, Z => n7385);
   U19061 : OAI21_X1 port map( B1 => n7378, B2 => n1466, A => n7377, ZN => 
                           n7380);
   U19062 : OAI21_X1 port map( B1 => n7382, B2 => n17219, A => n7380, ZN => 
                           n7383);
   U19063 : XOR2_X1 port map( A => n1901, B => n7383, Z => n7384);
   U19064 : XOR2_X1 port map( A => n1900, B => n7388, Z => n7396);
   U19065 : OAI21_X1 port map( B1 => n7390, B2 => n7391, A => n7389, ZN => 
                           n7392);
   U19066 : XOR2_X1 port map( A => n1900, B => n7394, Z => n7395);
   U19067 : OAI21_X1 port map( B1 => n7401, B2 => n1838, A => n7400, ZN => 
                           n7402);
   U19068 : OAI21_X1 port map( B1 => n7403, B2 => n7404, A => n7402, ZN => 
                           n7405);
   U19069 : XOR2_X1 port map( A => n1880, B => n7412, Z => n7422);
   U19070 : AOI21_X1 port map( B1 => n7415, B2 => n7414, A => n1831, ZN => 
                           n7416);
   U19071 : OAI22_X1 port map( A1 => n7418, A2 => n7417, B1 => n1502, B2 => 
                           n7416, ZN => n7419);
   U19072 : INV_X1 port map( A => n7426, ZN => n7429);
   U19073 : AOI21_X1 port map( B1 => n7427, B2 => n1401, A => n1832, ZN => 
                           n7428);
   U19074 : OAI22_X1 port map( A1 => n17221, A2 => n7430, B1 => n7429, B2 => 
                           n7428, ZN => n7431);
   U19075 : OAI21_X1 port map( B1 => n7433, B2 => n7432, A => n7431, ZN => 
                           n7434);
   U19076 : OAI22_X1 port map( A1 => n7443, A2 => n763, B1 => n1786, B2 => 
                           n7442, ZN => n7444);
   U19077 : XOR2_X1 port map( A => n1881, B => n7450, Z => n7455);
   U19078 : OAI21_X1 port map( B1 => n1418, B2 => n1717, A => n7451, ZN => 
                           n7452);
   U19079 : INV_X1 port map( A => n7458, ZN => n7462);
   U19080 : AOI21_X1 port map( B1 => n825, B2 => n7460, A => n1828, ZN => n7461
                           );
   U19081 : OAI22_X1 port map( A1 => n1726, A2 => n1420, B1 => n7462, B2 => 
                           n7461, ZN => n7463);
   U19082 : OAI21_X1 port map( B1 => n7465, B2 => n7464, A => n7463, ZN => 
                           n7466);
   U19083 : XOR2_X1 port map( A => n1882, B => n7466, Z => n7467);
   U19084 : OAI211_X1 port map( C1 => n7478, C2 => n7476, A => n7472, B => 
                           n7471, ZN => n7480);
   U19085 : OAI211_X1 port map( C1 => n7476, C2 => n7474, A => n7473, B => 
                           n7647, ZN => n7475);
   U19086 : NAND3_X1 port map( A1 => n7482, A2 => n7481, A3 => n7483, ZN => 
                           n7486);
   U19087 : NAND3_X1 port map( A1 => n7579, A2 => n7483, A3 => n7482, ZN => 
                           n7484);
   U19088 : OAI21_X1 port map( B1 => n1308, B2 => n7581, A => n7484, ZN => 
                           n7485);
   U19089 : NAND2_X1 port map( A1 => n7485, A2 => n7486, ZN => n7503);
   U19090 : OAI222_X1 port map( A1 => n7488, A2 => n7487, B1 => n1507, B2 => 
                           n7487, C1 => n1541, C2 => n587, ZN => n7490);
   U19091 : NAND2_X1 port map( A1 => n7491, A2 => n7581, ZN => n7504);
   U19092 : NAND3_X1 port map( A1 => n7550, A2 => n7495, A3 => n2258, ZN => 
                           n7507);
   U19093 : OAI22_X1 port map( A1 => n7499, A2 => n7498, B1 => n7979, B2 => 
                           n7497, ZN => n7500);
   U19094 : INV_X1 port map( A => n7500, ZN => n7502);
   U19095 : NAND3_X1 port map( A1 => n1130, A2 => n7503, A3 => n7502, ZN => 
                           n7505);
   U19096 : NAND2_X1 port map( A1 => n1235, A2 => n1548, ZN => n7546);
   U19097 : NAND3_X1 port map( A1 => n7513, A2 => n7512, A3 => n7511, ZN => 
                           n8660);
   U19098 : INV_X1 port map( A => n7514, ZN => n7746);
   U19099 : NAND2_X1 port map( A1 => n1907, A2 => n7746, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n150);
   U19100 : XOR2_X1 port map( A => n7516, B => n8058, Z => n7520);
   U19101 : INV_X1 port map( A => n7965, ZN => n7924);
   U19102 : NAND2_X1 port map( A1 => n7924, A2 => n7515, ZN => n7518);
   U19103 : INV_X1 port map( A => n7969, ZN => n7925);
   U19104 : NAND2_X1 port map( A1 => n7925, A2 => n8058, ZN => n7517);
   U19105 : INV_X1 port map( A => n7979, ZN => n8323);
   U19106 : NAND2_X1 port map( A1 => DRAM_ADDRESS_30_port, A2 => n8323, ZN => 
                           n7542);
   U19107 : OAI211_X1 port map( C1 => n7520, C2 => n2187, A => n7519, B => 
                           n7542, ZN => n7545);
   U19108 : XOR2_X1 port map( A => n7524, B => n7521, Z => n7541);
   U19109 : INV_X1 port map( A => n7522, ZN => n7523);
   U19110 : XOR2_X1 port map( A => n7524, B => n7523, Z => n7540);
   U19111 : INV_X1 port map( A => n7525, ZN => n7816);
   U19112 : OAI222_X1 port map( A1 => n4139, A2 => n8061, B1 => n2279, B2 => 
                           n7526, C1 => n266, C2 => n2238, ZN => n7527);
   U19113 : INV_X1 port map( A => n7527, ZN => n8055);
   U19114 : OAI22_X1 port map( A1 => n2277, A2 => n7528, B1 => n2273, B2 => 
                           n8055, ZN => n8012);
   U19115 : AOI222_X1 port map( A1 => n8116, A2 => n7530, B1 => n8034, B2 => 
                           n8012, C1 => n7529, C2 => n8073, ZN => n7531);
   U19116 : OAI221_X1 port map( B1 => n7816, B2 => n2134, C1 => n7532, C2 => 
                           n8037, A => n7531, ZN => n7754);
   U19117 : INV_X1 port map( A => n7754, ZN => n11491);
   U19118 : INV_X1 port map( A => n7533, ZN => n8308);
   U19119 : NAND3_X1 port map( A1 => n7746, A2 => n4135, A3 => n2130, ZN => 
                           n8099);
   U19120 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n150, A2 => 
                           n8030, ZN => n7727);
   U19121 : NAND3_X1 port map( A1 => n7746, A2 => n259, A3 => n2130, ZN => 
                           n8025);
   U19122 : NAND2_X1 port map( A1 => n1769, A2 => n8025, ZN => n7698);
   U19123 : AOI222_X1 port map( A1 => n7727, A2 => n7596, B1 => n7698, B2 => 
                           n7563, C1 => n7697, C2 => n7561, ZN => n7534);
   U19124 : OAI221_X1 port map( B1 => n2984, B2 => n11491, C1 => n8308, C2 => 
                           n8099, A => n7534, ZN => n7538);
   U19125 : INV_X1 port map( A => n7535, ZN => n8317);
   U19126 : INV_X1 port map( A => n7536, ZN => n8318);
   U19127 : OAI222_X1 port map( A1 => n8317, A2 => n8026, B1 => n8318, B2 => 
                           n2242, C1 => n8316, C2 => n8031, ZN => n7537);
   U19128 : NOR4_X1 port map( A1 => n7538, A2 => n7537, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n250, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n260, ZN => n7539);
   U19129 : OAI222_X1 port map( A1 => n7541, A2 => n7568, B1 => n7540, B2 => 
                           n7572, C1 => n7539, C2 => n8140, ZN => n7544);
   U19130 : INV_X1 port map( A => n7542, ZN => n7543);
   U19131 : OAI22_X1 port map( A1 => n7545, A2 => n7544, B1 => n7550, B2 => 
                           n7543, ZN => n7552);
   U19132 : OAI22_X1 port map( A1 => n590, A2 => n7548, B1 => n7546, B2 => 
                           n7547, ZN => n7549);
   U19133 : NAND2_X1 port map( A1 => n7551, A2 => n7552, ZN => n8661);
   U19134 : INV_X1 port map( A => n7553, ZN => n7848);
   U19135 : OAI222_X1 port map( A1 => n4139, A2 => n8070, B1 => n2279, B2 => 
                           n7554, C1 => n266, C2 => n2239, ZN => n7555);
   U19136 : INV_X1 port map( A => n7555, ZN => n8064);
   U19137 : OAI22_X1 port map( A1 => n2277, A2 => n7556, B1 => n2273, B2 => 
                           n8064, ZN => n8027);
   U19138 : AOI222_X1 port map( A1 => n8116, A2 => n7558, B1 => n8034, B2 => 
                           n8027, C1 => n7557, C2 => n8073, ZN => n7559);
   U19139 : OAI221_X1 port map( B1 => n7848, B2 => n2134, C1 => n7560, C2 => 
                           n8037, A => n7559, ZN => n7788);
   U19140 : INV_X1 port map( A => n7788, ZN => n7821);
   U19141 : AOI222_X1 port map( A1 => n7727, A2 => n7754, B1 => n7698, B2 => 
                           n7561, C1 => n7697, C2 => n7596, ZN => n7562);
   U19142 : OAI221_X1 port map( B1 => n2984, B2 => n7821, C1 => n8318, C2 => 
                           n8099, A => n7562, ZN => n7565);
   U19143 : INV_X1 port map( A => n7563, ZN => n8313);
   U19144 : OAI222_X1 port map( A1 => n8308, A2 => n8026, B1 => n8317, B2 => 
                           n8031, C1 => n8313, C2 => n2242, ZN => n7564);
   U19145 : NOR4_X1 port map( A1 => n7565, A2 => n7564, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n275, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n282, ZN => n7570);
   U19146 : INV_X1 port map( A => n7566, ZN => n7571);
   U19147 : XOR2_X1 port map( A => n7567, B => n7571, Z => n7569);
   U19148 : OAI22_X1 port map( A1 => n7570, A2 => n8140, B1 => n7569, B2 => 
                           n7568, ZN => n7585);
   U19149 : MUX2_X1 port map( A => n7965, B => n2187, S => n8067, Z => n7575);
   U19150 : MUX2_X1 port map( A => n2187, B => n7969, S => n8067, Z => n7574);
   U19151 : XOR2_X1 port map( A => n7571, B => n369, Z => n7573);
   U19152 : OAI222_X1 port map( A1 => n7581, A2 => n7575, B1 => n7579, B2 => 
                           n7574, C1 => n7573, C2 => n7572, ZN => n7584);
   U19153 : XOR2_X1 port map( A => n1800, B => n992, Z => n7582);
   U19154 : XOR2_X1 port map( A => n1800, B => n1808, Z => n7580);
   U19155 : OAI33_X1 port map( A1 => n7582, A2 => n7581, A3 => n2253, B1 => 
                           n7580, B2 => n7579, B3 => n2253, ZN => n7583);
   U19156 : NOR3_X1 port map( A1 => n7583, A2 => n7584, A3 => n7585, ZN => 
                           n7587);
   U19157 : OAI22_X1 port map( A1 => n7587, A2 => n7980, B1 => n7979, B2 => 
                           n7586, ZN => n8662);
   U19158 : XOR2_X1 port map( A => n7608, B => n8079, Z => n7602);
   U19159 : AOI21_X1 port map( B1 => n231, B2 => n7588, A => n433, ZN => n7601)
                           ;
   U19160 : INV_X1 port map( A => n7589, ZN => n7879);
   U19161 : OAI222_X1 port map( A1 => n8083, A2 => n4136, B1 => n7590, B2 => 
                           n7991, C1 => n2240, C2 => n266, ZN => n8016);
   U19162 : INV_X1 port map( A => n8016, ZN => n8076);
   U19163 : OAI22_X1 port map( A1 => n2277, A2 => n7591, B1 => n2273, B2 => 
                           n8076, ZN => n8015);
   U19164 : AOI222_X1 port map( A1 => n8116, A2 => n7593, B1 => n8034, B2 => 
                           n8015, C1 => n7592, C2 => n8073, ZN => n7594);
   U19165 : OAI221_X1 port map( B1 => n7879, B2 => n2134, C1 => n7595, C2 => 
                           n8037, A => n7594, ZN => n7819);
   U19166 : INV_X1 port map( A => n7819, ZN => n7853);
   U19167 : AOI222_X1 port map( A1 => n7727, A2 => n7788, B1 => n7698, B2 => 
                           n7596, C1 => n7697, C2 => n7754, ZN => n7597);
   U19168 : OAI221_X1 port map( B1 => n2984, B2 => n7853, C1 => n8313, C2 => 
                           n8099, A => n7597, ZN => n7599);
   U19169 : OAI222_X1 port map( A1 => n8308, A2 => n8031, B1 => n8318, B2 => 
                           n8026, C1 => n8319, C2 => n2242, ZN => n7598);
   U19170 : NOR4_X1 port map( A1 => n7599, A2 => n7598, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n289, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n296, ZN => n7600);
   U19171 : OAI222_X1 port map( A1 => n7602, A2 => n2186, B1 => n7601, B2 => 
                           n2252, C1 => n7600, C2 => n8140, ZN => n7614);
   U19172 : INV_X1 port map( A => n7603, ZN => n7604);
   U19173 : MUX2_X1 port map( A => n7606, B => n7605, S => n7604, Z => n7613);
   U19174 : NOR2_X1 port map( A1 => n8079, A2 => n7965, ZN => n7611);
   U19175 : NOR2_X1 port map( A1 => n7607, A2 => n7969, ZN => n7610);
   U19176 : INV_X1 port map( A => n7608, ZN => n7609);
   U19177 : MUX2_X1 port map( A => n7611, B => n7610, S => n7609, Z => n7612);
   U19178 : NOR3_X1 port map( A1 => n7614, A2 => n7613, A3 => n7612, ZN => 
                           n7616);
   U19179 : OAI22_X1 port map( A1 => n7616, A2 => n7980, B1 => n7979, B2 => 
                           n7615, ZN => n8663);
   U19180 : INV_X1 port map( A => n12931, ZN => n7617);
   U19181 : NAND2_X1 port map( A1 => n7618, A2 => n7702, ZN => n7687);
   U19182 : INV_X1 port map( A => n7687, ZN => n7619);
   U19183 : OAI21_X1 port map( B1 => n7637, B2 => n7619, A => n7636, ZN => 
                           n7655);
   U19184 : INV_X1 port map( A => n7655, ZN => n7621);
   U19185 : OAI21_X1 port map( B1 => n7622, B2 => n7621, A => n7620, ZN => 
                           n7623);
   U19186 : XOR2_X1 port map( A => n7623, B => n364, Z => n7652);
   U19187 : OAI222_X1 port map( A1 => n7626, A2 => n7991, B1 => n7625, B2 => 
                           n4135, C1 => n2227, C2 => n266, ZN => n8021);
   U19188 : INV_X1 port map( A => n8021, ZN => n8105);
   U19189 : OAI22_X1 port map( A1 => n2277, A2 => n7627, B1 => n2273, B2 => 
                           n8105, ZN => n8020);
   U19190 : AOI222_X1 port map( A1 => n8116, A2 => n7629, B1 => n8034, B2 => 
                           n8020, C1 => n7628, C2 => n8073, ZN => n7630);
   U19191 : OAI221_X1 port map( B1 => n7632, B2 => n2134, C1 => n7631, C2 => 
                           n8037, A => n7630, ZN => n7851);
   U19192 : INV_X1 port map( A => n7851, ZN => n11493);
   U19193 : AOI222_X1 port map( A1 => n7727, A2 => n7819, B1 => n7698, B2 => 
                           n7754, C1 => n7697, C2 => n7788, ZN => n7633);
   U19194 : OAI221_X1 port map( B1 => n2984, B2 => n11493, C1 => n8319, C2 => 
                           n8099, A => n7633, ZN => n7635);
   U19195 : OAI222_X1 port map( A1 => n8318, A2 => n8031, B1 => n8320, B2 => 
                           n2242, C1 => n8313, C2 => n8026, ZN => n7634);
   U19196 : NOR4_X1 port map( A1 => n7635, A2 => n7634, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n303, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n310, ZN => n7640);
   U19197 : OAI21_X1 port map( B1 => n7637, B2 => n7702, A => n7636, ZN => 
                           n7656);
   U19198 : AOI21_X1 port map( B1 => n7656, B2 => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_27_port, A 
                           => DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_0_0_27_port,
                           ZN => n7638);
   U19199 : XOR2_X1 port map( A => n364, B => n7638, Z => n7639);
   U19200 : NAND2_X1 port map( A1 => n12931, A2 => n2272, ZN => n7734);
   U19201 : OAI22_X1 port map( A1 => n7640, A2 => n8140, B1 => n7639, B2 => 
                           n7734, ZN => n7651);
   U19202 : XOR2_X1 port map( A => n434, B => n431, Z => n7643);
   U19203 : MUX2_X1 port map( A => n7965, B => n2186, S => n7644, Z => n7642);
   U19204 : OAI21_X1 port map( B1 => n7643, B2 => n2254, A => n7642, ZN => 
                           n7649);
   U19205 : XOR2_X1 port map( A => n1305, B => n1818, Z => n7646);
   U19206 : MUX2_X1 port map( A => n2186, B => n7969, S => n7644, Z => n7645);
   U19207 : OAI21_X1 port map( B1 => n7646, B2 => n2254, A => n7645, ZN => 
                           n7648);
   U19208 : MUX2_X1 port map( A => n7649, B => n7648, S => n7647, Z => n7650);
   U19209 : AOI211_X1 port map( C1 => n365, C2 => n7652, A => n7651, B => n7650
                           , ZN => n7654);
   U19210 : OAI22_X1 port map( A1 => n7654, A2 => n7980, B1 => n7979, B2 => 
                           n7653, ZN => n8664);
   U19211 : XOR2_X1 port map( A => n7655, B => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_27_port, Z 
                           => n7684);
   U19212 : INV_X1 port map( A => n7656, ZN => n7657);
   U19213 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_27_port, B 
                           => n7657, Z => n7676);
   U19214 : OAI222_X1 port map( A1 => n7660, A2 => n7991, B1 => n7659, B2 => 
                           n4135, C1 => n2229, C2 => n266, ZN => n8004);
   U19215 : INV_X1 port map( A => n8004, ZN => n8112);
   U19216 : OAI22_X1 port map( A1 => n2278, A2 => n7661, B1 => n2273, B2 => 
                           n8112, ZN => n8003);
   U19217 : AOI222_X1 port map( A1 => n8116, A2 => n7663, B1 => n8034, B2 => 
                           n8003, C1 => n7662, C2 => n8073, ZN => n7664);
   U19218 : OAI221_X1 port map( B1 => n7666, B2 => n2134, C1 => n7665, C2 => 
                           n8037, A => n7664, ZN => n7885);
   U19219 : INV_X1 port map( A => n7885, ZN => n8303);
   U19220 : AOI222_X1 port map( A1 => n7727, A2 => n7851, B1 => n7698, B2 => 
                           n7788, C1 => n7697, C2 => n7819, ZN => n7667);
   U19221 : OAI221_X1 port map( B1 => n2984, B2 => n8303, C1 => n11491, C2 => 
                           n2242, A => n7667, ZN => n7669);
   U19222 : OAI222_X1 port map( A1 => n8319, A2 => n8026, B1 => n8320, B2 => 
                           n8099, C1 => n8313, C2 => n8031, ZN => n7668);
   U19223 : NOR4_X1 port map( A1 => n7669, A2 => n7668, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n317, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n324, ZN => n7675);
   U19224 : NAND2_X1 port map( A1 => n7924, A2 => n7670, ZN => n7673);
   U19225 : NAND2_X1 port map( A1 => n7925, A2 => n7677, ZN => n7672);
   U19226 : INV_X1 port map( A => n7678, ZN => n7671);
   U19227 : MUX2_X1 port map( A => n7673, B => n7672, S => n7671, Z => n7674);
   U19228 : OAI221_X1 port map( B1 => n7676, B2 => n7734, C1 => n7675, C2 => 
                           n8140, A => n7674, ZN => n7683);
   U19229 : XOR2_X1 port map( A => n7678, B => n7677, Z => n7681);
   U19230 : AOI21_X1 port map( B1 => n1699, B2 => n7679, A => n1305, ZN => 
                           n7680);
   U19231 : OAI22_X1 port map( A1 => n7681, A2 => n2187, B1 => n7680, B2 => 
                           n2253, ZN => n7682);
   U19232 : AOI211_X1 port map( C1 => n365, C2 => n7684, A => n7683, B => n7682
                           , ZN => n7686);
   U19233 : OAI22_X1 port map( A1 => n7686, A2 => n7980, B1 => n7979, B2 => 
                           n7685, ZN => n8665);
   U19234 : XOR2_X1 port map( A => n7687, B => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_26_port, Z 
                           => n7717);
   U19235 : OAI222_X1 port map( A1 => n4139, A2 => n7690, B1 => n2279, B2 => 
                           n7689, C1 => n266, C2 => n2147, ZN => n8000);
   U19236 : INV_X1 port map( A => n8000, ZN => n8123);
   U19237 : OAI22_X1 port map( A1 => n2278, A2 => n7691, B1 => n2273, B2 => 
                           n8123, ZN => n7999);
   U19238 : AOI222_X1 port map( A1 => n8116, A2 => n7693, B1 => n8034, B2 => 
                           n7999, C1 => n7692, C2 => n8073, ZN => n7694);
   U19239 : OAI221_X1 port map( B1 => n7696, B2 => n2134, C1 => n7695, C2 => 
                           n8037, A => n7694, ZN => n7919);
   U19240 : INV_X1 port map( A => n7919, ZN => n8302);
   U19241 : AOI222_X1 port map( A1 => n7727, A2 => n7885, B1 => n7698, B2 => 
                           n7819, C1 => n7697, C2 => n7851, ZN => n7699);
   U19242 : OAI221_X1 port map( B1 => n2984, B2 => n8302, C1 => n7821, C2 => 
                           n2242, A => n7699, ZN => n7701);
   U19243 : OAI222_X1 port map( A1 => n8320, A2 => n8026, B1 => n11491, B2 => 
                           n8099, C1 => n8319, C2 => n8031, ZN => n7700);
   U19244 : NOR4_X1 port map( A1 => n7701, A2 => n7700, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n331, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n338, ZN => n7704);
   U19245 : XOR2_X1 port map( A => n7702, B => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_26_port, Z 
                           => n7703);
   U19246 : OAI22_X1 port map( A1 => n7704, A2 => n8140, B1 => n7703, B2 => 
                           n7734, ZN => n7716);
   U19247 : XOR2_X1 port map( A => n1781, B => n1819, Z => n7707);
   U19248 : MUX2_X1 port map( A => n7965, B => n2186, S => n7709, Z => n7706);
   U19249 : OAI21_X1 port map( B1 => n7707, B2 => n2254, A => n7706, ZN => 
                           n7714);
   U19250 : XOR2_X1 port map( A => n984, B => n1819, Z => n7711);
   U19251 : MUX2_X1 port map( A => n2186, B => n7969, S => n7709, Z => n7710);
   U19252 : OAI21_X1 port map( B1 => n7711, B2 => n2254, A => n7710, ZN => 
                           n7713);
   U19253 : MUX2_X1 port map( A => n7714, B => n7713, S => n7712, Z => n7715);
   U19254 : AOI211_X1 port map( C1 => n365, C2 => n7717, A => n7716, B => n7715
                           , ZN => n7719);
   U19255 : OAI22_X1 port map( A1 => n7719, A2 => n7980, B1 => n7979, B2 => 
                           n7718, ZN => n8666);
   U19256 : OAI222_X1 port map( A1 => n4139, A2 => n7721, B1 => n2279, B2 => 
                           n7720, C1 => n266, C2 => n771, ZN => n8097);
   U19257 : INV_X1 port map( A => n8097, ZN => n8039);
   U19258 : OAI22_X1 port map( A1 => n2278, A2 => n7725, B1 => n2273, B2 => 
                           n8039, ZN => n8035);
   U19259 : AOI222_X1 port map( A1 => n7723, A2 => n8073, B1 => n8034, B2 => 
                           n8035, C1 => n7994, C2 => n7722, ZN => n7724);
   U19260 : OAI221_X1 port map( B1 => n7725, B2 => n8089, C1 => n7987, C2 => 
                           n2134, A => n7724, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n344);
   U19261 : XOR2_X1 port map( A => n7737, B => n7736, Z => n7733);
   U19262 : AOI21_X1 port map( B1 => n916, B2 => n7726, A => n984, ZN => n7732)
                           ;
   U19263 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n191, A2 => 
                           n8099, ZN => n7954);
   U19264 : AOI222_X1 port map( A1 => n7727, A2 => n7919, B1 => n7788, B2 => 
                           n7954, C1 => n7953, C2 => n7754, ZN => n7728);
   U19265 : OAI221_X1 port map( B1 => n8303, B2 => n8032, C1 => n11493, C2 => 
                           n8025, A => n7728, ZN => n7730);
   U19266 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n344, ZN => n8301);
   U19267 : OAI222_X1 port map( A1 => n8320, A2 => n8031, B1 => n7853, B2 => 
                           n2242, C1 => n2984, C2 => n8301, ZN => n7729);
   U19268 : NOR4_X1 port map( A1 => n7730, A2 => n7729, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n345, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n354, ZN => n7731);
   U19269 : OAI222_X1 port map( A1 => n7733, A2 => n2186, B1 => n7732, B2 => 
                           n2252, C1 => n7731, C2 => n8140, ZN => n7743);
   U19270 : INV_X1 port map( A => n7734, ZN => n7735);
   U19271 : MUX2_X1 port map( A => n365, B => n7735, S => 
                           DataPath_ALUhw_ADDER_CARRYGEN_sigmtx_1_0_25_port, Z 
                           => n7742);
   U19272 : NOR2_X1 port map( A1 => n7736, A2 => n7965, ZN => n7740);
   U19273 : NOR2_X1 port map( A1 => n8094, A2 => n7969, ZN => n7739);
   U19274 : INV_X1 port map( A => n7737, ZN => n7738);
   U19275 : MUX2_X1 port map( A => n7740, B => n7739, S => n7738, Z => n7741);
   U19276 : NOR3_X1 port map( A1 => n7743, A2 => n7742, A3 => n7741, ZN => 
                           n7745);
   U19277 : OAI22_X1 port map( A1 => n7745, A2 => n7980, B1 => n7979, B2 => 
                           n7744, ZN => n8667);
   U19278 : INV_X1 port map( A => n12930, ZN => n7748);
   U19279 : NAND2_X1 port map( A1 => n7860, A2 => n7825, ZN => n7818);
   U19280 : INV_X1 port map( A => n7818, ZN => n7750);
   U19281 : OAI21_X1 port map( B1 => n7817, B2 => n7750, A => n7749, ZN => 
                           n7785);
   U19282 : INV_X1 port map( A => n7785, ZN => n7751);
   U19283 : OAI21_X1 port map( B1 => n7752, B2 => n7751, A => n7758, ZN => 
                           n7753);
   U19284 : XOR2_X1 port map( A => n7753, B => n7761, Z => n7776);
   U19285 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n182, A2 => 
                           n8031, ZN => n7955);
   U19286 : AOI222_X1 port map( A1 => n7955, A2 => n7754, B1 => n7819, B2 => 
                           n7954, C1 => n7788, C2 => n7953, ZN => n7755);
   U19287 : OAI221_X1 port map( B1 => n8302, B2 => n8032, C1 => n8303, C2 => 
                           n8025, A => n7755, ZN => n7757);
   U19288 : OAI222_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n181, A2 => 
                           n8320, B1 => n11493, B2 => n2242, C1 => n8301, C2 =>
                           n8030, ZN => n7756);
   U19289 : NOR4_X1 port map( A1 => n7757, A2 => n7756, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n360, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n367, ZN => n7763);
   U19290 : INV_X1 port map( A => n7758, ZN => n7759);
   U19291 : AOI21_X1 port map( B1 => n11529, B2 => n7787, A => n7759, ZN => 
                           n7760);
   U19292 : XOR2_X1 port map( A => n7761, B => n7760, Z => n7762);
   U19293 : NAND2_X1 port map( A1 => n12930, A2 => n2272, ZN => n7859);
   U19294 : OAI22_X1 port map( A1 => n7763, A2 => n8140, B1 => n7762, B2 => 
                           n7859, ZN => n7775);
   U19295 : XOR2_X1 port map( A => n1076, B => n1854, Z => n7766);
   U19296 : MUX2_X1 port map( A => n7965, B => n2187, S => n7768, Z => n7765);
   U19297 : OAI21_X1 port map( B1 => n7766, B2 => n2254, A => n7765, ZN => 
                           n7773);
   U19298 : INV_X1 port map( A => n7767, ZN => n7801);
   U19299 : XOR2_X1 port map( A => n7801, B => n1854, Z => n7770);
   U19300 : MUX2_X1 port map( A => n2187, B => n7969, S => n7768, Z => n7769);
   U19301 : OAI21_X1 port map( B1 => n7770, B2 => n2254, A => n7769, ZN => 
                           n7772);
   U19302 : MUX2_X1 port map( A => n7773, B => n7772, S => n7771, Z => n7774);
   U19303 : AOI211_X1 port map( C1 => n366, C2 => n7776, A => n7775, B => n7774
                           , ZN => n7778);
   U19304 : OAI22_X1 port map( A1 => n7778, A2 => n7980, B1 => n7979, B2 => 
                           n7777, ZN => n8668);
   U19305 : OAI21_X1 port map( B1 => n2278, B2 => n8010, A => n7779, ZN => 
                           n8040);
   U19306 : INV_X1 port map( A => n8040, ZN => n7780);
   U19307 : OAI22_X1 port map( A1 => n7784, A2 => n7991, B1 => n7780, B2 => 
                           n7989, ZN => n8041);
   U19308 : AOI222_X1 port map( A1 => n7781, A2 => n8073, B1 => n8034, B2 => 
                           n8041, C1 => n8043, C2 => n8007, ZN => n7782);
   U19309 : OAI221_X1 port map( B1 => n7784, B2 => n8089, C1 => n7783, C2 => 
                           n8037, A => n7782, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n380);
   U19310 : XOR2_X1 port map( A => n7785, B => n7787, Z => n7808);
   U19311 : INV_X1 port map( A => n11529, ZN => n7786);
   U19312 : XOR2_X1 port map( A => n7787, B => n7786, Z => n7798);
   U19313 : AOI222_X1 port map( A1 => n7788, A2 => n7955, B1 => n7954, B2 => 
                           n7851, C1 => n7819, C2 => n7953, ZN => n7789);
   U19314 : OAI221_X1 port map( B1 => n8302, B2 => n8025, C1 => n8303, C2 => 
                           n2242, A => n7789, ZN => n7791);
   U19315 : OAI222_X1 port map( A1 => n8301, A2 => n8032, B1 => 
                           DataPath_ALUhw_SHIFTER_HW_n181, B2 => n11491, C1 => 
                           n8298, C2 => n8030, ZN => n7790);
   U19316 : NOR4_X1 port map( A1 => n7791, A2 => n7790, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n373, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n378, ZN => n7797);
   U19317 : NAND2_X1 port map( A1 => n7924, A2 => n7792, ZN => n7795);
   U19318 : NAND2_X1 port map( A1 => n7925, A2 => n7799, ZN => n7794);
   U19319 : INV_X1 port map( A => n7800, ZN => n7793);
   U19320 : MUX2_X1 port map( A => n7795, B => n7794, S => n7793, Z => n7796);
   U19321 : OAI221_X1 port map( B1 => n7798, B2 => n7859, C1 => n7797, C2 => 
                           n8140, A => n7796, ZN => n7807);
   U19322 : XOR2_X1 port map( A => n7800, B => n7799, Z => n7805);
   U19323 : AOI21_X1 port map( B1 => n7803, B2 => n7802, A => n7801, ZN => 
                           n7804);
   U19324 : OAI22_X1 port map( A1 => n7805, A2 => n2186, B1 => n7804, B2 => 
                           n2252, ZN => n7806);
   U19325 : AOI211_X1 port map( C1 => n366, C2 => n7808, A => n7807, B => n7806
                           , ZN => n7810);
   U19326 : OAI22_X1 port map( A1 => n7810, A2 => n7980, B1 => n7979, B2 => 
                           n7809, ZN => n8669);
   U19327 : OAI21_X1 port map( B1 => n2278, B2 => n8014, A => n7811, ZN => 
                           n8053);
   U19328 : INV_X1 port map( A => n8053, ZN => n7812);
   U19329 : OAI22_X1 port map( A1 => n7815, A2 => n7991, B1 => n7812, B2 => 
                           n7989, ZN => n8054);
   U19330 : AOI222_X1 port map( A1 => n7994, A2 => n7813, B1 => n8034, B2 => 
                           n8054, C1 => n8043, C2 => n8012, ZN => n7814);
   U19331 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n600, B2 => 
                           n7816, C1 => n7815, C2 => n8089, A => n7814, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n392);
   U19332 : INV_X1 port map( A => n7817, ZN => n7824);
   U19333 : XOR2_X1 port map( A => n7818, B => n7824, Z => n7840);
   U19334 : AOI222_X1 port map( A1 => n7819, A2 => n7955, B1 => n7954, B2 => 
                           n7885, C1 => n7953, C2 => n7851, ZN => n7820);
   U19335 : OAI221_X1 port map( B1 => n8302, B2 => n2242, C1 => 
                           DataPath_ALUhw_SHIFTER_HW_n181, C2 => n7821, A => 
                           n7820, ZN => n7823);
   U19336 : OAI222_X1 port map( A1 => n8298, A2 => n8032, B1 => n8301, B2 => 
                           n8025, C1 => n8297, C2 => n8030, ZN => n7822);
   U19337 : NOR4_X1 port map( A1 => n7823, A2 => n7822, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n385, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n390, ZN => n7827);
   U19338 : XOR2_X1 port map( A => n7825, B => n7824, Z => n7826);
   U19339 : OAI22_X1 port map( A1 => n7827, A2 => n8140, B1 => n7826, B2 => 
                           n7859, ZN => n7839);
   U19340 : XOR2_X1 port map( A => n714, B => n1853, Z => n7830);
   U19341 : MUX2_X1 port map( A => n7965, B => n2187, S => n7832, Z => n7829);
   U19342 : OAI21_X1 port map( B1 => n7830, B2 => n2253, A => n7829, ZN => 
                           n7837);
   U19343 : INV_X1 port map( A => n7831, ZN => n7849);
   U19344 : XOR2_X1 port map( A => n7849, B => n1853, Z => n7834);
   U19345 : MUX2_X1 port map( A => n2187, B => n7969, S => n7832, Z => n7833);
   U19346 : OAI21_X1 port map( B1 => n7834, B2 => n2253, A => n7833, ZN => 
                           n7836);
   U19347 : MUX2_X1 port map( A => n7837, B => n7836, S => n7835, Z => n7838);
   U19348 : AOI211_X1 port map( C1 => n366, C2 => n7840, A => n7839, B => n7838
                           , ZN => n7842);
   U19349 : OAI22_X1 port map( A1 => n7842, A2 => n7980, B1 => n7979, B2 => 
                           n7841, ZN => n8670);
   U19350 : OAI21_X1 port map( B1 => n2278, B2 => n8029, A => n7843, ZN => 
                           n8062);
   U19351 : INV_X1 port map( A => n8062, ZN => n7844);
   U19352 : OAI22_X1 port map( A1 => n7847, A2 => n7991, B1 => n7844, B2 => 
                           n7989, ZN => n8063);
   U19353 : AOI222_X1 port map( A1 => n7994, A2 => n7845, B1 => n8034, B2 => 
                           n8063, C1 => n8043, C2 => n8027, ZN => n7846);
   U19354 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n600, B2 => 
                           n7848, C1 => n7847, C2 => n8089, A => n7846, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n405);
   U19355 : XOR2_X1 port map( A => n7865, B => n7863, Z => n7858);
   U19356 : AOI21_X1 port map( B1 => n1027, B2 => n7850, A => n7849, ZN => 
                           n7857);
   U19357 : AOI222_X1 port map( A1 => n7955, A2 => n7851, B1 => n7954, B2 => 
                           n7919, C1 => n7953, C2 => n7885, ZN => n7852);
   U19358 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n181, B2 => 
                           n7853, C1 => n8298, C2 => n8025, A => n7852, ZN => 
                           n7855);
   U19359 : OAI222_X1 port map( A1 => n8297, A2 => n8032, B1 => n8301, B2 => 
                           n2242, C1 => n8296, C2 => n8030, ZN => n7854);
   U19360 : NOR4_X1 port map( A1 => n7855, A2 => n7854, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n397, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n403, ZN => n7856);
   U19361 : OAI222_X1 port map( A1 => n7858, A2 => n2187, B1 => n7857, B2 => 
                           n2252, C1 => n7856, C2 => n8140, ZN => n7871);
   U19362 : INV_X1 port map( A => n7859, ZN => n7862);
   U19363 : INV_X1 port map( A => n7860, ZN => n7861);
   U19364 : MUX2_X1 port map( A => n366, B => n7862, S => n7861, Z => n7870);
   U19365 : NOR2_X1 port map( A1 => n7863, A2 => n7965, ZN => n7868);
   U19366 : NOR2_X1 port map( A1 => n7864, A2 => n7969, ZN => n7867);
   U19367 : INV_X1 port map( A => n7865, ZN => n7866);
   U19368 : MUX2_X1 port map( A => n7868, B => n7867, S => n7866, Z => n7869);
   U19369 : NOR3_X1 port map( A1 => n7871, A2 => n7870, A3 => n7869, ZN => 
                           n7873);
   U19370 : OAI22_X1 port map( A1 => n7873, A2 => n7980, B1 => n7979, B2 => 
                           n7872, ZN => n8671);
   U19371 : OAI21_X1 port map( B1 => n2278, B2 => n8018, A => n7874, ZN => 
                           n8072);
   U19372 : INV_X1 port map( A => n8072, ZN => n7875);
   U19373 : OAI22_X1 port map( A1 => n7878, A2 => n7991, B1 => n7875, B2 => 
                           n7989, ZN => n8074);
   U19374 : AOI222_X1 port map( A1 => n7994, A2 => n7876, B1 => n8034, B2 => 
                           n8074, C1 => n8043, C2 => n8015, ZN => n7877);
   U19375 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n600, B2 => 
                           n7879, C1 => n7878, C2 => n8089, A => n7877, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n432);
   U19376 : NAND2_X1 port map( A1 => n8222, A2 => n7960, ZN => n7952);
   U19377 : INV_X1 port map( A => n7952, ZN => n7881);
   U19378 : OAI21_X1 port map( B1 => n7951, B2 => n7881, A => n7880, ZN => 
                           n7916);
   U19379 : INV_X1 port map( A => n7916, ZN => n7882);
   U19380 : OAI21_X1 port map( B1 => n7883, B2 => n7882, A => n7889, ZN => 
                           n7884);
   U19381 : XOR2_X1 port map( A => n7884, B => n7892, Z => n7906);
   U19382 : AOI222_X1 port map( A1 => n7955, A2 => n7885, B1 => n7954, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n344, C1 => n7953, C2 => 
                           n7919, ZN => n7886);
   U19383 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n181, B2 => 
                           n11493, C1 => n8297, C2 => n8025, A => n7886, ZN => 
                           n7888);
   U19384 : OAI222_X1 port map( A1 => n8296, A2 => n8032, B1 => n8298, B2 => 
                           n2242, C1 => n8295, C2 => n8030, ZN => n7887);
   U19385 : NOR4_X1 port map( A1 => n7888, A2 => n7887, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n424, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n430, ZN => n7894);
   U19386 : INV_X1 port map( A => n7889, ZN => n7890);
   U19387 : AOI21_X1 port map( B1 => n11526, B2 => n7918, A => n7890, ZN => 
                           n7891);
   U19388 : XOR2_X1 port map( A => n7892, B => n7891, Z => n7893);
   U19389 : NAND2_X1 port map( A1 => n2272, A2 => n12929, ZN => n7961);
   U19390 : OAI22_X1 port map( A1 => n7894, A2 => n8140, B1 => n7893, B2 => 
                           n7961, ZN => n7905);
   U19391 : XOR2_X1 port map( A => n1783, B => n1857, Z => n7897);
   U19392 : MUX2_X1 port map( A => n7965, B => n2186, S => n7899, Z => n7896);
   U19393 : OAI21_X1 port map( B1 => n7897, B2 => n2254, A => n7896, ZN => 
                           n7903);
   U19394 : INV_X1 port map( A => n7898, ZN => n7934);
   U19395 : XOR2_X1 port map( A => n7934, B => n1857, Z => n7901);
   U19396 : MUX2_X1 port map( A => n2186, B => n7969, S => n7899, Z => n7900);
   U19397 : OAI21_X1 port map( B1 => n7901, B2 => n2255, A => n7900, ZN => 
                           n7902);
   U19398 : MUX2_X1 port map( A => n7903, B => n7902, S => n1702, Z => n7904);
   U19399 : AOI211_X1 port map( C1 => n367, C2 => n7906, A => n7905, B => n7904
                           , ZN => n7908);
   U19400 : OAI22_X1 port map( A1 => n7908, A2 => n7980, B1 => n7979, B2 => 
                           n7907, ZN => n8672);
   U19401 : OAI21_X1 port map( B1 => n2278, B2 => n8024, A => n7909, ZN => 
                           n8100);
   U19402 : INV_X1 port map( A => n8100, ZN => n7910);
   U19403 : OAI22_X1 port map( A1 => n7915, A2 => n7991, B1 => n7910, B2 => 
                           n7989, ZN => n7911);
   U19404 : INV_X1 port map( A => n7911, ZN => DataPath_ALUhw_SHIFTER_HW_n529);
   U19405 : AOI222_X1 port map( A1 => n7913, A2 => n8073, B1 => n8043, B2 => 
                           n8020, C1 => n7994, C2 => n7912, ZN => n7914);
   U19406 : OAI221_X1 port map( B1 => n7915, B2 => n8089, C1 => 
                           DataPath_ALUhw_SHIFTER_HW_n529, C2 => n7997, A => 
                           n7914, ZN => DataPath_ALUhw_SHIFTER_HW_n445);
   U19407 : XOR2_X1 port map( A => n7916, B => n7918, Z => n7941);
   U19408 : INV_X1 port map( A => n11526, ZN => n7917);
   U19409 : XOR2_X1 port map( A => n7918, B => n7917, Z => n7931);
   U19410 : AOI222_X1 port map( A1 => n7955, A2 => n7919, B1 => n7954, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n380, C1 => n7953, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n344, ZN => n7920);
   U19411 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n181, B2 => 
                           n8303, C1 => n8296, C2 => n8025, A => n7920, ZN => 
                           n7922);
   U19412 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n445, ZN => n8294);
   U19413 : OAI222_X1 port map( A1 => n8295, A2 => n8032, B1 => n8297, B2 => 
                           n2242, C1 => n8294, C2 => n8030, ZN => n7921);
   U19414 : NOR4_X1 port map( A1 => n7922, A2 => n7921, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n437, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n443, ZN => n7930);
   U19415 : NAND2_X1 port map( A1 => n7924, A2 => n7923, ZN => n7928);
   U19416 : NAND2_X1 port map( A1 => n7925, A2 => n7932, ZN => n7927);
   U19417 : INV_X1 port map( A => n7933, ZN => n7926);
   U19418 : MUX2_X1 port map( A => n7928, B => n7927, S => n7926, Z => n7929);
   U19419 : OAI221_X1 port map( B1 => n7931, B2 => n7961, C1 => n7930, C2 => 
                           n8140, A => n7929, ZN => n7940);
   U19420 : XOR2_X1 port map( A => n7933, B => n7932, Z => n7938);
   U19421 : AOI21_X1 port map( B1 => n7936, B2 => n7935, A => n7934, ZN => 
                           n7937);
   U19422 : OAI22_X1 port map( A1 => n7938, A2 => n2186, B1 => n7937, B2 => 
                           n2253, ZN => n7939);
   U19423 : AOI211_X1 port map( C1 => n367, C2 => n7941, A => n7940, B => n7939
                           , ZN => n7943);
   U19424 : OAI22_X1 port map( A1 => n7943, A2 => n7980, B1 => n7979, B2 => 
                           n7942, ZN => n8673);
   U19425 : OAI21_X1 port map( B1 => n2278, B2 => n8006, A => n7944, ZN => 
                           n8108);
   U19426 : INV_X1 port map( A => n8108, ZN => n7945);
   U19427 : OAI22_X1 port map( A1 => n7950, A2 => n7991, B1 => n7945, B2 => 
                           n7989, ZN => n7946);
   U19428 : INV_X1 port map( A => n7946, ZN => DataPath_ALUhw_SHIFTER_HW_n540);
   U19429 : AOI222_X1 port map( A1 => n7948, A2 => n8073, B1 => n8043, B2 => 
                           n8003, C1 => n7994, C2 => n7947, ZN => n7949);
   U19430 : OAI221_X1 port map( B1 => n7950, B2 => n8089, C1 => 
                           DataPath_ALUhw_SHIFTER_HW_n540, C2 => n7997, A => 
                           n7949, ZN => DataPath_ALUhw_SHIFTER_HW_n455);
   U19431 : INV_X1 port map( A => n7951, ZN => n7959);
   U19432 : XOR2_X1 port map( A => n7952, B => n7959, Z => n7978);
   U19433 : AOI222_X1 port map( A1 => n7955, A2 => 
                           DataPath_ALUhw_SHIFTER_HW_n344, B1 => n7954, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n392, C1 => n7953, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n380, ZN => n7956);
   U19434 : OAI221_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n181, B2 => 
                           n8302, C1 => n8295, C2 => n8025, A => n7956, ZN => 
                           n7958);
   U19435 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n455, ZN => n8293);
   U19436 : OAI222_X1 port map( A1 => n8294, A2 => n8032, B1 => n8296, B2 => 
                           n2242, C1 => n8293, C2 => n8030, ZN => n7957);
   U19437 : NOR4_X1 port map( A1 => n7958, A2 => n7957, A3 => 
                           DataPath_ALUhw_SHIFTER_HW_n450, A4 => 
                           DataPath_ALUhw_SHIFTER_HW_n453, ZN => n7963);
   U19438 : XOR2_X1 port map( A => n7960, B => n7959, Z => n7962);
   U19439 : OAI22_X1 port map( A1 => n7963, A2 => n8140, B1 => n7962, B2 => 
                           n7961, ZN => n7977);
   U19440 : XOR2_X1 port map( A => n773, B => n1856, Z => n7967);
   U19441 : MUX2_X1 port map( A => n7965, B => n2186, S => n7968, Z => n7966);
   U19442 : OAI21_X1 port map( B1 => n7967, B2 => n2255, A => n7966, ZN => 
                           n7975);
   U19443 : MUX2_X1 port map( A => n2186, B => n7969, S => n7968, Z => n7971);
   U19444 : OAI21_X1 port map( B1 => n7972, B2 => n2255, A => n7971, ZN => 
                           n7974);
   U19445 : MUX2_X1 port map( A => n7975, B => n7974, S => n7973, Z => n7976);
   U19446 : AOI211_X1 port map( C1 => n367, C2 => n7978, A => n7977, B => n7976
                           , ZN => n7981);
   U19447 : OAI22_X1 port map( A1 => n7981, A2 => n7980, B1 => n7979, B2 => 
                           n424, ZN => n8674);
   U19448 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n182, ZN => n8300);
   U19449 : OAI21_X1 port map( B1 => n2278, B2 => n8038, A => n7982, ZN => 
                           n7983);
   U19450 : INV_X1 port map( A => n7983, ZN => n8090);
   U19451 : OAI22_X1 port map( A1 => n2278, A2 => n7986, B1 => n2273, B2 => 
                           n8090, ZN => n8087);
   U19452 : AOI222_X1 port map( A1 => n7994, A2 => n7984, B1 => n8034, B2 => 
                           n8087, C1 => n8043, C2 => n8035, ZN => n7985);
   U19453 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n181, ZN => n8299);
   U19454 : OAI21_X1 port map( B1 => n2278, B2 => n8002, A => n7988, ZN => 
                           n8115);
   U19455 : INV_X1 port map( A => n8115, ZN => n7990);
   U19456 : OAI22_X1 port map( A1 => n7998, A2 => n7991, B1 => n7990, B2 => 
                           n7989, ZN => n7992);
   U19457 : INV_X1 port map( A => n7992, ZN => DataPath_ALUhw_SHIFTER_HW_n411);
   U19458 : AOI222_X1 port map( A1 => n7995, A2 => n8073, B1 => n8043, B2 => 
                           n7999, C1 => n7994, C2 => n7993, ZN => n7996);
   U19459 : AOI222_X1 port map( A1 => n8116, A2 => n8000, B1 => n8034, B2 => 
                           n8126, C1 => n7999, C2 => n8073, ZN => n8001);
   U19460 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n171, ZN => n8292);
   U19461 : AOI222_X1 port map( A1 => n8116, A2 => n8004, B1 => n8034, B2 => 
                           n8114, C1 => n8003, C2 => n8073, ZN => n8005);
   U19462 : OAI221_X1 port map( B1 => n8006, B2 => n8037, C1 => 
                           DataPath_ALUhw_SHIFTER_HW_n540, C2 => n2134, A => 
                           n8005, ZN => DataPath_ALUhw_SHIFTER_HW_n161);
   U19463 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n161, ZN => n8291);
   U19464 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n192, ZN => n8314);
   U19465 : INV_X1 port map( A => n8007, ZN => n8011);
   U19466 : AOI222_X1 port map( A1 => n8043, A2 => n8041, B1 => n8034, B2 => 
                           n8048, C1 => n8116, C2 => n8008, ZN => n8009);
   U19467 : AOI222_X1 port map( A1 => n8012, A2 => n8073, B1 => n8034, B2 => 
                           n8057, C1 => n8043, C2 => n8054, ZN => n8013);
   U19468 : OAI221_X1 port map( B1 => n8055, B2 => n8089, C1 => n8014, C2 => 
                           n8037, A => n8013, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n152);
   U19469 : INV_X1 port map( A => n8015, ZN => n8019);
   U19470 : AOI222_X1 port map( A1 => n8043, A2 => n8074, B1 => n8034, B2 => 
                           n8078, C1 => n8116, C2 => n8016, ZN => n8017);
   U19471 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n156, ZN => n8288);
   U19472 : AOI222_X1 port map( A1 => n8116, A2 => n8021, B1 => n8034, B2 => 
                           n8107, C1 => n8020, C2 => n8073, ZN => n8022);
   U19473 : OAI221_X1 port map( B1 => n8024, B2 => n8037, C1 => 
                           DataPath_ALUhw_SHIFTER_HW_n529, C2 => n2134, A => 
                           n8022, ZN => DataPath_ALUhw_SHIFTER_HW_n164);
   U19474 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n164, ZN => n8287);
   U19475 : AOI222_X1 port map( A1 => n8027, A2 => n8073, B1 => n8034, B2 => 
                           n8066, C1 => n8043, C2 => n8063, ZN => n8028);
   U19476 : OAI221_X1 port map( B1 => n8064, B2 => n8089, C1 => n8029, C2 => 
                           n8037, A => n8028, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n172);
   U19477 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n152, ZN => n8289);
   U19478 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n172, ZN => n8286);
   U19479 : OAI22_X1 port map( A1 => n8289, A2 => n8099, B1 => n8286, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n157);
   U19480 : AOI222_X1 port map( A1 => n8035, A2 => n8073, B1 => n8034, B2 => 
                           n8033, C1 => n8043, C2 => n8087, ZN => n8036);
   U19481 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n150, ZN => n8304);
   U19482 : OAI22_X1 port map( A1 => n8286, A2 => n8099, B1 => n8288, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n174);
   U19483 : AOI22_X1 port map( A1 => n8041, A2 => n8073, B1 => n8116, B2 => 
                           n8040, ZN => n8051);
   U19484 : NAND3_X1 port map( A1 => n11538, A2 => n8181, A3 => n2250, ZN => 
                           n8120);
   U19485 : INV_X1 port map( A => n8120, ZN => n8042);
   U19486 : NAND2_X1 port map( A1 => n11538, A2 => n8043, ZN => n8092);
   U19487 : INV_X1 port map( A => n8092, ZN => n8127);
   U19488 : NAND2_X1 port map( A1 => DataPath_ALUhw_SHIFTER_HW_n549, A2 => 
                           n8043, ZN => n8122);
   U19489 : OAI21_X1 port map( B1 => DataPath_ALUhw_SHIFTER_HW_n597, B2 => 
                           n8120, A => n8102, ZN => n8044);
   U19490 : INV_X1 port map( A => n8044, ZN => n8075);
   U19491 : OAI22_X1 port map( A1 => n8046, A2 => n8122, B1 => n17240, B2 => 
                           n8075, ZN => n8047);
   U19492 : AOI221_X1 port map( B1 => n282, B2 => n8049, C1 => n8127, C2 => 
                           n8048, A => n8047, ZN => n8050);
   U19493 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n151, ZN => n8290);
   U19494 : OAI22_X1 port map( A1 => n8288, A2 => n8099, B1 => n8287, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n184);
   U19495 : AOI22_X1 port map( A1 => n8054, A2 => n8073, B1 => n8116, B2 => 
                           n8053, ZN => n8060);
   U19496 : OAI22_X1 port map( A1 => n8055, A2 => n8122, B1 => n2238, B2 => 
                           n8075, ZN => n8056);
   U19497 : AOI221_X1 port map( B1 => n282, B2 => n8058, C1 => n8127, C2 => 
                           n8057, A => n8056, ZN => n8059);
   U19498 : OAI211_X1 port map( C1 => n8061, C2 => n8082, A => n8060, B => 
                           n8059, ZN => DataPath_ALUhw_SHIFTER_HW_n201);
   U19499 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n201, ZN => n8284);
   U19500 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n179, ZN => n8285);
   U19501 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n155, ZN => n8311);
   U19502 : OAI22_X1 port map( A1 => n8287, A2 => n8099, B1 => n8291, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n193);
   U19503 : AOI22_X1 port map( A1 => n8063, A2 => n8073, B1 => n8116, B2 => 
                           n8062, ZN => n8069);
   U19504 : OAI22_X1 port map( A1 => n8064, A2 => n8122, B1 => n2239, B2 => 
                           n8075, ZN => n8065);
   U19505 : AOI221_X1 port map( B1 => n282, B2 => n8067, C1 => n8127, C2 => 
                           n8066, A => n8065, ZN => n8068);
   U19506 : OAI211_X1 port map( C1 => n8070, C2 => n8082, A => n8069, B => 
                           n8068, ZN => DataPath_ALUhw_SHIFTER_HW_n211);
   U19507 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n211, ZN => n8283);
   U19508 : OAI22_X1 port map( A1 => n8291, A2 => n8099, B1 => n8292, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n200);
   U19509 : OAI22_X1 port map( A1 => n8292, A2 => n8099, B1 => n522, B2 => 
                           n2242, ZN => n8071);
   U19510 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n179, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n161, A => n8071, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n203);
   U19511 : AOI22_X1 port map( A1 => n8074, A2 => n8073, B1 => n8116, B2 => 
                           n8072, ZN => n8081);
   U19512 : OAI22_X1 port map( A1 => n8076, A2 => n8122, B1 => n2240, B2 => 
                           n8075, ZN => n8077);
   U19513 : AOI221_X1 port map( B1 => n282, B2 => n8079, C1 => n8127, C2 => 
                           n8078, A => n8077, ZN => n8080);
   U19514 : OAI211_X1 port map( C1 => n8083, C2 => n8082, A => n8081, B => 
                           n8080, ZN => DataPath_ALUhw_SHIFTER_HW_n219);
   U19515 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n219, ZN => n8282);
   U19516 : OAI22_X1 port map( A1 => n522, A2 => n8099, B1 => n8285, B2 => 
                           n2242, ZN => n8084);
   U19517 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n201, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n171, A => n8084, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n213);
   U19518 : OAI22_X1 port map( A1 => n8285, A2 => n8099, B1 => n8284, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n268);
   U19519 : OAI22_X1 port map( A1 => n8284, A2 => n8099, B1 => n8283, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n418);
   U19520 : INV_X1 port map( A => DataPath_ALUhw_SHIFTER_HW_n146, ZN => n11490)
                           ;
   U19521 : OAI22_X1 port map( A1 => n8296, A2 => n8099, B1 => n8295, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n467);
   U19522 : OAI22_X1 port map( A1 => n8295, A2 => n8099, B1 => n8294, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n482);
   U19523 : OAI22_X1 port map( A1 => n8294, A2 => n8099, B1 => n8293, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n495);
   U19524 : OAI22_X1 port map( A1 => n8293, A2 => n8099, B1 => n520, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n508);
   U19525 : OAI22_X1 port map( A1 => n11490, A2 => n2242, B1 => n520, B2 => 
                           n8099, ZN => n8085);
   U19526 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n151, C1 => n8315, C2 => 
                           DataPath_ALUhw_SHIFTER_HW_n455, A => n8085, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n510);
   U19527 : OAI22_X1 port map( A1 => n8290, A2 => n2242, B1 => n11490, B2 => 
                           n8099, ZN => n8086);
   U19528 : AOI221_X1 port map( B1 => n8305, B2 => 
                           DataPath_ALUhw_SHIFTER_HW_n152, C1 => n8315, C2 => 
                           n521, A => n8086, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n523);
   U19529 : OAI22_X1 port map( A1 => n8290, A2 => n8099, B1 => n8289, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n552);
   U19530 : INV_X1 port map( A => n8122, ZN => n8098);
   U19531 : INV_X1 port map( A => n8087, ZN => n8088);
   U19532 : OAI22_X1 port map( A1 => n8094, A2 => n8120, B1 => n8093, B2 => 
                           n8092, ZN => n8095);
   U19533 : AOI211_X1 port map( C1 => n8098, C2 => n8097, A => n8096, B => 
                           n8095, ZN => DataPath_ALUhw_SHIFTER_HW_n587);
   U19534 : OAI22_X1 port map( A1 => n8283, A2 => n8099, B1 => n8282, B2 => 
                           n2242, ZN => DataPath_ALUhw_SHIFTER_HW_n606);
   U19535 : AOI22_X1 port map( A1 => n8118, A2 => n8101, B1 => n8116, B2 => 
                           n8100, ZN => DataPath_ALUhw_SHIFTER_HW_n621);
   U19536 : INV_X1 port map( A => n8102, ZN => n8125);
   U19537 : INV_X1 port map( A => n8103, ZN => n8104);
   U19538 : OAI22_X1 port map( A1 => n8105, A2 => n8122, B1 => n8104, B2 => 
                           n8120, ZN => n8106);
   U19539 : AOI221_X1 port map( B1 => n8127, B2 => n8107, C1 => n8125, C2 => 
                           n2228, A => n8106, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n622);
   U19540 : AOI22_X1 port map( A1 => n8118, A2 => n8109, B1 => n8116, B2 => 
                           n8108, ZN => DataPath_ALUhw_SHIFTER_HW_n625);
   U19541 : INV_X1 port map( A => n8110, ZN => n8111);
   U19542 : OAI22_X1 port map( A1 => n8112, A2 => n8122, B1 => n8111, B2 => 
                           n8120, ZN => n8113);
   U19543 : AOI221_X1 port map( B1 => n8127, B2 => n8114, C1 => n8125, C2 => 
                           n2231, A => n8113, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n626);
   U19544 : AOI22_X1 port map( A1 => n8118, A2 => n8117, B1 => n8116, B2 => 
                           n8115, ZN => DataPath_ALUhw_SHIFTER_HW_n635);
   U19545 : INV_X1 port map( A => n8119, ZN => n8121);
   U19546 : OAI22_X1 port map( A1 => n8123, A2 => n8122, B1 => n8121, B2 => 
                           n8120, ZN => n8124);
   U19547 : AOI221_X1 port map( B1 => n8127, B2 => n8126, C1 => n8125, C2 => 
                           n2146, A => n8124, ZN => 
                           DataPath_ALUhw_SHIFTER_HW_n636);
   U19548 : XOR2_X1 port map( A => n1439, B => n8128, Z => n8132);
   U19549 : NAND2_X1 port map( A1 => n1872, A2 => n1090, ZN => n8141);
   U19550 : INV_X1 port map( A => n8141, ZN => n8131);
   U19551 : XOR2_X1 port map( A => n8132, B => n8131, Z => n8133);
   U19552 : MUX2_X1 port map( A => n8134, B => n8133, S => n2243, Z => n8139);
   U19553 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2987, S => 
                           n2243, Z => n8137);
   U19554 : MUX2_X1 port map( A => n2986, B => DataPath_ALUhw_BWISE_n72, S => 
                           n2243, Z => n8136);
   U19555 : MUX2_X1 port map( A => n8137, B => n8136, S => n797, Z => n8138);
   U19556 : AOI22_X1 port map( A1 => n2258, A2 => n8139, B1 => n8322, B2 => 
                           n8138, ZN => DataPath_ALUhw_MUXOUT_n3);
   U19557 : INV_X1 port map( A => n8140, ZN => n8321);
   U19558 : OAI21_X1 port map( B1 => n1872, B2 => n1090, A => n8141, ZN => 
                           n8148);
   U19559 : INV_X1 port map( A => n8143, ZN => n8144);
   U19560 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2987, S => 
                           n8144, Z => n8146);
   U19561 : MUX2_X1 port map( A => n2986, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8144, Z => n8145);
   U19562 : MUX2_X1 port map( A => n8146, B => n8145, S => n2202, Z => n8147);
   U19563 : AOI22_X1 port map( A1 => n2258, A2 => n8148, B1 => n8322, B2 => 
                           n8147, ZN => DataPath_ALUhw_MUXOUT_n9);
   U19564 : XOR2_X1 port map( A => n8149, B => n12927, Z => n11507);
   U19565 : XOR2_X1 port map( A => n1532, B => n8150, Z => n8155);
   U19566 : NOR2_X1 port map( A1 => n956, A2 => n8152, ZN => n8153);
   U19567 : XOR2_X1 port map( A => n8155, B => n8153, Z => n8157);
   U19568 : XOR2_X1 port map( A => n8154, B => n8155, Z => n8156);
   U19569 : MUX2_X1 port map( A => n8157, B => n8156, S => n2245, Z => n8162);
   U19570 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n1520, Z => n8160);
   U19571 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n1520, Z => n8159);
   U19572 : MUX2_X1 port map( A => n8160, B => n8159, S => n2245, Z => n8161);
   U19573 : AOI22_X1 port map( A1 => n2258, A2 => n8162, B1 => n8322, B2 => 
                           n8161, ZN => DataPath_ALUhw_MUXOUT_n11);
   U19574 : OAI21_X1 port map( B1 => n8165, B2 => n956, A => n1149, ZN => n8170
                           );
   U19575 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n8166, Z => n8168);
   U19576 : MUX2_X1 port map( A => n2986, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8166, Z => n8167);
   U19577 : MUX2_X1 port map( A => n8168, B => n8167, S => n1933, Z => n8169);
   U19578 : AOI22_X1 port map( A1 => n2258, A2 => n8170, B1 => n8322, B2 => 
                           n8169, ZN => DataPath_ALUhw_MUXOUT_n13);
   U19579 : XOR2_X1 port map( A => n8171, B => n1358, Z => n8172);
   U19580 : XOR2_X1 port map( A => n8172, B => n1237, Z => n8174);
   U19581 : XOR2_X1 port map( A => n8172, B => n17248, Z => n8173);
   U19582 : MUX2_X1 port map( A => n8174, B => n8173, S => n2247, Z => n8178);
   U19583 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n2247, Z => n8176);
   U19584 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n2248, Z => n8175);
   U19585 : MUX2_X1 port map( A => n8176, B => n8175, S => n788, Z => n8177);
   U19586 : AOI22_X1 port map( A1 => n2258, A2 => n8178, B1 => n8322, B2 => 
                           n8177, ZN => DataPath_ALUhw_MUXOUT_n15);
   U19587 : OAI21_X1 port map( B1 => n1875, B2 => n453, A => n17211, ZN => 
                           n8185);
   U19588 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n8181, Z => n8183);
   U19589 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8181, Z => n8182);
   U19590 : MUX2_X1 port map( A => n8183, B => n8182, S => n2241, Z => n8184);
   U19591 : AOI22_X1 port map( A1 => n2258, A2 => n8185, B1 => n8322, B2 => 
                           n8184, ZN => DataPath_ALUhw_MUXOUT_n17);
   U19592 : XOR2_X1 port map( A => n8186, B => n12926, Z => n11512);
   U19593 : XOR2_X1 port map( A => n1320, B => n1118, Z => n8191);
   U19594 : INV_X1 port map( A => n1246, ZN => n8190);
   U19595 : XOR2_X1 port map( A => n8191, B => n8190, Z => n8193);
   U19596 : XOR2_X1 port map( A => n8191, B => n1710, Z => n8192);
   U19597 : MUX2_X1 port map( A => n8193, B => n8192, S => n2250, Z => n8197);
   U19598 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n2228, Z => n8195);
   U19599 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n2228, Z => n8194);
   U19600 : MUX2_X1 port map( A => n8195, B => n8194, S => n804, Z => n8196);
   U19601 : AOI22_X1 port map( A1 => n2258, A2 => n8197, B1 => n8322, B2 => 
                           n8196, ZN => DataPath_ALUhw_MUXOUT_n19);
   U19602 : OAI21_X1 port map( B1 => n1878, B2 => n829, A => n598, ZN => n8203)
                           ;
   U19603 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n2130, Z => n8201);
   U19604 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n2130, Z => n8200);
   U19605 : MUX2_X1 port map( A => n8201, B => n8200, S => n2231, Z => n8202);
   U19606 : AOI22_X1 port map( A1 => n2258, A2 => n8203, B1 => n8322, B2 => 
                           n8202, ZN => DataPath_ALUhw_MUXOUT_n25);
   U19607 : INV_X1 port map( A => n777, ZN => n8207);
   U19608 : AOI21_X1 port map( B1 => n661, B2 => n8207, A => n2252, ZN => n8214
                           );
   U19609 : NAND2_X1 port map( A1 => n770, A2 => n2259, ZN => n8209);
   U19610 : MUX2_X1 port map( A => n8209, B => n2261, S => n8207, Z => n8213);
   U19611 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n71, S => 
                           n17161, Z => n8211);
   U19612 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n72, B => n2986, S => 
                           n2263, Z => n8210);
   U19613 : MUX2_X1 port map( A => n8211, B => n8210, S => n2146, Z => n8212);
   U19614 : AOI22_X1 port map( A1 => n8214, A2 => n8213, B1 => n8322, B2 => 
                           n8212, ZN => DataPath_ALUhw_MUXOUT_n47);
   U19615 : INV_X1 port map( A => n8215, ZN => n8216);
   U19616 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n8216, Z => n8219);
   U19617 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8216, Z => n8218);
   U19618 : MUX2_X1 port map( A => n8219, B => n8218, S => n8217, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_80_port);
   U19619 : OAI21_X1 port map( B1 => n1894, B2 => n853, A => n742, ZN => n11584
                           );
   U19620 : XOR2_X1 port map( A => n8222, B => n12929, Z => n11501);
   U19621 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n8223, Z => n8225);
   U19622 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8223, Z => n8224);
   U19623 : MUX2_X1 port map( A => n8225, B => n8224, S => n8229, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_79_port);
   U19624 : XOR2_X1 port map( A => n8227, B => n884, Z => n8228);
   U19625 : XOR2_X1 port map( A => n8228, B => n2166, Z => n8231);
   U19626 : XOR2_X1 port map( A => n8228, B => n1278, Z => n8230);
   U19627 : MUX2_X1 port map( A => n8231, B => n8230, S => n8229, Z => n11585);
   U19628 : INV_X1 port map( A => n8232, ZN => n8233);
   U19629 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n8233, Z => n8236);
   U19630 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8233, Z => n8235);
   U19631 : MUX2_X1 port map( A => n8236, B => n8235, S => n8234, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_78_port);
   U19632 : OAI21_X1 port map( B1 => n8239, B2 => n1581, A => n8237, ZN => 
                           n11586);
   U19633 : XOR2_X1 port map( A => n8240, B => n1715, Z => n8242);
   U19634 : XOR2_X1 port map( A => n8242, B => n1709, Z => n8244);
   U19635 : INV_X1 port map( A => n8254, ZN => n8241);
   U19636 : XOR2_X1 port map( A => n8242, B => n8241, Z => n8243);
   U19637 : MUX2_X1 port map( A => n8244, B => n8243, S => n2265, Z => n8249);
   U19638 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n2265, Z => n8247);
   U19639 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n2265, Z => n8246);
   U19640 : MUX2_X1 port map( A => n8247, B => n8246, S => n1935, Z => n8248);
   U19641 : AOI22_X1 port map( A1 => n2258, A2 => n8249, B1 => n8322, B2 => 
                           n8248, ZN => DataPath_ALUhw_MUXOUT_n61);
   U19642 : INV_X1 port map( A => n8250, ZN => n8251);
   U19643 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n8251, Z => n8253);
   U19644 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8251, Z => n8252);
   U19645 : MUX2_X1 port map( A => n8253, B => n8252, S => n1934, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_76_port);
   U19646 : OAI21_X1 port map( B1 => n1892, B2 => n1429, A => n1480, ZN => 
                           n11587);
   U19647 : XOR2_X1 port map( A => n8256, B => n12928, Z => n11502);
   U19648 : XOR2_X1 port map( A => n8258, B => n8257, Z => n8260);
   U19649 : XOR2_X1 port map( A => n8260, B => n1826, Z => n8262);
   U19650 : INV_X1 port map( A => n8268, ZN => n8259);
   U19651 : XOR2_X1 port map( A => n8260, B => n8259, Z => n8261);
   U19652 : MUX2_X1 port map( A => n8262, B => n8261, S => n2267, Z => n8267);
   U19653 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2986, S => 
                           n2207, Z => n8265);
   U19654 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n2207, Z => n8264);
   U19655 : MUX2_X1 port map( A => n8265, B => n8264, S => n2268, Z => n8266);
   U19656 : AOI22_X1 port map( A1 => n2258, A2 => n8267, B1 => n8322, B2 => 
                           n8266, ZN => DataPath_ALUhw_MUXOUT_n65);
   U19657 : OAI21_X1 port map( B1 => n1893, B2 => n8269, A => n8268, ZN => 
                           n8275);
   U19658 : INV_X1 port map( A => n8270, ZN => n8271);
   U19659 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n71, B => n2987, S => 
                           n8271, Z => n8273);
   U19660 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n72, S => 
                           n8271, Z => n8272);
   U19661 : MUX2_X1 port map( A => n8273, B => n8272, S => n2211, Z => n8274);
   U19662 : AOI22_X1 port map( A1 => n2258, A2 => n8275, B1 => n8322, B2 => 
                           n8274, ZN => DataPath_ALUhw_MUXOUT_n67);
   U19663 : MUX2_X1 port map( A => n2985, B => DataPath_ALUhw_BWISE_n71, S => 
                           n2269, Z => n8279);
   U19664 : MUX2_X1 port map( A => DataPath_ALUhw_BWISE_n72, B => n2987, S => 
                           n2269, Z => n8278);
   U19665 : MUX2_X1 port map( A => n8279, B => n8278, S => n2154, Z => n8281);
   U19666 : AOI22_X1 port map( A1 => n8322, A2 => n8281, B1 => n2258, B2 => 
                           n770, ZN => DataPath_ALUhw_MUXOUT_n69);
   U19667 : MUX2_X1 port map( A => n4132, B => n259, S => n1860, Z => n11488);
   U19668 : NAND4_X1 port map( A1 => n12883, A2 => n12884, A3 => n12885, A4 => 
                           n12886, ZN => n8345);
   U19669 : NAND4_X1 port map( A1 => n12879, A2 => n12880, A3 => n12881, A4 => 
                           n12882, ZN => n8346);
   U19670 : NAND4_X1 port map( A1 => n12843, A2 => n12844, A3 => n12845, A4 => 
                           n12846, ZN => n8343);
   U19671 : NAND4_X1 port map( A1 => n12839, A2 => n12840, A3 => n12841, A4 => 
                           n12842, ZN => n8344);
   U19672 : NAND4_X1 port map( A1 => n12803, A2 => n12804, A3 => n12805, A4 => 
                           n12806, ZN => n8341);
   U19673 : NAND4_X1 port map( A1 => n12799, A2 => n12800, A3 => n12801, A4 => 
                           n12802, ZN => n8342);
   U19674 : NAND4_X1 port map( A1 => n12763, A2 => n12764, A3 => n12765, A4 => 
                           n12766, ZN => n8339);
   U19675 : NAND4_X1 port map( A1 => n12759, A2 => n12760, A3 => n12761, A4 => 
                           n12762, ZN => n8340);
   U19676 : NAND4_X1 port map( A1 => n12723, A2 => n12724, A3 => n12725, A4 => 
                           n12726, ZN => n8337);
   U19677 : NAND4_X1 port map( A1 => n12719, A2 => n12720, A3 => n12721, A4 => 
                           n12722, ZN => n8338);
   U19678 : NAND4_X1 port map( A1 => n12683, A2 => n12684, A3 => n12685, A4 => 
                           n12686, ZN => n8335);
   U19679 : NAND4_X1 port map( A1 => n12679, A2 => n12680, A3 => n12681, A4 => 
                           n12682, ZN => n8336);
   U19680 : NAND4_X1 port map( A1 => n12643, A2 => n12644, A3 => n12645, A4 => 
                           n12646, ZN => n8333);
   U19681 : NAND4_X1 port map( A1 => n12639, A2 => n12640, A3 => n12641, A4 => 
                           n12642, ZN => n8334);
   U19682 : NAND4_X1 port map( A1 => n12603, A2 => n12604, A3 => n12605, A4 => 
                           n12606, ZN => n8389);
   U19683 : NAND4_X1 port map( A1 => n12599, A2 => n12600, A3 => n12601, A4 => 
                           n12602, ZN => n8390);
   U19684 : NAND4_X1 port map( A1 => n12563, A2 => n12564, A3 => n12565, A4 => 
                           n12566, ZN => n8387);
   U19685 : NAND4_X1 port map( A1 => n12559, A2 => n12560, A3 => n12561, A4 => 
                           n12562, ZN => n8388);
   U19686 : NAND4_X1 port map( A1 => n12523, A2 => n12524, A3 => n12525, A4 => 
                           n12526, ZN => n8331);
   U19687 : NAND4_X1 port map( A1 => n12519, A2 => n12520, A3 => n12521, A4 => 
                           n12522, ZN => n8332);
   U19688 : NAND4_X1 port map( A1 => n12483, A2 => n12484, A3 => n12485, A4 => 
                           n12486, ZN => n8385);
   U19689 : NAND4_X1 port map( A1 => n12479, A2 => n12480, A3 => n12481, A4 => 
                           n12482, ZN => n8386);
   U19690 : NAND4_X1 port map( A1 => n12443, A2 => n12444, A3 => n12445, A4 => 
                           n12446, ZN => n8383);
   U19691 : NAND4_X1 port map( A1 => n12439, A2 => n12440, A3 => n12441, A4 => 
                           n12442, ZN => n8384);
   U19692 : NAND4_X1 port map( A1 => n12403, A2 => n12404, A3 => n12405, A4 => 
                           n12406, ZN => n8381);
   U19693 : NAND4_X1 port map( A1 => n12399, A2 => n12400, A3 => n12401, A4 => 
                           n12402, ZN => n8382);
   U19694 : NAND4_X1 port map( A1 => n12363, A2 => n12364, A3 => n12365, A4 => 
                           n12366, ZN => n8379);
   U19695 : NAND4_X1 port map( A1 => n12359, A2 => n12360, A3 => n12361, A4 => 
                           n12362, ZN => n8380);
   U19696 : NAND4_X1 port map( A1 => n12323, A2 => n12324, A3 => n12325, A4 => 
                           n12326, ZN => n8377);
   U19697 : NAND4_X1 port map( A1 => n12319, A2 => n12320, A3 => n12321, A4 => 
                           n12322, ZN => n8378);
   U19698 : NAND4_X1 port map( A1 => n12283, A2 => n12284, A3 => n12285, A4 => 
                           n12286, ZN => n8375);
   U19699 : NAND4_X1 port map( A1 => n12279, A2 => n12280, A3 => n12281, A4 => 
                           n12282, ZN => n8376);
   U19700 : NAND4_X1 port map( A1 => n12243, A2 => n12244, A3 => n12245, A4 => 
                           n12246, ZN => n8373);
   U19701 : NAND4_X1 port map( A1 => n12239, A2 => n12240, A3 => n12241, A4 => 
                           n12242, ZN => n8374);
   U19702 : NAND4_X1 port map( A1 => n12203, A2 => n12204, A3 => n12205, A4 => 
                           n12206, ZN => n8371);
   U19703 : NAND4_X1 port map( A1 => n12199, A2 => n12200, A3 => n12201, A4 => 
                           n12202, ZN => n8372);
   U19704 : NAND4_X1 port map( A1 => n12163, A2 => n12164, A3 => n12165, A4 => 
                           n12166, ZN => n8369);
   U19705 : NAND4_X1 port map( A1 => n12159, A2 => n12160, A3 => n12161, A4 => 
                           n12162, ZN => n8370);
   U19706 : NAND4_X1 port map( A1 => n12123, A2 => n12124, A3 => n12125, A4 => 
                           n12126, ZN => n8367);
   U19707 : NAND4_X1 port map( A1 => n12119, A2 => n12120, A3 => n12121, A4 => 
                           n12122, ZN => n8368);
   U19708 : NAND4_X1 port map( A1 => n12083, A2 => n12084, A3 => n12085, A4 => 
                           n12086, ZN => n8329);
   U19709 : NAND4_X1 port map( A1 => n12079, A2 => n12080, A3 => n12081, A4 => 
                           n12082, ZN => n8330);
   U19710 : NAND4_X1 port map( A1 => n12043, A2 => n12044, A3 => n12045, A4 => 
                           n12046, ZN => n8365);
   U19711 : NAND4_X1 port map( A1 => n12039, A2 => n12040, A3 => n12041, A4 => 
                           n12042, ZN => n8366);
   U19712 : NAND4_X1 port map( A1 => n12003, A2 => n12004, A3 => n12005, A4 => 
                           n12006, ZN => n8363);
   U19713 : NAND4_X1 port map( A1 => n11999, A2 => n12000, A3 => n12001, A4 => 
                           n12002, ZN => n8364);
   U19714 : NAND4_X1 port map( A1 => n11963, A2 => n11964, A3 => n11965, A4 => 
                           n11966, ZN => n8361);
   U19715 : NAND4_X1 port map( A1 => n11959, A2 => n11960, A3 => n11961, A4 => 
                           n11962, ZN => n8362);
   U19716 : NAND4_X1 port map( A1 => n11923, A2 => n11924, A3 => n11925, A4 => 
                           n11926, ZN => n8359);
   U19717 : NAND4_X1 port map( A1 => n11919, A2 => n11920, A3 => n11921, A4 => 
                           n11922, ZN => n8360);
   U19718 : NAND4_X1 port map( A1 => n11883, A2 => n11884, A3 => n11885, A4 => 
                           n11886, ZN => n8357);
   U19719 : NAND4_X1 port map( A1 => n11879, A2 => n11880, A3 => n11881, A4 => 
                           n11882, ZN => n8358);
   U19720 : NAND4_X1 port map( A1 => n11843, A2 => n11844, A3 => n11845, A4 => 
                           n11846, ZN => n8355);
   U19721 : NAND4_X1 port map( A1 => n11839, A2 => n11840, A3 => n11841, A4 => 
                           n11842, ZN => n8356);
   U19722 : NAND4_X1 port map( A1 => n11803, A2 => n11804, A3 => n11805, A4 => 
                           n11806, ZN => n8353);
   U19723 : NAND4_X1 port map( A1 => n11799, A2 => n11800, A3 => n11801, A4 => 
                           n11802, ZN => n8354);
   U19724 : NAND4_X1 port map( A1 => n11763, A2 => n11764, A3 => n11765, A4 => 
                           n11766, ZN => n8351);
   U19725 : NAND4_X1 port map( A1 => n11759, A2 => n11760, A3 => n11761, A4 => 
                           n11762, ZN => n8352);
   U19726 : NAND4_X1 port map( A1 => n11723, A2 => n11724, A3 => n11725, A4 => 
                           n11726, ZN => n8349);
   U19727 : NAND4_X1 port map( A1 => n11719, A2 => n11720, A3 => n11721, A4 => 
                           n11722, ZN => n8350);
   U19728 : NAND4_X1 port map( A1 => n11683, A2 => n11684, A3 => n11685, A4 => 
                           n11686, ZN => n8347);
   U19729 : NAND4_X1 port map( A1 => n11679, A2 => n11680, A3 => n11681, A4 => 
                           n11682, ZN => n8348);
   U19730 : NAND4_X1 port map( A1 => n11643, A2 => n11644, A3 => n11645, A4 => 
                           n11646, ZN => n8327);
   U19731 : NAND4_X1 port map( A1 => n11639, A2 => n11640, A3 => n11641, A4 => 
                           n11642, ZN => n8328);
   U19732 : NAND4_X1 port map( A1 => n12875, A2 => n12876, A3 => n12877, A4 => 
                           n12878, ZN => n8409);
   U19733 : NAND4_X1 port map( A1 => n12871, A2 => n12872, A3 => n12873, A4 => 
                           n12874, ZN => n8410);
   U19734 : NAND4_X1 port map( A1 => n12835, A2 => n12836, A3 => n12837, A4 => 
                           n12838, ZN => n8407);
   U19735 : NAND4_X1 port map( A1 => n12831, A2 => n12832, A3 => n12833, A4 => 
                           n12834, ZN => n8408);
   U19736 : NAND4_X1 port map( A1 => n12795, A2 => n12796, A3 => n12797, A4 => 
                           n12798, ZN => n8405);
   U19737 : NAND4_X1 port map( A1 => n12791, A2 => n12792, A3 => n12793, A4 => 
                           n12794, ZN => n8406);
   U19738 : NAND4_X1 port map( A1 => n12755, A2 => n12756, A3 => n12757, A4 => 
                           n12758, ZN => n8403);
   U19739 : NAND4_X1 port map( A1 => n12751, A2 => n12752, A3 => n12753, A4 => 
                           n12754, ZN => n8404);
   U19740 : NAND4_X1 port map( A1 => n12715, A2 => n12716, A3 => n12717, A4 => 
                           n12718, ZN => n8401);
   U19741 : NAND4_X1 port map( A1 => n12711, A2 => n12712, A3 => n12713, A4 => 
                           n12714, ZN => n8402);
   U19742 : NAND4_X1 port map( A1 => n12675, A2 => n12676, A3 => n12677, A4 => 
                           n12678, ZN => n8399);
   U19743 : NAND4_X1 port map( A1 => n12671, A2 => n12672, A3 => n12673, A4 => 
                           n12674, ZN => n8400);
   U19744 : NAND4_X1 port map( A1 => n12635, A2 => n12636, A3 => n12637, A4 => 
                           n12638, ZN => n8397);
   U19745 : NAND4_X1 port map( A1 => n12631, A2 => n12632, A3 => n12633, A4 => 
                           n12634, ZN => n8398);
   U19746 : NAND4_X1 port map( A1 => n12595, A2 => n12596, A3 => n12597, A4 => 
                           n12598, ZN => n8453);
   U19747 : NAND4_X1 port map( A1 => n12591, A2 => n12592, A3 => n12593, A4 => 
                           n12594, ZN => n8454);
   U19748 : NAND4_X1 port map( A1 => n12555, A2 => n12556, A3 => n12557, A4 => 
                           n12558, ZN => n8451);
   U19749 : NAND4_X1 port map( A1 => n12551, A2 => n12552, A3 => n12553, A4 => 
                           n12554, ZN => n8452);
   U19750 : NAND4_X1 port map( A1 => n12515, A2 => n12516, A3 => n12517, A4 => 
                           n12518, ZN => n8395);
   U19751 : NAND4_X1 port map( A1 => n12511, A2 => n12512, A3 => n12513, A4 => 
                           n12514, ZN => n8396);
   U19752 : NAND4_X1 port map( A1 => n12475, A2 => n12476, A3 => n12477, A4 => 
                           n12478, ZN => n8449);
   U19753 : NAND4_X1 port map( A1 => n12471, A2 => n12472, A3 => n12473, A4 => 
                           n12474, ZN => n8450);
   U19754 : NAND4_X1 port map( A1 => n12435, A2 => n12436, A3 => n12437, A4 => 
                           n12438, ZN => n8447);
   U19755 : NAND4_X1 port map( A1 => n12431, A2 => n12432, A3 => n12433, A4 => 
                           n12434, ZN => n8448);
   U19756 : NAND4_X1 port map( A1 => n12395, A2 => n12396, A3 => n12397, A4 => 
                           n12398, ZN => n8445);
   U19757 : NAND4_X1 port map( A1 => n12391, A2 => n12392, A3 => n12393, A4 => 
                           n12394, ZN => n8446);
   U19758 : NAND4_X1 port map( A1 => n12355, A2 => n12356, A3 => n12357, A4 => 
                           n12358, ZN => n8443);
   U19759 : NAND4_X1 port map( A1 => n12351, A2 => n12352, A3 => n12353, A4 => 
                           n12354, ZN => n8444);
   U19760 : NAND4_X1 port map( A1 => n12315, A2 => n12316, A3 => n12317, A4 => 
                           n12318, ZN => n8441);
   U19761 : NAND4_X1 port map( A1 => n12311, A2 => n12312, A3 => n12313, A4 => 
                           n12314, ZN => n8442);
   U19762 : NAND4_X1 port map( A1 => n12275, A2 => n12276, A3 => n12277, A4 => 
                           n12278, ZN => n8439);
   U19763 : NAND4_X1 port map( A1 => n12271, A2 => n12272, A3 => n12273, A4 => 
                           n12274, ZN => n8440);
   U19764 : NAND4_X1 port map( A1 => n12235, A2 => n12236, A3 => n12237, A4 => 
                           n12238, ZN => n8437);
   U19765 : NAND4_X1 port map( A1 => n12231, A2 => n12232, A3 => n12233, A4 => 
                           n12234, ZN => n8438);
   U19766 : NAND4_X1 port map( A1 => n12195, A2 => n12196, A3 => n12197, A4 => 
                           n12198, ZN => n8435);
   U19767 : NAND4_X1 port map( A1 => n12191, A2 => n12192, A3 => n12193, A4 => 
                           n12194, ZN => n8436);
   U19768 : NAND4_X1 port map( A1 => n12155, A2 => n12156, A3 => n12157, A4 => 
                           n12158, ZN => n8433);
   U19769 : NAND4_X1 port map( A1 => n12151, A2 => n12152, A3 => n12153, A4 => 
                           n12154, ZN => n8434);
   U19770 : NAND4_X1 port map( A1 => n12115, A2 => n12116, A3 => n12117, A4 => 
                           n12118, ZN => n8431);
   U19771 : NAND4_X1 port map( A1 => n12111, A2 => n12112, A3 => n12113, A4 => 
                           n12114, ZN => n8432);
   U19772 : NAND4_X1 port map( A1 => n12075, A2 => n12076, A3 => n12077, A4 => 
                           n12078, ZN => n8393);
   U19773 : NAND4_X1 port map( A1 => n12071, A2 => n12072, A3 => n12073, A4 => 
                           n12074, ZN => n8394);
   U19774 : NAND4_X1 port map( A1 => n12035, A2 => n12036, A3 => n12037, A4 => 
                           n12038, ZN => n8429);
   U19775 : NAND4_X1 port map( A1 => n12031, A2 => n12032, A3 => n12033, A4 => 
                           n12034, ZN => n8430);
   U19776 : NAND4_X1 port map( A1 => n11995, A2 => n11996, A3 => n11997, A4 => 
                           n11998, ZN => n8427);
   U19777 : NAND4_X1 port map( A1 => n11991, A2 => n11992, A3 => n11993, A4 => 
                           n11994, ZN => n8428);
   U19778 : NAND4_X1 port map( A1 => n11955, A2 => n11956, A3 => n11957, A4 => 
                           n11958, ZN => n8425);
   U19779 : NAND4_X1 port map( A1 => n11951, A2 => n11952, A3 => n11953, A4 => 
                           n11954, ZN => n8426);
   U19780 : NAND4_X1 port map( A1 => n11915, A2 => n11916, A3 => n11917, A4 => 
                           n11918, ZN => n8423);
   U19781 : NAND4_X1 port map( A1 => n11911, A2 => n11912, A3 => n11913, A4 => 
                           n11914, ZN => n8424);
   U19782 : NAND4_X1 port map( A1 => n11875, A2 => n11876, A3 => n11877, A4 => 
                           n11878, ZN => n8421);
   U19783 : NAND4_X1 port map( A1 => n11871, A2 => n11872, A3 => n11873, A4 => 
                           n11874, ZN => n8422);
   U19784 : NAND4_X1 port map( A1 => n11835, A2 => n11836, A3 => n11837, A4 => 
                           n11838, ZN => n8419);
   U19785 : NAND4_X1 port map( A1 => n11831, A2 => n11832, A3 => n11833, A4 => 
                           n11834, ZN => n8420);
   U19786 : NAND4_X1 port map( A1 => n11795, A2 => n11796, A3 => n11797, A4 => 
                           n11798, ZN => n8417);
   U19787 : NAND4_X1 port map( A1 => n11791, A2 => n11792, A3 => n11793, A4 => 
                           n11794, ZN => n8418);
   U19788 : NAND4_X1 port map( A1 => n11755, A2 => n11756, A3 => n11757, A4 => 
                           n11758, ZN => n8415);
   U19789 : NAND4_X1 port map( A1 => n11751, A2 => n11752, A3 => n11753, A4 => 
                           n11754, ZN => n8416);
   U19790 : NAND4_X1 port map( A1 => n11715, A2 => n11716, A3 => n11717, A4 => 
                           n11718, ZN => n8413);
   U19791 : NAND4_X1 port map( A1 => n11711, A2 => n11712, A3 => n11713, A4 => 
                           n11714, ZN => n8414);
   U19792 : NAND4_X1 port map( A1 => n11675, A2 => n11676, A3 => n11677, A4 => 
                           n11678, ZN => n8411);
   U19793 : NAND4_X1 port map( A1 => n11671, A2 => n11672, A3 => n11673, A4 => 
                           n11674, ZN => n8412);
   U19794 : NAND4_X1 port map( A1 => n11635, A2 => n11636, A3 => n11637, A4 => 
                           n11638, ZN => n8391);
   U19795 : NAND4_X1 port map( A1 => n11631, A2 => n11632, A3 => n11633, A4 => 
                           n11634, ZN => n8392);
   U19796 : NAND4_X1 port map( A1 => n12867, A2 => n12868, A3 => n12869, A4 => 
                           n12870, ZN => n8473);
   U19797 : NAND4_X1 port map( A1 => n12863, A2 => n12864, A3 => n12865, A4 => 
                           n12866, ZN => n8474);
   U19798 : NAND4_X1 port map( A1 => n12827, A2 => n12828, A3 => n12829, A4 => 
                           n12830, ZN => n8471);
   U19799 : NAND4_X1 port map( A1 => n12823, A2 => n12824, A3 => n12825, A4 => 
                           n12826, ZN => n8472);
   U19800 : NAND4_X1 port map( A1 => n12787, A2 => n12788, A3 => n12789, A4 => 
                           n12790, ZN => n8469);
   U19801 : NAND4_X1 port map( A1 => n12783, A2 => n12784, A3 => n12785, A4 => 
                           n12786, ZN => n8470);
   U19802 : NAND4_X1 port map( A1 => n12747, A2 => n12748, A3 => n12749, A4 => 
                           n12750, ZN => n8467);
   U19803 : NAND4_X1 port map( A1 => n12743, A2 => n12744, A3 => n12745, A4 => 
                           n12746, ZN => n8468);
   U19804 : NAND4_X1 port map( A1 => n12707, A2 => n12708, A3 => n12709, A4 => 
                           n12710, ZN => n8465);
   U19805 : NAND4_X1 port map( A1 => n12703, A2 => n12704, A3 => n12705, A4 => 
                           n12706, ZN => n8466);
   U19806 : NAND4_X1 port map( A1 => n12667, A2 => n12668, A3 => n12669, A4 => 
                           n12670, ZN => n8463);
   U19807 : NAND4_X1 port map( A1 => n12663, A2 => n12664, A3 => n12665, A4 => 
                           n12666, ZN => n8464);
   U19808 : NAND4_X1 port map( A1 => n12627, A2 => n12628, A3 => n12629, A4 => 
                           n12630, ZN => n8461);
   U19809 : NAND4_X1 port map( A1 => n12623, A2 => n12624, A3 => n12625, A4 => 
                           n12626, ZN => n8462);
   U19810 : NAND4_X1 port map( A1 => n12587, A2 => n12588, A3 => n12589, A4 => 
                           n12590, ZN => n8517);
   U19811 : NAND4_X1 port map( A1 => n12583, A2 => n12584, A3 => n12585, A4 => 
                           n12586, ZN => n8518);
   U19812 : NAND4_X1 port map( A1 => n12547, A2 => n12548, A3 => n12549, A4 => 
                           n12550, ZN => n8515);
   U19813 : NAND4_X1 port map( A1 => n12543, A2 => n12544, A3 => n12545, A4 => 
                           n12546, ZN => n8516);
   U19814 : NAND4_X1 port map( A1 => n12507, A2 => n12508, A3 => n12509, A4 => 
                           n12510, ZN => n8459);
   U19815 : NAND4_X1 port map( A1 => n12503, A2 => n12504, A3 => n12505, A4 => 
                           n12506, ZN => n8460);
   U19816 : NAND4_X1 port map( A1 => n12467, A2 => n12468, A3 => n12469, A4 => 
                           n12470, ZN => n8513);
   U19817 : NAND4_X1 port map( A1 => n12463, A2 => n12464, A3 => n12465, A4 => 
                           n12466, ZN => n8514);
   U19818 : NAND4_X1 port map( A1 => n12427, A2 => n12428, A3 => n12429, A4 => 
                           n12430, ZN => n8511);
   U19819 : NAND4_X1 port map( A1 => n12423, A2 => n12424, A3 => n12425, A4 => 
                           n12426, ZN => n8512);
   U19820 : NAND4_X1 port map( A1 => n12387, A2 => n12388, A3 => n12389, A4 => 
                           n12390, ZN => n8509);
   U19821 : NAND4_X1 port map( A1 => n12383, A2 => n12384, A3 => n12385, A4 => 
                           n12386, ZN => n8510);
   U19822 : NAND4_X1 port map( A1 => n12347, A2 => n12348, A3 => n12349, A4 => 
                           n12350, ZN => n8507);
   U19823 : NAND4_X1 port map( A1 => n12343, A2 => n12344, A3 => n12345, A4 => 
                           n12346, ZN => n8508);
   U19824 : NAND4_X1 port map( A1 => n12307, A2 => n12308, A3 => n12309, A4 => 
                           n12310, ZN => n8505);
   U19825 : NAND4_X1 port map( A1 => n12303, A2 => n12304, A3 => n12305, A4 => 
                           n12306, ZN => n8506);
   U19826 : NAND4_X1 port map( A1 => n12267, A2 => n12268, A3 => n12269, A4 => 
                           n12270, ZN => n8503);
   U19827 : NAND4_X1 port map( A1 => n12263, A2 => n12264, A3 => n12265, A4 => 
                           n12266, ZN => n8504);
   U19828 : NAND4_X1 port map( A1 => n12227, A2 => n12228, A3 => n12229, A4 => 
                           n12230, ZN => n8501);
   U19829 : NAND4_X1 port map( A1 => n12223, A2 => n12224, A3 => n12225, A4 => 
                           n12226, ZN => n8502);
   U19830 : NAND4_X1 port map( A1 => n12187, A2 => n12188, A3 => n12189, A4 => 
                           n12190, ZN => n8499);
   U19831 : NAND4_X1 port map( A1 => n12183, A2 => n12184, A3 => n12185, A4 => 
                           n12186, ZN => n8500);
   U19832 : NAND4_X1 port map( A1 => n12147, A2 => n12148, A3 => n12149, A4 => 
                           n12150, ZN => n8497);
   U19833 : NAND4_X1 port map( A1 => n12143, A2 => n12144, A3 => n12145, A4 => 
                           n12146, ZN => n8498);
   U19834 : NAND4_X1 port map( A1 => n12107, A2 => n12108, A3 => n12109, A4 => 
                           n12110, ZN => n8495);
   U19835 : NAND4_X1 port map( A1 => n12103, A2 => n12104, A3 => n12105, A4 => 
                           n12106, ZN => n8496);
   U19836 : NAND4_X1 port map( A1 => n12067, A2 => n12068, A3 => n12069, A4 => 
                           n12070, ZN => n8457);
   U19837 : NAND4_X1 port map( A1 => n12063, A2 => n12064, A3 => n12065, A4 => 
                           n12066, ZN => n8458);
   U19838 : NAND4_X1 port map( A1 => n12027, A2 => n12028, A3 => n12029, A4 => 
                           n12030, ZN => n8493);
   U19839 : NAND4_X1 port map( A1 => n12023, A2 => n12024, A3 => n12025, A4 => 
                           n12026, ZN => n8494);
   U19840 : NAND4_X1 port map( A1 => n11987, A2 => n11988, A3 => n11989, A4 => 
                           n11990, ZN => n8491);
   U19841 : NAND4_X1 port map( A1 => n11983, A2 => n11984, A3 => n11985, A4 => 
                           n11986, ZN => n8492);
   U19842 : NAND4_X1 port map( A1 => n11947, A2 => n11948, A3 => n11949, A4 => 
                           n11950, ZN => n8489);
   U19843 : NAND4_X1 port map( A1 => n11943, A2 => n11944, A3 => n11945, A4 => 
                           n11946, ZN => n8490);
   U19844 : NAND4_X1 port map( A1 => n11907, A2 => n11908, A3 => n11909, A4 => 
                           n11910, ZN => n8487);
   U19845 : NAND4_X1 port map( A1 => n11903, A2 => n11904, A3 => n11905, A4 => 
                           n11906, ZN => n8488);
   U19846 : NAND4_X1 port map( A1 => n11867, A2 => n11868, A3 => n11869, A4 => 
                           n11870, ZN => n8485);
   U19847 : NAND4_X1 port map( A1 => n11863, A2 => n11864, A3 => n11865, A4 => 
                           n11866, ZN => n8486);
   U19848 : NAND4_X1 port map( A1 => n11827, A2 => n11828, A3 => n11829, A4 => 
                           n11830, ZN => n8483);
   U19849 : NAND4_X1 port map( A1 => n11823, A2 => n11824, A3 => n11825, A4 => 
                           n11826, ZN => n8484);
   U19850 : NAND4_X1 port map( A1 => n11787, A2 => n11788, A3 => n11789, A4 => 
                           n11790, ZN => n8481);
   U19851 : NAND4_X1 port map( A1 => n11783, A2 => n11784, A3 => n11785, A4 => 
                           n11786, ZN => n8482);
   U19852 : NAND4_X1 port map( A1 => n11747, A2 => n11748, A3 => n11749, A4 => 
                           n11750, ZN => n8479);
   U19853 : NAND4_X1 port map( A1 => n11743, A2 => n11744, A3 => n11745, A4 => 
                           n11746, ZN => n8480);
   U19854 : NAND4_X1 port map( A1 => n11707, A2 => n11708, A3 => n11709, A4 => 
                           n11710, ZN => n8477);
   U19855 : NAND4_X1 port map( A1 => n11703, A2 => n11704, A3 => n11705, A4 => 
                           n11706, ZN => n8478);
   U19856 : NAND4_X1 port map( A1 => n11667, A2 => n11668, A3 => n11669, A4 => 
                           n11670, ZN => n8475);
   U19857 : NAND4_X1 port map( A1 => n11663, A2 => n11664, A3 => n11665, A4 => 
                           n11666, ZN => n8476);
   U19858 : NAND4_X1 port map( A1 => n11627, A2 => n11628, A3 => n11629, A4 => 
                           n11630, ZN => n8455);
   U19859 : NAND4_X1 port map( A1 => n11623, A2 => n11624, A3 => n11625, A4 => 
                           n11626, ZN => n8456);
   U19860 : NAND4_X1 port map( A1 => n12859, A2 => n12860, A3 => n12861, A4 => 
                           n12862, ZN => n8537);
   U19861 : NAND4_X1 port map( A1 => n12855, A2 => n12856, A3 => n12857, A4 => 
                           n12858, ZN => n8538);
   U19862 : NAND4_X1 port map( A1 => n12819, A2 => n12820, A3 => n12821, A4 => 
                           n12822, ZN => n8535);
   U19863 : NAND4_X1 port map( A1 => n12815, A2 => n12816, A3 => n12817, A4 => 
                           n12818, ZN => n8536);
   U19864 : NAND4_X1 port map( A1 => n12779, A2 => n12780, A3 => n12781, A4 => 
                           n12782, ZN => n8533);
   U19865 : NAND4_X1 port map( A1 => n12775, A2 => n12776, A3 => n12777, A4 => 
                           n12778, ZN => n8534);
   U19866 : NAND4_X1 port map( A1 => n12739, A2 => n12740, A3 => n12741, A4 => 
                           n12742, ZN => n8531);
   U19867 : NAND4_X1 port map( A1 => n12735, A2 => n12736, A3 => n12737, A4 => 
                           n12738, ZN => n8532);
   U19868 : NAND4_X1 port map( A1 => n12699, A2 => n12700, A3 => n12701, A4 => 
                           n12702, ZN => n8529);
   U19869 : NAND4_X1 port map( A1 => n12695, A2 => n12696, A3 => n12697, A4 => 
                           n12698, ZN => n8530);
   U19870 : NAND4_X1 port map( A1 => n12659, A2 => n12660, A3 => n12661, A4 => 
                           n12662, ZN => n8527);
   U19871 : NAND4_X1 port map( A1 => n12655, A2 => n12656, A3 => n12657, A4 => 
                           n12658, ZN => n8528);
   U19872 : NAND4_X1 port map( A1 => n12619, A2 => n12620, A3 => n12621, A4 => 
                           n12622, ZN => n8525);
   U19873 : NAND4_X1 port map( A1 => n12615, A2 => n12616, A3 => n12617, A4 => 
                           n12618, ZN => n8526);
   U19874 : NAND4_X1 port map( A1 => n12579, A2 => n12580, A3 => n12581, A4 => 
                           n12582, ZN => n8581);
   U19875 : NAND4_X1 port map( A1 => n12575, A2 => n12576, A3 => n12577, A4 => 
                           n12578, ZN => n8582);
   U19876 : NAND4_X1 port map( A1 => n12539, A2 => n12540, A3 => n12541, A4 => 
                           n12542, ZN => n8579);
   U19877 : NAND4_X1 port map( A1 => n12535, A2 => n12536, A3 => n12537, A4 => 
                           n12538, ZN => n8580);
   U19878 : NAND4_X1 port map( A1 => n12499, A2 => n12500, A3 => n12501, A4 => 
                           n12502, ZN => n8523);
   U19879 : NAND4_X1 port map( A1 => n12495, A2 => n12496, A3 => n12497, A4 => 
                           n12498, ZN => n8524);
   U19880 : NAND4_X1 port map( A1 => n12459, A2 => n12460, A3 => n12461, A4 => 
                           n12462, ZN => n8577);
   U19881 : NAND4_X1 port map( A1 => n12455, A2 => n12456, A3 => n12457, A4 => 
                           n12458, ZN => n8578);
   U19882 : NAND4_X1 port map( A1 => n12419, A2 => n12420, A3 => n12421, A4 => 
                           n12422, ZN => n8575);
   U19883 : NAND4_X1 port map( A1 => n12415, A2 => n12416, A3 => n12417, A4 => 
                           n12418, ZN => n8576);
   U19884 : NAND4_X1 port map( A1 => n12379, A2 => n12380, A3 => n12381, A4 => 
                           n12382, ZN => n8573);
   U19885 : NAND4_X1 port map( A1 => n12375, A2 => n12376, A3 => n12377, A4 => 
                           n12378, ZN => n8574);
   U19886 : NAND4_X1 port map( A1 => n12339, A2 => n12340, A3 => n12341, A4 => 
                           n12342, ZN => n8571);
   U19887 : NAND4_X1 port map( A1 => n12335, A2 => n12336, A3 => n12337, A4 => 
                           n12338, ZN => n8572);
   U19888 : NAND4_X1 port map( A1 => n12299, A2 => n12300, A3 => n12301, A4 => 
                           n12302, ZN => n8569);
   U19889 : NAND4_X1 port map( A1 => n12295, A2 => n12296, A3 => n12297, A4 => 
                           n12298, ZN => n8570);
   U19890 : NAND4_X1 port map( A1 => n12259, A2 => n12260, A3 => n12261, A4 => 
                           n12262, ZN => n8567);
   U19891 : NAND4_X1 port map( A1 => n12255, A2 => n12256, A3 => n12257, A4 => 
                           n12258, ZN => n8568);
   U19892 : NAND4_X1 port map( A1 => n12219, A2 => n12220, A3 => n12221, A4 => 
                           n12222, ZN => n8565);
   U19893 : NAND4_X1 port map( A1 => n12215, A2 => n12216, A3 => n12217, A4 => 
                           n12218, ZN => n8566);
   U19894 : NAND4_X1 port map( A1 => n12179, A2 => n12180, A3 => n12181, A4 => 
                           n12182, ZN => n8563);
   U19895 : NAND4_X1 port map( A1 => n12175, A2 => n12176, A3 => n12177, A4 => 
                           n12178, ZN => n8564);
   U19896 : NAND4_X1 port map( A1 => n12139, A2 => n12140, A3 => n12141, A4 => 
                           n12142, ZN => n8561);
   U19897 : NAND4_X1 port map( A1 => n12135, A2 => n12136, A3 => n12137, A4 => 
                           n12138, ZN => n8562);
   U19898 : NAND4_X1 port map( A1 => n12099, A2 => n12100, A3 => n12101, A4 => 
                           n12102, ZN => n8559);
   U19899 : NAND4_X1 port map( A1 => n12095, A2 => n12096, A3 => n12097, A4 => 
                           n12098, ZN => n8560);
   U19900 : NAND4_X1 port map( A1 => n12059, A2 => n12060, A3 => n12061, A4 => 
                           n12062, ZN => n8521);
   U19901 : NAND4_X1 port map( A1 => n12055, A2 => n12056, A3 => n12057, A4 => 
                           n12058, ZN => n8522);
   U19902 : NAND4_X1 port map( A1 => n12019, A2 => n12020, A3 => n12021, A4 => 
                           n12022, ZN => n8557);
   U19903 : NAND4_X1 port map( A1 => n12015, A2 => n12016, A3 => n12017, A4 => 
                           n12018, ZN => n8558);
   U19904 : NAND4_X1 port map( A1 => n11979, A2 => n11980, A3 => n11981, A4 => 
                           n11982, ZN => n8555);
   U19905 : NAND4_X1 port map( A1 => n11975, A2 => n11976, A3 => n11977, A4 => 
                           n11978, ZN => n8556);
   U19906 : NAND4_X1 port map( A1 => n11939, A2 => n11940, A3 => n11941, A4 => 
                           n11942, ZN => n8553);
   U19907 : NAND4_X1 port map( A1 => n11935, A2 => n11936, A3 => n11937, A4 => 
                           n11938, ZN => n8554);
   U19908 : NAND4_X1 port map( A1 => n11899, A2 => n11900, A3 => n11901, A4 => 
                           n11902, ZN => n8551);
   U19909 : NAND4_X1 port map( A1 => n11895, A2 => n11896, A3 => n11897, A4 => 
                           n11898, ZN => n8552);
   U19910 : NAND4_X1 port map( A1 => n11859, A2 => n11860, A3 => n11861, A4 => 
                           n11862, ZN => n8549);
   U19911 : NAND4_X1 port map( A1 => n11855, A2 => n11856, A3 => n11857, A4 => 
                           n11858, ZN => n8550);
   U19912 : NAND4_X1 port map( A1 => n11819, A2 => n11820, A3 => n11821, A4 => 
                           n11822, ZN => n8547);
   U19913 : NAND4_X1 port map( A1 => n11815, A2 => n11816, A3 => n11817, A4 => 
                           n11818, ZN => n8548);
   U19914 : NAND4_X1 port map( A1 => n11779, A2 => n11780, A3 => n11781, A4 => 
                           n11782, ZN => n8545);
   U19915 : NAND4_X1 port map( A1 => n11775, A2 => n11776, A3 => n11777, A4 => 
                           n11778, ZN => n8546);
   U19916 : NAND4_X1 port map( A1 => n11739, A2 => n11740, A3 => n11741, A4 => 
                           n11742, ZN => n8543);
   U19917 : NAND4_X1 port map( A1 => n11735, A2 => n11736, A3 => n11737, A4 => 
                           n11738, ZN => n8544);
   U19918 : NAND4_X1 port map( A1 => n11699, A2 => n11700, A3 => n11701, A4 => 
                           n11702, ZN => n8541);
   U19919 : NAND4_X1 port map( A1 => n11695, A2 => n11696, A3 => n11697, A4 => 
                           n11698, ZN => n8542);
   U19920 : NAND4_X1 port map( A1 => n11659, A2 => n11660, A3 => n11661, A4 => 
                           n11662, ZN => n8539);
   U19921 : NAND4_X1 port map( A1 => n11655, A2 => n11656, A3 => n11657, A4 => 
                           n11658, ZN => n8540);
   U19922 : NAND4_X1 port map( A1 => n11619, A2 => n11620, A3 => n11621, A4 => 
                           n11622, ZN => n8519);
   U19923 : NAND4_X1 port map( A1 => n11615, A2 => n11616, A3 => n11617, A4 => 
                           n11618, ZN => n8520);
   U19924 : NAND4_X1 port map( A1 => n12852, A2 => n12853, A3 => n12854, A4 => 
                           n12887, ZN => n8601);
   U19925 : NAND4_X1 port map( A1 => n12848, A2 => n12849, A3 => n12850, A4 => 
                           n12851, ZN => n8602);
   U19926 : NAND4_X1 port map( A1 => n12812, A2 => n12813, A3 => n12814, A4 => 
                           n12847, ZN => n8599);
   U19927 : NAND4_X1 port map( A1 => n12808, A2 => n12809, A3 => n12810, A4 => 
                           n12811, ZN => n8600);
   U19928 : NAND4_X1 port map( A1 => n12772, A2 => n12773, A3 => n12774, A4 => 
                           n12807, ZN => n8597);
   U19929 : NAND4_X1 port map( A1 => n12768, A2 => n12769, A3 => n12770, A4 => 
                           n12771, ZN => n8598);
   U19930 : NAND4_X1 port map( A1 => n12732, A2 => n12733, A3 => n12734, A4 => 
                           n12767, ZN => n8595);
   U19931 : NAND4_X1 port map( A1 => n12728, A2 => n12729, A3 => n12730, A4 => 
                           n12731, ZN => n8596);
   U19932 : NAND4_X1 port map( A1 => n12692, A2 => n12693, A3 => n12694, A4 => 
                           n12727, ZN => n8593);
   U19933 : NAND4_X1 port map( A1 => n12688, A2 => n12689, A3 => n12690, A4 => 
                           n12691, ZN => n8594);
   U19934 : NAND4_X1 port map( A1 => n12652, A2 => n12653, A3 => n12654, A4 => 
                           n12687, ZN => n8591);
   U19935 : NAND4_X1 port map( A1 => n12648, A2 => n12649, A3 => n12650, A4 => 
                           n12651, ZN => n8592);
   U19936 : NAND4_X1 port map( A1 => n12612, A2 => n12613, A3 => n12614, A4 => 
                           n12647, ZN => n8589);
   U19937 : NAND4_X1 port map( A1 => n12608, A2 => n12609, A3 => n12610, A4 => 
                           n12611, ZN => n8590);
   U19938 : NAND4_X1 port map( A1 => n12572, A2 => n12573, A3 => n12574, A4 => 
                           n12607, ZN => n8645);
   U19939 : NAND4_X1 port map( A1 => n12568, A2 => n12569, A3 => n12570, A4 => 
                           n12571, ZN => n8646);
   U19940 : NAND4_X1 port map( A1 => n12532, A2 => n12533, A3 => n12534, A4 => 
                           n12567, ZN => n8643);
   U19941 : NAND4_X1 port map( A1 => n12528, A2 => n12529, A3 => n12530, A4 => 
                           n12531, ZN => n8644);
   U19942 : NAND4_X1 port map( A1 => n12492, A2 => n12493, A3 => n12494, A4 => 
                           n12527, ZN => n8587);
   U19943 : NAND4_X1 port map( A1 => n12488, A2 => n12489, A3 => n12490, A4 => 
                           n12491, ZN => n8588);
   U19944 : NAND4_X1 port map( A1 => n12452, A2 => n12453, A3 => n12454, A4 => 
                           n12487, ZN => n8641);
   U19945 : NAND4_X1 port map( A1 => n12448, A2 => n12449, A3 => n12450, A4 => 
                           n12451, ZN => n8642);
   U19946 : NAND4_X1 port map( A1 => n12412, A2 => n12413, A3 => n12414, A4 => 
                           n12447, ZN => n8639);
   U19947 : NAND4_X1 port map( A1 => n12408, A2 => n12409, A3 => n12410, A4 => 
                           n12411, ZN => n8640);
   U19948 : NAND4_X1 port map( A1 => n12372, A2 => n12373, A3 => n12374, A4 => 
                           n12407, ZN => n8637);
   U19949 : NAND4_X1 port map( A1 => n12368, A2 => n12369, A3 => n12370, A4 => 
                           n12371, ZN => n8638);
   U19950 : NAND4_X1 port map( A1 => n12332, A2 => n12333, A3 => n12334, A4 => 
                           n12367, ZN => n8635);
   U19951 : NAND4_X1 port map( A1 => n12328, A2 => n12329, A3 => n12330, A4 => 
                           n12331, ZN => n8636);
   U19952 : NAND4_X1 port map( A1 => n12292, A2 => n12293, A3 => n12294, A4 => 
                           n12327, ZN => n8633);
   U19953 : NAND4_X1 port map( A1 => n12288, A2 => n12289, A3 => n12290, A4 => 
                           n12291, ZN => n8634);
   U19954 : NAND4_X1 port map( A1 => n12252, A2 => n12253, A3 => n12254, A4 => 
                           n12287, ZN => n8631);
   U19955 : NAND4_X1 port map( A1 => n12248, A2 => n12249, A3 => n12250, A4 => 
                           n12251, ZN => n8632);
   U19956 : NAND4_X1 port map( A1 => n12212, A2 => n12213, A3 => n12214, A4 => 
                           n12247, ZN => n8629);
   U19957 : NAND4_X1 port map( A1 => n12208, A2 => n12209, A3 => n12210, A4 => 
                           n12211, ZN => n8630);
   U19958 : NAND4_X1 port map( A1 => n12172, A2 => n12173, A3 => n12174, A4 => 
                           n12207, ZN => n8627);
   U19959 : NAND4_X1 port map( A1 => n12168, A2 => n12169, A3 => n12170, A4 => 
                           n12171, ZN => n8628);
   U19960 : NAND4_X1 port map( A1 => n12132, A2 => n12133, A3 => n12134, A4 => 
                           n12167, ZN => n8625);
   U19961 : NAND4_X1 port map( A1 => n12128, A2 => n12129, A3 => n12130, A4 => 
                           n12131, ZN => n8626);
   U19962 : NAND4_X1 port map( A1 => n12092, A2 => n12093, A3 => n12094, A4 => 
                           n12127, ZN => n8623);
   U19963 : NAND4_X1 port map( A1 => n12088, A2 => n12089, A3 => n12090, A4 => 
                           n12091, ZN => n8624);
   U19964 : NAND4_X1 port map( A1 => n12052, A2 => n12053, A3 => n12054, A4 => 
                           n12087, ZN => n8585);
   U19965 : NAND4_X1 port map( A1 => n12048, A2 => n12049, A3 => n12050, A4 => 
                           n12051, ZN => n8586);
   U19966 : NAND4_X1 port map( A1 => n12012, A2 => n12013, A3 => n12014, A4 => 
                           n12047, ZN => n8621);
   U19967 : NAND4_X1 port map( A1 => n12008, A2 => n12009, A3 => n12010, A4 => 
                           n12011, ZN => n8622);
   U19968 : NAND4_X1 port map( A1 => n11972, A2 => n11973, A3 => n11974, A4 => 
                           n12007, ZN => n8619);
   U19969 : NAND4_X1 port map( A1 => n11968, A2 => n11969, A3 => n11970, A4 => 
                           n11971, ZN => n8620);
   U19970 : NAND4_X1 port map( A1 => n11932, A2 => n11933, A3 => n11934, A4 => 
                           n11967, ZN => n8617);
   U19971 : NAND4_X1 port map( A1 => n11928, A2 => n11929, A3 => n11930, A4 => 
                           n11931, ZN => n8618);
   U19972 : NAND4_X1 port map( A1 => n11892, A2 => n11893, A3 => n11894, A4 => 
                           n11927, ZN => n8615);
   U19973 : NAND4_X1 port map( A1 => n11888, A2 => n11889, A3 => n11890, A4 => 
                           n11891, ZN => n8616);
   U19974 : NAND4_X1 port map( A1 => n11852, A2 => n11853, A3 => n11854, A4 => 
                           n11887, ZN => n8613);
   U19975 : NAND4_X1 port map( A1 => n11848, A2 => n11849, A3 => n11850, A4 => 
                           n11851, ZN => n8614);
   U19976 : NAND4_X1 port map( A1 => n11812, A2 => n11813, A3 => n11814, A4 => 
                           n11847, ZN => n8611);
   U19977 : NAND4_X1 port map( A1 => n11808, A2 => n11809, A3 => n11810, A4 => 
                           n11811, ZN => n8612);
   U19978 : NAND4_X1 port map( A1 => n11772, A2 => n11773, A3 => n11774, A4 => 
                           n11807, ZN => n8609);
   U19979 : NAND4_X1 port map( A1 => n11768, A2 => n11769, A3 => n11770, A4 => 
                           n11771, ZN => n8610);
   U19980 : NAND4_X1 port map( A1 => n11732, A2 => n11733, A3 => n11734, A4 => 
                           n11767, ZN => n8607);
   U19981 : NAND4_X1 port map( A1 => n11728, A2 => n11729, A3 => n11730, A4 => 
                           n11731, ZN => n8608);
   U19982 : NAND4_X1 port map( A1 => n11692, A2 => n11693, A3 => n11694, A4 => 
                           n11727, ZN => n8605);
   U19983 : NAND4_X1 port map( A1 => n11688, A2 => n11689, A3 => n11690, A4 => 
                           n11691, ZN => n8606);
   U19984 : NAND4_X1 port map( A1 => n11652, A2 => n11653, A3 => n11654, A4 => 
                           n11687, ZN => n8603);
   U19985 : NAND4_X1 port map( A1 => n11648, A2 => n11649, A3 => n11650, A4 => 
                           n11651, ZN => n8604);
   U19986 : NAND4_X1 port map( A1 => n11612, A2 => n11613, A3 => n11614, A4 => 
                           n11647, ZN => n8583);
   U19987 : NAND4_X1 port map( A1 => n11608, A2 => n11609, A3 => n11610, A4 => 
                           n11611, ZN => n8584);
   RS2_4_port <= '0';
   DataPath_REG_IN1_Q_reg_8_inst : DFF_X1 port map( D => n2051, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_8_port, QN => n328);
   U146 : NAND2_X1 port map( A1 => n5524, A2 => n1508, ZN => n17146);
   U147 : OAI221_X4 port map( B1 => n5841, B2 => n5840, C1 => n5839, C2 => 
                           n6776, A => n5838, ZN => n17152);
   U149 : OR2_X1 port map( A1 => n6392, A2 => n17186, ZN => n17148);
   U150 : NAND2_X1 port map( A1 => n17148, A2 => n6340, ZN => n6372);
   U151 : AND2_X2 port map( A1 => n1404, A2 => n1405, ZN => n916);
   U152 : BUF_X1 port map( A => n5148, Z => n828);
   U153 : CLKBUF_X1 port map( A => n4580, Z => n17149);
   U154 : CLKBUF_X1 port map( A => n6103, Z => n17150);
   U156 : MUX2_X1 port map( A => n5607, B => n5606, S => n2244, Z => n1058);
   U157 : OR2_X2 port map( A1 => n4481, A2 => n4468, ZN => n4477);
   U158 : NAND2_X1 port map( A1 => n17216, A2 => n1483, ZN => n17153);
   U159 : XNOR2_X1 port map( A => n4695, B => n4690, ZN => n4698);
   U160 : CLKBUF_X1 port map( A => CU_I_n108, Z => n547);
   U161 : BUF_X1 port map( A => n6833, Z => n579);
   U162 : CLKBUF_X1 port map( A => n5291, Z => n639);
   U163 : XNOR2_X1 port map( A => n6296, B => n6202, ZN => n17154);
   U164 : XNOR2_X1 port map( A => n708, B => n6555, ZN => n17155);
   U166 : MUX2_X1 port map( A => n1666, B => n1665, S => n4436, Z => n1664);
   U167 : MUX2_X1 port map( A => n7017, B => n7018, S => n4436, Z => n17156);
   U168 : MUX2_X1 port map( A => n7017, B => n7018, S => n4436, Z => n7477);
   U169 : AND2_X1 port map( A1 => n644, A2 => n645, ZN => n17157);
   U170 : AND2_X1 port map( A1 => n5798, A2 => n5799, ZN => n5555);
   U171 : AND2_X1 port map( A1 => n4826, A2 => n4827, ZN => n1156);
   U172 : MUX2_X1 port map( A => n6239, B => n6240, S => n6839, Z => n1317);
   U173 : INV_X1 port map( A => n1058, ZN => n17158);
   U174 : MUX2_X2 port map( A => n5607, B => n5606, S => n2244, Z => n5879);
   U175 : CLKBUF_X1 port map( A => n1002, Z => n1237);
   U177 : OR2_X1 port map( A1 => n915, A2 => n8227, ZN => n17159);
   U184 : NAND2_X1 port map( A1 => n17159, A2 => n6207, ZN => n6329);
   U198 : INV_X1 port map( A => n2259, ZN => n17161);
   U217 : INV_X2 port map( A => n2263, ZN => n2259);
   U242 : CLKBUF_X1 port map( A => n6514, Z => n631);
   U251 : NAND2_X1 port map( A1 => n465, A2 => n466, ZN => n17162);
   U261 : MUX2_X1 port map( A => n6260, B => n6261, S => n859, Z => n1416);
   U269 : MUX2_X1 port map( A => n5918, B => n5917, S => n2268, Z => n17163);
   U276 : MUX2_X1 port map( A => n5918, B => n5917, S => n2268, Z => n6010);
   U315 : MUX2_X1 port map( A => n6675, B => n6676, S => n6594, Z => n1576);
   U333 : MUX2_X2 port map( A => n1719, B => n1720, S => n2265, Z => n17164);
   U336 : MUX2_X1 port map( A => n6257, B => n6256, S => n8229, Z => n855);
   U443 : CLKBUF_X1 port map( A => n4561, Z => n17165);
   U495 : INV_X1 port map( A => n6473, ZN => n17166);
   U566 : INV_X1 port map( A => n913, ZN => n17167);
   U730 : MUX2_X2 port map( A => n5901, B => n5902, S => n1211, Z => n17168);
   U733 : MUX2_X1 port map( A => n5901, B => n5902, S => n1211, Z => n6118);
   U879 : MUX2_X1 port map( A => n2174, B => n2173, S => n529, Z => n2172);
   U947 : CLKBUF_X1 port map( A => n8142, Z => n17169);
   U965 : AND2_X1 port map( A1 => n17249, A2 => n6176, ZN => n17170);
   U985 : AND2_X1 port map( A1 => n6175, A2 => n6176, ZN => n1775);
   U992 : NOR2_X1 port map( A1 => n6397, A2 => n6396, ZN => n17171);
   U996 : AND2_X1 port map( A1 => n644, A2 => n645, ZN => n813);
   U1082 : BUF_X1 port map( A => n6178, Z => n1481);
   U1092 : CLKBUF_X1 port map( A => n1131, Z => n17172);
   U1117 : INV_X1 port map( A => n1935, ZN => n2214);
   U1169 : AOI22_X1 port map( A1 => n4607, A2 => n1368, B1 => n4663, B2 => 
                           n17242, ZN => n17173);
   U1175 : NAND2_X2 port map( A1 => n4535, A2 => n4534, ZN => n4797);
   U1197 : AND2_X1 port map( A1 => n490, A2 => n217, ZN => n17174);
   U1209 : CLKBUF_X1 port map( A => n2149, Z => n17175);
   U1274 : MUX2_X2 port map( A => n6257, B => n6256, S => n8229, Z => n6397);
   U1283 : MUX2_X2 port map( A => n6117, B => n6116, S => n2266, Z => n1178);
   U1310 : AND3_X1 port map( A1 => n17177, A2 => n17178, A3 => n17176, ZN => 
                           n6058);
   U1340 : INV_X32 port map( A => n349, ZN => n17176);
   U1401 : NAND3_X1 port map( A1 => n6056, A2 => n851, A3 => n6055, ZN => 
                           n17177);
   U1452 : NAND2_X1 port map( A1 => n1131, A2 => n6070, ZN => n17178);
   U1469 : XNOR2_X1 port map( A => n17162, B => n6019, ZN => n1505);
   U1512 : CLKBUF_X1 port map( A => n17175, Z => n17179);
   U1526 : OAI211_X1 port map( C1 => n1064, C2 => n5072, A => n923, B => n5073,
                           ZN => n17180);
   U1599 : MUX2_X2 port map( A => n6394, B => n6395, S => n529, Z => n850);
   U1610 : MUX2_X2 port map( A => n6408, B => n6409, S => n754, Z => n1120);
   U1714 : OAI21_X1 port map( B1 => n6039, B2 => n6032, A => n5996, ZN => 
                           n17182);
   U1729 : MUX2_X1 port map( A => n5740, B => n5739, S => n2243, Z => n17183);
   U1745 : MUX2_X1 port map( A => n5740, B => n5739, S => n2243, Z => n5915);
   U1828 : INV_X1 port map( A => n5272, ZN => n17184);
   U1836 : OAI33_X1 port map( A1 => n449, A2 => n646, A3 => n472, B1 => n4810, 
                           B2 => n4803, B3 => n818, ZN => n17185);
   U1977 : MUX2_X1 port map( A => n6247, B => n6248, S => n859, Z => n6378);
   U2174 : INV_X1 port map( A => n8198, ZN => n17187);
   U2217 : AND2_X2 port map( A1 => n5968, A2 => n1648, ZN => n1607);
   U2225 : INV_X1 port map( A => n916, ZN => n17188);
   U2257 : CLKBUF_X1 port map( A => n237, Z => n17189);
   U2271 : CLKBUF_X1 port map( A => n766, Z => n17190);
   U2686 : NAND2_X1 port map( A1 => n496, A2 => n497, ZN => n17191);
   U2860 : AND2_X2 port map( A1 => n5338, A2 => n5337, ZN => n1780);
   U3807 : AND2_X1 port map( A1 => n6226, A2 => n1622, ZN => n17192);
   U16918 : AND2_X1 port map( A1 => n6226, A2 => n1622, ZN => n570);
   U16921 : MUX2_X1 port map( A => n4898, B => n4897, S => n2251, Z => n8180);
   U17159 : INV_X1 port map( A => n2136, ZN => n17193);
   U17577 : CLKBUF_X3 port map( A => n6858, Z => n2136);
   U17925 : INV_X1 port map( A => n2154, ZN => n17194);
   U18118 : BUF_X1 port map( A => n8091, Z => n2131);
   U18127 : CLKBUF_X1 port map( A => n7688, Z => n17195);
   U18194 : NAND2_X1 port map( A1 => n17196, A2 => n7069, ZN => n7578);
   U18221 : AND2_X1 port map( A1 => n963, A2 => n964, ZN => n17196);
   U19989 : INV_X1 port map( A => n8151, ZN => n17197);
   IRAM_ADDRESS_31_port <= '0';
   IRAM_ADDRESS_30_port <= '0';
   IRAM_ADDRESS_29_port <= '0';
   IRAM_ADDRESS_28_port <= '0';
   IRAM_ADDRESS_27_port <= '0';
   IRAM_ADDRESS_26_port <= '0';
   IRAM_ADDRESS_25_port <= '0';
   IRAM_ADDRESS_24_port <= '0';
   IRAM_ADDRESS_23_port <= '0';
   IRAM_ADDRESS_22_port <= '0';
   IRAM_ADDRESS_21_port <= '0';
   IRAM_ADDRESS_20_port <= '0';
   IRAM_ADDRESS_19_port <= '0';
   IRAM_ADDRESS_18_port <= '0';
   IRAM_ADDRESS_17_port <= '0';
   IRAM_ADDRESS_16_port <= '0';
   IRAM_ADDRESS_15_port <= '0';
   IRAM_ADDRESS_14_port <= '0';
   IRAM_ADDRESS_13_port <= '0';
   IRAM_ADDRESS_12_port <= '0';
   IRAM_ADDRESS_11_port <= '0';
   IRAM_ADDRESS_10_port <= '0';
   IRAM_ADDRESS_9_port <= '0';
   IRAM_ADDRESS_8_port <= '0';
   IRAM_ADDRESS_7_port <= '0';
   IRAM_ADDRESS_6_port <= '0';
   IRAM_ADDRESS_5_port <= '0';
   IRAM_ADDRESS_4_port <= '0';
   IRAM_ADDRESS_3_port <= '0';
   IRAM_ADDRESS_2_port <= '0';
   IRAM_ADDRESS_1_port <= '0';
   IRAM_ADDRESS_0_port <= '0';
   DataPath_REG_ALU_OUT_Q_reg_22_inst : DFF_X1 port map( D => n8669, CK => CLK,
                           Q => DRAM_ADDRESS_22_port, QN => n7809);
   DataPath_REG_ALU_OUT_Q_reg_23_inst : DFF_X1 port map( D => n8668, CK => CLK,
                           Q => DRAM_ADDRESS_23_port, QN => n7777);
   DataPath_REG_ALU_OUT_Q_reg_24_inst : DFF_X1 port map( D => n8667, CK => CLK,
                           Q => DRAM_ADDRESS_24_port, QN => n7744);
   DataPath_REG_ALU_OUT_Q_reg_25_inst : DFF_X1 port map( D => n8666, CK => CLK,
                           Q => DRAM_ADDRESS_25_port, QN => n7718);
   DataPath_REG_ALU_OUT_Q_reg_26_inst : DFF_X1 port map( D => n8665, CK => CLK,
                           Q => DRAM_ADDRESS_26_port, QN => n7685);
   DataPath_REG_ALU_OUT_Q_reg_27_inst : DFF_X1 port map( D => n8664, CK => CLK,
                           Q => DRAM_ADDRESS_27_port, QN => n7653);
   DataPath_REG_ALU_OUT_Q_reg_28_inst : DFF_X1 port map( D => n8663, CK => CLK,
                           Q => DRAM_ADDRESS_28_port, QN => n7615);
   DataPath_REG_IN1_Q_reg_5_inst : DFF_X1 port map( D => n2054, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN1_5_port, QN => n_3780);
   DataPath_REG_B_Q_reg_3_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_3_port, QN => n_3781);
   DataPath_REG_ALU_OUT_Q_reg_30_inst : DFF_X2 port map( D => n8661, CK => CLK,
                           Q => DRAM_ADDRESS_30_port, QN => n_3782);
   DataPath_REG_ALU_OUT_Q_reg_29_inst : DFF_X2 port map( D => n8662, CK => CLK,
                           Q => DRAM_ADDRESS_29_port, QN => n7586);
   U148 : MUX2_X2 port map( A => n6102, B => n6101, S => n2266, Z => n1003);
   U155 : MUX2_X1 port map( A => n6101, B => n6102, S => n17198, Z => n6262);
   U165 : INV_X32 port map( A => n2266, ZN => n17198);
   U176 : MUX2_X2 port map( A => n6116, B => n6117, S => n750, Z => n6288);
   U189 : OR2_X1 port map( A1 => n6734, A2 => n6733, ZN => n17199);
   U202 : NAND2_X1 port map( A1 => n17199, A2 => n6732, ZN => n6735);
   U211 : OR2_X1 port map( A1 => n4974, A2 => n4976, ZN => n17200);
   U223 : NAND2_X1 port map( A1 => n17200, A2 => n4927, ZN => n5014);
   U244 : NAND2_X1 port map( A1 => n17201, A2 => n17202, ZN => n17203);
   U250 : NAND2_X1 port map( A1 => n17203, A2 => n5768, ZN => n6732);
   U300 : INV_X1 port map( A => n5770, ZN => n17201);
   U301 : INV_X1 port map( A => n462, ZN => n17202);
   U302 : XNOR2_X1 port map( A => n7375, B => n7374, ZN => n17204);
   U305 : OR2_X1 port map( A1 => n4926, A2 => n5031, ZN => n17205);
   U306 : OR2_X1 port map( A1 => n5038, A2 => n5037, ZN => n17206);
   U344 : NAND3_X1 port map( A1 => n17205, A2 => n17206, A3 => n4925, ZN => 
                           n5021);
   U496 : OR2_X1 port map( A1 => n6883, A2 => n6882, ZN => n17207);
   U560 : NAND2_X1 port map( A1 => n17207, A2 => n6881, ZN => n7313);
   U600 : MUX2_X2 port map( A => n6729, B => n6728, S => n2250, Z => n6882);
   U622 : AND2_X1 port map( A1 => n6175, A2 => n6003, ZN => n17208);
   U636 : AND2_X1 port map( A1 => n6175, A2 => n6003, ZN => n1772);
   U656 : MUX2_X1 port map( A => n5891, B => n5890, S => n2268, Z => n6112);
   U668 : MUX2_X1 port map( A => n1349, B => n1348, S => n7712, Z => n756);
   U683 : CLKBUF_X1 port map( A => n6498, Z => n1475);
   U725 : BUF_X1 port map( A => n756, Z => n17209);
   U770 : MUX2_X1 port map( A => n5677, B => n5678, S => n1351, Z => n1352);
   U798 : MUX2_X1 port map( A => n2171, B => n2170, S => n6776, Z => n2169);
   U841 : NAND2_X1 port map( A1 => n6558, A2 => n6557, ZN => n17210);
   U846 : MUX2_X2 port map( A => n5636, B => n5635, S => n2244, Z => n620);
   U848 : INV_X1 port map( A => n17248, ZN => n17211);
   U855 : INV_X1 port map( A => n4636, ZN => n17212);
   U857 : AND2_X2 port map( A1 => n5880, A2 => n5881, ZN => n5883);
   U859 : XOR2_X1 port map( A => n1069, B => n6634, Z => n17213);
   U860 : MUX2_X2 port map( A => n6533, B => n6532, S => n1702, Z => n1580);
   U861 : MUX2_X2 port map( A => n5421, B => n5420, S => n2245, Z => n5657);
   U876 : MUX2_X2 port map( A => n5064, B => n5063, S => n2248, Z => n17214);
   U883 : MUX2_X1 port map( A => n5064, B => n5063, S => n2248, Z => n5397);
   U919 : NAND2_X1 port map( A1 => n6104, A2 => n1515, ZN => n17215);
   U1050 : OR2_X2 port map( A1 => n698, A2 => n5919, ZN => n690);
   U1085 : MUX2_X2 port map( A => n5947, B => n5946, S => n2267, Z => n5999);
   U1099 : OAI21_X1 port map( B1 => n1212, B2 => n5868, A => n5866, ZN => 
                           n17216);
   U1126 : CLKBUF_X1 port map( A => n4655, Z => n17217);
   U1134 : CLKBUF_X1 port map( A => n4557, Z => n835);
   U1136 : MUX2_X2 port map( A => n5947, B => n5946, S => n1706, Z => n776);
   U1141 : OAI33_X1 port map( A1 => n6912, A2 => n6911, A3 => n7365, B1 => 
                           n6910, B2 => n6909, B3 => n2244, ZN => n17218);
   U1195 : OR3_X1 port map( A1 => n6913, A2 => n447, A3 => n446, ZN => n17219);
   U1203 : INV_X1 port map( A => n5497, ZN => n17220);
   U1222 : CLKBUF_X1 port map( A => n1676, Z => n17221);
   U1263 : CLKBUF_X1 port map( A => n1469, Z => n17222);
   U1370 : CLKBUF_X1 port map( A => n1030, Z => n17223);
   U1371 : INV_X1 port map( A => n996, ZN => n17224);
   U1393 : MUX2_X2 port map( A => n6517, B => n6518, S => n6369, Z => n996);
   U1404 : BUF_X1 port map( A => n1729, Z => n565);
   U1409 : BUF_X1 port map( A => n727, Z => n17225);
   U1422 : OAI33_X1 port map( A1 => n4631, A2 => n2264, A3 => n4630, B1 => 
                           n4631, B2 => n2261, B3 => n450, ZN => n17226);
   U1509 : MUX2_X2 port map( A => n5885, B => n5886, S => n1211, Z => n6103);
   U1519 : OAI211_X1 port map( C1 => n5544, C2 => n5546, A => n5517, B => n5641
                           , ZN => n17227);
   U1558 : CLKBUF_X1 port map( A => n4639, Z => n17228);
   U1572 : XNOR2_X1 port map( A => n5359, B => n17229, ZN => n5362);
   U1606 : AND3_X1 port map( A1 => n888, A2 => n5207, A3 => n889, ZN => n17229)
                           ;
   U1687 : OR2_X2 port map( A1 => n6581, A2 => n6583, ZN => n1551);
   U1719 : AND2_X2 port map( A1 => n983, A2 => n4571, ZN => n555);
   U1875 : INV_X2 port map( A => n2167, ZN => n2141);
   U1928 : MUX2_X1 port map( A => n1719, B => n1720, S => n2265, Z => n1718);
   U2053 : MUX2_X1 port map( A => n6368, B => n6367, S => n986, Z => n1400);
   U2062 : MUX2_X1 port map( A => n5704, B => n5705, S => n6912, Z => n5815);
   U2069 : OR2_X2 port map( A1 => n6519, A2 => n6468, ZN => n6511);
   U2245 : NAND2_X1 port map( A1 => n4567, A2 => n1878, ZN => n17230);
   U2301 : BUF_X1 port map( A => n4864, Z => n1705);
   U2360 : MUX2_X2 port map( A => n5120, B => n5119, S => n2248, Z => n552);
   U2517 : OR2_X1 port map( A1 => n4499, A2 => n4463, ZN => n17231);
   U2550 : OR2_X2 port map( A1 => n17231, A2 => n17232, ZN => n4489);
   U2599 : OR2_X1 port map( A1 => n4465, A2 => n4464, ZN => n17232);
   U2615 : OR2_X1 port map( A1 => n1518, A2 => n1519, ZN => n17233);
   U2649 : OR2_X2 port map( A1 => n17233, A2 => n17234, ZN => n4512);
   U3825 : OR2_X1 port map( A1 => n4459, A2 => n4458, ZN => n17234);
   U6902 : BUF_X1 port map( A => n1228, Z => n17151);
   U16531 : NAND2_X1 port map( A1 => n1206, A2 => n4677, ZN => n17235);
   U16564 : OR2_X1 port map( A1 => n7370, A2 => n7369, ZN => n17236);
   U16579 : NAND2_X1 port map( A1 => n17236, A2 => n7368, ZN => n7371);
   U16880 : OR2_X2 port map( A1 => n4477, A2 => n4470, ZN => n5214);
   U16926 : INV_X2 port map( A => n2236, ZN => n17237);
   U16927 : INV_X1 port map( A => n17237, ZN => n17238);
   U16930 : INV_X2 port map( A => n17237, ZN => n17239);
   U17034 : INV_X1 port map( A => n17237, ZN => n17240);
   U17277 : MUX2_X1 port map( A => n6247, B => n6248, S => n6839, Z => n17186);
   U17299 : AND2_X2 port map( A1 => n983, A2 => n4571, ZN => n1467);
   U17300 : BUF_X1 port map( A => n4883, Z => n753);
   U17301 : AND2_X1 port map( A1 => n4871, A2 => n4870, ZN => n17241);
   U17304 : INV_X1 port map( A => n4783, ZN => n17242);
   U17316 : AND2_X2 port map( A1 => n1265, A2 => n1264, ZN => n1064);
   U17317 : BUF_X1 port map( A => n4948, Z => n734);
   U17426 : NAND2_X1 port map( A1 => n597, A2 => n2232, ZN => n17243);
   U17494 : XNOR2_X1 port map( A => n17244, B => n5877, ZN => n5886);
   U17520 : XOR2_X1 port map( A => n5879, B => n5878, Z => n17244);
   U17591 : AND2_X2 port map( A1 => n4490, A2 => n4489, ZN => n251);
   U17635 : INV_X1 port map( A => n251, ZN => n4681);
   U17681 : NAND2_X1 port map( A1 => n612, A2 => n6948, ZN => n17245);
   U17749 : CLKBUF_X1 port map( A => n6924, Z => n17246);
   U17840 : OR2_X1 port map( A1 => n4545, A2 => n4546, ZN => n17247);
   U17879 : OR2_X1 port map( A1 => n4545, A2 => n4546, ZN => n4652);
   U17952 : BUF_X1 port map( A => n548, Z => n597);
   U18265 : CLKBUF_X1 port map( A => n2155, Z => n609);
   U18266 : INV_X1 port map( A => n8179, ZN => n17248);
   U18411 : OR2_X1 port map( A1 => n6936, A2 => n6935, ZN => n6937);
   U18451 : INV_X1 port map( A => n776, ZN => n17249);
   U18500 : MUX2_X1 port map( A => n5727, B => n5726, S => n2243, Z => n17250);
   U18501 : MUX2_X1 port map( A => n5727, B => n5726, S => n2243, Z => n17251);
   U18571 : AND3_X1 port map( A1 => n4862, A2 => n17181, A3 => n1606, ZN => 
                           n17252);
   U18612 : MUX2_X1 port map( A => n5727, B => n5726, S => n2243, Z => n5821);
   U19017 : BUF_X1 port map( A => n4861, Z => n17181);
   U19058 : NAND2_X1 port map( A1 => n5018, A2 => n17253, ZN => n17254);
   U20022 : NAND2_X1 port map( A1 => n5017, A2 => n2248, ZN => n17255);
   U20023 : NAND2_X1 port map( A1 => n17254, A2 => n17255, ZN => n5357);
   U20024 : INV_X1 port map( A => n2248, ZN => n17253);
   U20025 : BUF_X4 port map( A => n799, Z => n2248);
   U20026 : MUX2_X1 port map( A => n5448, B => n5447, S => n2245, Z => n17256);
   U20027 : OAI21_X1 port map( B1 => n17258, B2 => n4944, A => n5165, ZN => 
                           n17257);
   U20028 : XNOR2_X1 port map( A => n513, B => n1817, ZN => n17258);
   U20029 : MUX2_X1 port map( A => n5448, B => n5447, S => n2245, Z => n1157);
   U20030 : MUX2_X1 port map( A => n5196, B => n5195, S => n2247, Z => n17259);
   U20031 : MUX2_X1 port map( A => n5196, B => n5195, S => n2247, Z => n5197);
   U20032 : OR2_X1 port map( A1 => n5385, A2 => n437, ZN => n17260);
   U20033 : OR2_X1 port map( A1 => n1600, A2 => n5387, ZN => n17261);
   U20034 : NAND3_X1 port map( A1 => n17260, A2 => n17261, A3 => n5288, ZN => 
                           n5380);
   U20035 : BUF_X1 port map( A => n5386, Z => n437);
   U20036 : BUF_X2 port map( A => n794, Z => n1358);
   U20037 : NAND2_X1 port map( A1 => n4873, A2 => n452, ZN => n17262);
   U20038 : XNOR2_X1 port map( A => n5858, B => n5857, ZN => n5863);
   U20039 : OR2_X1 port map( A1 => n6524, A2 => n17263, ZN => n6506);
   U20040 : INV_X1 port map( A => n6484, ZN => n17263);
   U20041 : XNOR2_X1 port map( A => n17168, B => n6016, ZN => n17264);
   U20042 : INV_X1 port map( A => n17264, ZN => n920);
   U20043 : MUX2_X2 port map( A => n6601, B => n6602, S => n6495, Z => n711);
   U20044 : XNOR2_X1 port map( A => n4981, B => n4988, ZN => n4995);
   U20045 : XNOR2_X1 port map( A => n5224, B => n5225, ZN => n4691);
   U20046 : OAI22_X1 port map( A1 => n2192, A2 => n7624, B1 => n2189, B2 => 
                           n1542, ZN => n4884);
   U20047 : XNOR2_X1 port map( A => n5254, B => n5255, ZN => n5226);
   U20048 : XNOR2_X1 port map( A => n489, B => n4773, ZN => n4774);
   U20049 : AOI22_X1 port map( A1 => n1368, A2 => n4607, B1 => n4663, B2 => 
                           n17242, ZN => n4778);
   U20050 : XOR2_X1 port map( A => n5069, B => n847, Z => n5070);
   U20051 : OAI211_X1 port map( C1 => n807, C2 => n4447, A => n4446, B => n4445
                           , ZN => n4576);
   U20052 : OAI222_X1 port map( A1 => n6947, A2 => n6946, B1 => n981, B2 => 
                           n1877, C1 => n6773, C2 => n6774, ZN => n6948);
   U20053 : OR2_X1 port map( A1 => n5122, A2 => n17265, ZN => n1288);
   U20054 : INV_X1 port map( A => n5145, ZN => n17265);
   U20055 : OAI33_X1 port map( A1 => n6698, A2 => n6697, A3 => n6699, B1 => 
                           n8229, B2 => n1154, B3 => n1846, ZN => n6791);
   U20056 : NAND3_X1 port map( A1 => n17266, A2 => n1875, A3 => n4943, ZN => 
                           n5148);
   U20057 : INV_X1 port map( A => n8180, ZN => n17266);
   U20058 : XNOR2_X1 port map( A => n896, B => n5523, ZN => n1766);
   U20059 : XNOR2_X1 port map( A => n5723, B => n5540, ZN => n5724);
   U20060 : AND3_X1 port map( A1 => n1899, A2 => n8164, A3 => n2154, ZN => 
                           n8154);
   U20061 : INV_X2 port map( A => n2131, ZN => n2154);
   U20062 : XNOR2_X1 port map( A => n908, B => n5336, ZN => n5340);
   U20063 : NAND2_X1 port map( A1 => n832, A2 => n1802, ZN => n5147);
   U20064 : AOI21_X1 port map( B1 => n4874, B2 => n4873, A => n1387, ZN => 
                           n4881);
   U20065 : AOI21_X1 port map( B1 => n4542, B2 => n17149, A => n2264, ZN => 
                           n4544);
   U20066 : NOR2_X1 port map( A1 => n17267, A2 => n1354, ZN => n1802);
   U20067 : INV_X1 port map( A => n1875, ZN => n17267);
   U20068 : OAI22_X1 port map( A1 => n1791, A2 => n5550, B1 => n5551, B2 => 
                           n5599, ZN => n5552);
   U20069 : OAI21_X1 port map( B1 => n6802, B2 => n1083, A => n6800, ZN => 
                           n17268);
   U20070 : INV_X1 port map( A => n17268, ZN => n7261);
   DataPath_REG_A_Q_reg_29_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_29_port, QN => n279);
   DataPath_REG_A_Q_reg_22_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_22_port, QN => n4411);
   DataPath_REG_A_Q_reg_24_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_24_port, QN => n4359);
   DataPath_REG_A_Q_reg_14_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_14_port, QN => n4334);
   DataPath_REG_A_Q_reg_7_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_7_port, QN => n4303);
   DataPath_REG_A_Q_reg_28_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_28_port, QN => n278);
   DataPath_REG_A_Q_reg_21_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_21_port, QN => n4417);
   DataPath_REG_A_Q_reg_18_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_18_port, QN => n4395);
   DataPath_REG_A_Q_reg_6_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_6_port, QN => n811);
   DataPath_REG_A_Q_reg_30_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_30_port, QN => n280);
   DataPath_REG_A_Q_reg_27_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_27_port, QN => n4367);
   DataPath_REG_A_Q_reg_23_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_23_port, QN => n4408);
   DataPath_REG_A_Q_reg_20_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_20_port, QN => n4414);
   DataPath_REG_A_Q_reg_17_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_17_port, QN => n4397);
   DataPath_REG_A_Q_reg_10_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_10_port, QN => n4314);
   DataPath_REG_A_Q_reg_25_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_25_port, QN => n4356);
   DataPath_REG_A_Q_reg_15_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_15_port, QN => n4343);
   DataPath_REG_A_Q_reg_8_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_8_port, QN => n4315);
   DataPath_REG_A_Q_reg_26_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_26_port, QN => n4370);
   DataPath_REG_A_Q_reg_19_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_19_port, QN => n4392);
   DataPath_REG_A_Q_reg_16_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_16_port, QN => n4396);
   DataPath_REG_A_Q_reg_31_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_31_port, QN => n7082);
   DataPath_REG_A_Q_reg_4_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_4_port, QN => n1544);
   DataPath_REG_A_Q_reg_0_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_0_port, QN => n4269);
   DataPath_REG_A_Q_reg_1_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_1_port, QN => n4267);
   DataPath_REG_A_Q_reg_2_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_2_port, QN => n4273);
   DataPath_REG_CMP_Q_reg_0_inst : DFF_X1 port map( D => n2032, CK => CLK, Q =>
                           DataPath_i_LGET_0_port, QN => n11591);
   CU_I_CW_WB_reg_1_inst : DFF_X1 port map( D => CU_I_N50, CK => CLK, Q => n256
                           , QN => n409);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N46_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n18);
   CU_I_aluOpcode1_reg_1_inst : DFF_X1 port map( D => CU_I_n154, CK => CLK, Q 
                           => i_ALU_OP_1_port, QN => n7080);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_14_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N60, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n4);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_13_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N59, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n5);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_12_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N58, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n6);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_11_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N57, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n7);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_10_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N56, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n8);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_9_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N55, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n9);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_8_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N54_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n10);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_7_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N53_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n11);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_6_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N52_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n12);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_5_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N51_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n13);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_4_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N50_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n14);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_3_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N49_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n15);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_2_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N48_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n16);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N47_port, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n17);
   CU_I_CW_EX_reg_18_inst : DFF_X1 port map( D => CU_I_n126, CK => CLK, Q => 
                           n4426, QN => CU_I_n109);
   CU_I_CW_EX_reg_17_inst : DFF_X1 port map( D => CU_I_n127, CK => CLK, Q => 
                           i_S1, QN => CU_I_n108);
   CU_I_CW_EX_reg_16_inst : DFF_X1 port map( D => CU_I_n128, CK => CLK, Q => 
                           i_S2, QN => CU_I_n107);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N61, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n1);
   CU_I_setcmp_1_reg_1_inst : DFF_X1 port map( D => CU_I_n146, CK => CLK, Q => 
                           i_SEL_LGET_1_port, QN => CU_I_n118);
   CU_I_setcmp_1_reg_0_inst : DFF_X1 port map( D => CU_I_n147, CK => CLK, Q => 
                           i_SEL_LGET_0_port, QN => n11483);
   CU_I_aluOpcode1_reg_2_inst : DFF_X1 port map( D => CU_I_n144, CK => CLK, Q 
                           => n259, QN => n4140);
   CU_I_sel_alu_setcmp_1_reg : DFF_X1 port map( D => CU_I_n152, CK => CLK, Q =>
                           i_SEL_ALU_SETCMP, QN => n8325);
   CU_I_aluOpcode1_reg_4_inst : DFF_X1 port map( D => CU_I_n156, CK => CLK, Q 
                           => i_ALU_OP_4_port, QN => n11540);
   CU_I_aluOpcode1_reg_3_inst : DFF_X1 port map( D => CU_I_n155, CK => CLK, Q 
                           => i_ALU_OP_3_port, QN => CU_I_n114);
   CU_I_aluOpcode1_reg_0_inst : DFF_X1 port map( D => CU_I_n153, CK => CLK, Q 
                           => i_ALU_OP_0_port, QN => n7081);
   CU_I_unsigned_2_reg : DFF_X1 port map( D => CU_I_n148, CK => CLK, Q => 
                           i_UNSIG_SIGN_N, QN => n11480);
   CU_I_CW_MEM_reg_5_inst : DFF_X1 port map( D => CU_I_n137, CK => CLK, Q => 
                           i_DATAMEM_RM, QN => CU_I_n104);
   CU_I_CW_MEM_reg_4_inst : DFF_X1 port map( D => CU_I_n138, CK => CLK, Q => 
                           DATA_SIZE_1_port, QN => CU_I_n102);
   CU_I_CW_MEM_reg_3_inst : DFF_X1 port map( D => CU_I_n139, CK => CLK, Q => 
                           DATA_SIZE_0_port, QN => n11579);
   DataPath_RF_CWP_Q_reg_0_inst : DFF_X1 port map( D => n429, CK => CLK, Q => 
                           DataPath_RF_c_win_0_port, QN => n11592);
   DataPath_RF_CWP_Q_reg_3_inst : DFF_X1 port map( D => n423, CK => CLK, Q => 
                           DataPath_RF_c_win_3_port, QN => n11595);
   DataPath_RF_CWP_Q_reg_1_inst : DFF_X1 port map( D => n421, CK => CLK, Q => 
                           DataPath_RF_c_win_1_port, QN => n11593);
   DataPath_RF_CWP_Q_reg_2_inst : DFF_X1 port map( D => n422, CK => CLK, Q => 
                           DataPath_RF_c_win_2_port, QN => n11594);
   DataPath_RF_PUSH_ADDRGEN_curr_state_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_n53, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_state_1_port, QN => 
                           DataPath_RF_PUSH_ADDRGEN_n20);

end SYN_dlx_rtl;
