
module hazard_table_N_REGS_LOG5 ( CLK, RST, WR1, WR2, ADD_WR1, ADD_WR2, 
        ADD_CHECK1, ADD_CHECK2, BUSY, BUSY_WINDOW );
  input [4:0] ADD_WR1;
  input [4:0] ADD_WR2;
  input [4:0] ADD_CHECK1;
  input [4:0] ADD_CHECK2;
  input CLK, RST, WR1, WR2;
  output BUSY, BUSY_WINDOW;
  wire   \Table[0][2] , \Table[0][1] , \Table[0][0] , \Table[1][2] ,
         \Table[1][1] , \Table[1][0] , \Table[2][2] , \Table[2][1] ,
         \Table[2][0] , \Table[3][2] , \Table[3][1] , \Table[3][0] ,
         \Table[4][2] , \Table[4][1] , \Table[4][0] , \Table[5][2] ,
         \Table[5][1] , \Table[5][0] , \Table[6][2] , \Table[6][1] ,
         \Table[6][0] , \Table[7][2] , \Table[7][1] , \Table[7][0] ,
         \Table[8][2] , \Table[8][1] , \Table[8][0] , \Table[9][2] ,
         \Table[9][1] , \Table[9][0] , \Table[10][2] , \Table[10][1] ,
         \Table[10][0] , \Table[11][2] , \Table[11][1] , \Table[11][0] ,
         \Table[12][2] , \Table[12][1] , \Table[12][0] , \Table[13][2] ,
         \Table[13][1] , \Table[13][0] , \Table[14][2] , \Table[14][1] ,
         \Table[14][0] , \Table[15][2] , \Table[15][1] , \Table[15][0] ,
         \Table[16][2] , \Table[16][1] , \Table[16][0] , \Table[17][2] ,
         \Table[17][1] , \Table[17][0] , \Table[18][2] , \Table[18][1] ,
         \Table[18][0] , \Table[19][2] , \Table[19][1] , \Table[19][0] ,
         \Table[20][2] , \Table[20][1] , \Table[20][0] , \Table[21][2] ,
         \Table[21][1] , \Table[21][0] , \Table[22][2] , \Table[22][1] ,
         \Table[22][0] , \Table[23][2] , \Table[23][1] , \Table[23][0] ,
         \Table[24][2] , \Table[24][1] , \Table[24][0] , \Table[25][2] ,
         \Table[25][1] , \Table[25][0] , \Table[26][2] , \Table[26][1] ,
         \Table[26][0] , \Table[27][2] , \Table[27][1] , \Table[27][0] ,
         \Table[28][2] , \Table[28][1] , \Table[28][0] , \Table[29][2] ,
         \Table[29][1] , \Table[29][0] , \Table[30][2] , \Table[30][1] ,
         \Table[30][0] , \Table[31][2] , \Table[31][1] , \Table[31][0] , N192,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671;
  assign BUSY = N192;

  DFF_X1 \Table_reg[19][0]  ( .D(n761), .CK(CLK), .Q(\Table[19][0] ), .QN(n50)
         );
  DFF_X1 \Table_reg[27][0]  ( .D(n785), .CK(CLK), .Q(\Table[27][0] ), .QN(n52)
         );
  DFF_X1 \Table_reg[19][2]  ( .D(n759), .CK(CLK), .Q(\Table[19][2] ), .QN(n51)
         );
  DFF_X1 \Table_reg[27][2]  ( .D(n783), .CK(CLK), .Q(\Table[27][2] ), .QN(n53)
         );
  DFF_X1 \Table_reg[30][2]  ( .D(n792), .CK(CLK), .Q(\Table[30][2] ), .QN(n54)
         );
  DFF_X1 \Table_reg[16][0]  ( .D(n752), .CK(CLK), .Q(\Table[16][0] ), .QN(n48)
         );
  DFF_X1 \Table_reg[15][0]  ( .D(n749), .CK(CLK), .Q(\Table[15][0] ), .QN(n521) );
  DFF_X1 \Table_reg[9][0]  ( .D(n731), .CK(CLK), .Q(\Table[9][0] ), .QN(n38)
         );
  DFF_X1 \Table_reg[8][0]  ( .D(n728), .CK(CLK), .Q(\Table[8][0] ), .QN(n589)
         );
  DFF_X1 \Table_reg[6][0]  ( .D(n722), .CK(CLK), .Q(\Table[6][0] ), .QN(n29)
         );
  DFF_X1 \Table_reg[5][0]  ( .D(n719), .CK(CLK), .Q(\Table[5][0] ), .QN(n39)
         );
  DFF_X1 \Table_reg[4][0]  ( .D(n716), .CK(CLK), .Q(\Table[4][0] ), .QN(n30)
         );
  DFF_X1 \Table_reg[3][0]  ( .D(n713), .CK(CLK), .Q(\Table[3][0] ), .QN(n19)
         );
  DFF_X1 \Table_reg[2][0]  ( .D(n710), .CK(CLK), .Q(\Table[2][0] ), .QN(n31)
         );
  DFF_X1 \Table_reg[1][0]  ( .D(n707), .CK(CLK), .Q(\Table[1][0] ), .QN(n40)
         );
  DFF_X1 \Table_reg[30][0]  ( .D(n794), .CK(CLK), .Q(\Table[30][0] ), .QN(n374) );
  DFF_X1 \Table_reg[29][0]  ( .D(n791), .CK(CLK), .Q(\Table[29][0] ), .QN(n384) );
  DFF_X1 \Table_reg[28][0]  ( .D(n788), .CK(CLK), .Q(\Table[28][0] ), .QN(n15)
         );
  DFF_X1 \Table_reg[26][0]  ( .D(n782), .CK(CLK), .Q(\Table[26][0] ), .QN(n413) );
  DFF_X1 \Table_reg[25][0]  ( .D(n779), .CK(CLK), .Q(\Table[25][0] ), .QN(n424) );
  DFF_X1 \Table_reg[24][0]  ( .D(n776), .CK(CLK), .Q(\Table[24][0] ), .QN(n20)
         );
  DFF_X1 \Table_reg[23][0]  ( .D(n773), .CK(CLK), .Q(\Table[23][0] ), .QN(n446) );
  DFF_X1 \Table_reg[22][0]  ( .D(n770), .CK(CLK), .Q(\Table[22][0] ), .QN(n456) );
  DFF_X1 \Table_reg[21][0]  ( .D(n767), .CK(CLK), .Q(\Table[21][0] ), .QN(n16)
         );
  DFF_X1 \Table_reg[20][0]  ( .D(n764), .CK(CLK), .Q(\Table[20][0] ), .QN(n474) );
  DFF_X1 \Table_reg[18][0]  ( .D(n758), .CK(CLK), .Q(\Table[18][0] ), .QN(n492) );
  DFF_X1 \Table_reg[17][0]  ( .D(n755), .CK(CLK), .Q(\Table[17][0] ), .QN(n502) );
  DFF_X1 \Table_reg[14][0]  ( .D(n746), .CK(CLK), .Q(\Table[14][0] ), .QN(n531) );
  DFF_X1 \Table_reg[13][0]  ( .D(n743), .CK(CLK), .Q(\Table[13][0] ), .QN(n541) );
  DFF_X1 \Table_reg[12][0]  ( .D(n740), .CK(CLK), .Q(\Table[12][0] ), .QN(n551) );
  DFF_X1 \Table_reg[11][0]  ( .D(n737), .CK(CLK), .Q(\Table[11][0] ), .QN(n561) );
  DFF_X1 \Table_reg[10][0]  ( .D(n734), .CK(CLK), .Q(\Table[10][0] ), .QN(n571) );
  DFF_X1 \Table_reg[7][0]  ( .D(n725), .CK(CLK), .Q(\Table[7][0] ), .QN(n18)
         );
  DFF_X1 \Table_reg[0][0]  ( .D(n704), .CK(CLK), .Q(\Table[0][0] ), .QN(n17)
         );
  DFF_X1 \Table_reg[31][0]  ( .D(n797), .CK(CLK), .Q(\Table[31][0] ), .QN(n261) );
  DFF_X1 \Table_reg[31][1]  ( .D(n796), .CK(CLK), .Q(\Table[31][1] ), .QN(n313) );
  DFF_X1 \Table_reg[30][1]  ( .D(n793), .CK(CLK), .Q(\Table[30][1] ), .QN(n376) );
  DFF_X1 \Table_reg[29][1]  ( .D(n790), .CK(CLK), .Q(\Table[29][1] ), .QN(n386) );
  DFF_X1 \Table_reg[28][1]  ( .D(n787), .CK(CLK), .Q(\Table[28][1] ), .QN(n21)
         );
  DFF_X1 \Table_reg[27][1]  ( .D(n784), .CK(CLK), .Q(\Table[27][1] ), .QN(n405) );
  DFF_X1 \Table_reg[26][1]  ( .D(n781), .CK(CLK), .Q(\Table[26][1] ), .QN(n415) );
  DFF_X1 \Table_reg[25][1]  ( .D(n778), .CK(CLK), .Q(\Table[25][1] ), .QN(n426) );
  DFF_X1 \Table_reg[24][1]  ( .D(n775), .CK(CLK), .Q(\Table[24][1] ), .QN(n437) );
  DFF_X1 \Table_reg[23][1]  ( .D(n772), .CK(CLK), .Q(\Table[23][1] ), .QN(n448) );
  DFF_X1 \Table_reg[22][1]  ( .D(n769), .CK(CLK), .Q(\Table[22][1] ), .QN(n458) );
  DFF_X1 \Table_reg[21][1]  ( .D(n766), .CK(CLK), .Q(\Table[21][1] ), .QN(n22)
         );
  DFF_X1 \Table_reg[20][1]  ( .D(n763), .CK(CLK), .Q(\Table[20][1] ), .QN(n476) );
  DFF_X1 \Table_reg[19][1]  ( .D(n760), .CK(CLK), .Q(\Table[19][1] ), .QN(n485) );
  DFF_X1 \Table_reg[18][1]  ( .D(n757), .CK(CLK), .Q(\Table[18][1] ), .QN(n494) );
  DFF_X1 \Table_reg[17][1]  ( .D(n754), .CK(CLK), .Q(\Table[17][1] ), .QN(n504) );
  DFF_X1 \Table_reg[16][1]  ( .D(n751), .CK(CLK), .Q(\Table[16][1] ), .QN(n5)
         );
  DFF_X1 \Table_reg[15][1]  ( .D(n748), .CK(CLK), .Q(\Table[15][1] ), .QN(n523) );
  DFF_X1 \Table_reg[14][1]  ( .D(n745), .CK(CLK), .Q(\Table[14][1] ), .QN(n533) );
  DFF_X1 \Table_reg[13][1]  ( .D(n742), .CK(CLK), .Q(\Table[13][1] ), .QN(n543) );
  DFF_X1 \Table_reg[12][1]  ( .D(n739), .CK(CLK), .Q(\Table[12][1] ), .QN(n553) );
  DFF_X1 \Table_reg[11][1]  ( .D(n736), .CK(CLK), .Q(\Table[11][1] ), .QN(n563) );
  DFF_X1 \Table_reg[10][1]  ( .D(n733), .CK(CLK), .Q(\Table[10][1] ), .QN(n573) );
  DFF_X1 \Table_reg[8][1]  ( .D(n727), .CK(CLK), .Q(\Table[8][1] ), .QN(n591)
         );
  DFF_X1 \Table_reg[7][1]  ( .D(n724), .CK(CLK), .Q(\Table[7][1] ), .QN(n24)
         );
  DFF_X1 \Table_reg[5][1]  ( .D(n718), .CK(CLK), .Q(\Table[5][1] ), .QN(n36)
         );
  DFF_X1 \Table_reg[3][1]  ( .D(n712), .CK(CLK), .Q(\Table[3][1] ), .QN(n25)
         );
  DFF_X1 \Table_reg[1][1]  ( .D(n706), .CK(CLK), .Q(\Table[1][1] ), .QN(n37)
         );
  DFF_X1 \Table_reg[0][1]  ( .D(n703), .CK(CLK), .Q(\Table[0][1] ), .QN(n23)
         );
  DFF_X1 \Table_reg[9][1]  ( .D(n730), .CK(CLK), .Q(\Table[9][1] ), .QN(n35)
         );
  DFF_X1 \Table_reg[6][1]  ( .D(n721), .CK(CLK), .Q(\Table[6][1] ), .QN(n26)
         );
  DFF_X1 \Table_reg[4][1]  ( .D(n715), .CK(CLK), .Q(\Table[4][1] ), .QN(n27)
         );
  DFF_X1 \Table_reg[2][1]  ( .D(n709), .CK(CLK), .Q(\Table[2][1] ), .QN(n28)
         );
  DFF_X1 \Table_reg[24][2]  ( .D(n774), .CK(CLK), .Q(\Table[24][2] ), .QN(n442) );
  DFF_X1 \Table_reg[9][2]  ( .D(n729), .CK(CLK), .Q(\Table[9][2] ), .QN(n41)
         );
  DFF_X1 \Table_reg[8][2]  ( .D(n726), .CK(CLK), .Q(\Table[8][2] ), .QN(n596)
         );
  DFF_X1 \Table_reg[7][2]  ( .D(n723), .CK(CLK), .Q(\Table[7][2] ), .QN(n13)
         );
  DFF_X1 \Table_reg[6][2]  ( .D(n720), .CK(CLK), .Q(\Table[6][2] ), .QN(n32)
         );
  DFF_X1 \Table_reg[5][2]  ( .D(n717), .CK(CLK), .Q(\Table[5][2] ), .QN(n42)
         );
  DFF_X1 \Table_reg[4][2]  ( .D(n714), .CK(CLK), .Q(\Table[4][2] ), .QN(n33)
         );
  DFF_X1 \Table_reg[3][2]  ( .D(n711), .CK(CLK), .Q(\Table[3][2] ), .QN(n14)
         );
  DFF_X1 \Table_reg[2][2]  ( .D(n708), .CK(CLK), .Q(\Table[2][2] ), .QN(n34)
         );
  DFF_X1 \Table_reg[1][2]  ( .D(n705), .CK(CLK), .Q(\Table[1][2] ), .QN(n43)
         );
  DFF_X1 \Table_reg[31][2]  ( .D(n795), .CK(CLK), .Q(\Table[31][2] ), .QN(n7)
         );
  DFF_X1 \Table_reg[29][2]  ( .D(n789), .CK(CLK), .Q(\Table[29][2] ), .QN(n391) );
  DFF_X1 \Table_reg[28][2]  ( .D(n786), .CK(CLK), .Q(\Table[28][2] ), .QN(n400) );
  DFF_X1 \Table_reg[26][2]  ( .D(n780), .CK(CLK), .Q(\Table[26][2] ), .QN(n420) );
  DFF_X1 \Table_reg[25][2]  ( .D(n777), .CK(CLK), .Q(\Table[25][2] ), .QN(n431) );
  DFF_X1 \Table_reg[23][2]  ( .D(n771), .CK(CLK), .Q(\Table[23][2] ), .QN(n453) );
  DFF_X1 \Table_reg[22][2]  ( .D(n768), .CK(CLK), .Q(\Table[22][2] ), .QN(n463) );
  DFF_X1 \Table_reg[21][2]  ( .D(n765), .CK(CLK), .Q(\Table[21][2] ), .QN(n471) );
  DFF_X1 \Table_reg[20][2]  ( .D(n762), .CK(CLK), .Q(\Table[20][2] ), .QN(n481) );
  DFF_X1 \Table_reg[18][2]  ( .D(n756), .CK(CLK), .Q(\Table[18][2] ), .QN(n499) );
  DFF_X1 \Table_reg[17][2]  ( .D(n753), .CK(CLK), .Q(\Table[17][2] ), .QN(n509) );
  DFF_X1 \Table_reg[16][2]  ( .D(n750), .CK(CLK), .Q(\Table[16][2] ), .QN(n49)
         );
  DFF_X1 \Table_reg[15][2]  ( .D(n747), .CK(CLK), .Q(\Table[15][2] ), .QN(n528) );
  DFF_X1 \Table_reg[14][2]  ( .D(n744), .CK(CLK), .Q(\Table[14][2] ), .QN(n538) );
  DFF_X1 \Table_reg[13][2]  ( .D(n741), .CK(CLK), .Q(\Table[13][2] ), .QN(n548) );
  DFF_X1 \Table_reg[12][2]  ( .D(n738), .CK(CLK), .Q(\Table[12][2] ), .QN(n558) );
  DFF_X1 \Table_reg[10][2]  ( .D(n732), .CK(CLK), .Q(\Table[10][2] ), .QN(n578) );
  DFF_X1 \Table_reg[0][2]  ( .D(n702), .CK(CLK), .Q(\Table[0][2] ), .QN(n12)
         );
  DFF_X1 \Table_reg[11][2]  ( .D(n735), .CK(CLK), .Q(\Table[11][2] ), .QN(n568) );
  AND2_X2 U3 ( .A1(n361), .A2(n284), .ZN(n660) );
  AOI21_X1 U4 ( .B1(n192), .B2(WR1), .A(n191), .ZN(n656) );
  AND3_X2 U5 ( .A1(n386), .A2(n391), .A3(n384), .ZN(n47) );
  BUF_X2 U6 ( .A(n663), .Z(n2) );
  BUF_X1 U7 ( .A(n656), .Z(n59) );
  BUF_X2 U8 ( .A(n668), .Z(n3) );
  BUF_X2 U9 ( .A(n662), .Z(n4) );
  INV_X1 U10 ( .A(ADD_WR1[2]), .ZN(n235) );
  INV_X1 U11 ( .A(ADD_WR1[1]), .ZN(n234) );
  AND3_X1 U12 ( .A1(n415), .A2(n413), .A3(n420), .ZN(n140) );
  AND3_X1 U13 ( .A1(n35), .A2(n38), .A3(n41), .ZN(n167) );
  AND3_X1 U14 ( .A1(n543), .A2(n541), .A3(n548), .ZN(n159) );
  AND3_X1 U15 ( .A1(n504), .A2(n502), .A3(n509), .ZN(n171) );
  AND3_X1 U16 ( .A1(n426), .A2(n424), .A3(n431), .ZN(n169) );
  BUF_X1 U17 ( .A(n665), .Z(n61) );
  NOR2_X2 U18 ( .A1(ADD_WR1[1]), .A2(n232), .ZN(n382) );
  NAND3_X1 U19 ( .A1(n553), .A2(n551), .A3(n558), .ZN(n6) );
  AND3_X1 U20 ( .A1(n448), .A2(n446), .A3(n453), .ZN(n8) );
  AND3_X1 U21 ( .A1(n376), .A2(n374), .A3(n54), .ZN(n148) );
  AND3_X1 U22 ( .A1(n563), .A2(n561), .A3(n568), .ZN(n136) );
  AND3_X1 U23 ( .A1(n573), .A2(n571), .A3(n578), .ZN(n9) );
  AND3_X1 U24 ( .A1(n533), .A2(n531), .A3(n538), .ZN(n10) );
  AND3_X1 U25 ( .A1(n405), .A2(n52), .A3(n53), .ZN(n137) );
  AND3_X1 U26 ( .A1(n591), .A2(n589), .A3(n596), .ZN(n96) );
  AND3_X1 U27 ( .A1(n485), .A2(n50), .A3(n51), .ZN(n141) );
  AND3_X1 U28 ( .A1(n523), .A2(n521), .A3(n528), .ZN(n145) );
  AND4_X1 U29 ( .A1(n140), .A2(n136), .A3(n137), .A4(n141), .ZN(n55) );
  AND2_X1 U30 ( .A1(n167), .A2(n67), .ZN(n11) );
  AND3_X1 U31 ( .A1(n313), .A2(n261), .A3(n7), .ZN(n146) );
  AND3_X1 U32 ( .A1(n553), .A2(n551), .A3(n558), .ZN(n97) );
  AND3_X1 U33 ( .A1(n448), .A2(n446), .A3(n453), .ZN(n149) );
  AND3_X1 U34 ( .A1(n573), .A2(n571), .A3(n578), .ZN(n91) );
  AND3_X1 U35 ( .A1(n533), .A2(n531), .A3(n538), .ZN(n92) );
  AND4_X1 U36 ( .A1(n148), .A2(n145), .A3(n146), .A4(n149), .ZN(n56) );
  AND4_X1 U37 ( .A1(n55), .A2(n56), .A3(n57), .A4(n58), .ZN(n65) );
  AND4_X1 U38 ( .A1(n97), .A2(n96), .A3(n91), .A4(n92), .ZN(n57) );
  NOR3_X1 U39 ( .A1(n64), .A2(n115), .A3(n163), .ZN(n66) );
  NAND3_X1 U40 ( .A1(n65), .A2(n11), .A3(n66), .ZN(BUSY_WINDOW) );
  BUF_X1 U41 ( .A(n659), .Z(n60) );
  INV_X1 U42 ( .A(ADD_WR1[0]), .ZN(n233) );
  INV_X1 U43 ( .A(ADD_CHECK2[4]), .ZN(n138) );
  INV_X1 U44 ( .A(n174), .ZN(n67) );
  AOI21_X1 U45 ( .B1(n364), .B2(n363), .A(n362), .ZN(n665) );
  NOR2_X1 U46 ( .A1(RST), .A2(n308), .ZN(n659) );
  NAND3_X1 U47 ( .A1(n437), .A2(n20), .A3(n442), .ZN(n174) );
  NAND3_X1 U48 ( .A1(n22), .A2(n16), .A3(n471), .ZN(n115) );
  NAND3_X1 U49 ( .A1(n21), .A2(n15), .A3(n400), .ZN(n163) );
  INV_X1 U50 ( .A(n393), .ZN(n624) );
  INV_X1 U51 ( .A(n422), .ZN(n648) );
  INV_X1 U52 ( .A(n402), .ZN(n632) );
  INV_X1 U53 ( .A(n433), .ZN(n658) );
  INV_X1 U54 ( .A(n411), .ZN(n640) );
  INV_X1 U55 ( .A(n370), .ZN(n608) );
  INV_X1 U56 ( .A(n328), .ZN(n600) );
  INV_X1 U57 ( .A(RST), .ZN(n62) );
  INV_X1 U58 ( .A(RST), .ZN(n63) );
  INV_X1 U59 ( .A(n382), .ZN(n616) );
  INV_X1 U60 ( .A(ADD_WR2[3]), .ZN(n213) );
  NOR3_X2 U61 ( .A1(n234), .A2(n235), .A3(n233), .ZN(n328) );
  NOR3_X2 U62 ( .A1(ADD_WR1[0]), .A2(n235), .A3(n234), .ZN(n370) );
  NOR3_X2 U63 ( .A1(ADD_WR1[1]), .A2(ADD_WR1[0]), .A3(n235), .ZN(n393) );
  NOR3_X2 U64 ( .A1(ADD_WR1[2]), .A2(n234), .A3(n233), .ZN(n402) );
  NOR3_X2 U65 ( .A1(ADD_WR1[2]), .A2(ADD_WR1[0]), .A3(n234), .ZN(n411) );
  NOR3_X2 U66 ( .A1(ADD_WR1[1]), .A2(ADD_WR1[2]), .A3(n233), .ZN(n422) );
  NOR3_X2 U67 ( .A1(ADD_WR1[1]), .A2(ADD_WR1[2]), .A3(ADD_WR1[0]), .ZN(n433)
         );
  INV_X1 U68 ( .A(ADD_WR2[2]), .ZN(n194) );
  INV_X1 U69 ( .A(ADD_WR2[4]), .ZN(n214) );
  OAI22_X1 U70 ( .A1(n170), .A2(n160), .B1(n47), .B2(n168), .ZN(n161) );
  OAI22_X1 U71 ( .A1(n123), .A2(n160), .B1(n47), .B2(n124), .ZN(n118) );
  AND3_X1 U72 ( .A1(n476), .A2(n474), .A3(n481), .ZN(n88) );
  AND3_X1 U73 ( .A1(n458), .A2(n456), .A3(n463), .ZN(n84) );
  AND3_X1 U74 ( .A1(n492), .A2(n494), .A3(n499), .ZN(n83) );
  NOR3_X1 U75 ( .A1(n45), .A2(n44), .A3(n46), .ZN(n58) );
  NAND4_X1 U76 ( .A1(n499), .A2(n456), .A3(n474), .A4(n463), .ZN(n44) );
  NAND4_X1 U77 ( .A1(n49), .A2(n48), .A3(n5), .A4(n481), .ZN(n45) );
  NAND4_X1 U78 ( .A1(n476), .A2(n492), .A3(n458), .A4(n494), .ZN(n46) );
  NAND4_X1 U79 ( .A1(n159), .A2(n171), .A3(n169), .A4(n47), .ZN(n64) );
  AOI221_X1 U80 ( .B1(n177), .B2(n83), .C1(ADD_CHECK2[2]), .C2(n84), .A(n69), 
        .ZN(n68) );
  NAND3_X1 U81 ( .A1(n5), .A2(n48), .A3(n49), .ZN(n86) );
  NOR2_X1 U82 ( .A1(ADD_CHECK2[1]), .A2(ADD_CHECK2[2]), .ZN(n71) );
  INV_X1 U83 ( .A(ADD_CHECK2[2]), .ZN(n177) );
  INV_X1 U84 ( .A(ADD_CHECK2[1]), .ZN(n69) );
  AOI211_X1 U85 ( .C1(n86), .C2(n71), .A(n138), .B(n68), .ZN(n76) );
  NAND2_X1 U86 ( .A1(n69), .A2(ADD_CHECK2[2]), .ZN(n75) );
  NOR3_X1 U87 ( .A1(\Table[4][1] ), .A2(\Table[4][0] ), .A3(\Table[4][2] ), 
        .ZN(n105) );
  NAND3_X1 U88 ( .A1(n23), .A2(n17), .A3(n12), .ZN(n102) );
  NOR3_X1 U89 ( .A1(\Table[2][1] ), .A2(\Table[2][0] ), .A3(\Table[2][2] ), 
        .ZN(n99) );
  NAND2_X1 U90 ( .A1(ADD_CHECK2[1]), .A2(n177), .ZN(n156) );
  NOR3_X1 U91 ( .A1(\Table[6][1] ), .A2(\Table[6][0] ), .A3(\Table[6][2] ), 
        .ZN(n100) );
  NAND2_X1 U92 ( .A1(ADD_CHECK2[1]), .A2(ADD_CHECK2[2]), .ZN(n154) );
  OAI22_X1 U93 ( .A1(n99), .A2(n156), .B1(n100), .B2(n154), .ZN(n70) );
  AOI211_X1 U94 ( .C1(n71), .C2(n102), .A(ADD_CHECK2[4]), .B(n70), .ZN(n72) );
  AOI221_X1 U95 ( .B1(n105), .B2(n72), .C1(n75), .C2(n72), .A(ADD_CHECK2[3]), 
        .ZN(n73) );
  INV_X1 U96 ( .A(n73), .ZN(n74) );
  AOI221_X1 U97 ( .B1(n76), .B2(n75), .C1(n76), .C2(n88), .A(n74), .ZN(n77) );
  INV_X1 U98 ( .A(n77), .ZN(n185) );
  OAI22_X1 U99 ( .A1(n9), .A2(n156), .B1(n10), .B2(n154), .ZN(n79) );
  AOI221_X1 U100 ( .B1(ADD_CHECK2[2]), .B2(n97), .C1(n177), .C2(n96), .A(
        ADD_CHECK2[1]), .ZN(n78) );
  OAI211_X1 U101 ( .C1(n79), .C2(n78), .A(ADD_CHECK2[3]), .B(n138), .ZN(n184)
         );
  NOR2_X1 U102 ( .A1(ADD_CHECK1[1]), .A2(ADD_CHECK1[2]), .ZN(n112) );
  INV_X1 U103 ( .A(ADD_CHECK1[3]), .ZN(n110) );
  NAND2_X1 U104 ( .A1(ADD_CHECK1[1]), .A2(ADD_CHECK1[2]), .ZN(n128) );
  INV_X1 U105 ( .A(ADD_CHECK1[1]), .ZN(n82) );
  NOR2_X1 U106 ( .A1(ADD_CHECK1[2]), .A2(n82), .ZN(n120) );
  INV_X1 U107 ( .A(n120), .ZN(n98) );
  OAI22_X1 U108 ( .A1(n128), .A2(n148), .B1(n140), .B2(n98), .ZN(n80) );
  AOI211_X1 U109 ( .C1(n174), .C2(n112), .A(n110), .B(n80), .ZN(n81) );
  INV_X1 U110 ( .A(n81), .ZN(n90) );
  NAND2_X1 U111 ( .A1(n82), .A2(ADD_CHECK1[2]), .ZN(n104) );
  INV_X1 U112 ( .A(n104), .ZN(n116) );
  OAI22_X1 U113 ( .A1(n84), .A2(n128), .B1(n83), .B2(n98), .ZN(n85) );
  AOI211_X1 U114 ( .C1(n112), .C2(n86), .A(ADD_CHECK1[3]), .B(n85), .ZN(n87)
         );
  OAI21_X1 U115 ( .B1(n88), .B2(n104), .A(n87), .ZN(n89) );
  OAI221_X1 U116 ( .B1(n90), .B2(n116), .C1(n90), .C2(n163), .A(n89), .ZN(n109) );
  INV_X1 U117 ( .A(ADD_CHECK1[4]), .ZN(n111) );
  INV_X1 U118 ( .A(n112), .ZN(n95) );
  OAI22_X1 U119 ( .A1(n128), .A2(n10), .B1(n98), .B2(n9), .ZN(n93) );
  INV_X1 U120 ( .A(n93), .ZN(n94) );
  OAI211_X1 U121 ( .C1(n96), .C2(n95), .A(ADD_CHECK1[3]), .B(n94), .ZN(n107)
         );
  OAI22_X1 U122 ( .A1(n100), .A2(n128), .B1(n99), .B2(n98), .ZN(n101) );
  AOI211_X1 U123 ( .C1(n112), .C2(n102), .A(ADD_CHECK1[3]), .B(n101), .ZN(n103) );
  OAI21_X1 U124 ( .B1(n105), .B2(n104), .A(n103), .ZN(n106) );
  OAI221_X1 U125 ( .B1(n107), .B2(n116), .C1(n107), .C2(n6), .A(n106), .ZN(
        n108) );
  AOI221_X1 U126 ( .B1(ADD_CHECK1[4]), .B2(n109), .C1(n111), .C2(n108), .A(
        ADD_CHECK1[0]), .ZN(n182) );
  NAND3_X1 U127 ( .A1(ADD_CHECK1[4]), .A2(ADD_CHECK1[0]), .A3(n110), .ZN(n123)
         );
  NAND3_X1 U128 ( .A1(ADD_CHECK1[0]), .A2(ADD_CHECK1[4]), .A3(ADD_CHECK1[3]), 
        .ZN(n124) );
  OAI22_X1 U129 ( .A1(n171), .A2(n123), .B1(n169), .B2(n124), .ZN(n114) );
  NAND3_X1 U130 ( .A1(ADD_CHECK1[0]), .A2(ADD_CHECK1[3]), .A3(n111), .ZN(n127)
         );
  NOR3_X1 U131 ( .A1(\Table[1][1] ), .A2(\Table[1][0] ), .A3(\Table[1][2] ), 
        .ZN(n165) );
  NAND3_X1 U132 ( .A1(ADD_CHECK1[0]), .A2(n111), .A3(n110), .ZN(n125) );
  OAI22_X1 U133 ( .A1(n167), .A2(n127), .B1(n165), .B2(n125), .ZN(n113) );
  OAI21_X1 U134 ( .B1(n114), .B2(n113), .A(n112), .ZN(n135) );
  INV_X1 U135 ( .A(n115), .ZN(n160) );
  NOR3_X1 U136 ( .A1(\Table[5][1] ), .A2(\Table[5][0] ), .A3(\Table[5][2] ), 
        .ZN(n158) );
  OAI22_X1 U137 ( .A1(n158), .A2(n125), .B1(n159), .B2(n127), .ZN(n117) );
  OAI21_X1 U138 ( .B1(n118), .B2(n117), .A(n116), .ZN(n134) );
  OAI22_X1 U139 ( .A1(n137), .A2(n124), .B1(n123), .B2(n141), .ZN(n122) );
  NAND3_X1 U140 ( .A1(n25), .A2(n19), .A3(n14), .ZN(n144) );
  INV_X1 U141 ( .A(n144), .ZN(n119) );
  OAI22_X1 U142 ( .A1(n136), .A2(n127), .B1(n119), .B2(n125), .ZN(n121) );
  OAI21_X1 U143 ( .B1(n122), .B2(n121), .A(n120), .ZN(n133) );
  OAI22_X1 U144 ( .A1(n146), .A2(n124), .B1(n123), .B2(n8), .ZN(n131) );
  NAND3_X1 U145 ( .A1(n24), .A2(n18), .A3(n13), .ZN(n152) );
  INV_X1 U146 ( .A(n152), .ZN(n126) );
  OAI22_X1 U147 ( .A1(n145), .A2(n127), .B1(n126), .B2(n125), .ZN(n130) );
  INV_X1 U148 ( .A(n128), .ZN(n129) );
  OAI21_X1 U149 ( .B1(n131), .B2(n130), .A(n129), .ZN(n132) );
  NAND4_X1 U150 ( .A1(n135), .A2(n134), .A3(n133), .A4(n132), .ZN(n181) );
  INV_X1 U151 ( .A(ADD_CHECK2[3]), .ZN(n139) );
  NAND3_X1 U152 ( .A1(n139), .A2(n138), .A3(ADD_CHECK2[0]), .ZN(n164) );
  INV_X1 U153 ( .A(n164), .ZN(n153) );
  NAND3_X1 U154 ( .A1(ADD_CHECK2[0]), .A2(ADD_CHECK2[3]), .A3(ADD_CHECK2[4]), 
        .ZN(n168) );
  NAND3_X1 U155 ( .A1(ADD_CHECK2[3]), .A2(ADD_CHECK2[0]), .A3(n138), .ZN(n166)
         );
  OAI22_X1 U156 ( .A1(n137), .A2(n168), .B1(n166), .B2(n136), .ZN(n143) );
  NAND3_X1 U157 ( .A1(ADD_CHECK2[0]), .A2(ADD_CHECK2[4]), .A3(n139), .ZN(n170)
         );
  NOR3_X1 U158 ( .A1(n139), .A2(n138), .A3(ADD_CHECK2[0]), .ZN(n175) );
  INV_X1 U159 ( .A(n175), .ZN(n147) );
  OAI22_X1 U160 ( .A1(n141), .A2(n170), .B1(n140), .B2(n147), .ZN(n142) );
  AOI211_X1 U161 ( .C1(n153), .C2(n144), .A(n143), .B(n142), .ZN(n157) );
  OAI22_X1 U162 ( .A1(n146), .A2(n168), .B1(n145), .B2(n166), .ZN(n151) );
  OAI22_X1 U163 ( .A1(n8), .A2(n170), .B1(n147), .B2(n148), .ZN(n150) );
  AOI211_X1 U164 ( .C1(n153), .C2(n152), .A(n151), .B(n150), .ZN(n155) );
  OAI22_X1 U165 ( .A1(n157), .A2(n156), .B1(n155), .B2(n154), .ZN(n180) );
  OAI22_X1 U166 ( .A1(n159), .A2(n166), .B1(n158), .B2(n164), .ZN(n162) );
  AOI211_X1 U167 ( .C1(n175), .C2(n163), .A(n162), .B(n161), .ZN(n178) );
  OAI22_X1 U168 ( .A1(n167), .A2(n166), .B1(n165), .B2(n164), .ZN(n173) );
  OAI22_X1 U169 ( .A1(n171), .A2(n170), .B1(n169), .B2(n168), .ZN(n172) );
  AOI211_X1 U170 ( .C1(n175), .C2(n174), .A(n173), .B(n172), .ZN(n176) );
  AOI221_X1 U171 ( .B1(ADD_CHECK2[2]), .B2(n178), .C1(n177), .C2(n176), .A(
        ADD_CHECK2[1]), .ZN(n179) );
  NOR4_X1 U172 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(n183) );
  OAI221_X1 U173 ( .B1(ADD_CHECK2[0]), .B2(n185), .C1(ADD_CHECK2[0]), .C2(n184), .A(n183), .ZN(N192) );
  NAND2_X1 U174 ( .A1(ADD_WR1[3]), .A2(ADD_WR1[4]), .ZN(n371) );
  NOR2_X1 U175 ( .A1(n600), .A2(n371), .ZN(n322) );
  INV_X1 U176 ( .A(ADD_WR1[4]), .ZN(n245) );
  INV_X1 U177 ( .A(ADD_WR2[0]), .ZN(n197) );
  INV_X1 U178 ( .A(ADD_WR1[3]), .ZN(n250) );
  AOI22_X1 U179 ( .A1(n234), .A2(ADD_WR2[1]), .B1(ADD_WR2[3]), .B2(n250), .ZN(
        n186) );
  OAI221_X1 U180 ( .B1(n234), .B2(ADD_WR2[1]), .C1(n250), .C2(ADD_WR2[3]), .A(
        n186), .ZN(n187) );
  AOI221_X1 U181 ( .B1(ADD_WR1[0]), .B2(n197), .C1(n233), .C2(ADD_WR2[0]), .A(
        n187), .ZN(n188) );
  OAI221_X1 U182 ( .B1(ADD_WR1[2]), .B2(n194), .C1(n235), .C2(ADD_WR2[2]), .A(
        n188), .ZN(n189) );
  AOI221_X1 U183 ( .B1(ADD_WR1[4]), .B2(n214), .C1(n245), .C2(ADD_WR2[4]), .A(
        n189), .ZN(n192) );
  INV_X1 U184 ( .A(WR1), .ZN(n190) );
  AOI21_X1 U185 ( .B1(n192), .B2(WR2), .A(n190), .ZN(n598) );
  INV_X1 U186 ( .A(WR2), .ZN(n191) );
  NAND2_X1 U187 ( .A1(ADD_WR2[4]), .A2(ADD_WR2[3]), .ZN(n198) );
  NAND3_X1 U188 ( .A1(ADD_WR2[2]), .A2(ADD_WR2[0]), .A3(ADD_WR2[1]), .ZN(n223)
         );
  NOR2_X1 U189 ( .A1(n198), .A2(n223), .ZN(n365) );
  NAND2_X1 U190 ( .A1(n59), .A2(n365), .ZN(n366) );
  INV_X1 U191 ( .A(n366), .ZN(n193) );
  AOI211_X1 U192 ( .C1(n322), .C2(n598), .A(RST), .B(n193), .ZN(n369) );
  NAND2_X1 U193 ( .A1(n63), .A2(n59), .ZN(n282) );
  INV_X1 U194 ( .A(n282), .ZN(n361) );
  NOR2_X1 U195 ( .A1(ADD_WR2[0]), .A2(ADD_WR2[1]), .ZN(n196) );
  NAND2_X1 U196 ( .A1(n196), .A2(n194), .ZN(n215) );
  NOR2_X1 U197 ( .A1(n198), .A2(n215), .ZN(n438) );
  INV_X1 U198 ( .A(ADD_WR2[1]), .ZN(n195) );
  NAND3_X1 U199 ( .A1(ADD_WR2[0]), .A2(n194), .A3(n195), .ZN(n216) );
  NOR2_X1 U200 ( .A1(n198), .A2(n216), .ZN(n427) );
  AOI22_X1 U201 ( .A1(\Table[24][0] ), .A2(n438), .B1(\Table[25][0] ), .B2(
        n427), .ZN(n202) );
  NAND3_X1 U202 ( .A1(ADD_WR2[1]), .A2(n194), .A3(n197), .ZN(n217) );
  NOR2_X1 U203 ( .A1(n198), .A2(n217), .ZN(n416) );
  NAND3_X1 U204 ( .A1(ADD_WR2[0]), .A2(ADD_WR2[1]), .A3(n194), .ZN(n218) );
  NOR2_X1 U205 ( .A1(n198), .A2(n218), .ZN(n406) );
  AOI22_X1 U206 ( .A1(\Table[26][0] ), .A2(n416), .B1(\Table[27][0] ), .B2(
        n406), .ZN(n201) );
  NAND3_X1 U207 ( .A1(ADD_WR2[0]), .A2(ADD_WR2[2]), .A3(n195), .ZN(n220) );
  NOR2_X1 U208 ( .A1(n198), .A2(n220), .ZN(n387) );
  NAND2_X1 U209 ( .A1(ADD_WR2[2]), .A2(n196), .ZN(n219) );
  NOR2_X1 U210 ( .A1(n198), .A2(n219), .ZN(n396) );
  AOI22_X1 U211 ( .A1(\Table[29][0] ), .A2(n387), .B1(\Table[28][0] ), .B2(
        n396), .ZN(n200) );
  NAND3_X1 U212 ( .A1(ADD_WR2[2]), .A2(ADD_WR2[1]), .A3(n197), .ZN(n221) );
  NOR2_X1 U213 ( .A1(n198), .A2(n221), .ZN(n377) );
  AOI22_X1 U214 ( .A1(\Table[30][0] ), .A2(n377), .B1(\Table[31][0] ), .B2(
        n365), .ZN(n199) );
  NAND4_X1 U215 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(n231) );
  NAND2_X1 U216 ( .A1(ADD_WR2[4]), .A2(n213), .ZN(n203) );
  NOR2_X1 U217 ( .A1(n215), .A2(n203), .ZN(n514) );
  NOR2_X1 U218 ( .A1(n216), .A2(n203), .ZN(n505) );
  AOI22_X1 U219 ( .A1(\Table[16][0] ), .A2(n514), .B1(\Table[17][0] ), .B2(
        n505), .ZN(n207) );
  NOR2_X1 U220 ( .A1(n217), .A2(n203), .ZN(n495) );
  NOR2_X1 U221 ( .A1(n218), .A2(n203), .ZN(n486) );
  AOI22_X1 U222 ( .A1(\Table[18][0] ), .A2(n495), .B1(\Table[19][0] ), .B2(
        n486), .ZN(n206) );
  NOR2_X1 U223 ( .A1(n219), .A2(n203), .ZN(n477) );
  NOR2_X1 U224 ( .A1(n220), .A2(n203), .ZN(n467) );
  AOI22_X1 U225 ( .A1(\Table[20][0] ), .A2(n477), .B1(\Table[21][0] ), .B2(
        n467), .ZN(n205) );
  NOR2_X1 U226 ( .A1(n221), .A2(n203), .ZN(n459) );
  NOR2_X1 U227 ( .A1(n223), .A2(n203), .ZN(n449) );
  AOI22_X1 U228 ( .A1(\Table[22][0] ), .A2(n459), .B1(\Table[23][0] ), .B2(
        n449), .ZN(n204) );
  NAND4_X1 U229 ( .A1(n207), .A2(n206), .A3(n205), .A4(n204), .ZN(n230) );
  NAND2_X1 U230 ( .A1(ADD_WR2[3]), .A2(n214), .ZN(n208) );
  NOR2_X1 U231 ( .A1(n215), .A2(n208), .ZN(n592) );
  NOR2_X1 U232 ( .A1(n216), .A2(n208), .ZN(n582) );
  AOI22_X1 U233 ( .A1(\Table[8][0] ), .A2(n592), .B1(\Table[9][0] ), .B2(n582), 
        .ZN(n212) );
  NOR2_X1 U234 ( .A1(n217), .A2(n208), .ZN(n574) );
  NOR2_X1 U235 ( .A1(n218), .A2(n208), .ZN(n564) );
  AOI22_X1 U236 ( .A1(\Table[10][0] ), .A2(n574), .B1(\Table[11][0] ), .B2(
        n564), .ZN(n211) );
  NOR2_X1 U237 ( .A1(n219), .A2(n208), .ZN(n554) );
  NOR2_X1 U238 ( .A1(n220), .A2(n208), .ZN(n544) );
  AOI22_X1 U239 ( .A1(\Table[12][0] ), .A2(n554), .B1(\Table[13][0] ), .B2(
        n544), .ZN(n210) );
  NOR2_X1 U240 ( .A1(n221), .A2(n208), .ZN(n534) );
  NOR2_X1 U241 ( .A1(n223), .A2(n208), .ZN(n524) );
  AOI22_X1 U242 ( .A1(\Table[14][0] ), .A2(n534), .B1(\Table[15][0] ), .B2(
        n524), .ZN(n209) );
  NAND4_X1 U243 ( .A1(n212), .A2(n211), .A3(n210), .A4(n209), .ZN(n229) );
  NAND2_X1 U244 ( .A1(n214), .A2(n213), .ZN(n222) );
  NOR2_X1 U245 ( .A1(n215), .A2(n222), .ZN(n666) );
  NOR2_X1 U246 ( .A1(n216), .A2(n222), .ZN(n651) );
  AOI22_X1 U247 ( .A1(\Table[0][0] ), .A2(n666), .B1(\Table[1][0] ), .B2(n651), 
        .ZN(n227) );
  NOR2_X1 U248 ( .A1(n217), .A2(n222), .ZN(n643) );
  NOR2_X1 U249 ( .A1(n218), .A2(n222), .ZN(n635) );
  AOI22_X1 U250 ( .A1(\Table[2][0] ), .A2(n643), .B1(\Table[3][0] ), .B2(n635), 
        .ZN(n226) );
  NOR2_X1 U251 ( .A1(n219), .A2(n222), .ZN(n627) );
  NOR2_X1 U252 ( .A1(n220), .A2(n222), .ZN(n619) );
  AOI22_X1 U253 ( .A1(\Table[4][0] ), .A2(n627), .B1(\Table[5][0] ), .B2(n619), 
        .ZN(n225) );
  NOR2_X1 U254 ( .A1(n221), .A2(n222), .ZN(n611) );
  NOR2_X1 U255 ( .A1(n223), .A2(n222), .ZN(n603) );
  AOI22_X1 U256 ( .A1(\Table[6][0] ), .A2(n611), .B1(\Table[7][0] ), .B2(n603), 
        .ZN(n224) );
  NAND4_X1 U257 ( .A1(n227), .A2(n226), .A3(n225), .A4(n224), .ZN(n228) );
  NOR4_X1 U258 ( .A1(n231), .A2(n230), .A3(n229), .A4(n228), .ZN(n284) );
  NAND2_X1 U259 ( .A1(ADD_WR1[2]), .A2(ADD_WR1[0]), .ZN(n232) );
  AOI22_X1 U260 ( .A1(n433), .A2(\Table[24][0] ), .B1(n422), .B2(
        \Table[25][0] ), .ZN(n238) );
  AOI22_X1 U261 ( .A1(n411), .A2(\Table[26][0] ), .B1(n402), .B2(
        \Table[27][0] ), .ZN(n237) );
  AOI22_X1 U262 ( .A1(n393), .A2(\Table[28][0] ), .B1(n370), .B2(
        \Table[30][0] ), .ZN(n236) );
  NAND3_X1 U263 ( .A1(n238), .A2(n237), .A3(n236), .ZN(n239) );
  AOI21_X1 U264 ( .B1(n382), .B2(\Table[29][0] ), .A(n239), .ZN(n259) );
  NOR2_X1 U265 ( .A1(ADD_WR1[3]), .A2(ADD_WR1[4]), .ZN(n599) );
  AOI22_X1 U266 ( .A1(n433), .A2(\Table[0][0] ), .B1(n422), .B2(\Table[1][0] ), 
        .ZN(n243) );
  AOI22_X1 U267 ( .A1(n411), .A2(\Table[2][0] ), .B1(n402), .B2(\Table[3][0] ), 
        .ZN(n242) );
  AOI22_X1 U268 ( .A1(n393), .A2(\Table[4][0] ), .B1(n382), .B2(\Table[5][0] ), 
        .ZN(n241) );
  AOI22_X1 U269 ( .A1(n370), .A2(\Table[6][0] ), .B1(n328), .B2(\Table[7][0] ), 
        .ZN(n240) );
  NAND4_X1 U270 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(n244) );
  AOI22_X1 U271 ( .A1(n599), .A2(n244), .B1(n322), .B2(\Table[31][0] ), .ZN(
        n258) );
  NOR2_X1 U272 ( .A1(ADD_WR1[3]), .A2(n245), .ZN(n444) );
  AOI22_X1 U273 ( .A1(n433), .A2(\Table[16][0] ), .B1(n422), .B2(
        \Table[17][0] ), .ZN(n249) );
  AOI22_X1 U274 ( .A1(n411), .A2(\Table[18][0] ), .B1(n402), .B2(
        \Table[19][0] ), .ZN(n248) );
  AOI22_X1 U275 ( .A1(n393), .A2(\Table[20][0] ), .B1(n382), .B2(
        \Table[21][0] ), .ZN(n247) );
  AOI22_X1 U276 ( .A1(n370), .A2(\Table[22][0] ), .B1(n328), .B2(
        \Table[23][0] ), .ZN(n246) );
  NAND4_X1 U277 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(n256) );
  NOR2_X1 U278 ( .A1(ADD_WR1[4]), .A2(n250), .ZN(n519) );
  AOI22_X1 U279 ( .A1(n433), .A2(\Table[8][0] ), .B1(n422), .B2(\Table[9][0] ), 
        .ZN(n254) );
  AOI22_X1 U280 ( .A1(n411), .A2(\Table[10][0] ), .B1(n402), .B2(
        \Table[11][0] ), .ZN(n253) );
  AOI22_X1 U281 ( .A1(n393), .A2(\Table[12][0] ), .B1(n382), .B2(
        \Table[13][0] ), .ZN(n252) );
  AOI22_X1 U282 ( .A1(n370), .A2(\Table[14][0] ), .B1(n328), .B2(
        \Table[15][0] ), .ZN(n251) );
  NAND4_X1 U283 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(n255) );
  AOI22_X1 U284 ( .A1(n444), .A2(n256), .B1(n519), .B2(n255), .ZN(n257) );
  OAI211_X1 U285 ( .C1(n259), .C2(n371), .A(n258), .B(n257), .ZN(n308) );
  AOI22_X1 U286 ( .A1(n365), .A2(n660), .B1(n60), .B2(n366), .ZN(n260) );
  INV_X1 U287 ( .A(n369), .ZN(n311) );
  AOI22_X1 U288 ( .A1(n369), .A2(n261), .B1(n260), .B2(n311), .ZN(n797) );
  AOI22_X1 U289 ( .A1(\Table[24][1] ), .A2(n438), .B1(\Table[25][1] ), .B2(
        n427), .ZN(n265) );
  AOI22_X1 U290 ( .A1(\Table[26][1] ), .A2(n416), .B1(\Table[27][1] ), .B2(
        n406), .ZN(n264) );
  AOI22_X1 U291 ( .A1(\Table[29][1] ), .A2(n387), .B1(\Table[28][1] ), .B2(
        n396), .ZN(n263) );
  AOI22_X1 U292 ( .A1(\Table[30][1] ), .A2(n377), .B1(\Table[31][1] ), .B2(
        n365), .ZN(n262) );
  NAND4_X1 U293 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(n281) );
  AOI22_X1 U294 ( .A1(\Table[16][1] ), .A2(n514), .B1(\Table[17][1] ), .B2(
        n505), .ZN(n269) );
  AOI22_X1 U295 ( .A1(\Table[18][1] ), .A2(n495), .B1(\Table[19][1] ), .B2(
        n486), .ZN(n268) );
  AOI22_X1 U296 ( .A1(\Table[20][1] ), .A2(n477), .B1(\Table[21][1] ), .B2(
        n467), .ZN(n267) );
  AOI22_X1 U297 ( .A1(\Table[22][1] ), .A2(n459), .B1(\Table[23][1] ), .B2(
        n449), .ZN(n266) );
  NAND4_X1 U298 ( .A1(n269), .A2(n268), .A3(n267), .A4(n266), .ZN(n280) );
  AOI22_X1 U299 ( .A1(\Table[8][1] ), .A2(n592), .B1(\Table[9][1] ), .B2(n582), 
        .ZN(n273) );
  AOI22_X1 U300 ( .A1(\Table[10][1] ), .A2(n574), .B1(\Table[11][1] ), .B2(
        n564), .ZN(n272) );
  AOI22_X1 U301 ( .A1(\Table[12][1] ), .A2(n554), .B1(\Table[13][1] ), .B2(
        n544), .ZN(n271) );
  AOI22_X1 U302 ( .A1(\Table[14][1] ), .A2(n534), .B1(\Table[15][1] ), .B2(
        n524), .ZN(n270) );
  NAND4_X1 U303 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .ZN(n279) );
  AOI22_X1 U304 ( .A1(\Table[0][1] ), .A2(n666), .B1(\Table[1][1] ), .B2(n651), 
        .ZN(n277) );
  AOI22_X1 U305 ( .A1(\Table[2][1] ), .A2(n643), .B1(\Table[3][1] ), .B2(n635), 
        .ZN(n276) );
  AOI22_X1 U306 ( .A1(\Table[4][1] ), .A2(n627), .B1(\Table[5][1] ), .B2(n619), 
        .ZN(n275) );
  AOI22_X1 U307 ( .A1(\Table[6][1] ), .A2(n611), .B1(\Table[7][1] ), .B2(n603), 
        .ZN(n274) );
  NAND4_X1 U308 ( .A1(n277), .A2(n276), .A3(n275), .A4(n274), .ZN(n278) );
  NOR4_X1 U309 ( .A1(n281), .A2(n280), .A3(n279), .A4(n278), .ZN(n283) );
  NAND2_X1 U310 ( .A1(n283), .A2(n284), .ZN(n363) );
  AOI221_X1 U311 ( .B1(n284), .B2(n363), .C1(n283), .C2(n363), .A(n282), .ZN(
        n663) );
  AOI22_X1 U312 ( .A1(n433), .A2(\Table[24][1] ), .B1(n422), .B2(
        \Table[25][1] ), .ZN(n287) );
  AOI22_X1 U313 ( .A1(n411), .A2(\Table[26][1] ), .B1(n402), .B2(
        \Table[27][1] ), .ZN(n286) );
  AOI22_X1 U314 ( .A1(n393), .A2(\Table[28][1] ), .B1(n370), .B2(
        \Table[30][1] ), .ZN(n285) );
  NAND3_X1 U315 ( .A1(n287), .A2(n286), .A3(n285), .ZN(n288) );
  AOI21_X1 U316 ( .B1(n382), .B2(\Table[29][1] ), .A(n288), .ZN(n306) );
  AOI22_X1 U317 ( .A1(n433), .A2(\Table[0][1] ), .B1(n422), .B2(\Table[1][1] ), 
        .ZN(n292) );
  AOI22_X1 U318 ( .A1(n411), .A2(\Table[2][1] ), .B1(n402), .B2(\Table[3][1] ), 
        .ZN(n291) );
  AOI22_X1 U319 ( .A1(n393), .A2(\Table[4][1] ), .B1(n382), .B2(\Table[5][1] ), 
        .ZN(n290) );
  AOI22_X1 U320 ( .A1(n370), .A2(\Table[6][1] ), .B1(n328), .B2(\Table[7][1] ), 
        .ZN(n289) );
  NAND4_X1 U321 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(n293) );
  AOI22_X1 U322 ( .A1(\Table[31][1] ), .A2(n322), .B1(n599), .B2(n293), .ZN(
        n305) );
  AOI22_X1 U323 ( .A1(n433), .A2(\Table[8][1] ), .B1(n422), .B2(\Table[9][1] ), 
        .ZN(n297) );
  AOI22_X1 U324 ( .A1(n411), .A2(\Table[10][1] ), .B1(n402), .B2(
        \Table[11][1] ), .ZN(n296) );
  AOI22_X1 U325 ( .A1(n393), .A2(\Table[12][1] ), .B1(n382), .B2(
        \Table[13][1] ), .ZN(n295) );
  AOI22_X1 U326 ( .A1(n370), .A2(\Table[14][1] ), .B1(n328), .B2(
        \Table[15][1] ), .ZN(n294) );
  NAND4_X1 U327 ( .A1(n297), .A2(n296), .A3(n295), .A4(n294), .ZN(n303) );
  AOI22_X1 U328 ( .A1(n433), .A2(\Table[16][1] ), .B1(n422), .B2(
        \Table[17][1] ), .ZN(n301) );
  AOI22_X1 U329 ( .A1(n411), .A2(\Table[18][1] ), .B1(n402), .B2(
        \Table[19][1] ), .ZN(n300) );
  AOI22_X1 U330 ( .A1(n393), .A2(\Table[20][1] ), .B1(n382), .B2(
        \Table[21][1] ), .ZN(n299) );
  AOI22_X1 U331 ( .A1(n370), .A2(\Table[22][1] ), .B1(n328), .B2(
        \Table[23][1] ), .ZN(n298) );
  NAND4_X1 U332 ( .A1(n301), .A2(n300), .A3(n299), .A4(n298), .ZN(n302) );
  AOI22_X1 U333 ( .A1(n519), .A2(n303), .B1(n444), .B2(n302), .ZN(n304) );
  OAI211_X1 U334 ( .C1(n306), .C2(n371), .A(n305), .B(n304), .ZN(n307) );
  INV_X1 U335 ( .A(n307), .ZN(n310) );
  INV_X1 U336 ( .A(n308), .ZN(n309) );
  NOR2_X1 U337 ( .A1(n310), .A2(n309), .ZN(n340) );
  AOI211_X1 U338 ( .C1(n310), .C2(n309), .A(RST), .B(n340), .ZN(n662) );
  AOI22_X1 U339 ( .A1(n365), .A2(n2), .B1(n4), .B2(n366), .ZN(n312) );
  AOI22_X1 U340 ( .A1(n369), .A2(n313), .B1(n312), .B2(n311), .ZN(n796) );
  AOI22_X1 U341 ( .A1(n433), .A2(\Table[24][2] ), .B1(n422), .B2(
        \Table[25][2] ), .ZN(n316) );
  AOI22_X1 U342 ( .A1(n411), .A2(\Table[26][2] ), .B1(n402), .B2(
        \Table[27][2] ), .ZN(n315) );
  AOI22_X1 U343 ( .A1(n393), .A2(\Table[28][2] ), .B1(n370), .B2(
        \Table[30][2] ), .ZN(n314) );
  NAND3_X1 U344 ( .A1(n316), .A2(n315), .A3(n314), .ZN(n317) );
  AOI21_X1 U345 ( .B1(n382), .B2(\Table[29][2] ), .A(n317), .ZN(n337) );
  AOI22_X1 U346 ( .A1(n433), .A2(\Table[0][2] ), .B1(n422), .B2(\Table[1][2] ), 
        .ZN(n321) );
  AOI22_X1 U347 ( .A1(n411), .A2(\Table[2][2] ), .B1(n402), .B2(\Table[3][2] ), 
        .ZN(n320) );
  AOI22_X1 U348 ( .A1(n393), .A2(\Table[4][2] ), .B1(n382), .B2(\Table[5][2] ), 
        .ZN(n319) );
  AOI22_X1 U349 ( .A1(n370), .A2(\Table[6][2] ), .B1(n328), .B2(\Table[7][2] ), 
        .ZN(n318) );
  NAND4_X1 U350 ( .A1(n321), .A2(n320), .A3(n319), .A4(n318), .ZN(n323) );
  AOI22_X1 U351 ( .A1(n599), .A2(n323), .B1(n322), .B2(\Table[31][2] ), .ZN(
        n336) );
  AOI22_X1 U352 ( .A1(n433), .A2(\Table[16][2] ), .B1(n422), .B2(
        \Table[17][2] ), .ZN(n327) );
  AOI22_X1 U353 ( .A1(n411), .A2(\Table[18][2] ), .B1(n402), .B2(
        \Table[19][2] ), .ZN(n326) );
  AOI22_X1 U354 ( .A1(n393), .A2(\Table[20][2] ), .B1(n382), .B2(
        \Table[21][2] ), .ZN(n325) );
  AOI22_X1 U355 ( .A1(n370), .A2(\Table[22][2] ), .B1(n328), .B2(
        \Table[23][2] ), .ZN(n324) );
  NAND4_X1 U356 ( .A1(n327), .A2(n326), .A3(n325), .A4(n324), .ZN(n334) );
  AOI22_X1 U357 ( .A1(n433), .A2(\Table[8][2] ), .B1(n422), .B2(\Table[9][2] ), 
        .ZN(n332) );
  AOI22_X1 U358 ( .A1(n411), .A2(\Table[10][2] ), .B1(n402), .B2(
        \Table[11][2] ), .ZN(n331) );
  AOI22_X1 U359 ( .A1(n393), .A2(\Table[12][2] ), .B1(n382), .B2(
        \Table[13][2] ), .ZN(n330) );
  AOI22_X1 U360 ( .A1(n370), .A2(\Table[14][2] ), .B1(n328), .B2(
        \Table[15][2] ), .ZN(n329) );
  NAND4_X1 U361 ( .A1(n332), .A2(n331), .A3(n330), .A4(n329), .ZN(n333) );
  AOI22_X1 U362 ( .A1(n444), .A2(n334), .B1(n519), .B2(n333), .ZN(n335) );
  OAI211_X1 U363 ( .C1(n337), .C2(n371), .A(n336), .B(n335), .ZN(n339) );
  NOR2_X1 U364 ( .A1(n340), .A2(n339), .ZN(n338) );
  AOI211_X1 U365 ( .C1(n340), .C2(n339), .A(RST), .B(n338), .ZN(n668) );
  AOI22_X1 U366 ( .A1(\Table[24][2] ), .A2(n438), .B1(\Table[25][2] ), .B2(
        n427), .ZN(n344) );
  AOI22_X1 U367 ( .A1(\Table[26][2] ), .A2(n416), .B1(\Table[27][2] ), .B2(
        n406), .ZN(n343) );
  AOI22_X1 U368 ( .A1(\Table[29][2] ), .A2(n387), .B1(\Table[28][2] ), .B2(
        n396), .ZN(n342) );
  AOI22_X1 U369 ( .A1(\Table[30][2] ), .A2(n377), .B1(\Table[31][2] ), .B2(
        n365), .ZN(n341) );
  NAND4_X1 U370 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .ZN(n360) );
  AOI22_X1 U371 ( .A1(\Table[16][2] ), .A2(n514), .B1(\Table[17][2] ), .B2(
        n505), .ZN(n348) );
  AOI22_X1 U372 ( .A1(\Table[18][2] ), .A2(n495), .B1(\Table[19][2] ), .B2(
        n486), .ZN(n347) );
  AOI22_X1 U373 ( .A1(\Table[20][2] ), .A2(n477), .B1(\Table[21][2] ), .B2(
        n467), .ZN(n346) );
  AOI22_X1 U374 ( .A1(\Table[22][2] ), .A2(n459), .B1(\Table[23][2] ), .B2(
        n449), .ZN(n345) );
  NAND4_X1 U375 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .ZN(n359) );
  AOI22_X1 U376 ( .A1(\Table[8][2] ), .A2(n592), .B1(\Table[9][2] ), .B2(n582), 
        .ZN(n352) );
  AOI22_X1 U377 ( .A1(\Table[10][2] ), .A2(n574), .B1(\Table[11][2] ), .B2(
        n564), .ZN(n351) );
  AOI22_X1 U378 ( .A1(\Table[12][2] ), .A2(n554), .B1(\Table[13][2] ), .B2(
        n544), .ZN(n350) );
  AOI22_X1 U379 ( .A1(\Table[14][2] ), .A2(n534), .B1(\Table[15][2] ), .B2(
        n524), .ZN(n349) );
  NAND4_X1 U380 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .ZN(n358) );
  AOI22_X1 U381 ( .A1(\Table[0][2] ), .A2(n666), .B1(\Table[1][2] ), .B2(n651), 
        .ZN(n356) );
  AOI22_X1 U382 ( .A1(\Table[2][2] ), .A2(n643), .B1(\Table[3][2] ), .B2(n635), 
        .ZN(n355) );
  AOI22_X1 U383 ( .A1(\Table[4][2] ), .A2(n627), .B1(\Table[5][2] ), .B2(n619), 
        .ZN(n354) );
  AOI22_X1 U384 ( .A1(\Table[6][2] ), .A2(n611), .B1(\Table[7][2] ), .B2(n603), 
        .ZN(n353) );
  NAND4_X1 U385 ( .A1(n356), .A2(n355), .A3(n354), .A4(n353), .ZN(n357) );
  NOR4_X1 U386 ( .A1(n360), .A2(n359), .A3(n358), .A4(n357), .ZN(n364) );
  OAI21_X1 U387 ( .B1(n364), .B2(n363), .A(n361), .ZN(n362) );
  AOI22_X1 U388 ( .A1(n3), .A2(n366), .B1(n365), .B2(n61), .ZN(n368) );
  NAND2_X1 U389 ( .A1(n369), .A2(\Table[31][2] ), .ZN(n367) );
  OAI21_X1 U390 ( .B1(n369), .B2(n368), .A(n367), .ZN(n795) );
  INV_X1 U391 ( .A(n371), .ZN(n372) );
  NAND2_X1 U392 ( .A1(n372), .A2(n598), .ZN(n434) );
  NAND2_X1 U393 ( .A1(n656), .A2(n377), .ZN(n378) );
  OAI211_X1 U394 ( .C1(n608), .C2(n434), .A(n62), .B(n378), .ZN(n379) );
  INV_X1 U395 ( .A(n379), .ZN(n381) );
  AOI22_X1 U396 ( .A1(n377), .A2(n660), .B1(n60), .B2(n378), .ZN(n373) );
  AOI22_X1 U397 ( .A1(n381), .A2(n374), .B1(n373), .B2(n379), .ZN(n794) );
  AOI22_X1 U398 ( .A1(n377), .A2(n2), .B1(n4), .B2(n378), .ZN(n375) );
  AOI22_X1 U399 ( .A1(n381), .A2(n376), .B1(n375), .B2(n379), .ZN(n793) );
  AOI22_X1 U400 ( .A1(n3), .A2(n378), .B1(n377), .B2(n61), .ZN(n380) );
  AOI22_X1 U401 ( .A1(n381), .A2(n54), .B1(n380), .B2(n379), .ZN(n792) );
  NAND2_X1 U402 ( .A1(n656), .A2(n387), .ZN(n388) );
  OAI211_X1 U403 ( .C1(n616), .C2(n434), .A(n63), .B(n388), .ZN(n389) );
  INV_X1 U404 ( .A(n389), .ZN(n392) );
  AOI22_X1 U405 ( .A1(n387), .A2(n660), .B1(n60), .B2(n388), .ZN(n383) );
  AOI22_X1 U406 ( .A1(n392), .A2(n384), .B1(n383), .B2(n389), .ZN(n791) );
  AOI22_X1 U407 ( .A1(n387), .A2(n2), .B1(n4), .B2(n388), .ZN(n385) );
  AOI22_X1 U408 ( .A1(n392), .A2(n386), .B1(n385), .B2(n389), .ZN(n790) );
  AOI22_X1 U409 ( .A1(n3), .A2(n388), .B1(n387), .B2(n61), .ZN(n390) );
  AOI22_X1 U410 ( .A1(n392), .A2(n391), .B1(n390), .B2(n389), .ZN(n789) );
  NAND2_X1 U411 ( .A1(n656), .A2(n396), .ZN(n397) );
  OAI211_X1 U412 ( .C1(n624), .C2(n434), .A(n62), .B(n397), .ZN(n398) );
  INV_X1 U413 ( .A(n398), .ZN(n401) );
  AOI22_X1 U414 ( .A1(n396), .A2(n660), .B1(n60), .B2(n397), .ZN(n394) );
  AOI22_X1 U415 ( .A1(n401), .A2(n15), .B1(n394), .B2(n398), .ZN(n788) );
  AOI22_X1 U416 ( .A1(n396), .A2(n2), .B1(n4), .B2(n397), .ZN(n395) );
  AOI22_X1 U417 ( .A1(n401), .A2(n21), .B1(n395), .B2(n398), .ZN(n787) );
  AOI22_X1 U418 ( .A1(n3), .A2(n397), .B1(n396), .B2(n61), .ZN(n399) );
  AOI22_X1 U419 ( .A1(n401), .A2(n400), .B1(n399), .B2(n398), .ZN(n786) );
  NAND2_X1 U420 ( .A1(n656), .A2(n406), .ZN(n407) );
  OAI211_X1 U421 ( .C1(n632), .C2(n434), .A(n63), .B(n407), .ZN(n408) );
  INV_X1 U422 ( .A(n408), .ZN(n410) );
  AOI22_X1 U423 ( .A1(n406), .A2(n660), .B1(n60), .B2(n407), .ZN(n403) );
  AOI22_X1 U424 ( .A1(n410), .A2(n52), .B1(n403), .B2(n408), .ZN(n785) );
  AOI22_X1 U425 ( .A1(n406), .A2(n2), .B1(n4), .B2(n407), .ZN(n404) );
  AOI22_X1 U426 ( .A1(n410), .A2(n405), .B1(n404), .B2(n408), .ZN(n784) );
  AOI22_X1 U427 ( .A1(n3), .A2(n407), .B1(n406), .B2(n61), .ZN(n409) );
  AOI22_X1 U428 ( .A1(n410), .A2(n53), .B1(n409), .B2(n408), .ZN(n783) );
  NAND2_X1 U429 ( .A1(n656), .A2(n416), .ZN(n417) );
  OAI211_X1 U430 ( .C1(n640), .C2(n434), .A(n62), .B(n417), .ZN(n418) );
  INV_X1 U431 ( .A(n418), .ZN(n421) );
  AOI22_X1 U432 ( .A1(n416), .A2(n660), .B1(n60), .B2(n417), .ZN(n412) );
  AOI22_X1 U433 ( .A1(n421), .A2(n413), .B1(n412), .B2(n418), .ZN(n782) );
  AOI22_X1 U434 ( .A1(n416), .A2(n2), .B1(n4), .B2(n417), .ZN(n414) );
  AOI22_X1 U435 ( .A1(n421), .A2(n415), .B1(n414), .B2(n418), .ZN(n781) );
  AOI22_X1 U436 ( .A1(n3), .A2(n417), .B1(n416), .B2(n61), .ZN(n419) );
  AOI22_X1 U437 ( .A1(n421), .A2(n420), .B1(n419), .B2(n418), .ZN(n780) );
  NAND2_X1 U438 ( .A1(n656), .A2(n427), .ZN(n428) );
  OAI211_X1 U439 ( .C1(n648), .C2(n434), .A(n63), .B(n428), .ZN(n429) );
  INV_X1 U440 ( .A(n429), .ZN(n432) );
  AOI22_X1 U441 ( .A1(n427), .A2(n660), .B1(n60), .B2(n428), .ZN(n423) );
  AOI22_X1 U442 ( .A1(n432), .A2(n424), .B1(n423), .B2(n429), .ZN(n779) );
  AOI22_X1 U443 ( .A1(n427), .A2(n2), .B1(n4), .B2(n428), .ZN(n425) );
  AOI22_X1 U444 ( .A1(n432), .A2(n426), .B1(n425), .B2(n429), .ZN(n778) );
  AOI22_X1 U445 ( .A1(n3), .A2(n428), .B1(n427), .B2(n61), .ZN(n430) );
  AOI22_X1 U446 ( .A1(n432), .A2(n431), .B1(n430), .B2(n429), .ZN(n777) );
  NAND2_X1 U447 ( .A1(n656), .A2(n438), .ZN(n439) );
  OAI211_X1 U448 ( .C1(n658), .C2(n434), .A(n62), .B(n439), .ZN(n440) );
  INV_X1 U449 ( .A(n440), .ZN(n443) );
  AOI22_X1 U450 ( .A1(n438), .A2(n660), .B1(n60), .B2(n439), .ZN(n435) );
  AOI22_X1 U451 ( .A1(n443), .A2(n20), .B1(n435), .B2(n440), .ZN(n776) );
  AOI22_X1 U452 ( .A1(n438), .A2(n2), .B1(n4), .B2(n439), .ZN(n436) );
  AOI22_X1 U453 ( .A1(n443), .A2(n437), .B1(n436), .B2(n440), .ZN(n775) );
  AOI22_X1 U454 ( .A1(n3), .A2(n439), .B1(n438), .B2(n665), .ZN(n441) );
  AOI22_X1 U455 ( .A1(n443), .A2(n442), .B1(n441), .B2(n440), .ZN(n774) );
  NAND2_X1 U456 ( .A1(n444), .A2(n598), .ZN(n511) );
  NAND2_X1 U457 ( .A1(n59), .A2(n449), .ZN(n450) );
  OAI211_X1 U458 ( .C1(n600), .C2(n511), .A(n63), .B(n450), .ZN(n451) );
  INV_X1 U459 ( .A(n451), .ZN(n454) );
  AOI22_X1 U460 ( .A1(n449), .A2(n660), .B1(n60), .B2(n450), .ZN(n445) );
  AOI22_X1 U461 ( .A1(n454), .A2(n446), .B1(n445), .B2(n451), .ZN(n773) );
  AOI22_X1 U462 ( .A1(n449), .A2(n2), .B1(n4), .B2(n450), .ZN(n447) );
  AOI22_X1 U463 ( .A1(n454), .A2(n448), .B1(n447), .B2(n451), .ZN(n772) );
  AOI22_X1 U464 ( .A1(n3), .A2(n450), .B1(n449), .B2(n61), .ZN(n452) );
  AOI22_X1 U465 ( .A1(n454), .A2(n453), .B1(n452), .B2(n451), .ZN(n771) );
  NAND2_X1 U466 ( .A1(n656), .A2(n459), .ZN(n460) );
  OAI211_X1 U467 ( .C1(n608), .C2(n511), .A(n62), .B(n460), .ZN(n461) );
  INV_X1 U468 ( .A(n461), .ZN(n464) );
  AOI22_X1 U469 ( .A1(n459), .A2(n660), .B1(n60), .B2(n460), .ZN(n455) );
  AOI22_X1 U470 ( .A1(n464), .A2(n456), .B1(n455), .B2(n461), .ZN(n770) );
  AOI22_X1 U471 ( .A1(n459), .A2(n2), .B1(n4), .B2(n460), .ZN(n457) );
  AOI22_X1 U472 ( .A1(n464), .A2(n458), .B1(n457), .B2(n461), .ZN(n769) );
  AOI22_X1 U473 ( .A1(n3), .A2(n460), .B1(n459), .B2(n61), .ZN(n462) );
  AOI22_X1 U474 ( .A1(n464), .A2(n463), .B1(n462), .B2(n461), .ZN(n768) );
  NAND2_X1 U475 ( .A1(n59), .A2(n467), .ZN(n468) );
  OAI211_X1 U476 ( .C1(n616), .C2(n511), .A(n63), .B(n468), .ZN(n469) );
  INV_X1 U477 ( .A(n469), .ZN(n472) );
  AOI22_X1 U478 ( .A1(n467), .A2(n660), .B1(n60), .B2(n468), .ZN(n465) );
  AOI22_X1 U479 ( .A1(n472), .A2(n16), .B1(n465), .B2(n469), .ZN(n767) );
  AOI22_X1 U480 ( .A1(n467), .A2(n2), .B1(n4), .B2(n468), .ZN(n466) );
  AOI22_X1 U481 ( .A1(n472), .A2(n22), .B1(n466), .B2(n469), .ZN(n766) );
  AOI22_X1 U482 ( .A1(n3), .A2(n468), .B1(n467), .B2(n61), .ZN(n470) );
  AOI22_X1 U483 ( .A1(n472), .A2(n471), .B1(n470), .B2(n469), .ZN(n765) );
  NAND2_X1 U484 ( .A1(n59), .A2(n477), .ZN(n478) );
  OAI211_X1 U485 ( .C1(n624), .C2(n511), .A(n63), .B(n478), .ZN(n479) );
  INV_X1 U486 ( .A(n479), .ZN(n482) );
  AOI22_X1 U487 ( .A1(n477), .A2(n660), .B1(n60), .B2(n478), .ZN(n473) );
  AOI22_X1 U488 ( .A1(n482), .A2(n474), .B1(n473), .B2(n479), .ZN(n764) );
  AOI22_X1 U489 ( .A1(n477), .A2(n2), .B1(n4), .B2(n478), .ZN(n475) );
  AOI22_X1 U490 ( .A1(n482), .A2(n476), .B1(n475), .B2(n479), .ZN(n763) );
  AOI22_X1 U491 ( .A1(n3), .A2(n478), .B1(n477), .B2(n61), .ZN(n480) );
  AOI22_X1 U492 ( .A1(n482), .A2(n481), .B1(n480), .B2(n479), .ZN(n762) );
  NAND2_X1 U493 ( .A1(n59), .A2(n486), .ZN(n487) );
  OAI211_X1 U494 ( .C1(n632), .C2(n511), .A(n63), .B(n487), .ZN(n488) );
  INV_X1 U495 ( .A(n488), .ZN(n490) );
  AOI22_X1 U496 ( .A1(n486), .A2(n660), .B1(n60), .B2(n487), .ZN(n483) );
  AOI22_X1 U497 ( .A1(n490), .A2(n50), .B1(n483), .B2(n488), .ZN(n761) );
  AOI22_X1 U498 ( .A1(n486), .A2(n2), .B1(n4), .B2(n487), .ZN(n484) );
  AOI22_X1 U499 ( .A1(n490), .A2(n485), .B1(n484), .B2(n488), .ZN(n760) );
  AOI22_X1 U500 ( .A1(n3), .A2(n487), .B1(n486), .B2(n61), .ZN(n489) );
  AOI22_X1 U501 ( .A1(n490), .A2(n51), .B1(n489), .B2(n488), .ZN(n759) );
  NAND2_X1 U502 ( .A1(n59), .A2(n495), .ZN(n496) );
  OAI211_X1 U503 ( .C1(n640), .C2(n511), .A(n63), .B(n496), .ZN(n497) );
  INV_X1 U504 ( .A(n497), .ZN(n500) );
  AOI22_X1 U505 ( .A1(n495), .A2(n660), .B1(n60), .B2(n496), .ZN(n491) );
  AOI22_X1 U506 ( .A1(n500), .A2(n492), .B1(n491), .B2(n497), .ZN(n758) );
  AOI22_X1 U507 ( .A1(n495), .A2(n2), .B1(n4), .B2(n496), .ZN(n493) );
  AOI22_X1 U508 ( .A1(n500), .A2(n494), .B1(n493), .B2(n497), .ZN(n757) );
  AOI22_X1 U509 ( .A1(n3), .A2(n496), .B1(n495), .B2(n61), .ZN(n498) );
  AOI22_X1 U510 ( .A1(n500), .A2(n499), .B1(n498), .B2(n497), .ZN(n756) );
  NAND2_X1 U511 ( .A1(n59), .A2(n505), .ZN(n506) );
  OAI211_X1 U512 ( .C1(n648), .C2(n511), .A(n63), .B(n506), .ZN(n507) );
  INV_X1 U513 ( .A(n507), .ZN(n510) );
  AOI22_X1 U514 ( .A1(n505), .A2(n660), .B1(n60), .B2(n506), .ZN(n501) );
  AOI22_X1 U515 ( .A1(n510), .A2(n502), .B1(n501), .B2(n507), .ZN(n755) );
  AOI22_X1 U516 ( .A1(n505), .A2(n2), .B1(n4), .B2(n506), .ZN(n503) );
  AOI22_X1 U517 ( .A1(n510), .A2(n504), .B1(n503), .B2(n507), .ZN(n754) );
  AOI22_X1 U518 ( .A1(n3), .A2(n506), .B1(n505), .B2(n61), .ZN(n508) );
  AOI22_X1 U519 ( .A1(n510), .A2(n509), .B1(n508), .B2(n507), .ZN(n753) );
  NAND2_X1 U520 ( .A1(n656), .A2(n514), .ZN(n515) );
  OAI211_X1 U521 ( .C1(n658), .C2(n511), .A(n63), .B(n515), .ZN(n516) );
  INV_X1 U522 ( .A(n516), .ZN(n518) );
  AOI22_X1 U523 ( .A1(n514), .A2(n660), .B1(n659), .B2(n515), .ZN(n512) );
  AOI22_X1 U524 ( .A1(n518), .A2(n48), .B1(n512), .B2(n516), .ZN(n752) );
  AOI22_X1 U525 ( .A1(n514), .A2(n2), .B1(n4), .B2(n515), .ZN(n513) );
  AOI22_X1 U526 ( .A1(n518), .A2(n5), .B1(n513), .B2(n516), .ZN(n751) );
  AOI22_X1 U527 ( .A1(n3), .A2(n515), .B1(n514), .B2(n61), .ZN(n517) );
  AOI22_X1 U528 ( .A1(n518), .A2(n49), .B1(n517), .B2(n516), .ZN(n750) );
  NAND2_X1 U529 ( .A1(n519), .A2(n598), .ZN(n587) );
  NAND2_X1 U530 ( .A1(n59), .A2(n524), .ZN(n525) );
  OAI211_X1 U531 ( .C1(n600), .C2(n587), .A(n63), .B(n525), .ZN(n526) );
  INV_X1 U532 ( .A(n526), .ZN(n529) );
  AOI22_X1 U533 ( .A1(n524), .A2(n660), .B1(n659), .B2(n525), .ZN(n520) );
  AOI22_X1 U534 ( .A1(n529), .A2(n521), .B1(n520), .B2(n526), .ZN(n749) );
  AOI22_X1 U535 ( .A1(n524), .A2(n2), .B1(n4), .B2(n525), .ZN(n522) );
  AOI22_X1 U536 ( .A1(n529), .A2(n523), .B1(n522), .B2(n526), .ZN(n748) );
  AOI22_X1 U537 ( .A1(n3), .A2(n525), .B1(n524), .B2(n61), .ZN(n527) );
  AOI22_X1 U538 ( .A1(n529), .A2(n528), .B1(n527), .B2(n526), .ZN(n747) );
  NAND2_X1 U539 ( .A1(n59), .A2(n534), .ZN(n535) );
  OAI211_X1 U540 ( .C1(n608), .C2(n587), .A(n63), .B(n535), .ZN(n536) );
  INV_X1 U541 ( .A(n536), .ZN(n539) );
  AOI22_X1 U542 ( .A1(n534), .A2(n660), .B1(n60), .B2(n535), .ZN(n530) );
  AOI22_X1 U543 ( .A1(n539), .A2(n531), .B1(n530), .B2(n536), .ZN(n746) );
  AOI22_X1 U544 ( .A1(n534), .A2(n2), .B1(n4), .B2(n535), .ZN(n532) );
  AOI22_X1 U545 ( .A1(n539), .A2(n533), .B1(n532), .B2(n536), .ZN(n745) );
  AOI22_X1 U546 ( .A1(n3), .A2(n535), .B1(n534), .B2(n61), .ZN(n537) );
  AOI22_X1 U547 ( .A1(n539), .A2(n538), .B1(n537), .B2(n536), .ZN(n744) );
  NAND2_X1 U548 ( .A1(n59), .A2(n544), .ZN(n545) );
  OAI211_X1 U549 ( .C1(n616), .C2(n587), .A(n63), .B(n545), .ZN(n546) );
  INV_X1 U550 ( .A(n546), .ZN(n549) );
  AOI22_X1 U551 ( .A1(n544), .A2(n660), .B1(n60), .B2(n545), .ZN(n540) );
  AOI22_X1 U552 ( .A1(n549), .A2(n541), .B1(n540), .B2(n546), .ZN(n743) );
  AOI22_X1 U553 ( .A1(n544), .A2(n2), .B1(n4), .B2(n545), .ZN(n542) );
  AOI22_X1 U554 ( .A1(n549), .A2(n543), .B1(n542), .B2(n546), .ZN(n742) );
  AOI22_X1 U555 ( .A1(n3), .A2(n545), .B1(n544), .B2(n61), .ZN(n547) );
  AOI22_X1 U556 ( .A1(n549), .A2(n548), .B1(n547), .B2(n546), .ZN(n741) );
  NAND2_X1 U557 ( .A1(n59), .A2(n554), .ZN(n555) );
  OAI211_X1 U558 ( .C1(n624), .C2(n587), .A(n63), .B(n555), .ZN(n556) );
  INV_X1 U559 ( .A(n556), .ZN(n559) );
  AOI22_X1 U560 ( .A1(n554), .A2(n660), .B1(n60), .B2(n555), .ZN(n550) );
  AOI22_X1 U561 ( .A1(n559), .A2(n551), .B1(n550), .B2(n556), .ZN(n740) );
  AOI22_X1 U562 ( .A1(n554), .A2(n2), .B1(n4), .B2(n555), .ZN(n552) );
  AOI22_X1 U563 ( .A1(n559), .A2(n553), .B1(n552), .B2(n556), .ZN(n739) );
  AOI22_X1 U564 ( .A1(n3), .A2(n555), .B1(n554), .B2(n61), .ZN(n557) );
  AOI22_X1 U565 ( .A1(n559), .A2(n558), .B1(n557), .B2(n556), .ZN(n738) );
  NAND2_X1 U566 ( .A1(n59), .A2(n564), .ZN(n565) );
  OAI211_X1 U567 ( .C1(n632), .C2(n587), .A(n63), .B(n565), .ZN(n566) );
  INV_X1 U568 ( .A(n566), .ZN(n569) );
  AOI22_X1 U569 ( .A1(n564), .A2(n660), .B1(n60), .B2(n565), .ZN(n560) );
  AOI22_X1 U570 ( .A1(n569), .A2(n561), .B1(n560), .B2(n566), .ZN(n737) );
  AOI22_X1 U571 ( .A1(n564), .A2(n2), .B1(n4), .B2(n565), .ZN(n562) );
  AOI22_X1 U572 ( .A1(n569), .A2(n563), .B1(n562), .B2(n566), .ZN(n736) );
  AOI22_X1 U573 ( .A1(n3), .A2(n565), .B1(n564), .B2(n61), .ZN(n567) );
  AOI22_X1 U574 ( .A1(n569), .A2(n568), .B1(n567), .B2(n566), .ZN(n735) );
  NAND2_X1 U575 ( .A1(n59), .A2(n574), .ZN(n575) );
  OAI211_X1 U576 ( .C1(n640), .C2(n587), .A(n62), .B(n575), .ZN(n576) );
  INV_X1 U577 ( .A(n576), .ZN(n579) );
  AOI22_X1 U578 ( .A1(n574), .A2(n660), .B1(n60), .B2(n575), .ZN(n570) );
  AOI22_X1 U579 ( .A1(n579), .A2(n571), .B1(n570), .B2(n576), .ZN(n734) );
  AOI22_X1 U580 ( .A1(n574), .A2(n2), .B1(n4), .B2(n575), .ZN(n572) );
  AOI22_X1 U581 ( .A1(n579), .A2(n573), .B1(n572), .B2(n576), .ZN(n733) );
  AOI22_X1 U582 ( .A1(n3), .A2(n575), .B1(n574), .B2(n61), .ZN(n577) );
  AOI22_X1 U583 ( .A1(n579), .A2(n578), .B1(n577), .B2(n576), .ZN(n732) );
  NAND2_X1 U584 ( .A1(n59), .A2(n582), .ZN(n583) );
  OAI211_X1 U585 ( .C1(n648), .C2(n587), .A(n62), .B(n583), .ZN(n584) );
  INV_X1 U586 ( .A(n584), .ZN(n586) );
  AOI22_X1 U587 ( .A1(n582), .A2(n660), .B1(n659), .B2(n583), .ZN(n580) );
  AOI22_X1 U588 ( .A1(n586), .A2(n38), .B1(n580), .B2(n584), .ZN(n731) );
  AOI22_X1 U589 ( .A1(n582), .A2(n2), .B1(n662), .B2(n583), .ZN(n581) );
  AOI22_X1 U590 ( .A1(n586), .A2(n35), .B1(n581), .B2(n584), .ZN(n730) );
  AOI22_X1 U591 ( .A1(n3), .A2(n583), .B1(n582), .B2(n665), .ZN(n585) );
  AOI22_X1 U592 ( .A1(n586), .A2(n41), .B1(n585), .B2(n584), .ZN(n729) );
  NAND2_X1 U593 ( .A1(n59), .A2(n592), .ZN(n593) );
  OAI211_X1 U594 ( .C1(n658), .C2(n587), .A(n62), .B(n593), .ZN(n594) );
  INV_X1 U595 ( .A(n594), .ZN(n597) );
  AOI22_X1 U596 ( .A1(n592), .A2(n660), .B1(n659), .B2(n593), .ZN(n588) );
  AOI22_X1 U597 ( .A1(n597), .A2(n589), .B1(n588), .B2(n594), .ZN(n728) );
  AOI22_X1 U598 ( .A1(n592), .A2(n2), .B1(n4), .B2(n593), .ZN(n590) );
  AOI22_X1 U599 ( .A1(n597), .A2(n591), .B1(n590), .B2(n594), .ZN(n727) );
  AOI22_X1 U600 ( .A1(n3), .A2(n593), .B1(n592), .B2(n665), .ZN(n595) );
  AOI22_X1 U601 ( .A1(n597), .A2(n596), .B1(n595), .B2(n594), .ZN(n726) );
  NAND2_X1 U602 ( .A1(n599), .A2(n598), .ZN(n657) );
  NAND2_X1 U603 ( .A1(n59), .A2(n603), .ZN(n604) );
  OAI211_X1 U604 ( .C1(n600), .C2(n657), .A(n62), .B(n604), .ZN(n605) );
  INV_X1 U605 ( .A(n605), .ZN(n607) );
  AOI22_X1 U606 ( .A1(n603), .A2(n660), .B1(n60), .B2(n604), .ZN(n601) );
  AOI22_X1 U607 ( .A1(n607), .A2(n18), .B1(n601), .B2(n605), .ZN(n725) );
  AOI22_X1 U608 ( .A1(n603), .A2(n2), .B1(n4), .B2(n604), .ZN(n602) );
  AOI22_X1 U609 ( .A1(n607), .A2(n24), .B1(n602), .B2(n605), .ZN(n724) );
  AOI22_X1 U610 ( .A1(n3), .A2(n604), .B1(n603), .B2(n665), .ZN(n606) );
  AOI22_X1 U611 ( .A1(n607), .A2(n13), .B1(n606), .B2(n605), .ZN(n723) );
  NAND2_X1 U612 ( .A1(n59), .A2(n611), .ZN(n612) );
  OAI211_X1 U613 ( .C1(n608), .C2(n657), .A(n62), .B(n612), .ZN(n613) );
  INV_X1 U614 ( .A(n613), .ZN(n615) );
  AOI22_X1 U615 ( .A1(n611), .A2(n660), .B1(n659), .B2(n612), .ZN(n609) );
  AOI22_X1 U616 ( .A1(n615), .A2(n29), .B1(n609), .B2(n613), .ZN(n722) );
  AOI22_X1 U617 ( .A1(n611), .A2(n2), .B1(n662), .B2(n612), .ZN(n610) );
  AOI22_X1 U618 ( .A1(n615), .A2(n26), .B1(n610), .B2(n613), .ZN(n721) );
  AOI22_X1 U619 ( .A1(n3), .A2(n612), .B1(n611), .B2(n665), .ZN(n614) );
  AOI22_X1 U620 ( .A1(n615), .A2(n32), .B1(n614), .B2(n613), .ZN(n720) );
  NAND2_X1 U621 ( .A1(n59), .A2(n619), .ZN(n620) );
  OAI211_X1 U622 ( .C1(n616), .C2(n657), .A(n62), .B(n620), .ZN(n621) );
  INV_X1 U623 ( .A(n621), .ZN(n623) );
  AOI22_X1 U624 ( .A1(n619), .A2(n660), .B1(n659), .B2(n620), .ZN(n617) );
  AOI22_X1 U625 ( .A1(n623), .A2(n39), .B1(n617), .B2(n621), .ZN(n719) );
  AOI22_X1 U626 ( .A1(n619), .A2(n2), .B1(n4), .B2(n620), .ZN(n618) );
  AOI22_X1 U627 ( .A1(n623), .A2(n36), .B1(n618), .B2(n621), .ZN(n718) );
  AOI22_X1 U628 ( .A1(n3), .A2(n620), .B1(n619), .B2(n665), .ZN(n622) );
  AOI22_X1 U629 ( .A1(n623), .A2(n42), .B1(n622), .B2(n621), .ZN(n717) );
  NAND2_X1 U630 ( .A1(n59), .A2(n627), .ZN(n628) );
  OAI211_X1 U631 ( .C1(n624), .C2(n657), .A(n62), .B(n628), .ZN(n629) );
  INV_X1 U632 ( .A(n629), .ZN(n631) );
  AOI22_X1 U633 ( .A1(n627), .A2(n660), .B1(n659), .B2(n628), .ZN(n625) );
  AOI22_X1 U634 ( .A1(n631), .A2(n30), .B1(n625), .B2(n629), .ZN(n716) );
  AOI22_X1 U635 ( .A1(n627), .A2(n2), .B1(n662), .B2(n628), .ZN(n626) );
  AOI22_X1 U636 ( .A1(n631), .A2(n27), .B1(n626), .B2(n629), .ZN(n715) );
  AOI22_X1 U637 ( .A1(n3), .A2(n628), .B1(n627), .B2(n665), .ZN(n630) );
  AOI22_X1 U638 ( .A1(n631), .A2(n33), .B1(n630), .B2(n629), .ZN(n714) );
  NAND2_X1 U639 ( .A1(n59), .A2(n635), .ZN(n636) );
  OAI211_X1 U640 ( .C1(n632), .C2(n657), .A(n62), .B(n636), .ZN(n637) );
  INV_X1 U641 ( .A(n637), .ZN(n639) );
  AOI22_X1 U642 ( .A1(n635), .A2(n660), .B1(n659), .B2(n636), .ZN(n633) );
  AOI22_X1 U643 ( .A1(n639), .A2(n19), .B1(n633), .B2(n637), .ZN(n713) );
  AOI22_X1 U644 ( .A1(n635), .A2(n2), .B1(n4), .B2(n636), .ZN(n634) );
  AOI22_X1 U645 ( .A1(n639), .A2(n25), .B1(n634), .B2(n637), .ZN(n712) );
  AOI22_X1 U646 ( .A1(n3), .A2(n636), .B1(n635), .B2(n665), .ZN(n638) );
  AOI22_X1 U647 ( .A1(n639), .A2(n14), .B1(n638), .B2(n637), .ZN(n711) );
  NAND2_X1 U648 ( .A1(n59), .A2(n643), .ZN(n644) );
  OAI211_X1 U649 ( .C1(n640), .C2(n657), .A(n62), .B(n644), .ZN(n645) );
  INV_X1 U650 ( .A(n645), .ZN(n647) );
  AOI22_X1 U651 ( .A1(n643), .A2(n660), .B1(n659), .B2(n644), .ZN(n641) );
  AOI22_X1 U652 ( .A1(n647), .A2(n31), .B1(n641), .B2(n645), .ZN(n710) );
  AOI22_X1 U653 ( .A1(n643), .A2(n2), .B1(n662), .B2(n644), .ZN(n642) );
  AOI22_X1 U654 ( .A1(n647), .A2(n28), .B1(n642), .B2(n645), .ZN(n709) );
  AOI22_X1 U655 ( .A1(n3), .A2(n644), .B1(n643), .B2(n665), .ZN(n646) );
  AOI22_X1 U656 ( .A1(n647), .A2(n34), .B1(n646), .B2(n645), .ZN(n708) );
  NAND2_X1 U657 ( .A1(n59), .A2(n651), .ZN(n652) );
  OAI211_X1 U658 ( .C1(n648), .C2(n657), .A(n62), .B(n652), .ZN(n653) );
  INV_X1 U659 ( .A(n653), .ZN(n655) );
  AOI22_X1 U660 ( .A1(n651), .A2(n660), .B1(n659), .B2(n652), .ZN(n649) );
  AOI22_X1 U661 ( .A1(n655), .A2(n40), .B1(n649), .B2(n653), .ZN(n707) );
  AOI22_X1 U662 ( .A1(n651), .A2(n2), .B1(n4), .B2(n652), .ZN(n650) );
  AOI22_X1 U663 ( .A1(n655), .A2(n37), .B1(n650), .B2(n653), .ZN(n706) );
  AOI22_X1 U664 ( .A1(n3), .A2(n652), .B1(n651), .B2(n665), .ZN(n654) );
  AOI22_X1 U665 ( .A1(n655), .A2(n43), .B1(n654), .B2(n653), .ZN(n705) );
  NAND2_X1 U666 ( .A1(n656), .A2(n666), .ZN(n667) );
  OAI211_X1 U667 ( .C1(n658), .C2(n657), .A(n62), .B(n667), .ZN(n669) );
  INV_X1 U668 ( .A(n669), .ZN(n671) );
  AOI22_X1 U669 ( .A1(n666), .A2(n660), .B1(n60), .B2(n667), .ZN(n661) );
  AOI22_X1 U670 ( .A1(n671), .A2(n17), .B1(n661), .B2(n669), .ZN(n704) );
  AOI22_X1 U671 ( .A1(n666), .A2(n2), .B1(n4), .B2(n667), .ZN(n664) );
  AOI22_X1 U672 ( .A1(n671), .A2(n23), .B1(n664), .B2(n669), .ZN(n703) );
  AOI22_X1 U673 ( .A1(n3), .A2(n667), .B1(n666), .B2(n61), .ZN(n670) );
  AOI22_X1 U674 ( .A1(n671), .A2(n12), .B1(n670), .B2(n669), .ZN(n702) );
endmodule


module in_loc_selblock_NBIT_DATA32_N8_F5 ( regs, win, curr_proc_regs );
  input [2559:0] regs;
  input [4:0] win;
  output [511:0] curr_proc_regs;
  wire   n1, n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585;

  CLKBUF_X3 U2 ( .A(n41), .Z(n38) );
  BUF_X2 U3 ( .A(n13), .Z(n14) );
  BUF_X4 U4 ( .A(n11), .Z(n13) );
  BUF_X4 U5 ( .A(n24), .Z(n28) );
  BUF_X2 U6 ( .A(n10), .Z(n1) );
  BUF_X2 U7 ( .A(n9), .Z(n2) );
  BUF_X4 U8 ( .A(n17), .Z(n11) );
  CLKBUF_X3 U9 ( .A(n1582), .Z(n35) );
  CLKBUF_X3 U10 ( .A(n1582), .Z(n34) );
  BUF_X4 U11 ( .A(n1582), .Z(n3) );
  BUF_X2 U12 ( .A(n37), .Z(n4) );
  BUF_X4 U13 ( .A(n1580), .Z(n5) );
  BUF_X2 U14 ( .A(win[4]), .Z(n41) );
  BUF_X2 U15 ( .A(n19), .Z(n7) );
  BUF_X2 U16 ( .A(n7), .Z(n16) );
  BUF_X2 U17 ( .A(n2), .Z(n31) );
  BUF_X2 U18 ( .A(n1), .Z(n8) );
  BUF_X4 U19 ( .A(n1582), .Z(n9) );
  BUF_X2 U20 ( .A(n4), .Z(n10) );
  BUF_X4 U21 ( .A(n5), .Z(n12) );
  BUF_X2 U22 ( .A(n1579), .Z(n15) );
  BUF_X2 U23 ( .A(n41), .Z(n39) );
  BUF_X2 U24 ( .A(n41), .Z(n37) );
  AND2_X2 U25 ( .A1(n43), .A2(win[1]), .ZN(n1579) );
  AND3_X2 U26 ( .A1(n43), .A2(win[0]), .A3(n42), .ZN(n1580) );
  NOR3_X2 U27 ( .A1(win[3]), .A2(win[4]), .A3(n44), .ZN(n1581) );
  BUF_X32 U28 ( .A(n1581), .Z(n29) );
  BUF_X1 U29 ( .A(n12), .Z(n22) );
  BUF_X1 U30 ( .A(n14), .Z(n20) );
  BUF_X1 U31 ( .A(n17), .Z(n18) );
  BUF_X1 U32 ( .A(n9), .Z(n32) );
  BUF_X1 U33 ( .A(n5), .Z(n23) );
  BUF_X1 U34 ( .A(n26), .Z(n25) );
  BUF_X1 U35 ( .A(n1580), .Z(n26) );
  BUF_X1 U36 ( .A(n28), .Z(n21) );
  BUF_X1 U37 ( .A(n1582), .Z(n33) );
  BUF_X1 U38 ( .A(n9), .Z(n30) );
  BUF_X1 U39 ( .A(n28), .Z(n27) );
  BUF_X1 U40 ( .A(n11), .Z(n19) );
  BUF_X1 U41 ( .A(n1579), .Z(n17) );
  BUF_X2 U42 ( .A(n5), .Z(n24) );
  BUF_X1 U43 ( .A(n8), .Z(n36) );
  BUF_X1 U44 ( .A(n41), .Z(n40) );
  NOR3_X1 U45 ( .A1(win[2]), .A2(win[3]), .A3(win[4]), .ZN(n43) );
  INV_X1 U46 ( .A(win[1]), .ZN(n42) );
  NAND2_X1 U47 ( .A1(regs[0]), .A2(n1580), .ZN(n48) );
  INV_X1 U48 ( .A(win[2]), .ZN(n44) );
  AOI22_X1 U49 ( .A1(n11), .A2(regs[512]), .B1(n29), .B2(regs[1024]), .ZN(n47)
         );
  INV_X1 U50 ( .A(win[3]), .ZN(n45) );
  NOR2_X1 U51 ( .A1(n38), .A2(n45), .ZN(n1582) );
  AOI22_X1 U52 ( .A1(win[4]), .A2(regs[2048]), .B1(n3), .B2(regs[1536]), .ZN(
        n46) );
  NAND3_X1 U53 ( .A1(n48), .A2(n47), .A3(n46), .ZN(curr_proc_regs[0]) );
  NAND2_X1 U54 ( .A1(regs[612]), .A2(n11), .ZN(n51) );
  AOI22_X1 U55 ( .A1(n29), .A2(regs[1124]), .B1(n21), .B2(regs[100]), .ZN(n50)
         );
  AOI22_X1 U56 ( .A1(win[4]), .A2(regs[2148]), .B1(n34), .B2(regs[1636]), .ZN(
        n49) );
  NAND3_X1 U57 ( .A1(n51), .A2(n50), .A3(n49), .ZN(curr_proc_regs[100]) );
  NAND2_X1 U58 ( .A1(regs[613]), .A2(n18), .ZN(n54) );
  AOI22_X1 U59 ( .A1(n29), .A2(regs[1125]), .B1(n21), .B2(regs[101]), .ZN(n53)
         );
  AOI22_X1 U60 ( .A1(win[4]), .A2(regs[2149]), .B1(n33), .B2(regs[1637]), .ZN(
        n52) );
  NAND3_X1 U61 ( .A1(n54), .A2(n53), .A3(n52), .ZN(curr_proc_regs[101]) );
  NAND2_X1 U62 ( .A1(regs[614]), .A2(n11), .ZN(n57) );
  AOI22_X1 U63 ( .A1(n29), .A2(regs[1126]), .B1(n22), .B2(regs[102]), .ZN(n56)
         );
  AOI22_X1 U64 ( .A1(n39), .A2(regs[2150]), .B1(n34), .B2(regs[1638]), .ZN(n55) );
  NAND3_X1 U65 ( .A1(n57), .A2(n56), .A3(n55), .ZN(curr_proc_regs[102]) );
  NAND2_X1 U66 ( .A1(regs[615]), .A2(n18), .ZN(n60) );
  AOI22_X1 U67 ( .A1(n29), .A2(regs[1127]), .B1(n1580), .B2(regs[103]), .ZN(
        n59) );
  AOI22_X1 U68 ( .A1(win[4]), .A2(regs[2151]), .B1(n9), .B2(regs[1639]), .ZN(
        n58) );
  NAND3_X1 U69 ( .A1(n60), .A2(n59), .A3(n58), .ZN(curr_proc_regs[103]) );
  NAND2_X1 U70 ( .A1(regs[616]), .A2(n11), .ZN(n63) );
  AOI22_X1 U71 ( .A1(n29), .A2(regs[1128]), .B1(n1580), .B2(regs[104]), .ZN(
        n62) );
  AOI22_X1 U72 ( .A1(win[4]), .A2(regs[2152]), .B1(n9), .B2(regs[1640]), .ZN(
        n61) );
  NAND3_X1 U73 ( .A1(n63), .A2(n62), .A3(n61), .ZN(curr_proc_regs[104]) );
  NAND2_X1 U74 ( .A1(regs[617]), .A2(n11), .ZN(n66) );
  AOI22_X1 U75 ( .A1(n29), .A2(regs[1129]), .B1(n22), .B2(regs[105]), .ZN(n65)
         );
  AOI22_X1 U76 ( .A1(win[4]), .A2(regs[2153]), .B1(n35), .B2(regs[1641]), .ZN(
        n64) );
  NAND3_X1 U77 ( .A1(n66), .A2(n65), .A3(n64), .ZN(curr_proc_regs[105]) );
  NAND2_X1 U78 ( .A1(regs[618]), .A2(n11), .ZN(n69) );
  AOI22_X1 U79 ( .A1(n29), .A2(regs[1130]), .B1(n21), .B2(regs[106]), .ZN(n68)
         );
  AOI22_X1 U80 ( .A1(n36), .A2(regs[2154]), .B1(n3), .B2(regs[1642]), .ZN(n67)
         );
  NAND3_X1 U81 ( .A1(n69), .A2(n68), .A3(n67), .ZN(curr_proc_regs[106]) );
  NAND2_X1 U82 ( .A1(regs[619]), .A2(n15), .ZN(n72) );
  AOI22_X1 U83 ( .A1(n29), .A2(regs[1131]), .B1(n22), .B2(regs[107]), .ZN(n71)
         );
  AOI22_X1 U84 ( .A1(win[4]), .A2(regs[2155]), .B1(n3), .B2(regs[1643]), .ZN(
        n70) );
  NAND3_X1 U85 ( .A1(n72), .A2(n71), .A3(n70), .ZN(curr_proc_regs[107]) );
  NAND2_X1 U86 ( .A1(regs[620]), .A2(n11), .ZN(n75) );
  AOI22_X1 U87 ( .A1(n29), .A2(regs[1132]), .B1(n1580), .B2(regs[108]), .ZN(
        n74) );
  AOI22_X1 U88 ( .A1(win[4]), .A2(regs[2156]), .B1(n34), .B2(regs[1644]), .ZN(
        n73) );
  NAND3_X1 U89 ( .A1(n75), .A2(n74), .A3(n73), .ZN(curr_proc_regs[108]) );
  NAND2_X1 U90 ( .A1(regs[621]), .A2(n1579), .ZN(n78) );
  AOI22_X1 U91 ( .A1(n29), .A2(regs[1133]), .B1(n24), .B2(regs[109]), .ZN(n77)
         );
  AOI22_X1 U92 ( .A1(win[4]), .A2(regs[2157]), .B1(n33), .B2(regs[1645]), .ZN(
        n76) );
  NAND3_X1 U93 ( .A1(n78), .A2(n77), .A3(n76), .ZN(curr_proc_regs[109]) );
  NAND2_X1 U94 ( .A1(regs[522]), .A2(n16), .ZN(n81) );
  AOI22_X1 U95 ( .A1(n29), .A2(regs[1034]), .B1(n12), .B2(regs[10]), .ZN(n80)
         );
  AOI22_X1 U96 ( .A1(n38), .A2(regs[2058]), .B1(n30), .B2(regs[1546]), .ZN(n79) );
  NAND3_X1 U97 ( .A1(n81), .A2(n80), .A3(n79), .ZN(curr_proc_regs[10]) );
  NAND2_X1 U98 ( .A1(regs[622]), .A2(n15), .ZN(n84) );
  AOI22_X1 U99 ( .A1(n29), .A2(regs[1134]), .B1(n24), .B2(regs[110]), .ZN(n83)
         );
  AOI22_X1 U100 ( .A1(n38), .A2(regs[2158]), .B1(n30), .B2(regs[1646]), .ZN(
        n82) );
  NAND3_X1 U101 ( .A1(n84), .A2(n83), .A3(n82), .ZN(curr_proc_regs[110]) );
  NAND2_X1 U102 ( .A1(regs[623]), .A2(n1579), .ZN(n87) );
  AOI22_X1 U103 ( .A1(n29), .A2(regs[1135]), .B1(n12), .B2(regs[111]), .ZN(n86) );
  AOI22_X1 U104 ( .A1(n38), .A2(regs[2159]), .B1(n30), .B2(regs[1647]), .ZN(
        n85) );
  NAND3_X1 U105 ( .A1(n87), .A2(n86), .A3(n85), .ZN(curr_proc_regs[111]) );
  NAND2_X1 U106 ( .A1(regs[624]), .A2(n16), .ZN(n90) );
  AOI22_X1 U107 ( .A1(n29), .A2(regs[1136]), .B1(n12), .B2(regs[112]), .ZN(n89) );
  AOI22_X1 U108 ( .A1(n38), .A2(regs[2160]), .B1(n30), .B2(regs[1648]), .ZN(
        n88) );
  NAND3_X1 U109 ( .A1(n90), .A2(n89), .A3(n88), .ZN(curr_proc_regs[112]) );
  NAND2_X1 U110 ( .A1(regs[625]), .A2(n15), .ZN(n93) );
  AOI22_X1 U111 ( .A1(n29), .A2(regs[1137]), .B1(n5), .B2(regs[113]), .ZN(n92)
         );
  AOI22_X1 U112 ( .A1(n38), .A2(regs[2161]), .B1(n30), .B2(regs[1649]), .ZN(
        n91) );
  NAND3_X1 U113 ( .A1(n93), .A2(n92), .A3(n91), .ZN(curr_proc_regs[113]) );
  NAND2_X1 U114 ( .A1(regs[626]), .A2(n1579), .ZN(n96) );
  AOI22_X1 U115 ( .A1(n29), .A2(regs[1138]), .B1(n28), .B2(regs[114]), .ZN(n95) );
  AOI22_X1 U116 ( .A1(n38), .A2(regs[2162]), .B1(n30), .B2(regs[1650]), .ZN(
        n94) );
  NAND3_X1 U117 ( .A1(n96), .A2(n95), .A3(n94), .ZN(curr_proc_regs[114]) );
  NAND2_X1 U118 ( .A1(regs[627]), .A2(n16), .ZN(n99) );
  AOI22_X1 U119 ( .A1(n29), .A2(regs[1139]), .B1(n24), .B2(regs[115]), .ZN(n98) );
  AOI22_X1 U120 ( .A1(n38), .A2(regs[2163]), .B1(n30), .B2(regs[1651]), .ZN(
        n97) );
  NAND3_X1 U121 ( .A1(n99), .A2(n98), .A3(n97), .ZN(curr_proc_regs[115]) );
  NAND2_X1 U122 ( .A1(regs[628]), .A2(n15), .ZN(n102) );
  AOI22_X1 U123 ( .A1(n29), .A2(regs[1140]), .B1(n1580), .B2(regs[116]), .ZN(
        n101) );
  AOI22_X1 U124 ( .A1(n38), .A2(regs[2164]), .B1(n30), .B2(regs[1652]), .ZN(
        n100) );
  NAND3_X1 U125 ( .A1(n102), .A2(n101), .A3(n100), .ZN(curr_proc_regs[116]) );
  NAND2_X1 U126 ( .A1(regs[629]), .A2(n1579), .ZN(n105) );
  AOI22_X1 U127 ( .A1(n29), .A2(regs[1141]), .B1(n12), .B2(regs[117]), .ZN(
        n104) );
  AOI22_X1 U128 ( .A1(n38), .A2(regs[2165]), .B1(n30), .B2(regs[1653]), .ZN(
        n103) );
  NAND3_X1 U129 ( .A1(n105), .A2(n104), .A3(n103), .ZN(curr_proc_regs[117]) );
  NAND2_X1 U130 ( .A1(regs[630]), .A2(n16), .ZN(n108) );
  AOI22_X1 U131 ( .A1(n29), .A2(regs[1142]), .B1(n22), .B2(regs[118]), .ZN(
        n107) );
  AOI22_X1 U132 ( .A1(n38), .A2(regs[2166]), .B1(n30), .B2(regs[1654]), .ZN(
        n106) );
  NAND3_X1 U133 ( .A1(n108), .A2(n107), .A3(n106), .ZN(curr_proc_regs[118]) );
  NAND2_X1 U134 ( .A1(regs[631]), .A2(n15), .ZN(n111) );
  AOI22_X1 U135 ( .A1(n29), .A2(regs[1143]), .B1(n25), .B2(regs[119]), .ZN(
        n110) );
  AOI22_X1 U136 ( .A1(n38), .A2(regs[2167]), .B1(n30), .B2(regs[1655]), .ZN(
        n109) );
  NAND3_X1 U137 ( .A1(n111), .A2(n110), .A3(n109), .ZN(curr_proc_regs[119]) );
  NAND2_X1 U138 ( .A1(regs[523]), .A2(n13), .ZN(n114) );
  AOI22_X1 U139 ( .A1(n29), .A2(regs[1035]), .B1(n22), .B2(regs[11]), .ZN(n113) );
  AOI22_X1 U140 ( .A1(n39), .A2(regs[2059]), .B1(n35), .B2(regs[1547]), .ZN(
        n112) );
  NAND3_X1 U141 ( .A1(n114), .A2(n113), .A3(n112), .ZN(curr_proc_regs[11]) );
  NAND2_X1 U142 ( .A1(regs[632]), .A2(n13), .ZN(n117) );
  AOI22_X1 U143 ( .A1(n29), .A2(regs[1144]), .B1(n1580), .B2(regs[120]), .ZN(
        n116) );
  AOI22_X1 U144 ( .A1(n39), .A2(regs[2168]), .B1(n35), .B2(regs[1656]), .ZN(
        n115) );
  NAND3_X1 U145 ( .A1(n117), .A2(n116), .A3(n115), .ZN(curr_proc_regs[120]) );
  NAND2_X1 U146 ( .A1(regs[633]), .A2(n13), .ZN(n120) );
  AOI22_X1 U147 ( .A1(n29), .A2(regs[1145]), .B1(n12), .B2(regs[121]), .ZN(
        n119) );
  AOI22_X1 U148 ( .A1(n40), .A2(regs[2169]), .B1(n35), .B2(regs[1657]), .ZN(
        n118) );
  NAND3_X1 U149 ( .A1(n120), .A2(n119), .A3(n118), .ZN(curr_proc_regs[121]) );
  NAND2_X1 U150 ( .A1(regs[634]), .A2(n13), .ZN(n123) );
  AOI22_X1 U151 ( .A1(n29), .A2(regs[1146]), .B1(n21), .B2(regs[122]), .ZN(
        n122) );
  AOI22_X1 U152 ( .A1(n41), .A2(regs[2170]), .B1(n35), .B2(regs[1658]), .ZN(
        n121) );
  NAND3_X1 U153 ( .A1(n123), .A2(n122), .A3(n121), .ZN(curr_proc_regs[122]) );
  NAND2_X1 U154 ( .A1(regs[635]), .A2(n13), .ZN(n126) );
  AOI22_X1 U155 ( .A1(n29), .A2(regs[1147]), .B1(n22), .B2(regs[123]), .ZN(
        n125) );
  AOI22_X1 U156 ( .A1(n8), .A2(regs[2171]), .B1(n35), .B2(regs[1659]), .ZN(
        n124) );
  NAND3_X1 U157 ( .A1(n126), .A2(n125), .A3(n124), .ZN(curr_proc_regs[123]) );
  NAND2_X1 U158 ( .A1(regs[636]), .A2(n13), .ZN(n129) );
  AOI22_X1 U159 ( .A1(n29), .A2(regs[1148]), .B1(n1580), .B2(regs[124]), .ZN(
        n128) );
  AOI22_X1 U160 ( .A1(n36), .A2(regs[2172]), .B1(n35), .B2(regs[1660]), .ZN(
        n127) );
  NAND3_X1 U161 ( .A1(n129), .A2(n128), .A3(n127), .ZN(curr_proc_regs[124]) );
  NAND2_X1 U162 ( .A1(regs[637]), .A2(n13), .ZN(n132) );
  AOI22_X1 U163 ( .A1(n29), .A2(regs[1149]), .B1(n28), .B2(regs[125]), .ZN(
        n131) );
  AOI22_X1 U164 ( .A1(n38), .A2(regs[2173]), .B1(n35), .B2(regs[1661]), .ZN(
        n130) );
  NAND3_X1 U165 ( .A1(n132), .A2(n131), .A3(n130), .ZN(curr_proc_regs[125]) );
  NAND2_X1 U166 ( .A1(regs[638]), .A2(n13), .ZN(n135) );
  AOI22_X1 U167 ( .A1(n29), .A2(regs[1150]), .B1(n21), .B2(regs[126]), .ZN(
        n134) );
  AOI22_X1 U168 ( .A1(n39), .A2(regs[2174]), .B1(n35), .B2(regs[1662]), .ZN(
        n133) );
  NAND3_X1 U169 ( .A1(n135), .A2(n134), .A3(n133), .ZN(curr_proc_regs[126]) );
  NAND2_X1 U170 ( .A1(regs[639]), .A2(n13), .ZN(n138) );
  AOI22_X1 U171 ( .A1(n29), .A2(regs[1151]), .B1(n22), .B2(regs[127]), .ZN(
        n137) );
  AOI22_X1 U172 ( .A1(n37), .A2(regs[2175]), .B1(n35), .B2(regs[1663]), .ZN(
        n136) );
  NAND3_X1 U173 ( .A1(n138), .A2(n137), .A3(n136), .ZN(curr_proc_regs[127]) );
  NAND2_X1 U174 ( .A1(regs[640]), .A2(n13), .ZN(n141) );
  AOI22_X1 U175 ( .A1(n29), .A2(regs[1152]), .B1(n1580), .B2(regs[128]), .ZN(
        n140) );
  AOI22_X1 U176 ( .A1(n38), .A2(regs[2176]), .B1(n35), .B2(regs[1664]), .ZN(
        n139) );
  NAND3_X1 U177 ( .A1(n141), .A2(n140), .A3(n139), .ZN(curr_proc_regs[128]) );
  NAND2_X1 U178 ( .A1(regs[641]), .A2(n13), .ZN(n144) );
  AOI22_X1 U179 ( .A1(n29), .A2(regs[1153]), .B1(n12), .B2(regs[129]), .ZN(
        n143) );
  AOI22_X1 U180 ( .A1(n38), .A2(regs[2177]), .B1(n35), .B2(regs[1665]), .ZN(
        n142) );
  NAND3_X1 U181 ( .A1(n144), .A2(n143), .A3(n142), .ZN(curr_proc_regs[129]) );
  NAND2_X1 U182 ( .A1(regs[524]), .A2(n14), .ZN(n147) );
  AOI22_X1 U183 ( .A1(n29), .A2(regs[1036]), .B1(n5), .B2(regs[12]), .ZN(n146)
         );
  AOI22_X1 U184 ( .A1(n39), .A2(regs[2060]), .B1(n2), .B2(regs[1548]), .ZN(
        n145) );
  NAND3_X1 U185 ( .A1(n147), .A2(n146), .A3(n145), .ZN(curr_proc_regs[12]) );
  NAND2_X1 U186 ( .A1(regs[642]), .A2(n14), .ZN(n150) );
  AOI22_X1 U187 ( .A1(n29), .A2(regs[1154]), .B1(n12), .B2(regs[130]), .ZN(
        n149) );
  AOI22_X1 U188 ( .A1(n37), .A2(regs[2178]), .B1(n2), .B2(regs[1666]), .ZN(
        n148) );
  NAND3_X1 U189 ( .A1(n150), .A2(n149), .A3(n148), .ZN(curr_proc_regs[130]) );
  NAND2_X1 U190 ( .A1(regs[643]), .A2(n14), .ZN(n153) );
  AOI22_X1 U191 ( .A1(n29), .A2(regs[1155]), .B1(n12), .B2(regs[131]), .ZN(
        n152) );
  AOI22_X1 U192 ( .A1(n4), .A2(regs[2179]), .B1(n2), .B2(regs[1667]), .ZN(n151) );
  NAND3_X1 U193 ( .A1(n153), .A2(n152), .A3(n151), .ZN(curr_proc_regs[131]) );
  NAND2_X1 U194 ( .A1(regs[644]), .A2(n14), .ZN(n156) );
  AOI22_X1 U195 ( .A1(n29), .A2(regs[1156]), .B1(n28), .B2(regs[132]), .ZN(
        n155) );
  AOI22_X1 U196 ( .A1(n10), .A2(regs[2180]), .B1(n2), .B2(regs[1668]), .ZN(
        n154) );
  NAND3_X1 U197 ( .A1(n156), .A2(n155), .A3(n154), .ZN(curr_proc_regs[132]) );
  NAND2_X1 U198 ( .A1(regs[645]), .A2(n14), .ZN(n159) );
  AOI22_X1 U199 ( .A1(n29), .A2(regs[1157]), .B1(n24), .B2(regs[133]), .ZN(
        n158) );
  AOI22_X1 U200 ( .A1(n1), .A2(regs[2181]), .B1(n2), .B2(regs[1669]), .ZN(n157) );
  NAND3_X1 U201 ( .A1(n159), .A2(n158), .A3(n157), .ZN(curr_proc_regs[133]) );
  NAND2_X1 U202 ( .A1(regs[646]), .A2(n14), .ZN(n162) );
  AOI22_X1 U203 ( .A1(n29), .A2(regs[1158]), .B1(n12), .B2(regs[134]), .ZN(
        n161) );
  AOI22_X1 U204 ( .A1(n41), .A2(regs[2182]), .B1(n2), .B2(regs[1670]), .ZN(
        n160) );
  NAND3_X1 U205 ( .A1(n162), .A2(n161), .A3(n160), .ZN(curr_proc_regs[134]) );
  NAND2_X1 U206 ( .A1(regs[647]), .A2(n14), .ZN(n165) );
  AOI22_X1 U207 ( .A1(n29), .A2(regs[1159]), .B1(n12), .B2(regs[135]), .ZN(
        n164) );
  AOI22_X1 U208 ( .A1(n8), .A2(regs[2183]), .B1(n2), .B2(regs[1671]), .ZN(n163) );
  NAND3_X1 U209 ( .A1(n165), .A2(n164), .A3(n163), .ZN(curr_proc_regs[135]) );
  NAND2_X1 U210 ( .A1(regs[648]), .A2(n14), .ZN(n168) );
  AOI22_X1 U211 ( .A1(n29), .A2(regs[1160]), .B1(n5), .B2(regs[136]), .ZN(n167) );
  AOI22_X1 U212 ( .A1(n38), .A2(regs[2184]), .B1(n2), .B2(regs[1672]), .ZN(
        n166) );
  NAND3_X1 U213 ( .A1(n168), .A2(n167), .A3(n166), .ZN(curr_proc_regs[136]) );
  NAND2_X1 U214 ( .A1(regs[649]), .A2(n14), .ZN(n171) );
  AOI22_X1 U215 ( .A1(n29), .A2(regs[1161]), .B1(n24), .B2(regs[137]), .ZN(
        n170) );
  AOI22_X1 U216 ( .A1(n38), .A2(regs[2185]), .B1(n2), .B2(regs[1673]), .ZN(
        n169) );
  NAND3_X1 U217 ( .A1(n171), .A2(n170), .A3(n169), .ZN(curr_proc_regs[137]) );
  NAND2_X1 U218 ( .A1(regs[650]), .A2(n14), .ZN(n174) );
  AOI22_X1 U219 ( .A1(n29), .A2(regs[1162]), .B1(n12), .B2(regs[138]), .ZN(
        n173) );
  AOI22_X1 U220 ( .A1(n38), .A2(regs[2186]), .B1(n2), .B2(regs[1674]), .ZN(
        n172) );
  NAND3_X1 U221 ( .A1(n174), .A2(n173), .A3(n172), .ZN(curr_proc_regs[138]) );
  NAND2_X1 U222 ( .A1(regs[651]), .A2(n14), .ZN(n177) );
  AOI22_X1 U223 ( .A1(n29), .A2(regs[1163]), .B1(n24), .B2(regs[139]), .ZN(
        n176) );
  AOI22_X1 U224 ( .A1(n38), .A2(regs[2187]), .B1(n2), .B2(regs[1675]), .ZN(
        n175) );
  NAND3_X1 U225 ( .A1(n177), .A2(n176), .A3(n175), .ZN(curr_proc_regs[139]) );
  NAND2_X1 U226 ( .A1(regs[525]), .A2(n15), .ZN(n180) );
  AOI22_X1 U227 ( .A1(n29), .A2(regs[1037]), .B1(n21), .B2(regs[13]), .ZN(n179) );
  AOI22_X1 U228 ( .A1(n41), .A2(regs[2061]), .B1(n9), .B2(regs[1549]), .ZN(
        n178) );
  NAND3_X1 U229 ( .A1(n180), .A2(n179), .A3(n178), .ZN(curr_proc_regs[13]) );
  NAND2_X1 U230 ( .A1(regs[652]), .A2(n15), .ZN(n183) );
  AOI22_X1 U231 ( .A1(n29), .A2(regs[1164]), .B1(n21), .B2(regs[140]), .ZN(
        n182) );
  AOI22_X1 U232 ( .A1(win[4]), .A2(regs[2188]), .B1(n9), .B2(regs[1676]), .ZN(
        n181) );
  NAND3_X1 U233 ( .A1(n183), .A2(n182), .A3(n181), .ZN(curr_proc_regs[140]) );
  NAND2_X1 U234 ( .A1(regs[653]), .A2(n15), .ZN(n186) );
  AOI22_X1 U235 ( .A1(n29), .A2(regs[1165]), .B1(n21), .B2(regs[141]), .ZN(
        n185) );
  AOI22_X1 U236 ( .A1(n36), .A2(regs[2189]), .B1(n35), .B2(regs[1677]), .ZN(
        n184) );
  NAND3_X1 U237 ( .A1(n186), .A2(n185), .A3(n184), .ZN(curr_proc_regs[141]) );
  NAND2_X1 U238 ( .A1(regs[654]), .A2(n15), .ZN(n189) );
  AOI22_X1 U239 ( .A1(n29), .A2(regs[1166]), .B1(n21), .B2(regs[142]), .ZN(
        n188) );
  AOI22_X1 U240 ( .A1(n40), .A2(regs[2190]), .B1(n3), .B2(regs[1678]), .ZN(
        n187) );
  NAND3_X1 U241 ( .A1(n189), .A2(n188), .A3(n187), .ZN(curr_proc_regs[142]) );
  NAND2_X1 U242 ( .A1(regs[655]), .A2(n15), .ZN(n192) );
  AOI22_X1 U243 ( .A1(n29), .A2(regs[1167]), .B1(n21), .B2(regs[143]), .ZN(
        n191) );
  AOI22_X1 U244 ( .A1(n10), .A2(regs[2191]), .B1(n3), .B2(regs[1679]), .ZN(
        n190) );
  NAND3_X1 U245 ( .A1(n192), .A2(n191), .A3(n190), .ZN(curr_proc_regs[143]) );
  NAND2_X1 U246 ( .A1(regs[656]), .A2(n15), .ZN(n195) );
  AOI22_X1 U247 ( .A1(n29), .A2(regs[1168]), .B1(n21), .B2(regs[144]), .ZN(
        n194) );
  AOI22_X1 U248 ( .A1(n8), .A2(regs[2192]), .B1(n34), .B2(regs[1680]), .ZN(
        n193) );
  NAND3_X1 U249 ( .A1(n195), .A2(n194), .A3(n193), .ZN(curr_proc_regs[144]) );
  NAND2_X1 U250 ( .A1(regs[657]), .A2(n15), .ZN(n198) );
  AOI22_X1 U251 ( .A1(n29), .A2(regs[1169]), .B1(n21), .B2(regs[145]), .ZN(
        n197) );
  AOI22_X1 U252 ( .A1(win[4]), .A2(regs[2193]), .B1(n9), .B2(regs[1681]), .ZN(
        n196) );
  NAND3_X1 U253 ( .A1(n198), .A2(n197), .A3(n196), .ZN(curr_proc_regs[145]) );
  NAND2_X1 U254 ( .A1(regs[658]), .A2(n15), .ZN(n201) );
  AOI22_X1 U255 ( .A1(n29), .A2(regs[1170]), .B1(n21), .B2(regs[146]), .ZN(
        n200) );
  AOI22_X1 U256 ( .A1(n4), .A2(regs[2194]), .B1(n9), .B2(regs[1682]), .ZN(n199) );
  NAND3_X1 U257 ( .A1(n201), .A2(n200), .A3(n199), .ZN(curr_proc_regs[146]) );
  NAND2_X1 U258 ( .A1(regs[659]), .A2(n15), .ZN(n204) );
  AOI22_X1 U259 ( .A1(n29), .A2(regs[1171]), .B1(n21), .B2(regs[147]), .ZN(
        n203) );
  AOI22_X1 U260 ( .A1(n10), .A2(regs[2195]), .B1(n35), .B2(regs[1683]), .ZN(
        n202) );
  NAND3_X1 U261 ( .A1(n204), .A2(n203), .A3(n202), .ZN(curr_proc_regs[147]) );
  NAND2_X1 U262 ( .A1(regs[660]), .A2(n15), .ZN(n207) );
  AOI22_X1 U263 ( .A1(n29), .A2(regs[1172]), .B1(n21), .B2(regs[148]), .ZN(
        n206) );
  AOI22_X1 U264 ( .A1(n39), .A2(regs[2196]), .B1(n3), .B2(regs[1684]), .ZN(
        n205) );
  NAND3_X1 U265 ( .A1(n207), .A2(n206), .A3(n205), .ZN(curr_proc_regs[148]) );
  NAND2_X1 U266 ( .A1(regs[661]), .A2(n15), .ZN(n210) );
  AOI22_X1 U267 ( .A1(n29), .A2(regs[1173]), .B1(n21), .B2(regs[149]), .ZN(
        n209) );
  AOI22_X1 U268 ( .A1(n4), .A2(regs[2197]), .B1(n3), .B2(regs[1685]), .ZN(n208) );
  NAND3_X1 U269 ( .A1(n210), .A2(n209), .A3(n208), .ZN(curr_proc_regs[149]) );
  NAND2_X1 U270 ( .A1(regs[526]), .A2(n17), .ZN(n213) );
  AOI22_X1 U271 ( .A1(n29), .A2(regs[1038]), .B1(n22), .B2(regs[14]), .ZN(n212) );
  AOI22_X1 U272 ( .A1(n10), .A2(regs[2062]), .B1(n33), .B2(regs[1550]), .ZN(
        n211) );
  NAND3_X1 U273 ( .A1(n213), .A2(n212), .A3(n211), .ZN(curr_proc_regs[14]) );
  NAND2_X1 U274 ( .A1(regs[662]), .A2(n11), .ZN(n216) );
  AOI22_X1 U275 ( .A1(n29), .A2(regs[1174]), .B1(n1580), .B2(regs[150]), .ZN(
        n215) );
  AOI22_X1 U276 ( .A1(n10), .A2(regs[2198]), .B1(n9), .B2(regs[1686]), .ZN(
        n214) );
  NAND3_X1 U277 ( .A1(n216), .A2(n215), .A3(n214), .ZN(curr_proc_regs[150]) );
  NAND2_X1 U278 ( .A1(regs[663]), .A2(n17), .ZN(n219) );
  AOI22_X1 U279 ( .A1(n29), .A2(regs[1175]), .B1(n26), .B2(regs[151]), .ZN(
        n218) );
  AOI22_X1 U280 ( .A1(n10), .A2(regs[2199]), .B1(n9), .B2(regs[1687]), .ZN(
        n217) );
  NAND3_X1 U281 ( .A1(n219), .A2(n218), .A3(n217), .ZN(curr_proc_regs[151]) );
  NAND2_X1 U282 ( .A1(regs[664]), .A2(n11), .ZN(n222) );
  AOI22_X1 U283 ( .A1(n29), .A2(regs[1176]), .B1(n1580), .B2(regs[152]), .ZN(
        n221) );
  AOI22_X1 U284 ( .A1(n10), .A2(regs[2200]), .B1(n35), .B2(regs[1688]), .ZN(
        n220) );
  NAND3_X1 U285 ( .A1(n222), .A2(n221), .A3(n220), .ZN(curr_proc_regs[152]) );
  NAND2_X1 U286 ( .A1(regs[665]), .A2(n17), .ZN(n225) );
  AOI22_X1 U287 ( .A1(n29), .A2(regs[1177]), .B1(n24), .B2(regs[153]), .ZN(
        n224) );
  AOI22_X1 U288 ( .A1(n10), .A2(regs[2201]), .B1(n3), .B2(regs[1689]), .ZN(
        n223) );
  NAND3_X1 U289 ( .A1(n225), .A2(n224), .A3(n223), .ZN(curr_proc_regs[153]) );
  NAND2_X1 U290 ( .A1(regs[666]), .A2(n11), .ZN(n228) );
  AOI22_X1 U291 ( .A1(n29), .A2(regs[1178]), .B1(n21), .B2(regs[154]), .ZN(
        n227) );
  AOI22_X1 U292 ( .A1(n10), .A2(regs[2202]), .B1(n3), .B2(regs[1690]), .ZN(
        n226) );
  NAND3_X1 U293 ( .A1(n228), .A2(n227), .A3(n226), .ZN(curr_proc_regs[154]) );
  NAND2_X1 U294 ( .A1(regs[667]), .A2(n17), .ZN(n231) );
  AOI22_X1 U295 ( .A1(n29), .A2(regs[1179]), .B1(n22), .B2(regs[155]), .ZN(
        n230) );
  AOI22_X1 U296 ( .A1(n10), .A2(regs[2203]), .B1(n34), .B2(regs[1691]), .ZN(
        n229) );
  NAND3_X1 U297 ( .A1(n231), .A2(n230), .A3(n229), .ZN(curr_proc_regs[155]) );
  NAND2_X1 U298 ( .A1(regs[668]), .A2(n11), .ZN(n234) );
  AOI22_X1 U299 ( .A1(n29), .A2(regs[1180]), .B1(n1580), .B2(regs[156]), .ZN(
        n233) );
  AOI22_X1 U300 ( .A1(n39), .A2(regs[2204]), .B1(n33), .B2(regs[1692]), .ZN(
        n232) );
  NAND3_X1 U301 ( .A1(n234), .A2(n233), .A3(n232), .ZN(curr_proc_regs[156]) );
  NAND2_X1 U302 ( .A1(regs[669]), .A2(n17), .ZN(n237) );
  AOI22_X1 U303 ( .A1(n29), .A2(regs[1181]), .B1(n5), .B2(regs[157]), .ZN(n236) );
  AOI22_X1 U304 ( .A1(n10), .A2(regs[2205]), .B1(n34), .B2(regs[1693]), .ZN(
        n235) );
  NAND3_X1 U305 ( .A1(n237), .A2(n236), .A3(n235), .ZN(curr_proc_regs[157]) );
  NAND2_X1 U306 ( .A1(regs[670]), .A2(n11), .ZN(n240) );
  AOI22_X1 U307 ( .A1(n29), .A2(regs[1182]), .B1(n24), .B2(regs[158]), .ZN(
        n239) );
  AOI22_X1 U308 ( .A1(n10), .A2(regs[2206]), .B1(n9), .B2(regs[1694]), .ZN(
        n238) );
  NAND3_X1 U309 ( .A1(n240), .A2(n239), .A3(n238), .ZN(curr_proc_regs[158]) );
  NAND2_X1 U310 ( .A1(regs[671]), .A2(n16), .ZN(n243) );
  AOI22_X1 U311 ( .A1(n29), .A2(regs[1183]), .B1(n1580), .B2(regs[159]), .ZN(
        n242) );
  AOI22_X1 U312 ( .A1(n10), .A2(regs[2207]), .B1(n9), .B2(regs[1695]), .ZN(
        n241) );
  NAND3_X1 U313 ( .A1(n243), .A2(n242), .A3(n241), .ZN(curr_proc_regs[159]) );
  NAND2_X1 U314 ( .A1(regs[527]), .A2(n13), .ZN(n246) );
  AOI22_X1 U315 ( .A1(n29), .A2(regs[1039]), .B1(n22), .B2(regs[15]), .ZN(n245) );
  AOI22_X1 U316 ( .A1(n40), .A2(regs[2063]), .B1(n31), .B2(regs[1551]), .ZN(
        n244) );
  NAND3_X1 U317 ( .A1(n246), .A2(n245), .A3(n244), .ZN(curr_proc_regs[15]) );
  NAND2_X1 U318 ( .A1(regs[672]), .A2(n13), .ZN(n249) );
  AOI22_X1 U319 ( .A1(n29), .A2(regs[1184]), .B1(n22), .B2(regs[160]), .ZN(
        n248) );
  AOI22_X1 U320 ( .A1(n40), .A2(regs[2208]), .B1(n31), .B2(regs[1696]), .ZN(
        n247) );
  NAND3_X1 U321 ( .A1(n249), .A2(n248), .A3(n247), .ZN(curr_proc_regs[160]) );
  NAND2_X1 U322 ( .A1(regs[673]), .A2(n13), .ZN(n252) );
  AOI22_X1 U323 ( .A1(n29), .A2(regs[1185]), .B1(n22), .B2(regs[161]), .ZN(
        n251) );
  AOI22_X1 U324 ( .A1(n40), .A2(regs[2209]), .B1(n3), .B2(regs[1697]), .ZN(
        n250) );
  NAND3_X1 U325 ( .A1(n252), .A2(n251), .A3(n250), .ZN(curr_proc_regs[161]) );
  NAND2_X1 U326 ( .A1(regs[674]), .A2(n13), .ZN(n255) );
  AOI22_X1 U327 ( .A1(n29), .A2(regs[1186]), .B1(n22), .B2(regs[162]), .ZN(
        n254) );
  AOI22_X1 U328 ( .A1(n40), .A2(regs[2210]), .B1(n2), .B2(regs[1698]), .ZN(
        n253) );
  NAND3_X1 U329 ( .A1(n255), .A2(n254), .A3(n253), .ZN(curr_proc_regs[162]) );
  NAND2_X1 U330 ( .A1(regs[675]), .A2(n13), .ZN(n258) );
  AOI22_X1 U331 ( .A1(n29), .A2(regs[1187]), .B1(n22), .B2(regs[163]), .ZN(
        n257) );
  AOI22_X1 U332 ( .A1(n40), .A2(regs[2211]), .B1(n31), .B2(regs[1699]), .ZN(
        n256) );
  NAND3_X1 U333 ( .A1(n258), .A2(n257), .A3(n256), .ZN(curr_proc_regs[163]) );
  NAND2_X1 U334 ( .A1(regs[676]), .A2(n13), .ZN(n261) );
  AOI22_X1 U335 ( .A1(n29), .A2(regs[1188]), .B1(n22), .B2(regs[164]), .ZN(
        n260) );
  AOI22_X1 U336 ( .A1(n40), .A2(regs[2212]), .B1(n31), .B2(regs[1700]), .ZN(
        n259) );
  NAND3_X1 U337 ( .A1(n261), .A2(n260), .A3(n259), .ZN(curr_proc_regs[164]) );
  NAND2_X1 U338 ( .A1(regs[677]), .A2(n13), .ZN(n264) );
  AOI22_X1 U339 ( .A1(n29), .A2(regs[1189]), .B1(n22), .B2(regs[165]), .ZN(
        n263) );
  AOI22_X1 U340 ( .A1(n40), .A2(regs[2213]), .B1(n34), .B2(regs[1701]), .ZN(
        n262) );
  NAND3_X1 U341 ( .A1(n264), .A2(n263), .A3(n262), .ZN(curr_proc_regs[165]) );
  NAND2_X1 U342 ( .A1(regs[678]), .A2(n13), .ZN(n267) );
  AOI22_X1 U343 ( .A1(n29), .A2(regs[1190]), .B1(n22), .B2(regs[166]), .ZN(
        n266) );
  AOI22_X1 U344 ( .A1(n40), .A2(regs[2214]), .B1(n2), .B2(regs[1702]), .ZN(
        n265) );
  NAND3_X1 U345 ( .A1(n267), .A2(n266), .A3(n265), .ZN(curr_proc_regs[166]) );
  NAND2_X1 U346 ( .A1(regs[679]), .A2(n13), .ZN(n270) );
  AOI22_X1 U347 ( .A1(n29), .A2(regs[1191]), .B1(n22), .B2(regs[167]), .ZN(
        n269) );
  AOI22_X1 U348 ( .A1(n40), .A2(regs[2215]), .B1(n31), .B2(regs[1703]), .ZN(
        n268) );
  NAND3_X1 U349 ( .A1(n270), .A2(n269), .A3(n268), .ZN(curr_proc_regs[167]) );
  NAND2_X1 U350 ( .A1(regs[680]), .A2(n13), .ZN(n273) );
  AOI22_X1 U351 ( .A1(n29), .A2(regs[1192]), .B1(n22), .B2(regs[168]), .ZN(
        n272) );
  AOI22_X1 U352 ( .A1(n40), .A2(regs[2216]), .B1(n31), .B2(regs[1704]), .ZN(
        n271) );
  NAND3_X1 U353 ( .A1(n273), .A2(n272), .A3(n271), .ZN(curr_proc_regs[168]) );
  NAND2_X1 U354 ( .A1(regs[681]), .A2(n13), .ZN(n276) );
  AOI22_X1 U355 ( .A1(n29), .A2(regs[1193]), .B1(n22), .B2(regs[169]), .ZN(
        n275) );
  AOI22_X1 U356 ( .A1(n40), .A2(regs[2217]), .B1(n9), .B2(regs[1705]), .ZN(
        n274) );
  NAND3_X1 U357 ( .A1(n276), .A2(n275), .A3(n274), .ZN(curr_proc_regs[169]) );
  NAND2_X1 U358 ( .A1(regs[528]), .A2(n16), .ZN(n279) );
  AOI22_X1 U359 ( .A1(n29), .A2(regs[1040]), .B1(n28), .B2(regs[16]), .ZN(n278) );
  AOI22_X1 U360 ( .A1(n39), .A2(regs[2064]), .B1(n2), .B2(regs[1552]), .ZN(
        n277) );
  NAND3_X1 U361 ( .A1(n279), .A2(n278), .A3(n277), .ZN(curr_proc_regs[16]) );
  NAND2_X1 U362 ( .A1(regs[682]), .A2(n16), .ZN(n282) );
  AOI22_X1 U363 ( .A1(n29), .A2(regs[1194]), .B1(n1580), .B2(regs[170]), .ZN(
        n281) );
  AOI22_X1 U364 ( .A1(n39), .A2(regs[2218]), .B1(n2), .B2(regs[1706]), .ZN(
        n280) );
  NAND3_X1 U365 ( .A1(n282), .A2(n281), .A3(n280), .ZN(curr_proc_regs[170]) );
  NAND2_X1 U366 ( .A1(regs[683]), .A2(n16), .ZN(n285) );
  AOI22_X1 U367 ( .A1(n29), .A2(regs[1195]), .B1(n1580), .B2(regs[171]), .ZN(
        n284) );
  AOI22_X1 U368 ( .A1(n39), .A2(regs[2219]), .B1(n2), .B2(regs[1707]), .ZN(
        n283) );
  NAND3_X1 U369 ( .A1(n285), .A2(n284), .A3(n283), .ZN(curr_proc_regs[171]) );
  NAND2_X1 U370 ( .A1(regs[684]), .A2(n16), .ZN(n288) );
  AOI22_X1 U371 ( .A1(n29), .A2(regs[1196]), .B1(n12), .B2(regs[172]), .ZN(
        n287) );
  AOI22_X1 U372 ( .A1(n39), .A2(regs[2220]), .B1(n2), .B2(regs[1708]), .ZN(
        n286) );
  NAND3_X1 U373 ( .A1(n288), .A2(n287), .A3(n286), .ZN(curr_proc_regs[172]) );
  NAND2_X1 U374 ( .A1(regs[685]), .A2(n16), .ZN(n291) );
  AOI22_X1 U375 ( .A1(n29), .A2(regs[1197]), .B1(n22), .B2(regs[173]), .ZN(
        n290) );
  AOI22_X1 U376 ( .A1(n39), .A2(regs[2221]), .B1(n2), .B2(regs[1709]), .ZN(
        n289) );
  NAND3_X1 U377 ( .A1(n291), .A2(n290), .A3(n289), .ZN(curr_proc_regs[173]) );
  NAND2_X1 U378 ( .A1(regs[686]), .A2(n16), .ZN(n294) );
  AOI22_X1 U379 ( .A1(n29), .A2(regs[1198]), .B1(n25), .B2(regs[174]), .ZN(
        n293) );
  AOI22_X1 U380 ( .A1(n39), .A2(regs[2222]), .B1(n2), .B2(regs[1710]), .ZN(
        n292) );
  NAND3_X1 U381 ( .A1(n294), .A2(n293), .A3(n292), .ZN(curr_proc_regs[174]) );
  NAND2_X1 U382 ( .A1(regs[687]), .A2(n16), .ZN(n297) );
  AOI22_X1 U383 ( .A1(n29), .A2(regs[1199]), .B1(n12), .B2(regs[175]), .ZN(
        n296) );
  AOI22_X1 U384 ( .A1(n39), .A2(regs[2223]), .B1(n2), .B2(regs[1711]), .ZN(
        n295) );
  NAND3_X1 U385 ( .A1(n297), .A2(n296), .A3(n295), .ZN(curr_proc_regs[175]) );
  NAND2_X1 U386 ( .A1(regs[688]), .A2(n16), .ZN(n300) );
  AOI22_X1 U387 ( .A1(n29), .A2(regs[1200]), .B1(n28), .B2(regs[176]), .ZN(
        n299) );
  AOI22_X1 U388 ( .A1(n39), .A2(regs[2224]), .B1(n2), .B2(regs[1712]), .ZN(
        n298) );
  NAND3_X1 U389 ( .A1(n300), .A2(n299), .A3(n298), .ZN(curr_proc_regs[176]) );
  NAND2_X1 U390 ( .A1(regs[689]), .A2(n16), .ZN(n303) );
  AOI22_X1 U391 ( .A1(n29), .A2(regs[1201]), .B1(n28), .B2(regs[177]), .ZN(
        n302) );
  AOI22_X1 U392 ( .A1(n39), .A2(regs[2225]), .B1(n2), .B2(regs[1713]), .ZN(
        n301) );
  NAND3_X1 U393 ( .A1(n303), .A2(n302), .A3(n301), .ZN(curr_proc_regs[177]) );
  NAND2_X1 U394 ( .A1(regs[690]), .A2(n16), .ZN(n306) );
  AOI22_X1 U395 ( .A1(n29), .A2(regs[1202]), .B1(n21), .B2(regs[178]), .ZN(
        n305) );
  AOI22_X1 U396 ( .A1(n39), .A2(regs[2226]), .B1(n2), .B2(regs[1714]), .ZN(
        n304) );
  NAND3_X1 U397 ( .A1(n306), .A2(n305), .A3(n304), .ZN(curr_proc_regs[178]) );
  NAND2_X1 U398 ( .A1(regs[691]), .A2(n16), .ZN(n309) );
  AOI22_X1 U399 ( .A1(n29), .A2(regs[1203]), .B1(n28), .B2(regs[179]), .ZN(
        n308) );
  AOI22_X1 U400 ( .A1(n39), .A2(regs[2227]), .B1(n2), .B2(regs[1715]), .ZN(
        n307) );
  NAND3_X1 U401 ( .A1(n309), .A2(n308), .A3(n307), .ZN(curr_proc_regs[179]) );
  NAND2_X1 U402 ( .A1(regs[529]), .A2(n17), .ZN(n312) );
  AOI22_X1 U403 ( .A1(n29), .A2(regs[1041]), .B1(n21), .B2(regs[17]), .ZN(n311) );
  AOI22_X1 U404 ( .A1(n38), .A2(regs[2065]), .B1(n9), .B2(regs[1553]), .ZN(
        n310) );
  NAND3_X1 U405 ( .A1(n312), .A2(n311), .A3(n310), .ZN(curr_proc_regs[17]) );
  NAND2_X1 U406 ( .A1(regs[692]), .A2(n17), .ZN(n315) );
  AOI22_X1 U407 ( .A1(n29), .A2(regs[1204]), .B1(n25), .B2(regs[180]), .ZN(
        n314) );
  AOI22_X1 U408 ( .A1(n38), .A2(regs[2228]), .B1(n9), .B2(regs[1716]), .ZN(
        n313) );
  NAND3_X1 U409 ( .A1(n315), .A2(n314), .A3(n313), .ZN(curr_proc_regs[180]) );
  NAND2_X1 U410 ( .A1(regs[693]), .A2(n17), .ZN(n318) );
  AOI22_X1 U411 ( .A1(n29), .A2(regs[1205]), .B1(n12), .B2(regs[181]), .ZN(
        n317) );
  AOI22_X1 U412 ( .A1(n38), .A2(regs[2229]), .B1(n35), .B2(regs[1717]), .ZN(
        n316) );
  NAND3_X1 U413 ( .A1(n318), .A2(n317), .A3(n316), .ZN(curr_proc_regs[181]) );
  NAND2_X1 U414 ( .A1(regs[694]), .A2(n17), .ZN(n321) );
  AOI22_X1 U415 ( .A1(n29), .A2(regs[1206]), .B1(n21), .B2(regs[182]), .ZN(
        n320) );
  AOI22_X1 U416 ( .A1(n38), .A2(regs[2230]), .B1(n30), .B2(regs[1718]), .ZN(
        n319) );
  NAND3_X1 U417 ( .A1(n321), .A2(n320), .A3(n319), .ZN(curr_proc_regs[182]) );
  NAND2_X1 U418 ( .A1(regs[695]), .A2(n17), .ZN(n324) );
  AOI22_X1 U419 ( .A1(n29), .A2(regs[1207]), .B1(n22), .B2(regs[183]), .ZN(
        n323) );
  AOI22_X1 U420 ( .A1(n38), .A2(regs[2231]), .B1(n3), .B2(regs[1719]), .ZN(
        n322) );
  NAND3_X1 U421 ( .A1(n324), .A2(n323), .A3(n322), .ZN(curr_proc_regs[183]) );
  NAND2_X1 U422 ( .A1(regs[696]), .A2(n17), .ZN(n327) );
  AOI22_X1 U423 ( .A1(n29), .A2(regs[1208]), .B1(n1580), .B2(regs[184]), .ZN(
        n326) );
  AOI22_X1 U424 ( .A1(n38), .A2(regs[2232]), .B1(n30), .B2(regs[1720]), .ZN(
        n325) );
  NAND3_X1 U425 ( .A1(n327), .A2(n326), .A3(n325), .ZN(curr_proc_regs[184]) );
  NAND2_X1 U426 ( .A1(regs[697]), .A2(n17), .ZN(n330) );
  AOI22_X1 U427 ( .A1(n29), .A2(regs[1209]), .B1(n5), .B2(regs[185]), .ZN(n329) );
  AOI22_X1 U428 ( .A1(n38), .A2(regs[2233]), .B1(n3), .B2(regs[1721]), .ZN(
        n328) );
  NAND3_X1 U429 ( .A1(n330), .A2(n329), .A3(n328), .ZN(curr_proc_regs[185]) );
  NAND2_X1 U430 ( .A1(regs[698]), .A2(n17), .ZN(n333) );
  AOI22_X1 U431 ( .A1(n29), .A2(regs[1210]), .B1(n5), .B2(regs[186]), .ZN(n332) );
  AOI22_X1 U432 ( .A1(n38), .A2(regs[2234]), .B1(n30), .B2(regs[1722]), .ZN(
        n331) );
  NAND3_X1 U433 ( .A1(n333), .A2(n332), .A3(n331), .ZN(curr_proc_regs[186]) );
  NAND2_X1 U434 ( .A1(regs[699]), .A2(n17), .ZN(n336) );
  AOI22_X1 U435 ( .A1(n29), .A2(regs[1211]), .B1(n12), .B2(regs[187]), .ZN(
        n335) );
  AOI22_X1 U436 ( .A1(n38), .A2(regs[2235]), .B1(n34), .B2(regs[1723]), .ZN(
        n334) );
  NAND3_X1 U437 ( .A1(n336), .A2(n335), .A3(n334), .ZN(curr_proc_regs[187]) );
  NAND2_X1 U438 ( .A1(regs[700]), .A2(n17), .ZN(n339) );
  AOI22_X1 U439 ( .A1(n29), .A2(regs[1212]), .B1(n21), .B2(regs[188]), .ZN(
        n338) );
  AOI22_X1 U440 ( .A1(n38), .A2(regs[2236]), .B1(n30), .B2(regs[1724]), .ZN(
        n337) );
  NAND3_X1 U441 ( .A1(n339), .A2(n338), .A3(n337), .ZN(curr_proc_regs[188]) );
  NAND2_X1 U442 ( .A1(regs[701]), .A2(n17), .ZN(n342) );
  AOI22_X1 U443 ( .A1(n29), .A2(regs[1213]), .B1(n5), .B2(regs[189]), .ZN(n341) );
  AOI22_X1 U444 ( .A1(n38), .A2(regs[2237]), .B1(n33), .B2(regs[1725]), .ZN(
        n340) );
  NAND3_X1 U445 ( .A1(n342), .A2(n341), .A3(n340), .ZN(curr_proc_regs[189]) );
  NAND2_X1 U446 ( .A1(regs[530]), .A2(n18), .ZN(n345) );
  AOI22_X1 U447 ( .A1(n29), .A2(regs[1042]), .B1(n1580), .B2(regs[18]), .ZN(
        n344) );
  AOI22_X1 U448 ( .A1(n37), .A2(regs[2066]), .B1(n31), .B2(regs[1554]), .ZN(
        n343) );
  NAND3_X1 U449 ( .A1(n345), .A2(n344), .A3(n343), .ZN(curr_proc_regs[18]) );
  NAND2_X1 U450 ( .A1(regs[702]), .A2(n18), .ZN(n348) );
  AOI22_X1 U451 ( .A1(n29), .A2(regs[1214]), .B1(n12), .B2(regs[190]), .ZN(
        n347) );
  AOI22_X1 U452 ( .A1(n37), .A2(regs[2238]), .B1(n33), .B2(regs[1726]), .ZN(
        n346) );
  NAND3_X1 U453 ( .A1(n348), .A2(n347), .A3(n346), .ZN(curr_proc_regs[190]) );
  NAND2_X1 U454 ( .A1(regs[703]), .A2(n18), .ZN(n351) );
  AOI22_X1 U455 ( .A1(n29), .A2(regs[1215]), .B1(n22), .B2(regs[191]), .ZN(
        n350) );
  AOI22_X1 U456 ( .A1(n37), .A2(regs[2239]), .B1(n9), .B2(regs[1727]), .ZN(
        n349) );
  NAND3_X1 U457 ( .A1(n351), .A2(n350), .A3(n349), .ZN(curr_proc_regs[191]) );
  NAND2_X1 U458 ( .A1(regs[704]), .A2(n18), .ZN(n354) );
  AOI22_X1 U459 ( .A1(n29), .A2(regs[1216]), .B1(n25), .B2(regs[192]), .ZN(
        n353) );
  AOI22_X1 U460 ( .A1(n37), .A2(regs[2240]), .B1(n9), .B2(regs[1728]), .ZN(
        n352) );
  NAND3_X1 U461 ( .A1(n354), .A2(n353), .A3(n352), .ZN(curr_proc_regs[192]) );
  NAND2_X1 U462 ( .A1(regs[705]), .A2(n18), .ZN(n357) );
  AOI22_X1 U463 ( .A1(n29), .A2(regs[1217]), .B1(n12), .B2(regs[193]), .ZN(
        n356) );
  AOI22_X1 U464 ( .A1(n37), .A2(regs[2241]), .B1(n35), .B2(regs[1729]), .ZN(
        n355) );
  NAND3_X1 U465 ( .A1(n357), .A2(n356), .A3(n355), .ZN(curr_proc_regs[193]) );
  NAND2_X1 U466 ( .A1(regs[706]), .A2(n18), .ZN(n360) );
  AOI22_X1 U467 ( .A1(n29), .A2(regs[1218]), .B1(n28), .B2(regs[194]), .ZN(
        n359) );
  AOI22_X1 U468 ( .A1(n37), .A2(regs[2242]), .B1(n3), .B2(regs[1730]), .ZN(
        n358) );
  NAND3_X1 U469 ( .A1(n360), .A2(n359), .A3(n358), .ZN(curr_proc_regs[194]) );
  NAND2_X1 U470 ( .A1(regs[707]), .A2(n18), .ZN(n363) );
  AOI22_X1 U471 ( .A1(n29), .A2(regs[1219]), .B1(n21), .B2(regs[195]), .ZN(
        n362) );
  AOI22_X1 U472 ( .A1(n37), .A2(regs[2243]), .B1(n3), .B2(regs[1731]), .ZN(
        n361) );
  NAND3_X1 U473 ( .A1(n363), .A2(n362), .A3(n361), .ZN(curr_proc_regs[195]) );
  NAND2_X1 U474 ( .A1(regs[708]), .A2(n18), .ZN(n366) );
  AOI22_X1 U475 ( .A1(n29), .A2(regs[1220]), .B1(n24), .B2(regs[196]), .ZN(
        n365) );
  AOI22_X1 U476 ( .A1(n37), .A2(regs[2244]), .B1(n34), .B2(regs[1732]), .ZN(
        n364) );
  NAND3_X1 U477 ( .A1(n366), .A2(n365), .A3(n364), .ZN(curr_proc_regs[196]) );
  NAND2_X1 U478 ( .A1(regs[709]), .A2(n18), .ZN(n369) );
  AOI22_X1 U479 ( .A1(n29), .A2(regs[1221]), .B1(n28), .B2(regs[197]), .ZN(
        n368) );
  AOI22_X1 U480 ( .A1(n37), .A2(regs[2245]), .B1(n2), .B2(regs[1733]), .ZN(
        n367) );
  NAND3_X1 U481 ( .A1(n369), .A2(n368), .A3(n367), .ZN(curr_proc_regs[197]) );
  NAND2_X1 U482 ( .A1(regs[710]), .A2(n18), .ZN(n372) );
  AOI22_X1 U483 ( .A1(n29), .A2(regs[1222]), .B1(n12), .B2(regs[198]), .ZN(
        n371) );
  AOI22_X1 U484 ( .A1(n37), .A2(regs[2246]), .B1(n33), .B2(regs[1734]), .ZN(
        n370) );
  NAND3_X1 U485 ( .A1(n372), .A2(n371), .A3(n370), .ZN(curr_proc_regs[198]) );
  NAND2_X1 U486 ( .A1(regs[711]), .A2(n18), .ZN(n375) );
  AOI22_X1 U487 ( .A1(n29), .A2(regs[1223]), .B1(n5), .B2(regs[199]), .ZN(n374) );
  AOI22_X1 U488 ( .A1(n37), .A2(regs[2247]), .B1(n9), .B2(regs[1735]), .ZN(
        n373) );
  NAND3_X1 U489 ( .A1(n375), .A2(n374), .A3(n373), .ZN(curr_proc_regs[199]) );
  NAND2_X1 U490 ( .A1(regs[531]), .A2(n19), .ZN(n378) );
  AOI22_X1 U491 ( .A1(n29), .A2(regs[1043]), .B1(n25), .B2(regs[19]), .ZN(n377) );
  AOI22_X1 U492 ( .A1(n41), .A2(regs[2067]), .B1(n32), .B2(regs[1555]), .ZN(
        n376) );
  NAND3_X1 U493 ( .A1(n378), .A2(n377), .A3(n376), .ZN(curr_proc_regs[19]) );
  NAND2_X1 U494 ( .A1(regs[513]), .A2(n19), .ZN(n381) );
  AOI22_X1 U495 ( .A1(n29), .A2(regs[1025]), .B1(n24), .B2(regs[1]), .ZN(n380)
         );
  AOI22_X1 U496 ( .A1(n1), .A2(regs[2049]), .B1(n9), .B2(regs[1537]), .ZN(n379) );
  NAND3_X1 U497 ( .A1(n381), .A2(n380), .A3(n379), .ZN(curr_proc_regs[1]) );
  NAND2_X1 U498 ( .A1(regs[712]), .A2(n19), .ZN(n384) );
  AOI22_X1 U499 ( .A1(n29), .A2(regs[1224]), .B1(n21), .B2(regs[200]), .ZN(
        n383) );
  AOI22_X1 U500 ( .A1(n10), .A2(regs[2248]), .B1(n32), .B2(regs[1736]), .ZN(
        n382) );
  NAND3_X1 U501 ( .A1(n384), .A2(n383), .A3(n382), .ZN(curr_proc_regs[200]) );
  NAND2_X1 U502 ( .A1(regs[713]), .A2(n19), .ZN(n387) );
  AOI22_X1 U503 ( .A1(n29), .A2(regs[1225]), .B1(n12), .B2(regs[201]), .ZN(
        n386) );
  AOI22_X1 U504 ( .A1(n4), .A2(regs[2249]), .B1(n9), .B2(regs[1737]), .ZN(n385) );
  NAND3_X1 U505 ( .A1(n387), .A2(n386), .A3(n385), .ZN(curr_proc_regs[201]) );
  NAND2_X1 U506 ( .A1(regs[714]), .A2(n19), .ZN(n390) );
  AOI22_X1 U507 ( .A1(n29), .A2(regs[1226]), .B1(n5), .B2(regs[202]), .ZN(n389) );
  AOI22_X1 U508 ( .A1(n37), .A2(regs[2250]), .B1(n32), .B2(regs[1738]), .ZN(
        n388) );
  NAND3_X1 U509 ( .A1(n390), .A2(n389), .A3(n388), .ZN(curr_proc_regs[202]) );
  NAND2_X1 U510 ( .A1(regs[715]), .A2(n19), .ZN(n393) );
  AOI22_X1 U511 ( .A1(n29), .A2(regs[1227]), .B1(n28), .B2(regs[203]), .ZN(
        n392) );
  AOI22_X1 U512 ( .A1(n39), .A2(regs[2251]), .B1(n35), .B2(regs[1739]), .ZN(
        n391) );
  NAND3_X1 U513 ( .A1(n393), .A2(n392), .A3(n391), .ZN(curr_proc_regs[203]) );
  NAND2_X1 U514 ( .A1(regs[716]), .A2(n19), .ZN(n396) );
  AOI22_X1 U515 ( .A1(n29), .A2(regs[1228]), .B1(n24), .B2(regs[204]), .ZN(
        n395) );
  AOI22_X1 U516 ( .A1(n8), .A2(regs[2252]), .B1(n32), .B2(regs[1740]), .ZN(
        n394) );
  NAND3_X1 U517 ( .A1(n396), .A2(n395), .A3(n394), .ZN(curr_proc_regs[204]) );
  NAND2_X1 U518 ( .A1(regs[717]), .A2(n19), .ZN(n399) );
  AOI22_X1 U519 ( .A1(n29), .A2(regs[1229]), .B1(n5), .B2(regs[205]), .ZN(n398) );
  AOI22_X1 U520 ( .A1(n41), .A2(regs[2253]), .B1(n3), .B2(regs[1741]), .ZN(
        n397) );
  NAND3_X1 U521 ( .A1(n399), .A2(n398), .A3(n397), .ZN(curr_proc_regs[205]) );
  NAND2_X1 U522 ( .A1(regs[718]), .A2(n19), .ZN(n402) );
  AOI22_X1 U523 ( .A1(n29), .A2(regs[1230]), .B1(n12), .B2(regs[206]), .ZN(
        n401) );
  AOI22_X1 U524 ( .A1(n1), .A2(regs[2254]), .B1(n32), .B2(regs[1742]), .ZN(
        n400) );
  NAND3_X1 U525 ( .A1(n402), .A2(n401), .A3(n400), .ZN(curr_proc_regs[206]) );
  NAND2_X1 U526 ( .A1(regs[719]), .A2(n19), .ZN(n405) );
  AOI22_X1 U527 ( .A1(n29), .A2(regs[1231]), .B1(n5), .B2(regs[207]), .ZN(n404) );
  AOI22_X1 U528 ( .A1(n10), .A2(regs[2255]), .B1(n3), .B2(regs[1743]), .ZN(
        n403) );
  NAND3_X1 U529 ( .A1(n405), .A2(n404), .A3(n403), .ZN(curr_proc_regs[207]) );
  NAND2_X1 U530 ( .A1(regs[720]), .A2(n19), .ZN(n408) );
  AOI22_X1 U531 ( .A1(n29), .A2(regs[1232]), .B1(n12), .B2(regs[208]), .ZN(
        n407) );
  AOI22_X1 U532 ( .A1(n4), .A2(regs[2256]), .B1(n32), .B2(regs[1744]), .ZN(
        n406) );
  NAND3_X1 U533 ( .A1(n408), .A2(n407), .A3(n406), .ZN(curr_proc_regs[208]) );
  NAND2_X1 U534 ( .A1(regs[721]), .A2(n11), .ZN(n411) );
  AOI22_X1 U535 ( .A1(n29), .A2(regs[1233]), .B1(n28), .B2(regs[209]), .ZN(
        n410) );
  AOI22_X1 U536 ( .A1(n41), .A2(regs[2257]), .B1(n34), .B2(regs[1745]), .ZN(
        n409) );
  NAND3_X1 U537 ( .A1(n411), .A2(n410), .A3(n409), .ZN(curr_proc_regs[209]) );
  NAND2_X1 U538 ( .A1(regs[532]), .A2(n11), .ZN(n414) );
  AOI22_X1 U539 ( .A1(n29), .A2(regs[1044]), .B1(n28), .B2(regs[20]), .ZN(n413) );
  AOI22_X1 U540 ( .A1(n41), .A2(regs[2068]), .B1(n9), .B2(regs[1556]), .ZN(
        n412) );
  NAND3_X1 U541 ( .A1(n414), .A2(n413), .A3(n412), .ZN(curr_proc_regs[20]) );
  NAND2_X1 U542 ( .A1(regs[722]), .A2(n11), .ZN(n417) );
  AOI22_X1 U543 ( .A1(n29), .A2(regs[1234]), .B1(n28), .B2(regs[210]), .ZN(
        n416) );
  AOI22_X1 U544 ( .A1(n41), .A2(regs[2258]), .B1(n9), .B2(regs[1746]), .ZN(
        n415) );
  NAND3_X1 U545 ( .A1(n417), .A2(n416), .A3(n415), .ZN(curr_proc_regs[210]) );
  NAND2_X1 U546 ( .A1(regs[723]), .A2(n11), .ZN(n420) );
  AOI22_X1 U547 ( .A1(n29), .A2(regs[1235]), .B1(n28), .B2(regs[211]), .ZN(
        n419) );
  AOI22_X1 U548 ( .A1(n41), .A2(regs[2259]), .B1(n3), .B2(regs[1747]), .ZN(
        n418) );
  NAND3_X1 U549 ( .A1(n420), .A2(n419), .A3(n418), .ZN(curr_proc_regs[211]) );
  NAND2_X1 U550 ( .A1(regs[724]), .A2(n11), .ZN(n423) );
  AOI22_X1 U551 ( .A1(n29), .A2(regs[1236]), .B1(n28), .B2(regs[212]), .ZN(
        n422) );
  AOI22_X1 U552 ( .A1(n41), .A2(regs[2260]), .B1(n9), .B2(regs[1748]), .ZN(
        n421) );
  NAND3_X1 U553 ( .A1(n423), .A2(n422), .A3(n421), .ZN(curr_proc_regs[212]) );
  NAND2_X1 U554 ( .A1(regs[725]), .A2(n11), .ZN(n426) );
  AOI22_X1 U555 ( .A1(n29), .A2(regs[1237]), .B1(n28), .B2(regs[213]), .ZN(
        n425) );
  AOI22_X1 U556 ( .A1(n41), .A2(regs[2261]), .B1(n34), .B2(regs[1749]), .ZN(
        n424) );
  NAND3_X1 U557 ( .A1(n426), .A2(n425), .A3(n424), .ZN(curr_proc_regs[213]) );
  NAND2_X1 U558 ( .A1(regs[726]), .A2(n11), .ZN(n429) );
  AOI22_X1 U559 ( .A1(n29), .A2(regs[1238]), .B1(n28), .B2(regs[214]), .ZN(
        n428) );
  AOI22_X1 U560 ( .A1(n10), .A2(regs[2262]), .B1(n3), .B2(regs[1750]), .ZN(
        n427) );
  NAND3_X1 U561 ( .A1(n429), .A2(n428), .A3(n427), .ZN(curr_proc_regs[214]) );
  NAND2_X1 U562 ( .A1(regs[727]), .A2(n11), .ZN(n432) );
  AOI22_X1 U563 ( .A1(n29), .A2(regs[1239]), .B1(n28), .B2(regs[215]), .ZN(
        n431) );
  AOI22_X1 U564 ( .A1(win[4]), .A2(regs[2263]), .B1(n35), .B2(regs[1751]), 
        .ZN(n430) );
  NAND3_X1 U565 ( .A1(n432), .A2(n431), .A3(n430), .ZN(curr_proc_regs[215]) );
  NAND2_X1 U566 ( .A1(regs[728]), .A2(n11), .ZN(n435) );
  AOI22_X1 U567 ( .A1(n29), .A2(regs[1240]), .B1(n28), .B2(regs[216]), .ZN(
        n434) );
  AOI22_X1 U568 ( .A1(win[4]), .A2(regs[2264]), .B1(n34), .B2(regs[1752]), 
        .ZN(n433) );
  NAND3_X1 U569 ( .A1(n435), .A2(n434), .A3(n433), .ZN(curr_proc_regs[216]) );
  NAND2_X1 U570 ( .A1(regs[729]), .A2(n11), .ZN(n438) );
  AOI22_X1 U571 ( .A1(n29), .A2(regs[1241]), .B1(n28), .B2(regs[217]), .ZN(
        n437) );
  AOI22_X1 U572 ( .A1(win[4]), .A2(regs[2265]), .B1(n9), .B2(regs[1753]), .ZN(
        n436) );
  NAND3_X1 U573 ( .A1(n438), .A2(n437), .A3(n436), .ZN(curr_proc_regs[217]) );
  NAND2_X1 U574 ( .A1(regs[730]), .A2(n11), .ZN(n441) );
  AOI22_X1 U575 ( .A1(n29), .A2(regs[1242]), .B1(n28), .B2(regs[218]), .ZN(
        n440) );
  AOI22_X1 U576 ( .A1(win[4]), .A2(regs[2266]), .B1(n9), .B2(regs[1754]), .ZN(
        n439) );
  NAND3_X1 U577 ( .A1(n441), .A2(n440), .A3(n439), .ZN(curr_proc_regs[218]) );
  NAND2_X1 U578 ( .A1(regs[731]), .A2(n7), .ZN(n444) );
  AOI22_X1 U579 ( .A1(n29), .A2(regs[1243]), .B1(n28), .B2(regs[219]), .ZN(
        n443) );
  AOI22_X1 U580 ( .A1(win[4]), .A2(regs[2267]), .B1(n31), .B2(regs[1755]), 
        .ZN(n442) );
  NAND3_X1 U581 ( .A1(n444), .A2(n443), .A3(n442), .ZN(curr_proc_regs[219]) );
  NAND2_X1 U582 ( .A1(regs[533]), .A2(n16), .ZN(n447) );
  AOI22_X1 U583 ( .A1(n29), .A2(regs[1045]), .B1(n28), .B2(regs[21]), .ZN(n446) );
  AOI22_X1 U584 ( .A1(win[4]), .A2(regs[2069]), .B1(n31), .B2(regs[1557]), 
        .ZN(n445) );
  NAND3_X1 U585 ( .A1(n447), .A2(n446), .A3(n445), .ZN(curr_proc_regs[21]) );
  NAND2_X1 U586 ( .A1(regs[732]), .A2(n13), .ZN(n450) );
  AOI22_X1 U587 ( .A1(n29), .A2(regs[1244]), .B1(n28), .B2(regs[220]), .ZN(
        n449) );
  AOI22_X1 U588 ( .A1(win[4]), .A2(regs[2268]), .B1(n31), .B2(regs[1756]), 
        .ZN(n448) );
  NAND3_X1 U589 ( .A1(n450), .A2(n449), .A3(n448), .ZN(curr_proc_regs[220]) );
  NAND2_X1 U590 ( .A1(regs[733]), .A2(n11), .ZN(n453) );
  AOI22_X1 U591 ( .A1(n29), .A2(regs[1245]), .B1(n28), .B2(regs[221]), .ZN(
        n452) );
  AOI22_X1 U592 ( .A1(n1), .A2(regs[2269]), .B1(n31), .B2(regs[1757]), .ZN(
        n451) );
  NAND3_X1 U593 ( .A1(n453), .A2(n452), .A3(n451), .ZN(curr_proc_regs[221]) );
  NAND2_X1 U594 ( .A1(regs[734]), .A2(n11), .ZN(n456) );
  AOI22_X1 U595 ( .A1(n29), .A2(regs[1246]), .B1(n28), .B2(regs[222]), .ZN(
        n455) );
  AOI22_X1 U596 ( .A1(n41), .A2(regs[2270]), .B1(n31), .B2(regs[1758]), .ZN(
        n454) );
  NAND3_X1 U597 ( .A1(n456), .A2(n455), .A3(n454), .ZN(curr_proc_regs[222]) );
  NAND2_X1 U598 ( .A1(regs[735]), .A2(n1579), .ZN(n459) );
  AOI22_X1 U599 ( .A1(n29), .A2(regs[1247]), .B1(n28), .B2(regs[223]), .ZN(
        n458) );
  AOI22_X1 U600 ( .A1(n4), .A2(regs[2271]), .B1(n31), .B2(regs[1759]), .ZN(
        n457) );
  NAND3_X1 U601 ( .A1(n459), .A2(n458), .A3(n457), .ZN(curr_proc_regs[223]) );
  NAND2_X1 U602 ( .A1(regs[736]), .A2(n1579), .ZN(n462) );
  AOI22_X1 U603 ( .A1(n29), .A2(regs[1248]), .B1(n28), .B2(regs[224]), .ZN(
        n461) );
  AOI22_X1 U604 ( .A1(n10), .A2(regs[2272]), .B1(n31), .B2(regs[1760]), .ZN(
        n460) );
  NAND3_X1 U605 ( .A1(n462), .A2(n461), .A3(n460), .ZN(curr_proc_regs[224]) );
  NAND2_X1 U606 ( .A1(regs[737]), .A2(n13), .ZN(n465) );
  AOI22_X1 U607 ( .A1(n29), .A2(regs[1249]), .B1(n28), .B2(regs[225]), .ZN(
        n464) );
  AOI22_X1 U608 ( .A1(n39), .A2(regs[2273]), .B1(n31), .B2(regs[1761]), .ZN(
        n463) );
  NAND3_X1 U609 ( .A1(n465), .A2(n464), .A3(n463), .ZN(curr_proc_regs[225]) );
  NAND2_X1 U610 ( .A1(regs[738]), .A2(n1579), .ZN(n468) );
  AOI22_X1 U611 ( .A1(n29), .A2(regs[1250]), .B1(n28), .B2(regs[226]), .ZN(
        n467) );
  AOI22_X1 U612 ( .A1(n37), .A2(regs[2274]), .B1(n31), .B2(regs[1762]), .ZN(
        n466) );
  NAND3_X1 U613 ( .A1(n468), .A2(n467), .A3(n466), .ZN(curr_proc_regs[226]) );
  NAND2_X1 U614 ( .A1(regs[739]), .A2(n14), .ZN(n471) );
  AOI22_X1 U615 ( .A1(n29), .A2(regs[1251]), .B1(n28), .B2(regs[227]), .ZN(
        n470) );
  AOI22_X1 U616 ( .A1(n41), .A2(regs[2275]), .B1(n31), .B2(regs[1763]), .ZN(
        n469) );
  NAND3_X1 U617 ( .A1(n471), .A2(n470), .A3(n469), .ZN(curr_proc_regs[227]) );
  NAND2_X1 U618 ( .A1(regs[740]), .A2(n13), .ZN(n474) );
  AOI22_X1 U619 ( .A1(n29), .A2(regs[1252]), .B1(n28), .B2(regs[228]), .ZN(
        n473) );
  AOI22_X1 U620 ( .A1(n8), .A2(regs[2276]), .B1(n31), .B2(regs[1764]), .ZN(
        n472) );
  NAND3_X1 U621 ( .A1(n474), .A2(n473), .A3(n472), .ZN(curr_proc_regs[228]) );
  NAND2_X1 U622 ( .A1(regs[741]), .A2(n15), .ZN(n477) );
  AOI22_X1 U623 ( .A1(n29), .A2(regs[1253]), .B1(n28), .B2(regs[229]), .ZN(
        n476) );
  AOI22_X1 U624 ( .A1(n41), .A2(regs[2277]), .B1(n3), .B2(regs[1765]), .ZN(
        n475) );
  NAND3_X1 U625 ( .A1(n477), .A2(n476), .A3(n475), .ZN(curr_proc_regs[229]) );
  NAND2_X1 U626 ( .A1(regs[534]), .A2(n15), .ZN(n480) );
  AOI22_X1 U627 ( .A1(n29), .A2(regs[1046]), .B1(n28), .B2(regs[22]), .ZN(n479) );
  AOI22_X1 U628 ( .A1(n1), .A2(regs[2070]), .B1(n3), .B2(regs[1558]), .ZN(n478) );
  NAND3_X1 U629 ( .A1(n480), .A2(n479), .A3(n478), .ZN(curr_proc_regs[22]) );
  NAND2_X1 U630 ( .A1(regs[742]), .A2(n15), .ZN(n483) );
  AOI22_X1 U631 ( .A1(n29), .A2(regs[1254]), .B1(n28), .B2(regs[230]), .ZN(
        n482) );
  AOI22_X1 U632 ( .A1(n1), .A2(regs[2278]), .B1(n34), .B2(regs[1766]), .ZN(
        n481) );
  NAND3_X1 U633 ( .A1(n483), .A2(n482), .A3(n481), .ZN(curr_proc_regs[230]) );
  NAND2_X1 U634 ( .A1(regs[743]), .A2(n15), .ZN(n486) );
  AOI22_X1 U635 ( .A1(n29), .A2(regs[1255]), .B1(n28), .B2(regs[231]), .ZN(
        n485) );
  AOI22_X1 U636 ( .A1(n41), .A2(regs[2279]), .B1(n1582), .B2(regs[1767]), .ZN(
        n484) );
  NAND3_X1 U637 ( .A1(n486), .A2(n485), .A3(n484), .ZN(curr_proc_regs[231]) );
  NAND2_X1 U638 ( .A1(regs[744]), .A2(n15), .ZN(n489) );
  AOI22_X1 U639 ( .A1(n29), .A2(regs[1256]), .B1(n28), .B2(regs[232]), .ZN(
        n488) );
  AOI22_X1 U640 ( .A1(n1), .A2(regs[2280]), .B1(n33), .B2(regs[1768]), .ZN(
        n487) );
  NAND3_X1 U641 ( .A1(n489), .A2(n488), .A3(n487), .ZN(curr_proc_regs[232]) );
  NAND2_X1 U642 ( .A1(regs[745]), .A2(n15), .ZN(n492) );
  AOI22_X1 U643 ( .A1(n29), .A2(regs[1257]), .B1(n28), .B2(regs[233]), .ZN(
        n491) );
  AOI22_X1 U644 ( .A1(n1), .A2(regs[2281]), .B1(n9), .B2(regs[1769]), .ZN(n490) );
  NAND3_X1 U645 ( .A1(n492), .A2(n491), .A3(n490), .ZN(curr_proc_regs[233]) );
  NAND2_X1 U646 ( .A1(regs[746]), .A2(n15), .ZN(n495) );
  AOI22_X1 U647 ( .A1(n29), .A2(regs[1258]), .B1(n28), .B2(regs[234]), .ZN(
        n494) );
  AOI22_X1 U648 ( .A1(n1), .A2(regs[2282]), .B1(n9), .B2(regs[1770]), .ZN(n493) );
  NAND3_X1 U649 ( .A1(n495), .A2(n494), .A3(n493), .ZN(curr_proc_regs[234]) );
  NAND2_X1 U650 ( .A1(regs[747]), .A2(n15), .ZN(n498) );
  AOI22_X1 U651 ( .A1(n29), .A2(regs[1259]), .B1(n28), .B2(regs[235]), .ZN(
        n497) );
  AOI22_X1 U652 ( .A1(n1), .A2(regs[2283]), .B1(n35), .B2(regs[1771]), .ZN(
        n496) );
  NAND3_X1 U653 ( .A1(n498), .A2(n497), .A3(n496), .ZN(curr_proc_regs[235]) );
  NAND2_X1 U654 ( .A1(regs[748]), .A2(n15), .ZN(n501) );
  AOI22_X1 U655 ( .A1(n29), .A2(regs[1260]), .B1(n28), .B2(regs[236]), .ZN(
        n500) );
  AOI22_X1 U656 ( .A1(n1), .A2(regs[2284]), .B1(n3), .B2(regs[1772]), .ZN(n499) );
  NAND3_X1 U657 ( .A1(n501), .A2(n500), .A3(n499), .ZN(curr_proc_regs[236]) );
  NAND2_X1 U658 ( .A1(regs[749]), .A2(n15), .ZN(n504) );
  AOI22_X1 U659 ( .A1(n29), .A2(regs[1261]), .B1(n28), .B2(regs[237]), .ZN(
        n503) );
  AOI22_X1 U660 ( .A1(n1), .A2(regs[2285]), .B1(n3), .B2(regs[1773]), .ZN(n502) );
  NAND3_X1 U661 ( .A1(n504), .A2(n503), .A3(n502), .ZN(curr_proc_regs[237]) );
  NAND2_X1 U662 ( .A1(regs[750]), .A2(n15), .ZN(n507) );
  AOI22_X1 U663 ( .A1(n29), .A2(regs[1262]), .B1(n28), .B2(regs[238]), .ZN(
        n506) );
  AOI22_X1 U664 ( .A1(n1), .A2(regs[2286]), .B1(n34), .B2(regs[1774]), .ZN(
        n505) );
  NAND3_X1 U665 ( .A1(n507), .A2(n506), .A3(n505), .ZN(curr_proc_regs[238]) );
  NAND2_X1 U666 ( .A1(regs[751]), .A2(n11), .ZN(n510) );
  AOI22_X1 U667 ( .A1(n29), .A2(regs[1263]), .B1(n28), .B2(regs[239]), .ZN(
        n509) );
  AOI22_X1 U668 ( .A1(n1), .A2(regs[2287]), .B1(n9), .B2(regs[1775]), .ZN(n508) );
  NAND3_X1 U669 ( .A1(n510), .A2(n509), .A3(n508), .ZN(curr_proc_regs[239]) );
  NAND2_X1 U670 ( .A1(regs[535]), .A2(n13), .ZN(n513) );
  AOI22_X1 U671 ( .A1(n29), .A2(regs[1047]), .B1(n28), .B2(regs[23]), .ZN(n512) );
  AOI22_X1 U672 ( .A1(n1), .A2(regs[2071]), .B1(n9), .B2(regs[1559]), .ZN(n511) );
  NAND3_X1 U673 ( .A1(n513), .A2(n512), .A3(n511), .ZN(curr_proc_regs[23]) );
  NAND2_X1 U674 ( .A1(regs[752]), .A2(n11), .ZN(n516) );
  AOI22_X1 U675 ( .A1(n29), .A2(regs[1264]), .B1(n28), .B2(regs[240]), .ZN(
        n515) );
  AOI22_X1 U676 ( .A1(n1), .A2(regs[2288]), .B1(n35), .B2(regs[1776]), .ZN(
        n514) );
  NAND3_X1 U677 ( .A1(n516), .A2(n515), .A3(n514), .ZN(curr_proc_regs[240]) );
  NAND2_X1 U678 ( .A1(regs[753]), .A2(n13), .ZN(n519) );
  AOI22_X1 U679 ( .A1(n29), .A2(regs[1265]), .B1(n28), .B2(regs[241]), .ZN(
        n518) );
  AOI22_X1 U680 ( .A1(n4), .A2(regs[2289]), .B1(n31), .B2(regs[1777]), .ZN(
        n517) );
  NAND3_X1 U681 ( .A1(n519), .A2(n518), .A3(n517), .ZN(curr_proc_regs[241]) );
  NAND2_X1 U682 ( .A1(regs[754]), .A2(n11), .ZN(n522) );
  AOI22_X1 U683 ( .A1(n29), .A2(regs[1266]), .B1(n28), .B2(regs[242]), .ZN(
        n521) );
  AOI22_X1 U684 ( .A1(n4), .A2(regs[2290]), .B1(n3), .B2(regs[1778]), .ZN(n520) );
  NAND3_X1 U685 ( .A1(n522), .A2(n521), .A3(n520), .ZN(curr_proc_regs[242]) );
  NAND2_X1 U686 ( .A1(regs[755]), .A2(n13), .ZN(n525) );
  AOI22_X1 U687 ( .A1(n29), .A2(regs[1267]), .B1(n28), .B2(regs[243]), .ZN(
        n524) );
  AOI22_X1 U688 ( .A1(n4), .A2(regs[2291]), .B1(n2), .B2(regs[1779]), .ZN(n523) );
  NAND3_X1 U689 ( .A1(n525), .A2(n524), .A3(n523), .ZN(curr_proc_regs[243]) );
  NAND2_X1 U690 ( .A1(regs[756]), .A2(n11), .ZN(n528) );
  AOI22_X1 U691 ( .A1(n29), .A2(regs[1268]), .B1(n28), .B2(regs[244]), .ZN(
        n527) );
  AOI22_X1 U692 ( .A1(n4), .A2(regs[2292]), .B1(n2), .B2(regs[1780]), .ZN(n526) );
  NAND3_X1 U693 ( .A1(n528), .A2(n527), .A3(n526), .ZN(curr_proc_regs[244]) );
  NAND2_X1 U694 ( .A1(regs[757]), .A2(n13), .ZN(n531) );
  AOI22_X1 U695 ( .A1(n29), .A2(regs[1269]), .B1(n28), .B2(regs[245]), .ZN(
        n530) );
  AOI22_X1 U696 ( .A1(n4), .A2(regs[2293]), .B1(n2), .B2(regs[1781]), .ZN(n529) );
  NAND3_X1 U697 ( .A1(n531), .A2(n530), .A3(n529), .ZN(curr_proc_regs[245]) );
  NAND2_X1 U698 ( .A1(regs[758]), .A2(n11), .ZN(n534) );
  AOI22_X1 U699 ( .A1(n29), .A2(regs[1270]), .B1(n28), .B2(regs[246]), .ZN(
        n533) );
  AOI22_X1 U700 ( .A1(n4), .A2(regs[2294]), .B1(n2), .B2(regs[1782]), .ZN(n532) );
  NAND3_X1 U701 ( .A1(n534), .A2(n533), .A3(n532), .ZN(curr_proc_regs[246]) );
  NAND2_X1 U702 ( .A1(regs[759]), .A2(n13), .ZN(n537) );
  AOI22_X1 U703 ( .A1(n29), .A2(regs[1271]), .B1(n28), .B2(regs[247]), .ZN(
        n536) );
  AOI22_X1 U704 ( .A1(n4), .A2(regs[2295]), .B1(n2), .B2(regs[1783]), .ZN(n535) );
  NAND3_X1 U705 ( .A1(n537), .A2(n536), .A3(n535), .ZN(curr_proc_regs[247]) );
  NAND2_X1 U706 ( .A1(regs[760]), .A2(n11), .ZN(n540) );
  AOI22_X1 U707 ( .A1(n29), .A2(regs[1272]), .B1(n28), .B2(regs[248]), .ZN(
        n539) );
  AOI22_X1 U708 ( .A1(n4), .A2(regs[2296]), .B1(n2), .B2(regs[1784]), .ZN(n538) );
  NAND3_X1 U709 ( .A1(n540), .A2(n539), .A3(n538), .ZN(curr_proc_regs[248]) );
  NAND2_X1 U710 ( .A1(regs[761]), .A2(n16), .ZN(n543) );
  AOI22_X1 U711 ( .A1(n29), .A2(regs[1273]), .B1(n28), .B2(regs[249]), .ZN(
        n542) );
  AOI22_X1 U712 ( .A1(n4), .A2(regs[2297]), .B1(n30), .B2(regs[1785]), .ZN(
        n541) );
  NAND3_X1 U713 ( .A1(n543), .A2(n542), .A3(n541), .ZN(curr_proc_regs[249]) );
  NAND2_X1 U714 ( .A1(regs[536]), .A2(n16), .ZN(n546) );
  AOI22_X1 U715 ( .A1(n29), .A2(regs[1048]), .B1(n28), .B2(regs[24]), .ZN(n545) );
  AOI22_X1 U716 ( .A1(n4), .A2(regs[2072]), .B1(n34), .B2(regs[1560]), .ZN(
        n544) );
  NAND3_X1 U717 ( .A1(n546), .A2(n545), .A3(n544), .ZN(curr_proc_regs[24]) );
  NAND2_X1 U718 ( .A1(regs[762]), .A2(n16), .ZN(n549) );
  AOI22_X1 U719 ( .A1(n29), .A2(regs[1274]), .B1(n28), .B2(regs[250]), .ZN(
        n548) );
  AOI22_X1 U720 ( .A1(n1), .A2(regs[2298]), .B1(n2), .B2(regs[1786]), .ZN(n547) );
  NAND3_X1 U721 ( .A1(n549), .A2(n548), .A3(n547), .ZN(curr_proc_regs[250]) );
  NAND2_X1 U722 ( .A1(regs[763]), .A2(n16), .ZN(n552) );
  AOI22_X1 U723 ( .A1(n29), .A2(regs[1275]), .B1(n28), .B2(regs[251]), .ZN(
        n551) );
  AOI22_X1 U724 ( .A1(n4), .A2(regs[2299]), .B1(n34), .B2(regs[1787]), .ZN(
        n550) );
  NAND3_X1 U725 ( .A1(n552), .A2(n551), .A3(n550), .ZN(curr_proc_regs[251]) );
  NAND2_X1 U726 ( .A1(regs[764]), .A2(n16), .ZN(n555) );
  AOI22_X1 U727 ( .A1(n29), .A2(regs[1276]), .B1(n28), .B2(regs[252]), .ZN(
        n554) );
  AOI22_X1 U728 ( .A1(n1), .A2(regs[2300]), .B1(n30), .B2(regs[1788]), .ZN(
        n553) );
  NAND3_X1 U729 ( .A1(n555), .A2(n554), .A3(n553), .ZN(curr_proc_regs[252]) );
  NAND2_X1 U730 ( .A1(regs[765]), .A2(n16), .ZN(n558) );
  AOI22_X1 U731 ( .A1(n29), .A2(regs[1277]), .B1(n28), .B2(regs[253]), .ZN(
        n557) );
  AOI22_X1 U732 ( .A1(n1), .A2(regs[2301]), .B1(n34), .B2(regs[1789]), .ZN(
        n556) );
  NAND3_X1 U733 ( .A1(n558), .A2(n557), .A3(n556), .ZN(curr_proc_regs[253]) );
  NAND2_X1 U734 ( .A1(regs[766]), .A2(n16), .ZN(n561) );
  AOI22_X1 U735 ( .A1(n29), .A2(regs[1278]), .B1(n28), .B2(regs[254]), .ZN(
        n560) );
  AOI22_X1 U736 ( .A1(n1), .A2(regs[2302]), .B1(n30), .B2(regs[1790]), .ZN(
        n559) );
  NAND3_X1 U737 ( .A1(n561), .A2(n560), .A3(n559), .ZN(curr_proc_regs[254]) );
  NAND2_X1 U738 ( .A1(regs[767]), .A2(n16), .ZN(n564) );
  AOI22_X1 U739 ( .A1(n29), .A2(regs[1279]), .B1(n28), .B2(regs[255]), .ZN(
        n563) );
  AOI22_X1 U740 ( .A1(n1), .A2(regs[2303]), .B1(n34), .B2(regs[1791]), .ZN(
        n562) );
  NAND3_X1 U741 ( .A1(n564), .A2(n563), .A3(n562), .ZN(curr_proc_regs[255]) );
  NAND2_X1 U742 ( .A1(regs[768]), .A2(n16), .ZN(n567) );
  AOI22_X1 U743 ( .A1(n29), .A2(regs[1280]), .B1(n28), .B2(regs[256]), .ZN(
        n566) );
  AOI22_X1 U744 ( .A1(n1), .A2(regs[2304]), .B1(n30), .B2(regs[1792]), .ZN(
        n565) );
  NAND3_X1 U745 ( .A1(n567), .A2(n566), .A3(n565), .ZN(curr_proc_regs[256]) );
  NAND2_X1 U746 ( .A1(regs[769]), .A2(n16), .ZN(n570) );
  AOI22_X1 U747 ( .A1(n29), .A2(regs[1281]), .B1(n28), .B2(regs[257]), .ZN(
        n569) );
  AOI22_X1 U748 ( .A1(n1), .A2(regs[2305]), .B1(n34), .B2(regs[1793]), .ZN(
        n568) );
  NAND3_X1 U749 ( .A1(n570), .A2(n569), .A3(n568), .ZN(curr_proc_regs[257]) );
  NAND2_X1 U750 ( .A1(regs[770]), .A2(n16), .ZN(n573) );
  AOI22_X1 U751 ( .A1(n29), .A2(regs[1282]), .B1(n28), .B2(regs[258]), .ZN(
        n572) );
  AOI22_X1 U752 ( .A1(n1), .A2(regs[2306]), .B1(n34), .B2(regs[1794]), .ZN(
        n571) );
  NAND3_X1 U753 ( .A1(n573), .A2(n572), .A3(n571), .ZN(curr_proc_regs[258]) );
  NAND2_X1 U754 ( .A1(regs[771]), .A2(n11), .ZN(n576) );
  AOI22_X1 U755 ( .A1(n29), .A2(regs[1283]), .B1(n28), .B2(regs[259]), .ZN(
        n575) );
  AOI22_X1 U756 ( .A1(n1), .A2(regs[2307]), .B1(n32), .B2(regs[1795]), .ZN(
        n574) );
  NAND3_X1 U757 ( .A1(n576), .A2(n575), .A3(n574), .ZN(curr_proc_regs[259]) );
  NAND2_X1 U758 ( .A1(regs[537]), .A2(n11), .ZN(n579) );
  AOI22_X1 U759 ( .A1(n29), .A2(regs[1049]), .B1(n28), .B2(regs[25]), .ZN(n578) );
  AOI22_X1 U760 ( .A1(n1), .A2(regs[2073]), .B1(n32), .B2(regs[1561]), .ZN(
        n577) );
  NAND3_X1 U761 ( .A1(n579), .A2(n578), .A3(n577), .ZN(curr_proc_regs[25]) );
  NAND2_X1 U762 ( .A1(regs[772]), .A2(n11), .ZN(n582) );
  AOI22_X1 U763 ( .A1(n29), .A2(regs[1284]), .B1(n28), .B2(regs[260]), .ZN(
        n581) );
  AOI22_X1 U764 ( .A1(n1), .A2(regs[2308]), .B1(n32), .B2(regs[1796]), .ZN(
        n580) );
  NAND3_X1 U765 ( .A1(n582), .A2(n581), .A3(n580), .ZN(curr_proc_regs[260]) );
  NAND2_X1 U766 ( .A1(regs[773]), .A2(n11), .ZN(n585) );
  AOI22_X1 U767 ( .A1(n29), .A2(regs[1285]), .B1(n28), .B2(regs[261]), .ZN(
        n584) );
  AOI22_X1 U768 ( .A1(n39), .A2(regs[2309]), .B1(n32), .B2(regs[1797]), .ZN(
        n583) );
  NAND3_X1 U769 ( .A1(n585), .A2(n584), .A3(n583), .ZN(curr_proc_regs[261]) );
  NAND2_X1 U770 ( .A1(regs[774]), .A2(n11), .ZN(n588) );
  AOI22_X1 U771 ( .A1(n29), .A2(regs[1286]), .B1(n28), .B2(regs[262]), .ZN(
        n587) );
  AOI22_X1 U772 ( .A1(n40), .A2(regs[2310]), .B1(n32), .B2(regs[1798]), .ZN(
        n586) );
  NAND3_X1 U773 ( .A1(n588), .A2(n587), .A3(n586), .ZN(curr_proc_regs[262]) );
  NAND2_X1 U774 ( .A1(regs[775]), .A2(n11), .ZN(n591) );
  AOI22_X1 U775 ( .A1(n29), .A2(regs[1287]), .B1(n28), .B2(regs[263]), .ZN(
        n590) );
  AOI22_X1 U776 ( .A1(n36), .A2(regs[2311]), .B1(n32), .B2(regs[1799]), .ZN(
        n589) );
  NAND3_X1 U777 ( .A1(n591), .A2(n590), .A3(n589), .ZN(curr_proc_regs[263]) );
  NAND2_X1 U778 ( .A1(regs[776]), .A2(n11), .ZN(n594) );
  AOI22_X1 U779 ( .A1(n29), .A2(regs[1288]), .B1(n28), .B2(regs[264]), .ZN(
        n593) );
  AOI22_X1 U780 ( .A1(win[4]), .A2(regs[2312]), .B1(n32), .B2(regs[1800]), 
        .ZN(n592) );
  NAND3_X1 U781 ( .A1(n594), .A2(n593), .A3(n592), .ZN(curr_proc_regs[264]) );
  NAND2_X1 U782 ( .A1(regs[777]), .A2(n11), .ZN(n597) );
  AOI22_X1 U783 ( .A1(n29), .A2(regs[1289]), .B1(n28), .B2(regs[265]), .ZN(
        n596) );
  AOI22_X1 U784 ( .A1(n8), .A2(regs[2313]), .B1(n32), .B2(regs[1801]), .ZN(
        n595) );
  NAND3_X1 U785 ( .A1(n597), .A2(n596), .A3(n595), .ZN(curr_proc_regs[265]) );
  NAND2_X1 U786 ( .A1(regs[778]), .A2(n11), .ZN(n600) );
  AOI22_X1 U787 ( .A1(n29), .A2(regs[1290]), .B1(n28), .B2(regs[266]), .ZN(
        n599) );
  AOI22_X1 U788 ( .A1(win[4]), .A2(regs[2314]), .B1(n32), .B2(regs[1802]), 
        .ZN(n598) );
  NAND3_X1 U789 ( .A1(n600), .A2(n599), .A3(n598), .ZN(curr_proc_regs[266]) );
  NAND2_X1 U790 ( .A1(regs[779]), .A2(n11), .ZN(n603) );
  AOI22_X1 U791 ( .A1(n29), .A2(regs[1291]), .B1(n28), .B2(regs[267]), .ZN(
        n602) );
  AOI22_X1 U792 ( .A1(n38), .A2(regs[2315]), .B1(n32), .B2(regs[1803]), .ZN(
        n601) );
  NAND3_X1 U793 ( .A1(n603), .A2(n602), .A3(n601), .ZN(curr_proc_regs[267]) );
  NAND2_X1 U794 ( .A1(regs[780]), .A2(n11), .ZN(n606) );
  AOI22_X1 U795 ( .A1(n29), .A2(regs[1292]), .B1(n28), .B2(regs[268]), .ZN(
        n605) );
  AOI22_X1 U796 ( .A1(win[4]), .A2(regs[2316]), .B1(n32), .B2(regs[1804]), 
        .ZN(n604) );
  NAND3_X1 U797 ( .A1(n606), .A2(n605), .A3(n604), .ZN(curr_proc_regs[268]) );
  NAND2_X1 U798 ( .A1(regs[781]), .A2(n13), .ZN(n609) );
  AOI22_X1 U799 ( .A1(n29), .A2(regs[1293]), .B1(n21), .B2(regs[269]), .ZN(
        n608) );
  AOI22_X1 U800 ( .A1(n41), .A2(regs[2317]), .B1(n31), .B2(regs[1805]), .ZN(
        n607) );
  NAND3_X1 U801 ( .A1(n609), .A2(n608), .A3(n607), .ZN(curr_proc_regs[269]) );
  NAND2_X1 U802 ( .A1(regs[538]), .A2(n13), .ZN(n612) );
  AOI22_X1 U803 ( .A1(n29), .A2(regs[1050]), .B1(n1580), .B2(regs[26]), .ZN(
        n611) );
  AOI22_X1 U804 ( .A1(win[4]), .A2(regs[2074]), .B1(n31), .B2(regs[1562]), 
        .ZN(n610) );
  NAND3_X1 U805 ( .A1(n612), .A2(n611), .A3(n610), .ZN(curr_proc_regs[26]) );
  NAND2_X1 U806 ( .A1(regs[782]), .A2(n13), .ZN(n615) );
  AOI22_X1 U807 ( .A1(n29), .A2(regs[1294]), .B1(n1580), .B2(regs[270]), .ZN(
        n614) );
  AOI22_X1 U808 ( .A1(n10), .A2(regs[2318]), .B1(n31), .B2(regs[1806]), .ZN(
        n613) );
  NAND3_X1 U809 ( .A1(n615), .A2(n614), .A3(n613), .ZN(curr_proc_regs[270]) );
  NAND2_X1 U810 ( .A1(regs[783]), .A2(n13), .ZN(n618) );
  AOI22_X1 U811 ( .A1(n29), .A2(regs[1295]), .B1(n1580), .B2(regs[271]), .ZN(
        n617) );
  AOI22_X1 U812 ( .A1(win[4]), .A2(regs[2319]), .B1(n31), .B2(regs[1807]), 
        .ZN(n616) );
  NAND3_X1 U813 ( .A1(n618), .A2(n617), .A3(n616), .ZN(curr_proc_regs[271]) );
  NAND2_X1 U814 ( .A1(regs[784]), .A2(n13), .ZN(n621) );
  AOI22_X1 U815 ( .A1(n29), .A2(regs[1296]), .B1(n1580), .B2(regs[272]), .ZN(
        n620) );
  AOI22_X1 U816 ( .A1(n41), .A2(regs[2320]), .B1(n31), .B2(regs[1808]), .ZN(
        n619) );
  NAND3_X1 U817 ( .A1(n621), .A2(n620), .A3(n619), .ZN(curr_proc_regs[272]) );
  NAND2_X1 U818 ( .A1(regs[785]), .A2(n13), .ZN(n624) );
  AOI22_X1 U819 ( .A1(n29), .A2(regs[1297]), .B1(n1580), .B2(regs[273]), .ZN(
        n623) );
  AOI22_X1 U820 ( .A1(n8), .A2(regs[2321]), .B1(n31), .B2(regs[1809]), .ZN(
        n622) );
  NAND3_X1 U821 ( .A1(n624), .A2(n623), .A3(n622), .ZN(curr_proc_regs[273]) );
  NAND2_X1 U822 ( .A1(regs[786]), .A2(n13), .ZN(n627) );
  AOI22_X1 U823 ( .A1(n29), .A2(regs[1298]), .B1(n23), .B2(regs[274]), .ZN(
        n626) );
  AOI22_X1 U824 ( .A1(n39), .A2(regs[2322]), .B1(n31), .B2(regs[1810]), .ZN(
        n625) );
  NAND3_X1 U825 ( .A1(n627), .A2(n626), .A3(n625), .ZN(curr_proc_regs[274]) );
  NAND2_X1 U826 ( .A1(regs[787]), .A2(n13), .ZN(n630) );
  AOI22_X1 U827 ( .A1(n29), .A2(regs[1299]), .B1(n5), .B2(regs[275]), .ZN(n629) );
  AOI22_X1 U828 ( .A1(n37), .A2(regs[2323]), .B1(n31), .B2(regs[1811]), .ZN(
        n628) );
  NAND3_X1 U829 ( .A1(n630), .A2(n629), .A3(n628), .ZN(curr_proc_regs[275]) );
  NAND2_X1 U830 ( .A1(regs[788]), .A2(n13), .ZN(n633) );
  AOI22_X1 U831 ( .A1(n29), .A2(regs[1300]), .B1(n23), .B2(regs[276]), .ZN(
        n632) );
  AOI22_X1 U832 ( .A1(n4), .A2(regs[2324]), .B1(n31), .B2(regs[1812]), .ZN(
        n631) );
  NAND3_X1 U833 ( .A1(n633), .A2(n632), .A3(n631), .ZN(curr_proc_regs[276]) );
  NAND2_X1 U834 ( .A1(regs[789]), .A2(n13), .ZN(n636) );
  AOI22_X1 U835 ( .A1(n29), .A2(regs[1301]), .B1(n5), .B2(regs[277]), .ZN(n635) );
  AOI22_X1 U836 ( .A1(n10), .A2(regs[2325]), .B1(n31), .B2(regs[1813]), .ZN(
        n634) );
  NAND3_X1 U837 ( .A1(n636), .A2(n635), .A3(n634), .ZN(curr_proc_regs[277]) );
  NAND2_X1 U838 ( .A1(regs[790]), .A2(n13), .ZN(n639) );
  AOI22_X1 U839 ( .A1(n29), .A2(regs[1302]), .B1(n5), .B2(regs[278]), .ZN(n638) );
  AOI22_X1 U840 ( .A1(n1), .A2(regs[2326]), .B1(n31), .B2(regs[1814]), .ZN(
        n637) );
  NAND3_X1 U841 ( .A1(n639), .A2(n638), .A3(n637), .ZN(curr_proc_regs[278]) );
  NAND2_X1 U842 ( .A1(regs[791]), .A2(n13), .ZN(n642) );
  AOI22_X1 U843 ( .A1(n29), .A2(regs[1303]), .B1(n23), .B2(regs[279]), .ZN(
        n641) );
  AOI22_X1 U844 ( .A1(n41), .A2(regs[2327]), .B1(n3), .B2(regs[1815]), .ZN(
        n640) );
  NAND3_X1 U845 ( .A1(n642), .A2(n641), .A3(n640), .ZN(curr_proc_regs[279]) );
  NAND2_X1 U846 ( .A1(regs[539]), .A2(n13), .ZN(n645) );
  AOI22_X1 U847 ( .A1(n29), .A2(regs[1051]), .B1(n5), .B2(regs[27]), .ZN(n644)
         );
  AOI22_X1 U848 ( .A1(n8), .A2(regs[2075]), .B1(n2), .B2(regs[1563]), .ZN(n643) );
  NAND3_X1 U849 ( .A1(n645), .A2(n644), .A3(n643), .ZN(curr_proc_regs[27]) );
  NAND2_X1 U850 ( .A1(regs[792]), .A2(n13), .ZN(n648) );
  AOI22_X1 U851 ( .A1(n29), .A2(regs[1304]), .B1(n28), .B2(regs[280]), .ZN(
        n647) );
  AOI22_X1 U852 ( .A1(n36), .A2(regs[2328]), .B1(n34), .B2(regs[1816]), .ZN(
        n646) );
  NAND3_X1 U853 ( .A1(n648), .A2(n647), .A3(n646), .ZN(curr_proc_regs[280]) );
  NAND2_X1 U854 ( .A1(regs[793]), .A2(n13), .ZN(n651) );
  AOI22_X1 U855 ( .A1(n29), .A2(regs[1305]), .B1(n23), .B2(regs[281]), .ZN(
        n650) );
  AOI22_X1 U856 ( .A1(n40), .A2(regs[2329]), .B1(n2), .B2(regs[1817]), .ZN(
        n649) );
  NAND3_X1 U857 ( .A1(n651), .A2(n650), .A3(n649), .ZN(curr_proc_regs[281]) );
  NAND2_X1 U858 ( .A1(regs[794]), .A2(n13), .ZN(n654) );
  AOI22_X1 U859 ( .A1(n29), .A2(regs[1306]), .B1(n5), .B2(regs[282]), .ZN(n653) );
  AOI22_X1 U860 ( .A1(n36), .A2(regs[2330]), .B1(n31), .B2(regs[1818]), .ZN(
        n652) );
  NAND3_X1 U861 ( .A1(n654), .A2(n653), .A3(n652), .ZN(curr_proc_regs[282]) );
  NAND2_X1 U862 ( .A1(regs[795]), .A2(n13), .ZN(n657) );
  AOI22_X1 U863 ( .A1(n29), .A2(regs[1307]), .B1(n1580), .B2(regs[283]), .ZN(
        n656) );
  AOI22_X1 U864 ( .A1(n40), .A2(regs[2331]), .B1(n2), .B2(regs[1819]), .ZN(
        n655) );
  NAND3_X1 U865 ( .A1(n657), .A2(n656), .A3(n655), .ZN(curr_proc_regs[283]) );
  NAND2_X1 U866 ( .A1(regs[796]), .A2(n13), .ZN(n660) );
  AOI22_X1 U867 ( .A1(n29), .A2(regs[1308]), .B1(n23), .B2(regs[284]), .ZN(
        n659) );
  AOI22_X1 U868 ( .A1(n36), .A2(regs[2332]), .B1(n2), .B2(regs[1820]), .ZN(
        n658) );
  NAND3_X1 U869 ( .A1(n660), .A2(n659), .A3(n658), .ZN(curr_proc_regs[284]) );
  NAND2_X1 U870 ( .A1(regs[797]), .A2(n13), .ZN(n663) );
  AOI22_X1 U871 ( .A1(n29), .A2(regs[1309]), .B1(n5), .B2(regs[285]), .ZN(n662) );
  AOI22_X1 U872 ( .A1(n40), .A2(regs[2333]), .B1(n2), .B2(regs[1821]), .ZN(
        n661) );
  NAND3_X1 U873 ( .A1(n663), .A2(n662), .A3(n661), .ZN(curr_proc_regs[285]) );
  NAND2_X1 U874 ( .A1(regs[798]), .A2(n13), .ZN(n666) );
  AOI22_X1 U875 ( .A1(n29), .A2(regs[1310]), .B1(n26), .B2(regs[286]), .ZN(
        n665) );
  AOI22_X1 U876 ( .A1(n36), .A2(regs[2334]), .B1(n2), .B2(regs[1822]), .ZN(
        n664) );
  NAND3_X1 U877 ( .A1(n666), .A2(n665), .A3(n664), .ZN(curr_proc_regs[286]) );
  NAND2_X1 U878 ( .A1(regs[799]), .A2(n13), .ZN(n669) );
  AOI22_X1 U879 ( .A1(n29), .A2(regs[1311]), .B1(n23), .B2(regs[287]), .ZN(
        n668) );
  AOI22_X1 U880 ( .A1(n40), .A2(regs[2335]), .B1(n2), .B2(regs[1823]), .ZN(
        n667) );
  NAND3_X1 U881 ( .A1(n669), .A2(n668), .A3(n667), .ZN(curr_proc_regs[287]) );
  NAND2_X1 U882 ( .A1(regs[800]), .A2(n13), .ZN(n672) );
  AOI22_X1 U883 ( .A1(n29), .A2(regs[1312]), .B1(n5), .B2(regs[288]), .ZN(n671) );
  AOI22_X1 U884 ( .A1(n36), .A2(regs[2336]), .B1(n2), .B2(regs[1824]), .ZN(
        n670) );
  NAND3_X1 U885 ( .A1(n672), .A2(n671), .A3(n670), .ZN(curr_proc_regs[288]) );
  NAND2_X1 U886 ( .A1(regs[801]), .A2(n13), .ZN(n675) );
  AOI22_X1 U887 ( .A1(n29), .A2(regs[1313]), .B1(n23), .B2(regs[289]), .ZN(
        n674) );
  AOI22_X1 U888 ( .A1(n40), .A2(regs[2337]), .B1(n34), .B2(regs[1825]), .ZN(
        n673) );
  NAND3_X1 U889 ( .A1(n675), .A2(n674), .A3(n673), .ZN(curr_proc_regs[289]) );
  NAND2_X1 U890 ( .A1(regs[540]), .A2(n16), .ZN(n678) );
  AOI22_X1 U891 ( .A1(n29), .A2(regs[1052]), .B1(n23), .B2(regs[28]), .ZN(n677) );
  AOI22_X1 U892 ( .A1(n36), .A2(regs[2076]), .B1(n34), .B2(regs[1564]), .ZN(
        n676) );
  NAND3_X1 U893 ( .A1(n678), .A2(n677), .A3(n676), .ZN(curr_proc_regs[28]) );
  NAND2_X1 U894 ( .A1(regs[802]), .A2(n11), .ZN(n681) );
  AOI22_X1 U895 ( .A1(n29), .A2(regs[1314]), .B1(n23), .B2(regs[290]), .ZN(
        n680) );
  AOI22_X1 U896 ( .A1(n1), .A2(regs[2338]), .B1(n34), .B2(regs[1826]), .ZN(
        n679) );
  NAND3_X1 U897 ( .A1(n681), .A2(n680), .A3(n679), .ZN(curr_proc_regs[290]) );
  NAND2_X1 U898 ( .A1(regs[803]), .A2(n16), .ZN(n684) );
  AOI22_X1 U899 ( .A1(n29), .A2(regs[1315]), .B1(n23), .B2(regs[291]), .ZN(
        n683) );
  AOI22_X1 U900 ( .A1(n10), .A2(regs[2339]), .B1(n34), .B2(regs[1827]), .ZN(
        n682) );
  NAND3_X1 U901 ( .A1(n684), .A2(n683), .A3(n682), .ZN(curr_proc_regs[291]) );
  NAND2_X1 U902 ( .A1(regs[804]), .A2(n13), .ZN(n687) );
  AOI22_X1 U903 ( .A1(n29), .A2(regs[1316]), .B1(n23), .B2(regs[292]), .ZN(
        n686) );
  AOI22_X1 U904 ( .A1(n1), .A2(regs[2340]), .B1(n34), .B2(regs[1828]), .ZN(
        n685) );
  NAND3_X1 U905 ( .A1(n687), .A2(n686), .A3(n685), .ZN(curr_proc_regs[292]) );
  NAND2_X1 U906 ( .A1(regs[805]), .A2(n16), .ZN(n690) );
  AOI22_X1 U907 ( .A1(n29), .A2(regs[1317]), .B1(n23), .B2(regs[293]), .ZN(
        n689) );
  AOI22_X1 U908 ( .A1(n10), .A2(regs[2341]), .B1(n34), .B2(regs[1829]), .ZN(
        n688) );
  NAND3_X1 U909 ( .A1(n690), .A2(n689), .A3(n688), .ZN(curr_proc_regs[293]) );
  NAND2_X1 U910 ( .A1(regs[806]), .A2(n14), .ZN(n693) );
  AOI22_X1 U911 ( .A1(n29), .A2(regs[1318]), .B1(n23), .B2(regs[294]), .ZN(
        n692) );
  AOI22_X1 U912 ( .A1(n1), .A2(regs[2342]), .B1(n34), .B2(regs[1830]), .ZN(
        n691) );
  NAND3_X1 U913 ( .A1(n693), .A2(n692), .A3(n691), .ZN(curr_proc_regs[294]) );
  NAND2_X1 U914 ( .A1(regs[807]), .A2(n16), .ZN(n696) );
  AOI22_X1 U915 ( .A1(n29), .A2(regs[1319]), .B1(n23), .B2(regs[295]), .ZN(
        n695) );
  AOI22_X1 U916 ( .A1(n10), .A2(regs[2343]), .B1(n34), .B2(regs[1831]), .ZN(
        n694) );
  NAND3_X1 U917 ( .A1(n696), .A2(n695), .A3(n694), .ZN(curr_proc_regs[295]) );
  NAND2_X1 U918 ( .A1(regs[808]), .A2(n13), .ZN(n699) );
  AOI22_X1 U919 ( .A1(n29), .A2(regs[1320]), .B1(n23), .B2(regs[296]), .ZN(
        n698) );
  AOI22_X1 U920 ( .A1(n1), .A2(regs[2344]), .B1(n34), .B2(regs[1832]), .ZN(
        n697) );
  NAND3_X1 U921 ( .A1(n699), .A2(n698), .A3(n697), .ZN(curr_proc_regs[296]) );
  NAND2_X1 U922 ( .A1(regs[809]), .A2(n16), .ZN(n702) );
  AOI22_X1 U923 ( .A1(n29), .A2(regs[1321]), .B1(n23), .B2(regs[297]), .ZN(
        n701) );
  AOI22_X1 U924 ( .A1(n10), .A2(regs[2345]), .B1(n34), .B2(regs[1833]), .ZN(
        n700) );
  NAND3_X1 U925 ( .A1(n702), .A2(n701), .A3(n700), .ZN(curr_proc_regs[297]) );
  NAND2_X1 U926 ( .A1(regs[810]), .A2(n16), .ZN(n705) );
  AOI22_X1 U927 ( .A1(n29), .A2(regs[1322]), .B1(n23), .B2(regs[298]), .ZN(
        n704) );
  AOI22_X1 U928 ( .A1(n1), .A2(regs[2346]), .B1(n34), .B2(regs[1834]), .ZN(
        n703) );
  NAND3_X1 U929 ( .A1(n705), .A2(n704), .A3(n703), .ZN(curr_proc_regs[298]) );
  NAND2_X1 U930 ( .A1(regs[811]), .A2(n11), .ZN(n708) );
  AOI22_X1 U931 ( .A1(n29), .A2(regs[1323]), .B1(n5), .B2(regs[299]), .ZN(n707) );
  AOI22_X1 U932 ( .A1(n10), .A2(regs[2347]), .B1(n3), .B2(regs[1835]), .ZN(
        n706) );
  NAND3_X1 U933 ( .A1(n708), .A2(n707), .A3(n706), .ZN(curr_proc_regs[299]) );
  NAND2_X1 U934 ( .A1(regs[541]), .A2(n11), .ZN(n711) );
  AOI22_X1 U935 ( .A1(n29), .A2(regs[1053]), .B1(n12), .B2(regs[29]), .ZN(n710) );
  AOI22_X1 U936 ( .A1(n1), .A2(regs[2077]), .B1(n33), .B2(regs[1565]), .ZN(
        n709) );
  NAND3_X1 U937 ( .A1(n711), .A2(n710), .A3(n709), .ZN(curr_proc_regs[29]) );
  NAND2_X1 U938 ( .A1(regs[514]), .A2(n11), .ZN(n714) );
  AOI22_X1 U939 ( .A1(n29), .A2(regs[1026]), .B1(n1580), .B2(regs[2]), .ZN(
        n713) );
  AOI22_X1 U940 ( .A1(n4), .A2(regs[2050]), .B1(n34), .B2(regs[1538]), .ZN(
        n712) );
  NAND3_X1 U941 ( .A1(n714), .A2(n713), .A3(n712), .ZN(curr_proc_regs[2]) );
  NAND2_X1 U942 ( .A1(regs[812]), .A2(n11), .ZN(n717) );
  AOI22_X1 U943 ( .A1(n29), .A2(regs[1324]), .B1(n23), .B2(regs[300]), .ZN(
        n716) );
  AOI22_X1 U944 ( .A1(win[4]), .A2(regs[2348]), .B1(n9), .B2(regs[1836]), .ZN(
        n715) );
  NAND3_X1 U945 ( .A1(n717), .A2(n716), .A3(n715), .ZN(curr_proc_regs[300]) );
  NAND2_X1 U946 ( .A1(regs[813]), .A2(n11), .ZN(n720) );
  AOI22_X1 U947 ( .A1(n29), .A2(regs[1325]), .B1(n5), .B2(regs[301]), .ZN(n719) );
  AOI22_X1 U948 ( .A1(n4), .A2(regs[2349]), .B1(n9), .B2(regs[1837]), .ZN(n718) );
  NAND3_X1 U949 ( .A1(n720), .A2(n719), .A3(n718), .ZN(curr_proc_regs[301]) );
  NAND2_X1 U950 ( .A1(regs[814]), .A2(n11), .ZN(n723) );
  AOI22_X1 U951 ( .A1(n29), .A2(regs[1326]), .B1(n23), .B2(regs[302]), .ZN(
        n722) );
  AOI22_X1 U952 ( .A1(n10), .A2(regs[2350]), .B1(n35), .B2(regs[1838]), .ZN(
        n721) );
  NAND3_X1 U953 ( .A1(n723), .A2(n722), .A3(n721), .ZN(curr_proc_regs[302]) );
  NAND2_X1 U954 ( .A1(regs[815]), .A2(n11), .ZN(n726) );
  AOI22_X1 U955 ( .A1(n29), .A2(regs[1327]), .B1(n22), .B2(regs[303]), .ZN(
        n725) );
  AOI22_X1 U956 ( .A1(n4), .A2(regs[2351]), .B1(n3), .B2(regs[1839]), .ZN(n724) );
  NAND3_X1 U957 ( .A1(n726), .A2(n725), .A3(n724), .ZN(curr_proc_regs[303]) );
  NAND2_X1 U958 ( .A1(regs[816]), .A2(n11), .ZN(n729) );
  AOI22_X1 U959 ( .A1(n29), .A2(regs[1328]), .B1(n23), .B2(regs[304]), .ZN(
        n728) );
  AOI22_X1 U960 ( .A1(win[4]), .A2(regs[2352]), .B1(n3), .B2(regs[1840]), .ZN(
        n727) );
  NAND3_X1 U961 ( .A1(n729), .A2(n728), .A3(n727), .ZN(curr_proc_regs[304]) );
  NAND2_X1 U962 ( .A1(regs[817]), .A2(n11), .ZN(n732) );
  AOI22_X1 U963 ( .A1(n29), .A2(regs[1329]), .B1(n5), .B2(regs[305]), .ZN(n731) );
  AOI22_X1 U964 ( .A1(n4), .A2(regs[2353]), .B1(n34), .B2(regs[1841]), .ZN(
        n730) );
  NAND3_X1 U965 ( .A1(n732), .A2(n731), .A3(n730), .ZN(curr_proc_regs[305]) );
  NAND2_X1 U966 ( .A1(regs[818]), .A2(n11), .ZN(n735) );
  AOI22_X1 U967 ( .A1(n29), .A2(regs[1330]), .B1(n5), .B2(regs[306]), .ZN(n734) );
  AOI22_X1 U968 ( .A1(n39), .A2(regs[2354]), .B1(n31), .B2(regs[1842]), .ZN(
        n733) );
  NAND3_X1 U969 ( .A1(n735), .A2(n734), .A3(n733), .ZN(curr_proc_regs[306]) );
  NAND2_X1 U970 ( .A1(regs[819]), .A2(n11), .ZN(n738) );
  AOI22_X1 U971 ( .A1(n29), .A2(regs[1331]), .B1(n1580), .B2(regs[307]), .ZN(
        n737) );
  AOI22_X1 U972 ( .A1(n4), .A2(regs[2355]), .B1(n33), .B2(regs[1843]), .ZN(
        n736) );
  NAND3_X1 U973 ( .A1(n738), .A2(n737), .A3(n736), .ZN(curr_proc_regs[307]) );
  NAND2_X1 U974 ( .A1(regs[820]), .A2(n14), .ZN(n741) );
  AOI22_X1 U975 ( .A1(n29), .A2(regs[1332]), .B1(n23), .B2(regs[308]), .ZN(
        n740) );
  AOI22_X1 U976 ( .A1(win[4]), .A2(regs[2356]), .B1(n9), .B2(regs[1844]), .ZN(
        n739) );
  NAND3_X1 U977 ( .A1(n741), .A2(n740), .A3(n739), .ZN(curr_proc_regs[308]) );
  NAND2_X1 U978 ( .A1(regs[821]), .A2(n1579), .ZN(n744) );
  AOI22_X1 U979 ( .A1(n29), .A2(regs[1333]), .B1(n1580), .B2(regs[309]), .ZN(
        n743) );
  AOI22_X1 U980 ( .A1(n4), .A2(regs[2357]), .B1(n9), .B2(regs[1845]), .ZN(n742) );
  NAND3_X1 U981 ( .A1(n744), .A2(n743), .A3(n742), .ZN(curr_proc_regs[309]) );
  NAND2_X1 U982 ( .A1(regs[542]), .A2(n16), .ZN(n747) );
  AOI22_X1 U983 ( .A1(n29), .A2(regs[1054]), .B1(n24), .B2(regs[30]), .ZN(n746) );
  AOI22_X1 U984 ( .A1(n41), .A2(regs[2078]), .B1(n35), .B2(regs[1566]), .ZN(
        n745) );
  NAND3_X1 U985 ( .A1(n747), .A2(n746), .A3(n745), .ZN(curr_proc_regs[30]) );
  NAND2_X1 U986 ( .A1(regs[822]), .A2(n15), .ZN(n750) );
  AOI22_X1 U987 ( .A1(n29), .A2(regs[1334]), .B1(n23), .B2(regs[310]), .ZN(
        n749) );
  AOI22_X1 U988 ( .A1(win[4]), .A2(regs[2358]), .B1(n3), .B2(regs[1846]), .ZN(
        n748) );
  NAND3_X1 U989 ( .A1(n750), .A2(n749), .A3(n748), .ZN(curr_proc_regs[310]) );
  NAND2_X1 U990 ( .A1(regs[823]), .A2(n14), .ZN(n753) );
  AOI22_X1 U991 ( .A1(n29), .A2(regs[1335]), .B1(n5), .B2(regs[311]), .ZN(n752) );
  AOI22_X1 U992 ( .A1(win[4]), .A2(regs[2359]), .B1(n3), .B2(regs[1847]), .ZN(
        n751) );
  NAND3_X1 U993 ( .A1(n753), .A2(n752), .A3(n751), .ZN(curr_proc_regs[311]) );
  NAND2_X1 U994 ( .A1(regs[824]), .A2(n1579), .ZN(n756) );
  AOI22_X1 U995 ( .A1(n29), .A2(regs[1336]), .B1(n5), .B2(regs[312]), .ZN(n755) );
  AOI22_X1 U996 ( .A1(n37), .A2(regs[2360]), .B1(n34), .B2(regs[1848]), .ZN(
        n754) );
  NAND3_X1 U997 ( .A1(n756), .A2(n755), .A3(n754), .ZN(curr_proc_regs[312]) );
  NAND2_X1 U998 ( .A1(regs[825]), .A2(n16), .ZN(n759) );
  AOI22_X1 U999 ( .A1(n29), .A2(regs[1337]), .B1(n23), .B2(regs[313]), .ZN(
        n758) );
  AOI22_X1 U1000 ( .A1(win[4]), .A2(regs[2361]), .B1(n31), .B2(regs[1849]), 
        .ZN(n757) );
  NAND3_X1 U1001 ( .A1(n759), .A2(n758), .A3(n757), .ZN(curr_proc_regs[313])
         );
  NAND2_X1 U1002 ( .A1(regs[826]), .A2(n15), .ZN(n762) );
  AOI22_X1 U1003 ( .A1(n29), .A2(regs[1338]), .B1(n5), .B2(regs[314]), .ZN(
        n761) );
  AOI22_X1 U1004 ( .A1(win[4]), .A2(regs[2362]), .B1(n33), .B2(regs[1850]), 
        .ZN(n760) );
  NAND3_X1 U1005 ( .A1(n762), .A2(n761), .A3(n760), .ZN(curr_proc_regs[314])
         );
  NAND2_X1 U1006 ( .A1(regs[827]), .A2(n7), .ZN(n765) );
  AOI22_X1 U1007 ( .A1(n29), .A2(regs[1339]), .B1(n5), .B2(regs[315]), .ZN(
        n764) );
  AOI22_X1 U1008 ( .A1(n38), .A2(regs[2363]), .B1(n9), .B2(regs[1851]), .ZN(
        n763) );
  NAND3_X1 U1009 ( .A1(n765), .A2(n764), .A3(n763), .ZN(curr_proc_regs[315])
         );
  NAND2_X1 U1010 ( .A1(regs[828]), .A2(n18), .ZN(n768) );
  AOI22_X1 U1011 ( .A1(n29), .A2(regs[1340]), .B1(n5), .B2(regs[316]), .ZN(
        n767) );
  AOI22_X1 U1012 ( .A1(win[4]), .A2(regs[2364]), .B1(n9), .B2(regs[1852]), 
        .ZN(n766) );
  NAND3_X1 U1013 ( .A1(n768), .A2(n767), .A3(n766), .ZN(curr_proc_regs[316])
         );
  NAND2_X1 U1014 ( .A1(regs[829]), .A2(n19), .ZN(n771) );
  AOI22_X1 U1015 ( .A1(n29), .A2(regs[1341]), .B1(n5), .B2(regs[317]), .ZN(
        n770) );
  AOI22_X1 U1016 ( .A1(win[4]), .A2(regs[2365]), .B1(n35), .B2(regs[1853]), 
        .ZN(n769) );
  NAND3_X1 U1017 ( .A1(n771), .A2(n770), .A3(n769), .ZN(curr_proc_regs[317])
         );
  NAND2_X1 U1018 ( .A1(regs[830]), .A2(n7), .ZN(n774) );
  AOI22_X1 U1019 ( .A1(n29), .A2(regs[1342]), .B1(n23), .B2(regs[318]), .ZN(
        n773) );
  AOI22_X1 U1020 ( .A1(n38), .A2(regs[2366]), .B1(n32), .B2(regs[1854]), .ZN(
        n772) );
  NAND3_X1 U1021 ( .A1(n774), .A2(n773), .A3(n772), .ZN(curr_proc_regs[318])
         );
  NAND2_X1 U1022 ( .A1(regs[831]), .A2(n7), .ZN(n777) );
  AOI22_X1 U1023 ( .A1(n29), .A2(regs[1343]), .B1(n5), .B2(regs[319]), .ZN(
        n776) );
  AOI22_X1 U1024 ( .A1(win[4]), .A2(regs[2367]), .B1(n34), .B2(regs[1855]), 
        .ZN(n775) );
  NAND3_X1 U1025 ( .A1(n777), .A2(n776), .A3(n775), .ZN(curr_proc_regs[319])
         );
  NAND2_X1 U1026 ( .A1(regs[543]), .A2(n7), .ZN(n780) );
  AOI22_X1 U1027 ( .A1(n29), .A2(regs[1055]), .B1(n5), .B2(regs[31]), .ZN(n779) );
  AOI22_X1 U1028 ( .A1(n39), .A2(regs[2079]), .B1(n32), .B2(regs[1567]), .ZN(
        n778) );
  NAND3_X1 U1029 ( .A1(n780), .A2(n779), .A3(n778), .ZN(curr_proc_regs[31]) );
  NAND2_X1 U1030 ( .A1(regs[832]), .A2(n7), .ZN(n783) );
  AOI22_X1 U1031 ( .A1(n29), .A2(regs[1344]), .B1(n5), .B2(regs[320]), .ZN(
        n782) );
  AOI22_X1 U1032 ( .A1(n39), .A2(regs[2368]), .B1(n31), .B2(regs[1856]), .ZN(
        n781) );
  NAND3_X1 U1033 ( .A1(n783), .A2(n782), .A3(n781), .ZN(curr_proc_regs[320])
         );
  NAND2_X1 U1034 ( .A1(regs[833]), .A2(n7), .ZN(n786) );
  AOI22_X1 U1035 ( .A1(n29), .A2(regs[1345]), .B1(n5), .B2(regs[321]), .ZN(
        n785) );
  AOI22_X1 U1036 ( .A1(n39), .A2(regs[2369]), .B1(n32), .B2(regs[1857]), .ZN(
        n784) );
  NAND3_X1 U1037 ( .A1(n786), .A2(n785), .A3(n784), .ZN(curr_proc_regs[321])
         );
  NAND2_X1 U1038 ( .A1(regs[834]), .A2(n7), .ZN(n789) );
  AOI22_X1 U1039 ( .A1(n29), .A2(regs[1346]), .B1(n12), .B2(regs[322]), .ZN(
        n788) );
  AOI22_X1 U1040 ( .A1(n39), .A2(regs[2370]), .B1(n33), .B2(regs[1858]), .ZN(
        n787) );
  NAND3_X1 U1041 ( .A1(n789), .A2(n788), .A3(n787), .ZN(curr_proc_regs[322])
         );
  NAND2_X1 U1042 ( .A1(regs[835]), .A2(n7), .ZN(n792) );
  AOI22_X1 U1043 ( .A1(n29), .A2(regs[1347]), .B1(n23), .B2(regs[323]), .ZN(
        n791) );
  AOI22_X1 U1044 ( .A1(n39), .A2(regs[2371]), .B1(n32), .B2(regs[1859]), .ZN(
        n790) );
  NAND3_X1 U1045 ( .A1(n792), .A2(n791), .A3(n790), .ZN(curr_proc_regs[323])
         );
  NAND2_X1 U1046 ( .A1(regs[836]), .A2(n7), .ZN(n795) );
  AOI22_X1 U1047 ( .A1(n29), .A2(regs[1348]), .B1(n5), .B2(regs[324]), .ZN(
        n794) );
  AOI22_X1 U1048 ( .A1(n39), .A2(regs[2372]), .B1(n9), .B2(regs[1860]), .ZN(
        n793) );
  NAND3_X1 U1049 ( .A1(n795), .A2(n794), .A3(n793), .ZN(curr_proc_regs[324])
         );
  NAND2_X1 U1050 ( .A1(regs[837]), .A2(n7), .ZN(n798) );
  AOI22_X1 U1051 ( .A1(n29), .A2(regs[1349]), .B1(n5), .B2(regs[325]), .ZN(
        n797) );
  AOI22_X1 U1052 ( .A1(n39), .A2(regs[2373]), .B1(n32), .B2(regs[1861]), .ZN(
        n796) );
  NAND3_X1 U1053 ( .A1(n798), .A2(n797), .A3(n796), .ZN(curr_proc_regs[325])
         );
  NAND2_X1 U1054 ( .A1(regs[838]), .A2(n7), .ZN(n801) );
  AOI22_X1 U1055 ( .A1(n29), .A2(regs[1350]), .B1(n5), .B2(regs[326]), .ZN(
        n800) );
  AOI22_X1 U1056 ( .A1(n39), .A2(regs[2374]), .B1(n9), .B2(regs[1862]), .ZN(
        n799) );
  NAND3_X1 U1057 ( .A1(n801), .A2(n800), .A3(n799), .ZN(curr_proc_regs[326])
         );
  NAND2_X1 U1058 ( .A1(regs[839]), .A2(n7), .ZN(n804) );
  AOI22_X1 U1059 ( .A1(n29), .A2(regs[1351]), .B1(n5), .B2(regs[327]), .ZN(
        n803) );
  AOI22_X1 U1060 ( .A1(n39), .A2(regs[2375]), .B1(n32), .B2(regs[1863]), .ZN(
        n802) );
  NAND3_X1 U1061 ( .A1(n804), .A2(n803), .A3(n802), .ZN(curr_proc_regs[327])
         );
  NAND2_X1 U1062 ( .A1(regs[840]), .A2(n15), .ZN(n807) );
  AOI22_X1 U1063 ( .A1(n29), .A2(regs[1352]), .B1(n1580), .B2(regs[328]), .ZN(
        n806) );
  AOI22_X1 U1064 ( .A1(n39), .A2(regs[2376]), .B1(n3), .B2(regs[1864]), .ZN(
        n805) );
  NAND3_X1 U1065 ( .A1(n807), .A2(n806), .A3(n805), .ZN(curr_proc_regs[328])
         );
  NAND2_X1 U1066 ( .A1(regs[841]), .A2(n19), .ZN(n810) );
  AOI22_X1 U1067 ( .A1(n29), .A2(regs[1353]), .B1(n12), .B2(regs[329]), .ZN(
        n809) );
  AOI22_X1 U1068 ( .A1(n1), .A2(regs[2377]), .B1(n34), .B2(regs[1865]), .ZN(
        n808) );
  NAND3_X1 U1069 ( .A1(n810), .A2(n809), .A3(n808), .ZN(curr_proc_regs[329])
         );
  NAND2_X1 U1070 ( .A1(regs[544]), .A2(n18), .ZN(n813) );
  AOI22_X1 U1071 ( .A1(n29), .A2(regs[1056]), .B1(n27), .B2(regs[32]), .ZN(
        n812) );
  AOI22_X1 U1072 ( .A1(n8), .A2(regs[2080]), .B1(n1582), .B2(regs[1568]), .ZN(
        n811) );
  NAND3_X1 U1073 ( .A1(n813), .A2(n812), .A3(n811), .ZN(curr_proc_regs[32]) );
  NAND2_X1 U1074 ( .A1(regs[842]), .A2(n15), .ZN(n816) );
  AOI22_X1 U1075 ( .A1(n29), .A2(regs[1354]), .B1(n28), .B2(regs[330]), .ZN(
        n815) );
  AOI22_X1 U1076 ( .A1(n38), .A2(regs[2378]), .B1(n33), .B2(regs[1866]), .ZN(
        n814) );
  NAND3_X1 U1077 ( .A1(n816), .A2(n815), .A3(n814), .ZN(curr_proc_regs[330])
         );
  NAND2_X1 U1078 ( .A1(regs[843]), .A2(n11), .ZN(n819) );
  AOI22_X1 U1079 ( .A1(n29), .A2(regs[1355]), .B1(n27), .B2(regs[331]), .ZN(
        n818) );
  AOI22_X1 U1080 ( .A1(n41), .A2(regs[2379]), .B1(n9), .B2(regs[1867]), .ZN(
        n817) );
  NAND3_X1 U1081 ( .A1(n819), .A2(n818), .A3(n817), .ZN(curr_proc_regs[331])
         );
  NAND2_X1 U1082 ( .A1(regs[844]), .A2(n7), .ZN(n822) );
  AOI22_X1 U1083 ( .A1(n29), .A2(regs[1356]), .B1(n27), .B2(regs[332]), .ZN(
        n821) );
  AOI22_X1 U1084 ( .A1(n37), .A2(regs[2380]), .B1(n9), .B2(regs[1868]), .ZN(
        n820) );
  NAND3_X1 U1085 ( .A1(n822), .A2(n821), .A3(n820), .ZN(curr_proc_regs[332])
         );
  NAND2_X1 U1086 ( .A1(regs[845]), .A2(n1579), .ZN(n825) );
  AOI22_X1 U1087 ( .A1(n29), .A2(regs[1357]), .B1(n5), .B2(regs[333]), .ZN(
        n824) );
  AOI22_X1 U1088 ( .A1(n37), .A2(regs[2381]), .B1(n35), .B2(regs[1869]), .ZN(
        n823) );
  NAND3_X1 U1089 ( .A1(n825), .A2(n824), .A3(n823), .ZN(curr_proc_regs[333])
         );
  NAND2_X1 U1090 ( .A1(regs[846]), .A2(n1579), .ZN(n828) );
  AOI22_X1 U1091 ( .A1(n29), .A2(regs[1358]), .B1(n27), .B2(regs[334]), .ZN(
        n827) );
  AOI22_X1 U1092 ( .A1(n38), .A2(regs[2382]), .B1(n3), .B2(regs[1870]), .ZN(
        n826) );
  NAND3_X1 U1093 ( .A1(n828), .A2(n827), .A3(n826), .ZN(curr_proc_regs[334])
         );
  NAND2_X1 U1094 ( .A1(regs[847]), .A2(n15), .ZN(n831) );
  AOI22_X1 U1095 ( .A1(n29), .A2(regs[1359]), .B1(n27), .B2(regs[335]), .ZN(
        n830) );
  AOI22_X1 U1096 ( .A1(n38), .A2(regs[2383]), .B1(n3), .B2(regs[1871]), .ZN(
        n829) );
  NAND3_X1 U1097 ( .A1(n831), .A2(n830), .A3(n829), .ZN(curr_proc_regs[335])
         );
  NAND2_X1 U1098 ( .A1(regs[848]), .A2(n19), .ZN(n834) );
  AOI22_X1 U1099 ( .A1(n29), .A2(regs[1360]), .B1(n28), .B2(regs[336]), .ZN(
        n833) );
  AOI22_X1 U1100 ( .A1(n41), .A2(regs[2384]), .B1(n34), .B2(regs[1872]), .ZN(
        n832) );
  NAND3_X1 U1101 ( .A1(n834), .A2(n833), .A3(n832), .ZN(curr_proc_regs[336])
         );
  NAND2_X1 U1102 ( .A1(regs[849]), .A2(n7), .ZN(n837) );
  AOI22_X1 U1103 ( .A1(n29), .A2(regs[1361]), .B1(n27), .B2(regs[337]), .ZN(
        n836) );
  AOI22_X1 U1104 ( .A1(n39), .A2(regs[2385]), .B1(n1582), .B2(regs[1873]), 
        .ZN(n835) );
  NAND3_X1 U1105 ( .A1(n837), .A2(n836), .A3(n835), .ZN(curr_proc_regs[337])
         );
  NAND2_X1 U1106 ( .A1(regs[850]), .A2(n20), .ZN(n840) );
  AOI22_X1 U1107 ( .A1(n29), .A2(regs[1362]), .B1(n24), .B2(regs[338]), .ZN(
        n839) );
  AOI22_X1 U1108 ( .A1(win[4]), .A2(regs[2386]), .B1(n3), .B2(regs[1874]), 
        .ZN(n838) );
  NAND3_X1 U1109 ( .A1(n840), .A2(n839), .A3(n838), .ZN(curr_proc_regs[338])
         );
  NAND2_X1 U1110 ( .A1(regs[851]), .A2(n14), .ZN(n843) );
  AOI22_X1 U1111 ( .A1(n29), .A2(regs[1363]), .B1(n5), .B2(regs[339]), .ZN(
        n842) );
  AOI22_X1 U1112 ( .A1(win[4]), .A2(regs[2387]), .B1(n35), .B2(regs[1875]), 
        .ZN(n841) );
  NAND3_X1 U1113 ( .A1(n843), .A2(n842), .A3(n841), .ZN(curr_proc_regs[339])
         );
  NAND2_X1 U1114 ( .A1(regs[545]), .A2(n20), .ZN(n846) );
  AOI22_X1 U1115 ( .A1(n29), .A2(regs[1057]), .B1(n27), .B2(regs[33]), .ZN(
        n845) );
  AOI22_X1 U1116 ( .A1(n37), .A2(regs[2081]), .B1(n9), .B2(regs[1569]), .ZN(
        n844) );
  NAND3_X1 U1117 ( .A1(n846), .A2(n845), .A3(n844), .ZN(curr_proc_regs[33]) );
  NAND2_X1 U1118 ( .A1(regs[852]), .A2(n20), .ZN(n849) );
  AOI22_X1 U1119 ( .A1(n29), .A2(regs[1364]), .B1(n12), .B2(regs[340]), .ZN(
        n848) );
  AOI22_X1 U1120 ( .A1(win[4]), .A2(regs[2388]), .B1(n3), .B2(regs[1876]), 
        .ZN(n847) );
  NAND3_X1 U1121 ( .A1(n849), .A2(n848), .A3(n847), .ZN(curr_proc_regs[340])
         );
  NAND2_X1 U1122 ( .A1(regs[853]), .A2(n14), .ZN(n852) );
  AOI22_X1 U1123 ( .A1(n29), .A2(regs[1365]), .B1(n12), .B2(regs[341]), .ZN(
        n851) );
  AOI22_X1 U1124 ( .A1(n39), .A2(regs[2389]), .B1(n3), .B2(regs[1877]), .ZN(
        n850) );
  NAND3_X1 U1125 ( .A1(n852), .A2(n851), .A3(n850), .ZN(curr_proc_regs[341])
         );
  NAND2_X1 U1126 ( .A1(regs[854]), .A2(n20), .ZN(n855) );
  AOI22_X1 U1127 ( .A1(n29), .A2(regs[1366]), .B1(n12), .B2(regs[342]), .ZN(
        n854) );
  AOI22_X1 U1128 ( .A1(n40), .A2(regs[2390]), .B1(n35), .B2(regs[1878]), .ZN(
        n853) );
  NAND3_X1 U1129 ( .A1(n855), .A2(n854), .A3(n853), .ZN(curr_proc_regs[342])
         );
  NAND2_X1 U1130 ( .A1(regs[855]), .A2(n20), .ZN(n858) );
  AOI22_X1 U1131 ( .A1(n29), .A2(regs[1367]), .B1(n27), .B2(regs[343]), .ZN(
        n857) );
  AOI22_X1 U1132 ( .A1(n41), .A2(regs[2391]), .B1(n35), .B2(regs[1879]), .ZN(
        n856) );
  NAND3_X1 U1133 ( .A1(n858), .A2(n857), .A3(n856), .ZN(curr_proc_regs[343])
         );
  NAND2_X1 U1134 ( .A1(regs[856]), .A2(n14), .ZN(n861) );
  AOI22_X1 U1135 ( .A1(n29), .A2(regs[1368]), .B1(n1580), .B2(regs[344]), .ZN(
        n860) );
  AOI22_X1 U1136 ( .A1(n8), .A2(regs[2392]), .B1(n34), .B2(regs[1880]), .ZN(
        n859) );
  NAND3_X1 U1137 ( .A1(n861), .A2(n860), .A3(n859), .ZN(curr_proc_regs[344])
         );
  NAND2_X1 U1138 ( .A1(regs[857]), .A2(n20), .ZN(n864) );
  AOI22_X1 U1139 ( .A1(n29), .A2(regs[1369]), .B1(n26), .B2(regs[345]), .ZN(
        n863) );
  AOI22_X1 U1140 ( .A1(n38), .A2(regs[2393]), .B1(n9), .B2(regs[1881]), .ZN(
        n862) );
  NAND3_X1 U1141 ( .A1(n864), .A2(n863), .A3(n862), .ZN(curr_proc_regs[345])
         );
  NAND2_X1 U1142 ( .A1(regs[858]), .A2(n20), .ZN(n867) );
  AOI22_X1 U1143 ( .A1(n29), .A2(regs[1370]), .B1(n24), .B2(regs[346]), .ZN(
        n866) );
  AOI22_X1 U1144 ( .A1(n39), .A2(regs[2394]), .B1(n35), .B2(regs[1882]), .ZN(
        n865) );
  NAND3_X1 U1145 ( .A1(n867), .A2(n866), .A3(n865), .ZN(curr_proc_regs[346])
         );
  NAND2_X1 U1146 ( .A1(regs[859]), .A2(n20), .ZN(n870) );
  AOI22_X1 U1147 ( .A1(n29), .A2(regs[1371]), .B1(n27), .B2(regs[347]), .ZN(
        n869) );
  AOI22_X1 U1148 ( .A1(n1), .A2(regs[2395]), .B1(n3), .B2(regs[1883]), .ZN(
        n868) );
  NAND3_X1 U1149 ( .A1(n870), .A2(n869), .A3(n868), .ZN(curr_proc_regs[347])
         );
  NAND2_X1 U1150 ( .A1(regs[860]), .A2(n13), .ZN(n873) );
  AOI22_X1 U1151 ( .A1(n29), .A2(regs[1372]), .B1(n26), .B2(regs[348]), .ZN(
        n872) );
  AOI22_X1 U1152 ( .A1(n41), .A2(regs[2396]), .B1(n31), .B2(regs[1884]), .ZN(
        n871) );
  NAND3_X1 U1153 ( .A1(n873), .A2(n872), .A3(n871), .ZN(curr_proc_regs[348])
         );
  NAND2_X1 U1154 ( .A1(regs[861]), .A2(n13), .ZN(n876) );
  AOI22_X1 U1155 ( .A1(n29), .A2(regs[1373]), .B1(n24), .B2(regs[349]), .ZN(
        n875) );
  AOI22_X1 U1156 ( .A1(n36), .A2(regs[2397]), .B1(n31), .B2(regs[1885]), .ZN(
        n874) );
  NAND3_X1 U1157 ( .A1(n876), .A2(n875), .A3(n874), .ZN(curr_proc_regs[349])
         );
  NAND2_X1 U1158 ( .A1(regs[546]), .A2(n13), .ZN(n879) );
  AOI22_X1 U1159 ( .A1(n29), .A2(regs[1058]), .B1(n12), .B2(regs[34]), .ZN(
        n878) );
  AOI22_X1 U1160 ( .A1(n1), .A2(regs[2082]), .B1(n31), .B2(regs[1570]), .ZN(
        n877) );
  NAND3_X1 U1161 ( .A1(n879), .A2(n878), .A3(n877), .ZN(curr_proc_regs[34]) );
  NAND2_X1 U1162 ( .A1(regs[862]), .A2(n13), .ZN(n882) );
  AOI22_X1 U1163 ( .A1(n29), .A2(regs[1374]), .B1(n24), .B2(regs[350]), .ZN(
        n881) );
  AOI22_X1 U1164 ( .A1(n41), .A2(regs[2398]), .B1(n31), .B2(regs[1886]), .ZN(
        n880) );
  NAND3_X1 U1165 ( .A1(n882), .A2(n881), .A3(n880), .ZN(curr_proc_regs[350])
         );
  NAND2_X1 U1166 ( .A1(regs[863]), .A2(n13), .ZN(n885) );
  AOI22_X1 U1167 ( .A1(n29), .A2(regs[1375]), .B1(n22), .B2(regs[351]), .ZN(
        n884) );
  AOI22_X1 U1168 ( .A1(n41), .A2(regs[2399]), .B1(n31), .B2(regs[1887]), .ZN(
        n883) );
  NAND3_X1 U1169 ( .A1(n885), .A2(n884), .A3(n883), .ZN(curr_proc_regs[351])
         );
  NAND2_X1 U1170 ( .A1(regs[864]), .A2(n13), .ZN(n888) );
  AOI22_X1 U1171 ( .A1(n29), .A2(regs[1376]), .B1(n1580), .B2(regs[352]), .ZN(
        n887) );
  AOI22_X1 U1172 ( .A1(n1), .A2(regs[2400]), .B1(n31), .B2(regs[1888]), .ZN(
        n886) );
  NAND3_X1 U1173 ( .A1(n888), .A2(n887), .A3(n886), .ZN(curr_proc_regs[352])
         );
  NAND2_X1 U1174 ( .A1(regs[865]), .A2(n13), .ZN(n891) );
  AOI22_X1 U1175 ( .A1(n29), .A2(regs[1377]), .B1(n28), .B2(regs[353]), .ZN(
        n890) );
  AOI22_X1 U1176 ( .A1(win[4]), .A2(regs[2401]), .B1(n31), .B2(regs[1889]), 
        .ZN(n889) );
  NAND3_X1 U1177 ( .A1(n891), .A2(n890), .A3(n889), .ZN(curr_proc_regs[353])
         );
  NAND2_X1 U1178 ( .A1(regs[866]), .A2(n13), .ZN(n894) );
  AOI22_X1 U1179 ( .A1(n29), .A2(regs[1378]), .B1(n5), .B2(regs[354]), .ZN(
        n893) );
  AOI22_X1 U1180 ( .A1(n38), .A2(regs[2402]), .B1(n31), .B2(regs[1890]), .ZN(
        n892) );
  NAND3_X1 U1181 ( .A1(n894), .A2(n893), .A3(n892), .ZN(curr_proc_regs[354])
         );
  NAND2_X1 U1182 ( .A1(regs[867]), .A2(n13), .ZN(n897) );
  AOI22_X1 U1183 ( .A1(n29), .A2(regs[1379]), .B1(n12), .B2(regs[355]), .ZN(
        n896) );
  AOI22_X1 U1184 ( .A1(win[4]), .A2(regs[2403]), .B1(n31), .B2(regs[1891]), 
        .ZN(n895) );
  NAND3_X1 U1185 ( .A1(n897), .A2(n896), .A3(n895), .ZN(curr_proc_regs[355])
         );
  NAND2_X1 U1186 ( .A1(regs[868]), .A2(n13), .ZN(n900) );
  AOI22_X1 U1187 ( .A1(n29), .A2(regs[1380]), .B1(n12), .B2(regs[356]), .ZN(
        n899) );
  AOI22_X1 U1188 ( .A1(n41), .A2(regs[2404]), .B1(n31), .B2(regs[1892]), .ZN(
        n898) );
  NAND3_X1 U1189 ( .A1(n900), .A2(n899), .A3(n898), .ZN(curr_proc_regs[356])
         );
  NAND2_X1 U1190 ( .A1(regs[869]), .A2(n13), .ZN(n903) );
  AOI22_X1 U1191 ( .A1(n29), .A2(regs[1381]), .B1(n21), .B2(regs[357]), .ZN(
        n902) );
  AOI22_X1 U1192 ( .A1(n41), .A2(regs[2405]), .B1(n31), .B2(regs[1893]), .ZN(
        n901) );
  NAND3_X1 U1193 ( .A1(n903), .A2(n902), .A3(n901), .ZN(curr_proc_regs[357])
         );
  NAND2_X1 U1194 ( .A1(regs[870]), .A2(n11), .ZN(n906) );
  AOI22_X1 U1195 ( .A1(n29), .A2(regs[1382]), .B1(n12), .B2(regs[358]), .ZN(
        n905) );
  AOI22_X1 U1196 ( .A1(n41), .A2(regs[2406]), .B1(n34), .B2(regs[1894]), .ZN(
        n904) );
  NAND3_X1 U1197 ( .A1(n906), .A2(n905), .A3(n904), .ZN(curr_proc_regs[358])
         );
  NAND2_X1 U1198 ( .A1(regs[871]), .A2(n11), .ZN(n909) );
  AOI22_X1 U1199 ( .A1(n29), .A2(regs[1383]), .B1(n27), .B2(regs[359]), .ZN(
        n908) );
  AOI22_X1 U1200 ( .A1(n39), .A2(regs[2407]), .B1(n9), .B2(regs[1895]), .ZN(
        n907) );
  NAND3_X1 U1201 ( .A1(n909), .A2(n908), .A3(n907), .ZN(curr_proc_regs[359])
         );
  NAND2_X1 U1202 ( .A1(regs[547]), .A2(n11), .ZN(n912) );
  AOI22_X1 U1203 ( .A1(n29), .A2(regs[1059]), .B1(n27), .B2(regs[35]), .ZN(
        n911) );
  AOI22_X1 U1204 ( .A1(n38), .A2(regs[2083]), .B1(n9), .B2(regs[1571]), .ZN(
        n910) );
  NAND3_X1 U1205 ( .A1(n912), .A2(n911), .A3(n910), .ZN(curr_proc_regs[35]) );
  NAND2_X1 U1206 ( .A1(regs[872]), .A2(n11), .ZN(n915) );
  AOI22_X1 U1207 ( .A1(n29), .A2(regs[1384]), .B1(n24), .B2(regs[360]), .ZN(
        n914) );
  AOI22_X1 U1208 ( .A1(win[4]), .A2(regs[2408]), .B1(n35), .B2(regs[1896]), 
        .ZN(n913) );
  NAND3_X1 U1209 ( .A1(n915), .A2(n914), .A3(n913), .ZN(curr_proc_regs[360])
         );
  NAND2_X1 U1210 ( .A1(regs[873]), .A2(n11), .ZN(n918) );
  AOI22_X1 U1211 ( .A1(n29), .A2(regs[1385]), .B1(n12), .B2(regs[361]), .ZN(
        n917) );
  AOI22_X1 U1212 ( .A1(win[4]), .A2(regs[2409]), .B1(n3), .B2(regs[1897]), 
        .ZN(n916) );
  NAND3_X1 U1213 ( .A1(n918), .A2(n917), .A3(n916), .ZN(curr_proc_regs[361])
         );
  NAND2_X1 U1214 ( .A1(regs[874]), .A2(n11), .ZN(n921) );
  AOI22_X1 U1215 ( .A1(n29), .A2(regs[1386]), .B1(n12), .B2(regs[362]), .ZN(
        n920) );
  AOI22_X1 U1216 ( .A1(win[4]), .A2(regs[2410]), .B1(n3), .B2(regs[1898]), 
        .ZN(n919) );
  NAND3_X1 U1217 ( .A1(n921), .A2(n920), .A3(n919), .ZN(curr_proc_regs[362])
         );
  NAND2_X1 U1218 ( .A1(regs[875]), .A2(n11), .ZN(n924) );
  AOI22_X1 U1219 ( .A1(n29), .A2(regs[1387]), .B1(n27), .B2(regs[363]), .ZN(
        n923) );
  AOI22_X1 U1220 ( .A1(n1), .A2(regs[2411]), .B1(n34), .B2(regs[1899]), .ZN(
        n922) );
  NAND3_X1 U1221 ( .A1(n924), .A2(n923), .A3(n922), .ZN(curr_proc_regs[363])
         );
  NAND2_X1 U1222 ( .A1(regs[876]), .A2(n11), .ZN(n927) );
  AOI22_X1 U1223 ( .A1(n29), .A2(regs[1388]), .B1(n1580), .B2(regs[364]), .ZN(
        n926) );
  AOI22_X1 U1224 ( .A1(n39), .A2(regs[2412]), .B1(n33), .B2(regs[1900]), .ZN(
        n925) );
  NAND3_X1 U1225 ( .A1(n927), .A2(n926), .A3(n925), .ZN(curr_proc_regs[364])
         );
  NAND2_X1 U1226 ( .A1(regs[877]), .A2(n11), .ZN(n930) );
  AOI22_X1 U1227 ( .A1(n29), .A2(regs[1389]), .B1(n27), .B2(regs[365]), .ZN(
        n929) );
  AOI22_X1 U1228 ( .A1(n39), .A2(regs[2413]), .B1(n34), .B2(regs[1901]), .ZN(
        n928) );
  NAND3_X1 U1229 ( .A1(n930), .A2(n929), .A3(n928), .ZN(curr_proc_regs[365])
         );
  NAND2_X1 U1230 ( .A1(regs[878]), .A2(n11), .ZN(n933) );
  AOI22_X1 U1231 ( .A1(n29), .A2(regs[1390]), .B1(n27), .B2(regs[366]), .ZN(
        n932) );
  AOI22_X1 U1232 ( .A1(n41), .A2(regs[2414]), .B1(n9), .B2(regs[1902]), .ZN(
        n931) );
  NAND3_X1 U1233 ( .A1(n933), .A2(n932), .A3(n931), .ZN(curr_proc_regs[366])
         );
  NAND2_X1 U1234 ( .A1(regs[879]), .A2(n11), .ZN(n936) );
  AOI22_X1 U1235 ( .A1(n29), .A2(regs[1391]), .B1(n27), .B2(regs[367]), .ZN(
        n935) );
  AOI22_X1 U1236 ( .A1(n40), .A2(regs[2415]), .B1(n9), .B2(regs[1903]), .ZN(
        n934) );
  NAND3_X1 U1237 ( .A1(n936), .A2(n935), .A3(n934), .ZN(curr_proc_regs[367])
         );
  NAND2_X1 U1238 ( .A1(regs[880]), .A2(n16), .ZN(n939) );
  AOI22_X1 U1239 ( .A1(n29), .A2(regs[1392]), .B1(n26), .B2(regs[368]), .ZN(
        n938) );
  AOI22_X1 U1240 ( .A1(n36), .A2(regs[2416]), .B1(n33), .B2(regs[1904]), .ZN(
        n937) );
  NAND3_X1 U1241 ( .A1(n939), .A2(n938), .A3(n937), .ZN(curr_proc_regs[368])
         );
  NAND2_X1 U1242 ( .A1(regs[881]), .A2(n1579), .ZN(n942) );
  AOI22_X1 U1243 ( .A1(n29), .A2(regs[1393]), .B1(n5), .B2(regs[369]), .ZN(
        n941) );
  AOI22_X1 U1244 ( .A1(n37), .A2(regs[2417]), .B1(n9), .B2(regs[1905]), .ZN(
        n940) );
  NAND3_X1 U1245 ( .A1(n942), .A2(n941), .A3(n940), .ZN(curr_proc_regs[369])
         );
  NAND2_X1 U1246 ( .A1(regs[548]), .A2(n11), .ZN(n945) );
  AOI22_X1 U1247 ( .A1(n29), .A2(regs[1060]), .B1(n5), .B2(regs[36]), .ZN(n944) );
  AOI22_X1 U1248 ( .A1(n39), .A2(regs[2084]), .B1(n9), .B2(regs[1572]), .ZN(
        n943) );
  NAND3_X1 U1249 ( .A1(n945), .A2(n944), .A3(n943), .ZN(curr_proc_regs[36]) );
  NAND2_X1 U1250 ( .A1(regs[882]), .A2(n1579), .ZN(n948) );
  AOI22_X1 U1251 ( .A1(n29), .A2(regs[1394]), .B1(n27), .B2(regs[370]), .ZN(
        n947) );
  AOI22_X1 U1252 ( .A1(n40), .A2(regs[2418]), .B1(n35), .B2(regs[1906]), .ZN(
        n946) );
  NAND3_X1 U1253 ( .A1(n948), .A2(n947), .A3(n946), .ZN(curr_proc_regs[370])
         );
  NAND2_X1 U1254 ( .A1(regs[883]), .A2(n13), .ZN(n951) );
  AOI22_X1 U1255 ( .A1(n29), .A2(regs[1395]), .B1(n27), .B2(regs[371]), .ZN(
        n950) );
  AOI22_X1 U1256 ( .A1(n41), .A2(regs[2419]), .B1(n31), .B2(regs[1907]), .ZN(
        n949) );
  NAND3_X1 U1257 ( .A1(n951), .A2(n950), .A3(n949), .ZN(curr_proc_regs[371])
         );
  NAND2_X1 U1258 ( .A1(regs[884]), .A2(n11), .ZN(n954) );
  AOI22_X1 U1259 ( .A1(n29), .A2(regs[1396]), .B1(n27), .B2(regs[372]), .ZN(
        n953) );
  AOI22_X1 U1260 ( .A1(n38), .A2(regs[2420]), .B1(n3), .B2(regs[1908]), .ZN(
        n952) );
  NAND3_X1 U1261 ( .A1(n954), .A2(n953), .A3(n952), .ZN(curr_proc_regs[372])
         );
  NAND2_X1 U1262 ( .A1(regs[885]), .A2(n13), .ZN(n957) );
  AOI22_X1 U1263 ( .A1(n29), .A2(regs[1397]), .B1(n27), .B2(regs[373]), .ZN(
        n956) );
  AOI22_X1 U1264 ( .A1(n8), .A2(regs[2421]), .B1(n3), .B2(regs[1909]), .ZN(
        n955) );
  NAND3_X1 U1265 ( .A1(n957), .A2(n956), .A3(n955), .ZN(curr_proc_regs[373])
         );
  NAND2_X1 U1266 ( .A1(regs[886]), .A2(n17), .ZN(n960) );
  AOI22_X1 U1267 ( .A1(n29), .A2(regs[1398]), .B1(n27), .B2(regs[374]), .ZN(
        n959) );
  AOI22_X1 U1268 ( .A1(n37), .A2(regs[2422]), .B1(n33), .B2(regs[1910]), .ZN(
        n958) );
  NAND3_X1 U1269 ( .A1(n960), .A2(n959), .A3(n958), .ZN(curr_proc_regs[374])
         );
  NAND2_X1 U1270 ( .A1(regs[887]), .A2(n14), .ZN(n963) );
  AOI22_X1 U1271 ( .A1(n29), .A2(regs[1399]), .B1(n5), .B2(regs[375]), .ZN(
        n962) );
  AOI22_X1 U1272 ( .A1(n38), .A2(regs[2423]), .B1(n34), .B2(regs[1911]), .ZN(
        n961) );
  NAND3_X1 U1273 ( .A1(n963), .A2(n962), .A3(n961), .ZN(curr_proc_regs[375])
         );
  NAND2_X1 U1274 ( .A1(regs[888]), .A2(n13), .ZN(n966) );
  AOI22_X1 U1275 ( .A1(n29), .A2(regs[1400]), .B1(n27), .B2(regs[376]), .ZN(
        n965) );
  AOI22_X1 U1276 ( .A1(n38), .A2(regs[2424]), .B1(n9), .B2(regs[1912]), .ZN(
        n964) );
  NAND3_X1 U1277 ( .A1(n966), .A2(n965), .A3(n964), .ZN(curr_proc_regs[376])
         );
  NAND2_X1 U1278 ( .A1(regs[889]), .A2(n1579), .ZN(n969) );
  AOI22_X1 U1279 ( .A1(n29), .A2(regs[1401]), .B1(n27), .B2(regs[377]), .ZN(
        n968) );
  AOI22_X1 U1280 ( .A1(n41), .A2(regs[2425]), .B1(n9), .B2(regs[1913]), .ZN(
        n967) );
  NAND3_X1 U1281 ( .A1(n969), .A2(n968), .A3(n967), .ZN(curr_proc_regs[377])
         );
  NAND2_X1 U1282 ( .A1(regs[890]), .A2(n18), .ZN(n972) );
  AOI22_X1 U1283 ( .A1(n29), .A2(regs[1402]), .B1(n12), .B2(regs[378]), .ZN(
        n971) );
  AOI22_X1 U1284 ( .A1(n37), .A2(regs[2426]), .B1(n35), .B2(regs[1914]), .ZN(
        n970) );
  NAND3_X1 U1285 ( .A1(n972), .A2(n971), .A3(n970), .ZN(curr_proc_regs[378])
         );
  NAND2_X1 U1286 ( .A1(regs[891]), .A2(n7), .ZN(n975) );
  AOI22_X1 U1287 ( .A1(n29), .A2(regs[1403]), .B1(n27), .B2(regs[379]), .ZN(
        n974) );
  AOI22_X1 U1288 ( .A1(n8), .A2(regs[2427]), .B1(n35), .B2(regs[1915]), .ZN(
        n973) );
  NAND3_X1 U1289 ( .A1(n975), .A2(n974), .A3(n973), .ZN(curr_proc_regs[379])
         );
  NAND2_X1 U1290 ( .A1(regs[549]), .A2(n7), .ZN(n978) );
  AOI22_X1 U1291 ( .A1(n29), .A2(regs[1061]), .B1(n12), .B2(regs[37]), .ZN(
        n977) );
  AOI22_X1 U1292 ( .A1(n36), .A2(regs[2085]), .B1(n3), .B2(regs[1573]), .ZN(
        n976) );
  NAND3_X1 U1293 ( .A1(n978), .A2(n977), .A3(n976), .ZN(curr_proc_regs[37]) );
  NAND2_X1 U1294 ( .A1(regs[892]), .A2(n15), .ZN(n981) );
  AOI22_X1 U1295 ( .A1(n29), .A2(regs[1404]), .B1(n27), .B2(regs[380]), .ZN(
        n980) );
  AOI22_X1 U1296 ( .A1(n1), .A2(regs[2428]), .B1(n3), .B2(regs[1916]), .ZN(
        n979) );
  NAND3_X1 U1297 ( .A1(n981), .A2(n980), .A3(n979), .ZN(curr_proc_regs[380])
         );
  NAND2_X1 U1298 ( .A1(regs[893]), .A2(n18), .ZN(n984) );
  AOI22_X1 U1299 ( .A1(n29), .A2(regs[1405]), .B1(n5), .B2(regs[381]), .ZN(
        n983) );
  AOI22_X1 U1300 ( .A1(n1), .A2(regs[2429]), .B1(n3), .B2(regs[1917]), .ZN(
        n982) );
  NAND3_X1 U1301 ( .A1(n984), .A2(n983), .A3(n982), .ZN(curr_proc_regs[381])
         );
  NAND2_X1 U1302 ( .A1(regs[894]), .A2(n19), .ZN(n987) );
  AOI22_X1 U1303 ( .A1(n29), .A2(regs[1406]), .B1(n27), .B2(regs[382]), .ZN(
        n986) );
  AOI22_X1 U1304 ( .A1(n8), .A2(regs[2430]), .B1(n3), .B2(regs[1918]), .ZN(
        n985) );
  NAND3_X1 U1305 ( .A1(n987), .A2(n986), .A3(n985), .ZN(curr_proc_regs[382])
         );
  NAND2_X1 U1306 ( .A1(regs[895]), .A2(n7), .ZN(n990) );
  AOI22_X1 U1307 ( .A1(n29), .A2(regs[1407]), .B1(n25), .B2(regs[383]), .ZN(
        n989) );
  AOI22_X1 U1308 ( .A1(n10), .A2(regs[2431]), .B1(n34), .B2(regs[1919]), .ZN(
        n988) );
  NAND3_X1 U1309 ( .A1(n990), .A2(n989), .A3(n988), .ZN(curr_proc_regs[383])
         );
  NAND2_X1 U1310 ( .A1(regs[896]), .A2(n16), .ZN(n993) );
  AOI22_X1 U1311 ( .A1(n29), .A2(regs[1408]), .B1(n28), .B2(regs[384]), .ZN(
        n992) );
  AOI22_X1 U1312 ( .A1(n8), .A2(regs[2432]), .B1(n34), .B2(regs[1920]), .ZN(
        n991) );
  NAND3_X1 U1313 ( .A1(n993), .A2(n992), .A3(n991), .ZN(curr_proc_regs[384])
         );
  NAND2_X1 U1314 ( .A1(regs[897]), .A2(n18), .ZN(n996) );
  AOI22_X1 U1315 ( .A1(n29), .A2(regs[1409]), .B1(n5), .B2(regs[385]), .ZN(
        n995) );
  AOI22_X1 U1316 ( .A1(n8), .A2(regs[2433]), .B1(n33), .B2(regs[1921]), .ZN(
        n994) );
  NAND3_X1 U1317 ( .A1(n996), .A2(n995), .A3(n994), .ZN(curr_proc_regs[385])
         );
  NAND2_X1 U1318 ( .A1(regs[898]), .A2(n7), .ZN(n999) );
  AOI22_X1 U1319 ( .A1(n29), .A2(regs[1410]), .B1(n26), .B2(regs[386]), .ZN(
        n998) );
  AOI22_X1 U1320 ( .A1(n4), .A2(regs[2434]), .B1(n34), .B2(regs[1922]), .ZN(
        n997) );
  NAND3_X1 U1321 ( .A1(n999), .A2(n998), .A3(n997), .ZN(curr_proc_regs[386])
         );
  NAND2_X1 U1322 ( .A1(regs[899]), .A2(n7), .ZN(n1002) );
  AOI22_X1 U1323 ( .A1(n29), .A2(regs[1411]), .B1(n1580), .B2(regs[387]), .ZN(
        n1001) );
  AOI22_X1 U1324 ( .A1(n41), .A2(regs[2435]), .B1(n34), .B2(regs[1923]), .ZN(
        n1000) );
  NAND3_X1 U1325 ( .A1(n1002), .A2(n1001), .A3(n1000), .ZN(curr_proc_regs[387]) );
  NAND2_X1 U1326 ( .A1(regs[900]), .A2(n11), .ZN(n1005) );
  AOI22_X1 U1327 ( .A1(n29), .A2(regs[1412]), .B1(n5), .B2(regs[388]), .ZN(
        n1004) );
  AOI22_X1 U1328 ( .A1(n8), .A2(regs[2436]), .B1(n3), .B2(regs[1924]), .ZN(
        n1003) );
  NAND3_X1 U1329 ( .A1(n1005), .A2(n1004), .A3(n1003), .ZN(curr_proc_regs[388]) );
  NAND2_X1 U1330 ( .A1(regs[901]), .A2(n15), .ZN(n1008) );
  AOI22_X1 U1331 ( .A1(n29), .A2(regs[1413]), .B1(n25), .B2(regs[389]), .ZN(
        n1007) );
  AOI22_X1 U1332 ( .A1(win[4]), .A2(regs[2437]), .B1(n35), .B2(regs[1925]), 
        .ZN(n1006) );
  NAND3_X1 U1333 ( .A1(n1008), .A2(n1007), .A3(n1006), .ZN(curr_proc_regs[389]) );
  NAND2_X1 U1334 ( .A1(regs[550]), .A2(n13), .ZN(n1011) );
  AOI22_X1 U1335 ( .A1(n29), .A2(regs[1062]), .B1(n5), .B2(regs[38]), .ZN(
        n1010) );
  AOI22_X1 U1336 ( .A1(win[4]), .A2(regs[2086]), .B1(n34), .B2(regs[1574]), 
        .ZN(n1009) );
  NAND3_X1 U1337 ( .A1(n1011), .A2(n1010), .A3(n1009), .ZN(curr_proc_regs[38])
         );
  NAND2_X1 U1338 ( .A1(regs[902]), .A2(n11), .ZN(n1014) );
  AOI22_X1 U1339 ( .A1(n29), .A2(regs[1414]), .B1(n24), .B2(regs[390]), .ZN(
        n1013) );
  AOI22_X1 U1340 ( .A1(win[4]), .A2(regs[2438]), .B1(n3), .B2(regs[1926]), 
        .ZN(n1012) );
  NAND3_X1 U1341 ( .A1(n1014), .A2(n1013), .A3(n1012), .ZN(curr_proc_regs[390]) );
  NAND2_X1 U1342 ( .A1(regs[903]), .A2(n11), .ZN(n1017) );
  AOI22_X1 U1343 ( .A1(n29), .A2(regs[1415]), .B1(n1580), .B2(regs[391]), .ZN(
        n1016) );
  AOI22_X1 U1344 ( .A1(n4), .A2(regs[2439]), .B1(n3), .B2(regs[1927]), .ZN(
        n1015) );
  NAND3_X1 U1345 ( .A1(n1017), .A2(n1016), .A3(n1015), .ZN(curr_proc_regs[391]) );
  NAND2_X1 U1346 ( .A1(regs[904]), .A2(n7), .ZN(n1020) );
  AOI22_X1 U1347 ( .A1(n29), .A2(regs[1416]), .B1(n24), .B2(regs[392]), .ZN(
        n1019) );
  AOI22_X1 U1348 ( .A1(n4), .A2(regs[2440]), .B1(n34), .B2(regs[1928]), .ZN(
        n1018) );
  NAND3_X1 U1349 ( .A1(n1020), .A2(n1019), .A3(n1018), .ZN(curr_proc_regs[392]) );
  NAND2_X1 U1350 ( .A1(regs[905]), .A2(n15), .ZN(n1023) );
  AOI22_X1 U1351 ( .A1(n29), .A2(regs[1417]), .B1(n12), .B2(regs[393]), .ZN(
        n1022) );
  AOI22_X1 U1352 ( .A1(n8), .A2(regs[2441]), .B1(n9), .B2(regs[1929]), .ZN(
        n1021) );
  NAND3_X1 U1353 ( .A1(n1023), .A2(n1022), .A3(n1021), .ZN(curr_proc_regs[393]) );
  NAND2_X1 U1354 ( .A1(regs[906]), .A2(n1579), .ZN(n1026) );
  AOI22_X1 U1355 ( .A1(n29), .A2(regs[1418]), .B1(n12), .B2(regs[394]), .ZN(
        n1025) );
  AOI22_X1 U1356 ( .A1(n10), .A2(regs[2442]), .B1(n9), .B2(regs[1930]), .ZN(
        n1024) );
  NAND3_X1 U1357 ( .A1(n1026), .A2(n1025), .A3(n1024), .ZN(curr_proc_regs[394]) );
  NAND2_X1 U1358 ( .A1(regs[907]), .A2(n16), .ZN(n1029) );
  AOI22_X1 U1359 ( .A1(n29), .A2(regs[1419]), .B1(n26), .B2(regs[395]), .ZN(
        n1028) );
  AOI22_X1 U1360 ( .A1(n40), .A2(regs[2443]), .B1(n35), .B2(regs[1931]), .ZN(
        n1027) );
  NAND3_X1 U1361 ( .A1(n1029), .A2(n1028), .A3(n1027), .ZN(curr_proc_regs[395]) );
  NAND2_X1 U1362 ( .A1(regs[908]), .A2(n13), .ZN(n1032) );
  AOI22_X1 U1363 ( .A1(n29), .A2(regs[1420]), .B1(n5), .B2(regs[396]), .ZN(
        n1031) );
  AOI22_X1 U1364 ( .A1(n37), .A2(regs[2444]), .B1(n3), .B2(regs[1932]), .ZN(
        n1030) );
  NAND3_X1 U1365 ( .A1(n1032), .A2(n1031), .A3(n1030), .ZN(curr_proc_regs[396]) );
  NAND2_X1 U1366 ( .A1(regs[909]), .A2(n1579), .ZN(n1035) );
  AOI22_X1 U1367 ( .A1(n29), .A2(regs[1421]), .B1(n24), .B2(regs[397]), .ZN(
        n1034) );
  AOI22_X1 U1368 ( .A1(win[4]), .A2(regs[2445]), .B1(n3), .B2(regs[1933]), 
        .ZN(n1033) );
  NAND3_X1 U1369 ( .A1(n1035), .A2(n1034), .A3(n1033), .ZN(curr_proc_regs[397]) );
  NAND2_X1 U1370 ( .A1(regs[910]), .A2(n15), .ZN(n1038) );
  AOI22_X1 U1371 ( .A1(n29), .A2(regs[1422]), .B1(n12), .B2(regs[398]), .ZN(
        n1037) );
  AOI22_X1 U1372 ( .A1(win[4]), .A2(regs[2446]), .B1(n1582), .B2(regs[1934]), 
        .ZN(n1036) );
  NAND3_X1 U1373 ( .A1(n1038), .A2(n1037), .A3(n1036), .ZN(curr_proc_regs[398]) );
  NAND2_X1 U1374 ( .A1(regs[911]), .A2(n15), .ZN(n1041) );
  AOI22_X1 U1375 ( .A1(n29), .A2(regs[1423]), .B1(n28), .B2(regs[399]), .ZN(
        n1040) );
  AOI22_X1 U1376 ( .A1(win[4]), .A2(regs[2447]), .B1(n34), .B2(regs[1935]), 
        .ZN(n1039) );
  NAND3_X1 U1377 ( .A1(n1041), .A2(n1040), .A3(n1039), .ZN(curr_proc_regs[399]) );
  NAND2_X1 U1378 ( .A1(regs[551]), .A2(n15), .ZN(n1044) );
  AOI22_X1 U1379 ( .A1(n29), .A2(regs[1063]), .B1(n25), .B2(regs[39]), .ZN(
        n1043) );
  AOI22_X1 U1380 ( .A1(win[4]), .A2(regs[2087]), .B1(n33), .B2(regs[1575]), 
        .ZN(n1042) );
  NAND3_X1 U1381 ( .A1(n1044), .A2(n1043), .A3(n1042), .ZN(curr_proc_regs[39])
         );
  NAND2_X1 U1382 ( .A1(regs[515]), .A2(n15), .ZN(n1047) );
  AOI22_X1 U1383 ( .A1(n29), .A2(regs[1027]), .B1(n5), .B2(regs[3]), .ZN(n1046) );
  AOI22_X1 U1384 ( .A1(win[4]), .A2(regs[2051]), .B1(n9), .B2(regs[1539]), 
        .ZN(n1045) );
  NAND3_X1 U1385 ( .A1(n1047), .A2(n1046), .A3(n1045), .ZN(curr_proc_regs[3])
         );
  NAND2_X1 U1386 ( .A1(regs[912]), .A2(n15), .ZN(n1050) );
  AOI22_X1 U1387 ( .A1(n29), .A2(regs[1424]), .B1(n5), .B2(regs[400]), .ZN(
        n1049) );
  AOI22_X1 U1388 ( .A1(win[4]), .A2(regs[2448]), .B1(n9), .B2(regs[1936]), 
        .ZN(n1048) );
  NAND3_X1 U1389 ( .A1(n1050), .A2(n1049), .A3(n1048), .ZN(curr_proc_regs[400]) );
  NAND2_X1 U1390 ( .A1(regs[913]), .A2(n15), .ZN(n1053) );
  AOI22_X1 U1391 ( .A1(n29), .A2(regs[1425]), .B1(n26), .B2(regs[401]), .ZN(
        n1052) );
  AOI22_X1 U1392 ( .A1(win[4]), .A2(regs[2449]), .B1(n9), .B2(regs[1937]), 
        .ZN(n1051) );
  NAND3_X1 U1393 ( .A1(n1053), .A2(n1052), .A3(n1051), .ZN(curr_proc_regs[401]) );
  NAND2_X1 U1394 ( .A1(regs[914]), .A2(n15), .ZN(n1056) );
  AOI22_X1 U1395 ( .A1(n29), .A2(regs[1426]), .B1(n1580), .B2(regs[402]), .ZN(
        n1055) );
  AOI22_X1 U1396 ( .A1(win[4]), .A2(regs[2450]), .B1(n9), .B2(regs[1938]), 
        .ZN(n1054) );
  NAND3_X1 U1397 ( .A1(n1056), .A2(n1055), .A3(n1054), .ZN(curr_proc_regs[402]) );
  NAND2_X1 U1398 ( .A1(regs[915]), .A2(n15), .ZN(n1059) );
  AOI22_X1 U1399 ( .A1(n29), .A2(regs[1427]), .B1(n24), .B2(regs[403]), .ZN(
        n1058) );
  AOI22_X1 U1400 ( .A1(win[4]), .A2(regs[2451]), .B1(n35), .B2(regs[1939]), 
        .ZN(n1057) );
  NAND3_X1 U1401 ( .A1(n1059), .A2(n1058), .A3(n1057), .ZN(curr_proc_regs[403]) );
  NAND2_X1 U1402 ( .A1(regs[916]), .A2(n15), .ZN(n1062) );
  AOI22_X1 U1403 ( .A1(n29), .A2(regs[1428]), .B1(n12), .B2(regs[404]), .ZN(
        n1061) );
  AOI22_X1 U1404 ( .A1(win[4]), .A2(regs[2452]), .B1(n35), .B2(regs[1940]), 
        .ZN(n1060) );
  NAND3_X1 U1405 ( .A1(n1062), .A2(n1061), .A3(n1060), .ZN(curr_proc_regs[404]) );
  NAND2_X1 U1406 ( .A1(regs[917]), .A2(n15), .ZN(n1065) );
  AOI22_X1 U1407 ( .A1(n29), .A2(regs[1429]), .B1(n12), .B2(regs[405]), .ZN(
        n1064) );
  AOI22_X1 U1408 ( .A1(win[4]), .A2(regs[2453]), .B1(n1582), .B2(regs[1941]), 
        .ZN(n1063) );
  NAND3_X1 U1409 ( .A1(n1065), .A2(n1064), .A3(n1063), .ZN(curr_proc_regs[405]) );
  NAND2_X1 U1410 ( .A1(regs[918]), .A2(n15), .ZN(n1068) );
  AOI22_X1 U1411 ( .A1(n29), .A2(regs[1430]), .B1(n5), .B2(regs[406]), .ZN(
        n1067) );
  AOI22_X1 U1412 ( .A1(n38), .A2(regs[2454]), .B1(n3), .B2(regs[1942]), .ZN(
        n1066) );
  NAND3_X1 U1413 ( .A1(n1068), .A2(n1067), .A3(n1066), .ZN(curr_proc_regs[406]) );
  NAND2_X1 U1414 ( .A1(regs[919]), .A2(n11), .ZN(n1071) );
  AOI22_X1 U1415 ( .A1(n29), .A2(regs[1431]), .B1(n12), .B2(regs[407]), .ZN(
        n1070) );
  AOI22_X1 U1416 ( .A1(n38), .A2(regs[2455]), .B1(n35), .B2(regs[1943]), .ZN(
        n1069) );
  NAND3_X1 U1417 ( .A1(n1071), .A2(n1070), .A3(n1069), .ZN(curr_proc_regs[407]) );
  NAND2_X1 U1418 ( .A1(regs[920]), .A2(n17), .ZN(n1074) );
  AOI22_X1 U1419 ( .A1(n29), .A2(regs[1432]), .B1(n12), .B2(regs[408]), .ZN(
        n1073) );
  AOI22_X1 U1420 ( .A1(n38), .A2(regs[2456]), .B1(n33), .B2(regs[1944]), .ZN(
        n1072) );
  NAND3_X1 U1421 ( .A1(n1074), .A2(n1073), .A3(n1072), .ZN(curr_proc_regs[408]) );
  NAND2_X1 U1422 ( .A1(regs[921]), .A2(n1579), .ZN(n1077) );
  AOI22_X1 U1423 ( .A1(n29), .A2(regs[1433]), .B1(n12), .B2(regs[409]), .ZN(
        n1076) );
  AOI22_X1 U1424 ( .A1(n38), .A2(regs[2457]), .B1(n31), .B2(regs[1945]), .ZN(
        n1075) );
  NAND3_X1 U1425 ( .A1(n1077), .A2(n1076), .A3(n1075), .ZN(curr_proc_regs[409]) );
  NAND2_X1 U1426 ( .A1(regs[552]), .A2(n7), .ZN(n1080) );
  AOI22_X1 U1427 ( .A1(n29), .A2(regs[1064]), .B1(n12), .B2(regs[40]), .ZN(
        n1079) );
  AOI22_X1 U1428 ( .A1(n38), .A2(regs[2088]), .B1(n9), .B2(regs[1576]), .ZN(
        n1078) );
  NAND3_X1 U1429 ( .A1(n1080), .A2(n1079), .A3(n1078), .ZN(curr_proc_regs[40])
         );
  NAND2_X1 U1430 ( .A1(regs[922]), .A2(n7), .ZN(n1083) );
  AOI22_X1 U1431 ( .A1(n29), .A2(regs[1434]), .B1(n12), .B2(regs[410]), .ZN(
        n1082) );
  AOI22_X1 U1432 ( .A1(n38), .A2(regs[2458]), .B1(n3), .B2(regs[1946]), .ZN(
        n1081) );
  NAND3_X1 U1433 ( .A1(n1083), .A2(n1082), .A3(n1081), .ZN(curr_proc_regs[410]) );
  NAND2_X1 U1434 ( .A1(regs[923]), .A2(n14), .ZN(n1086) );
  AOI22_X1 U1435 ( .A1(n29), .A2(regs[1435]), .B1(n12), .B2(regs[411]), .ZN(
        n1085) );
  AOI22_X1 U1436 ( .A1(n38), .A2(regs[2459]), .B1(n9), .B2(regs[1947]), .ZN(
        n1084) );
  NAND3_X1 U1437 ( .A1(n1086), .A2(n1085), .A3(n1084), .ZN(curr_proc_regs[411]) );
  NAND2_X1 U1438 ( .A1(regs[924]), .A2(n18), .ZN(n1089) );
  AOI22_X1 U1439 ( .A1(n29), .A2(regs[1436]), .B1(n12), .B2(regs[412]), .ZN(
        n1088) );
  AOI22_X1 U1440 ( .A1(n38), .A2(regs[2460]), .B1(n3), .B2(regs[1948]), .ZN(
        n1087) );
  NAND3_X1 U1441 ( .A1(n1089), .A2(n1088), .A3(n1087), .ZN(curr_proc_regs[412]) );
  NAND2_X1 U1442 ( .A1(regs[925]), .A2(n11), .ZN(n1092) );
  AOI22_X1 U1443 ( .A1(n29), .A2(regs[1437]), .B1(n12), .B2(regs[413]), .ZN(
        n1091) );
  AOI22_X1 U1444 ( .A1(n38), .A2(regs[2461]), .B1(n35), .B2(regs[1949]), .ZN(
        n1090) );
  NAND3_X1 U1445 ( .A1(n1092), .A2(n1091), .A3(n1090), .ZN(curr_proc_regs[413]) );
  NAND2_X1 U1446 ( .A1(regs[926]), .A2(n1579), .ZN(n1095) );
  AOI22_X1 U1447 ( .A1(n29), .A2(regs[1438]), .B1(n12), .B2(regs[414]), .ZN(
        n1094) );
  AOI22_X1 U1448 ( .A1(n38), .A2(regs[2462]), .B1(n33), .B2(regs[1950]), .ZN(
        n1093) );
  NAND3_X1 U1449 ( .A1(n1095), .A2(n1094), .A3(n1093), .ZN(curr_proc_regs[414]) );
  NAND2_X1 U1450 ( .A1(regs[927]), .A2(n16), .ZN(n1098) );
  AOI22_X1 U1451 ( .A1(n29), .A2(regs[1439]), .B1(n12), .B2(regs[415]), .ZN(
        n1097) );
  AOI22_X1 U1452 ( .A1(n38), .A2(regs[2463]), .B1(n3), .B2(regs[1951]), .ZN(
        n1096) );
  NAND3_X1 U1453 ( .A1(n1098), .A2(n1097), .A3(n1096), .ZN(curr_proc_regs[415]) );
  NAND2_X1 U1454 ( .A1(regs[928]), .A2(n7), .ZN(n1101) );
  AOI22_X1 U1455 ( .A1(n29), .A2(regs[1440]), .B1(n12), .B2(regs[416]), .ZN(
        n1100) );
  AOI22_X1 U1456 ( .A1(n8), .A2(regs[2464]), .B1(n34), .B2(regs[1952]), .ZN(
        n1099) );
  NAND3_X1 U1457 ( .A1(n1101), .A2(n1100), .A3(n1099), .ZN(curr_proc_regs[416]) );
  NAND2_X1 U1458 ( .A1(regs[929]), .A2(n7), .ZN(n1104) );
  AOI22_X1 U1459 ( .A1(n29), .A2(regs[1441]), .B1(n24), .B2(regs[417]), .ZN(
        n1103) );
  AOI22_X1 U1460 ( .A1(n8), .A2(regs[2465]), .B1(n35), .B2(regs[1953]), .ZN(
        n1102) );
  NAND3_X1 U1461 ( .A1(n1104), .A2(n1103), .A3(n1102), .ZN(curr_proc_regs[417]) );
  NAND2_X1 U1462 ( .A1(regs[930]), .A2(n7), .ZN(n1107) );
  AOI22_X1 U1463 ( .A1(n29), .A2(regs[1442]), .B1(n12), .B2(regs[418]), .ZN(
        n1106) );
  AOI22_X1 U1464 ( .A1(n8), .A2(regs[2466]), .B1(n35), .B2(regs[1954]), .ZN(
        n1105) );
  NAND3_X1 U1465 ( .A1(n1107), .A2(n1106), .A3(n1105), .ZN(curr_proc_regs[418]) );
  NAND2_X1 U1466 ( .A1(regs[931]), .A2(n7), .ZN(n1110) );
  AOI22_X1 U1467 ( .A1(n29), .A2(regs[1443]), .B1(n24), .B2(regs[419]), .ZN(
        n1109) );
  AOI22_X1 U1468 ( .A1(n8), .A2(regs[2467]), .B1(n3), .B2(regs[1955]), .ZN(
        n1108) );
  NAND3_X1 U1469 ( .A1(n1110), .A2(n1109), .A3(n1108), .ZN(curr_proc_regs[419]) );
  NAND2_X1 U1470 ( .A1(regs[553]), .A2(n7), .ZN(n1113) );
  AOI22_X1 U1471 ( .A1(n29), .A2(regs[1065]), .B1(n12), .B2(regs[41]), .ZN(
        n1112) );
  AOI22_X1 U1472 ( .A1(n8), .A2(regs[2089]), .B1(n3), .B2(regs[1577]), .ZN(
        n1111) );
  NAND3_X1 U1473 ( .A1(n1113), .A2(n1112), .A3(n1111), .ZN(curr_proc_regs[41])
         );
  NAND2_X1 U1474 ( .A1(regs[932]), .A2(n7), .ZN(n1116) );
  AOI22_X1 U1475 ( .A1(n29), .A2(regs[1444]), .B1(n1580), .B2(regs[420]), .ZN(
        n1115) );
  AOI22_X1 U1476 ( .A1(n8), .A2(regs[2468]), .B1(n35), .B2(regs[1956]), .ZN(
        n1114) );
  NAND3_X1 U1477 ( .A1(n1116), .A2(n1115), .A3(n1114), .ZN(curr_proc_regs[420]) );
  NAND2_X1 U1478 ( .A1(regs[933]), .A2(n7), .ZN(n1119) );
  AOI22_X1 U1479 ( .A1(n29), .A2(regs[1445]), .B1(n12), .B2(regs[421]), .ZN(
        n1118) );
  AOI22_X1 U1480 ( .A1(n8), .A2(regs[2469]), .B1(n35), .B2(regs[1957]), .ZN(
        n1117) );
  NAND3_X1 U1481 ( .A1(n1119), .A2(n1118), .A3(n1117), .ZN(curr_proc_regs[421]) );
  NAND2_X1 U1482 ( .A1(regs[934]), .A2(n7), .ZN(n1122) );
  AOI22_X1 U1483 ( .A1(n29), .A2(regs[1446]), .B1(n12), .B2(regs[422]), .ZN(
        n1121) );
  AOI22_X1 U1484 ( .A1(n8), .A2(regs[2470]), .B1(n9), .B2(regs[1958]), .ZN(
        n1120) );
  NAND3_X1 U1485 ( .A1(n1122), .A2(n1121), .A3(n1120), .ZN(curr_proc_regs[422]) );
  NAND2_X1 U1486 ( .A1(regs[935]), .A2(n7), .ZN(n1125) );
  AOI22_X1 U1487 ( .A1(n29), .A2(regs[1447]), .B1(n24), .B2(regs[423]), .ZN(
        n1124) );
  AOI22_X1 U1488 ( .A1(n8), .A2(regs[2471]), .B1(n9), .B2(regs[1959]), .ZN(
        n1123) );
  NAND3_X1 U1489 ( .A1(n1125), .A2(n1124), .A3(n1123), .ZN(curr_proc_regs[423]) );
  NAND2_X1 U1490 ( .A1(regs[936]), .A2(n7), .ZN(n1128) );
  AOI22_X1 U1491 ( .A1(n29), .A2(regs[1448]), .B1(n24), .B2(regs[424]), .ZN(
        n1127) );
  AOI22_X1 U1492 ( .A1(n8), .A2(regs[2472]), .B1(n34), .B2(regs[1960]), .ZN(
        n1126) );
  NAND3_X1 U1493 ( .A1(n1128), .A2(n1127), .A3(n1126), .ZN(curr_proc_regs[424]) );
  NAND2_X1 U1494 ( .A1(regs[937]), .A2(n7), .ZN(n1131) );
  AOI22_X1 U1495 ( .A1(n29), .A2(regs[1449]), .B1(n12), .B2(regs[425]), .ZN(
        n1130) );
  AOI22_X1 U1496 ( .A1(n8), .A2(regs[2473]), .B1(n9), .B2(regs[1961]), .ZN(
        n1129) );
  NAND3_X1 U1497 ( .A1(n1131), .A2(n1130), .A3(n1129), .ZN(curr_proc_regs[425]) );
  NAND2_X1 U1498 ( .A1(regs[938]), .A2(n7), .ZN(n1134) );
  AOI22_X1 U1499 ( .A1(n29), .A2(regs[1450]), .B1(n12), .B2(regs[426]), .ZN(
        n1133) );
  AOI22_X1 U1500 ( .A1(n10), .A2(regs[2474]), .B1(n35), .B2(regs[1962]), .ZN(
        n1132) );
  NAND3_X1 U1501 ( .A1(n1134), .A2(n1133), .A3(n1132), .ZN(curr_proc_regs[426]) );
  NAND2_X1 U1502 ( .A1(regs[939]), .A2(n13), .ZN(n1137) );
  AOI22_X1 U1503 ( .A1(n29), .A2(regs[1451]), .B1(n25), .B2(regs[427]), .ZN(
        n1136) );
  AOI22_X1 U1504 ( .A1(n10), .A2(regs[2475]), .B1(n3), .B2(regs[1963]), .ZN(
        n1135) );
  NAND3_X1 U1505 ( .A1(n1137), .A2(n1136), .A3(n1135), .ZN(curr_proc_regs[427]) );
  NAND2_X1 U1506 ( .A1(regs[940]), .A2(n13), .ZN(n1140) );
  AOI22_X1 U1507 ( .A1(n29), .A2(regs[1452]), .B1(n5), .B2(regs[428]), .ZN(
        n1139) );
  AOI22_X1 U1508 ( .A1(n10), .A2(regs[2476]), .B1(n9), .B2(regs[1964]), .ZN(
        n1138) );
  NAND3_X1 U1509 ( .A1(n1140), .A2(n1139), .A3(n1138), .ZN(curr_proc_regs[428]) );
  NAND2_X1 U1510 ( .A1(regs[941]), .A2(n13), .ZN(n1143) );
  AOI22_X1 U1511 ( .A1(n29), .A2(regs[1453]), .B1(n5), .B2(regs[429]), .ZN(
        n1142) );
  AOI22_X1 U1512 ( .A1(n10), .A2(regs[2477]), .B1(n3), .B2(regs[1965]), .ZN(
        n1141) );
  NAND3_X1 U1513 ( .A1(n1143), .A2(n1142), .A3(n1141), .ZN(curr_proc_regs[429]) );
  NAND2_X1 U1514 ( .A1(regs[554]), .A2(n13), .ZN(n1146) );
  AOI22_X1 U1515 ( .A1(n29), .A2(regs[1066]), .B1(n26), .B2(regs[42]), .ZN(
        n1145) );
  AOI22_X1 U1516 ( .A1(n10), .A2(regs[2090]), .B1(n35), .B2(regs[1578]), .ZN(
        n1144) );
  NAND3_X1 U1517 ( .A1(n1146), .A2(n1145), .A3(n1144), .ZN(curr_proc_regs[42])
         );
  NAND2_X1 U1518 ( .A1(regs[942]), .A2(n13), .ZN(n1149) );
  AOI22_X1 U1519 ( .A1(n29), .A2(regs[1454]), .B1(n1580), .B2(regs[430]), .ZN(
        n1148) );
  AOI22_X1 U1520 ( .A1(n10), .A2(regs[2478]), .B1(n33), .B2(regs[1966]), .ZN(
        n1147) );
  NAND3_X1 U1521 ( .A1(n1149), .A2(n1148), .A3(n1147), .ZN(curr_proc_regs[430]) );
  NAND2_X1 U1522 ( .A1(regs[943]), .A2(n13), .ZN(n1152) );
  AOI22_X1 U1523 ( .A1(n29), .A2(regs[1455]), .B1(n24), .B2(regs[431]), .ZN(
        n1151) );
  AOI22_X1 U1524 ( .A1(n10), .A2(regs[2479]), .B1(n31), .B2(regs[1967]), .ZN(
        n1150) );
  NAND3_X1 U1525 ( .A1(n1152), .A2(n1151), .A3(n1150), .ZN(curr_proc_regs[431]) );
  NAND2_X1 U1526 ( .A1(regs[944]), .A2(n13), .ZN(n1155) );
  AOI22_X1 U1527 ( .A1(n29), .A2(regs[1456]), .B1(n12), .B2(regs[432]), .ZN(
        n1154) );
  AOI22_X1 U1528 ( .A1(n10), .A2(regs[2480]), .B1(n34), .B2(regs[1968]), .ZN(
        n1153) );
  NAND3_X1 U1529 ( .A1(n1155), .A2(n1154), .A3(n1153), .ZN(curr_proc_regs[432]) );
  NAND2_X1 U1530 ( .A1(regs[945]), .A2(n13), .ZN(n1158) );
  AOI22_X1 U1531 ( .A1(n29), .A2(regs[1457]), .B1(n12), .B2(regs[433]), .ZN(
        n1157) );
  AOI22_X1 U1532 ( .A1(n10), .A2(regs[2481]), .B1(n3), .B2(regs[1969]), .ZN(
        n1156) );
  NAND3_X1 U1533 ( .A1(n1158), .A2(n1157), .A3(n1156), .ZN(curr_proc_regs[433]) );
  NAND2_X1 U1534 ( .A1(regs[946]), .A2(n13), .ZN(n1161) );
  AOI22_X1 U1535 ( .A1(n29), .A2(regs[1458]), .B1(n28), .B2(regs[434]), .ZN(
        n1160) );
  AOI22_X1 U1536 ( .A1(n10), .A2(regs[2482]), .B1(n2), .B2(regs[1970]), .ZN(
        n1159) );
  NAND3_X1 U1537 ( .A1(n1161), .A2(n1160), .A3(n1159), .ZN(curr_proc_regs[434]) );
  NAND2_X1 U1538 ( .A1(regs[947]), .A2(n13), .ZN(n1164) );
  AOI22_X1 U1539 ( .A1(n29), .A2(regs[1459]), .B1(n25), .B2(regs[435]), .ZN(
        n1163) );
  AOI22_X1 U1540 ( .A1(n10), .A2(regs[2483]), .B1(n3), .B2(regs[1971]), .ZN(
        n1162) );
  NAND3_X1 U1541 ( .A1(n1164), .A2(n1163), .A3(n1162), .ZN(curr_proc_regs[435]) );
  NAND2_X1 U1542 ( .A1(regs[948]), .A2(n13), .ZN(n1167) );
  AOI22_X1 U1543 ( .A1(n29), .A2(regs[1460]), .B1(n1580), .B2(regs[436]), .ZN(
        n1166) );
  AOI22_X1 U1544 ( .A1(n4), .A2(regs[2484]), .B1(n9), .B2(regs[1972]), .ZN(
        n1165) );
  NAND3_X1 U1545 ( .A1(n1167), .A2(n1166), .A3(n1165), .ZN(curr_proc_regs[436]) );
  NAND2_X1 U1546 ( .A1(regs[949]), .A2(n13), .ZN(n1170) );
  AOI22_X1 U1547 ( .A1(n29), .A2(regs[1461]), .B1(n5), .B2(regs[437]), .ZN(
        n1169) );
  AOI22_X1 U1548 ( .A1(n1), .A2(regs[2485]), .B1(n33), .B2(regs[1973]), .ZN(
        n1168) );
  NAND3_X1 U1549 ( .A1(n1170), .A2(n1169), .A3(n1168), .ZN(curr_proc_regs[437]) );
  NAND2_X1 U1550 ( .A1(regs[950]), .A2(n11), .ZN(n1173) );
  AOI22_X1 U1551 ( .A1(n29), .A2(regs[1462]), .B1(n1580), .B2(regs[438]), .ZN(
        n1172) );
  AOI22_X1 U1552 ( .A1(n37), .A2(regs[2486]), .B1(n30), .B2(regs[1974]), .ZN(
        n1171) );
  NAND3_X1 U1553 ( .A1(n1173), .A2(n1172), .A3(n1171), .ZN(curr_proc_regs[438]) );
  NAND2_X1 U1554 ( .A1(regs[951]), .A2(n13), .ZN(n1176) );
  AOI22_X1 U1555 ( .A1(n29), .A2(regs[1463]), .B1(n24), .B2(regs[439]), .ZN(
        n1175) );
  AOI22_X1 U1556 ( .A1(n41), .A2(regs[2487]), .B1(n9), .B2(regs[1975]), .ZN(
        n1174) );
  NAND3_X1 U1557 ( .A1(n1176), .A2(n1175), .A3(n1174), .ZN(curr_proc_regs[439]) );
  NAND2_X1 U1558 ( .A1(regs[555]), .A2(n14), .ZN(n1179) );
  AOI22_X1 U1559 ( .A1(n29), .A2(regs[1067]), .B1(n12), .B2(regs[43]), .ZN(
        n1178) );
  AOI22_X1 U1560 ( .A1(n39), .A2(regs[2091]), .B1(n30), .B2(regs[1579]), .ZN(
        n1177) );
  NAND3_X1 U1561 ( .A1(n1179), .A2(n1178), .A3(n1177), .ZN(curr_proc_regs[43])
         );
  NAND2_X1 U1562 ( .A1(regs[952]), .A2(n13), .ZN(n1182) );
  AOI22_X1 U1563 ( .A1(n29), .A2(regs[1464]), .B1(n24), .B2(regs[440]), .ZN(
        n1181) );
  AOI22_X1 U1564 ( .A1(n10), .A2(regs[2488]), .B1(n34), .B2(regs[1976]), .ZN(
        n1180) );
  NAND3_X1 U1565 ( .A1(n1182), .A2(n1181), .A3(n1180), .ZN(curr_proc_regs[440]) );
  NAND2_X1 U1566 ( .A1(regs[953]), .A2(n11), .ZN(n1185) );
  AOI22_X1 U1567 ( .A1(n29), .A2(regs[1465]), .B1(n12), .B2(regs[441]), .ZN(
        n1184) );
  AOI22_X1 U1568 ( .A1(n8), .A2(regs[2489]), .B1(n30), .B2(regs[1977]), .ZN(
        n1183) );
  NAND3_X1 U1569 ( .A1(n1185), .A2(n1184), .A3(n1183), .ZN(curr_proc_regs[441]) );
  NAND2_X1 U1570 ( .A1(regs[954]), .A2(n17), .ZN(n1188) );
  AOI22_X1 U1571 ( .A1(n29), .A2(regs[1466]), .B1(n28), .B2(regs[442]), .ZN(
        n1187) );
  AOI22_X1 U1572 ( .A1(n10), .A2(regs[2490]), .B1(n35), .B2(regs[1978]), .ZN(
        n1186) );
  NAND3_X1 U1573 ( .A1(n1188), .A2(n1187), .A3(n1186), .ZN(curr_proc_regs[442]) );
  NAND2_X1 U1574 ( .A1(regs[955]), .A2(n18), .ZN(n1191) );
  AOI22_X1 U1575 ( .A1(n29), .A2(regs[1467]), .B1(n12), .B2(regs[443]), .ZN(
        n1190) );
  AOI22_X1 U1576 ( .A1(n37), .A2(regs[2491]), .B1(n30), .B2(regs[1979]), .ZN(
        n1189) );
  NAND3_X1 U1577 ( .A1(n1191), .A2(n1190), .A3(n1189), .ZN(curr_proc_regs[443]) );
  NAND2_X1 U1578 ( .A1(regs[956]), .A2(n19), .ZN(n1194) );
  AOI22_X1 U1579 ( .A1(n29), .A2(regs[1468]), .B1(n24), .B2(regs[444]), .ZN(
        n1193) );
  AOI22_X1 U1580 ( .A1(n38), .A2(regs[2492]), .B1(n3), .B2(regs[1980]), .ZN(
        n1192) );
  NAND3_X1 U1581 ( .A1(n1194), .A2(n1193), .A3(n1192), .ZN(curr_proc_regs[444]) );
  NAND2_X1 U1582 ( .A1(regs[957]), .A2(n1579), .ZN(n1197) );
  AOI22_X1 U1583 ( .A1(n29), .A2(regs[1469]), .B1(n12), .B2(regs[445]), .ZN(
        n1196) );
  AOI22_X1 U1584 ( .A1(n41), .A2(regs[2493]), .B1(n30), .B2(regs[1981]), .ZN(
        n1195) );
  NAND3_X1 U1585 ( .A1(n1197), .A2(n1196), .A3(n1195), .ZN(curr_proc_regs[445]) );
  NAND2_X1 U1586 ( .A1(regs[958]), .A2(n11), .ZN(n1200) );
  AOI22_X1 U1587 ( .A1(n29), .A2(regs[1470]), .B1(n5), .B2(regs[446]), .ZN(
        n1199) );
  AOI22_X1 U1588 ( .A1(n41), .A2(regs[2494]), .B1(n30), .B2(regs[1982]), .ZN(
        n1198) );
  NAND3_X1 U1589 ( .A1(n1200), .A2(n1199), .A3(n1198), .ZN(curr_proc_regs[446]) );
  NAND2_X1 U1590 ( .A1(regs[959]), .A2(n20), .ZN(n1203) );
  AOI22_X1 U1591 ( .A1(n29), .A2(regs[1471]), .B1(n5), .B2(regs[447]), .ZN(
        n1202) );
  AOI22_X1 U1592 ( .A1(n41), .A2(regs[2495]), .B1(n9), .B2(regs[1983]), .ZN(
        n1201) );
  NAND3_X1 U1593 ( .A1(n1203), .A2(n1202), .A3(n1201), .ZN(curr_proc_regs[447]) );
  NAND2_X1 U1594 ( .A1(regs[960]), .A2(n14), .ZN(n1206) );
  AOI22_X1 U1595 ( .A1(n29), .A2(regs[1472]), .B1(n25), .B2(regs[448]), .ZN(
        n1205) );
  AOI22_X1 U1596 ( .A1(n41), .A2(regs[2496]), .B1(n9), .B2(regs[1984]), .ZN(
        n1204) );
  NAND3_X1 U1597 ( .A1(n1206), .A2(n1205), .A3(n1204), .ZN(curr_proc_regs[448]) );
  NAND2_X1 U1598 ( .A1(regs[961]), .A2(n20), .ZN(n1209) );
  AOI22_X1 U1599 ( .A1(n29), .A2(regs[1473]), .B1(n5), .B2(regs[449]), .ZN(
        n1208) );
  AOI22_X1 U1600 ( .A1(n41), .A2(regs[2497]), .B1(n35), .B2(regs[1985]), .ZN(
        n1207) );
  NAND3_X1 U1601 ( .A1(n1209), .A2(n1208), .A3(n1207), .ZN(curr_proc_regs[449]) );
  NAND2_X1 U1602 ( .A1(regs[556]), .A2(n14), .ZN(n1212) );
  AOI22_X1 U1603 ( .A1(n29), .A2(regs[1068]), .B1(n5), .B2(regs[44]), .ZN(
        n1211) );
  AOI22_X1 U1604 ( .A1(n10), .A2(regs[2092]), .B1(n9), .B2(regs[1580]), .ZN(
        n1210) );
  NAND3_X1 U1605 ( .A1(n1212), .A2(n1211), .A3(n1210), .ZN(curr_proc_regs[44])
         );
  NAND2_X1 U1606 ( .A1(regs[962]), .A2(n14), .ZN(n1215) );
  AOI22_X1 U1607 ( .A1(n29), .A2(regs[1474]), .B1(n12), .B2(regs[450]), .ZN(
        n1214) );
  AOI22_X1 U1608 ( .A1(n8), .A2(regs[2498]), .B1(n9), .B2(regs[1986]), .ZN(
        n1213) );
  NAND3_X1 U1609 ( .A1(n1215), .A2(n1214), .A3(n1213), .ZN(curr_proc_regs[450]) );
  NAND2_X1 U1610 ( .A1(regs[963]), .A2(n14), .ZN(n1218) );
  AOI22_X1 U1611 ( .A1(n29), .A2(regs[1475]), .B1(n12), .B2(regs[451]), .ZN(
        n1217) );
  AOI22_X1 U1612 ( .A1(n4), .A2(regs[2499]), .B1(n34), .B2(regs[1987]), .ZN(
        n1216) );
  NAND3_X1 U1613 ( .A1(n1218), .A2(n1217), .A3(n1216), .ZN(curr_proc_regs[451]) );
  NAND2_X1 U1614 ( .A1(regs[964]), .A2(n20), .ZN(n1221) );
  AOI22_X1 U1615 ( .A1(n29), .A2(regs[1476]), .B1(n1580), .B2(regs[452]), .ZN(
        n1220) );
  AOI22_X1 U1616 ( .A1(n8), .A2(regs[2500]), .B1(n3), .B2(regs[1988]), .ZN(
        n1219) );
  NAND3_X1 U1617 ( .A1(n1221), .A2(n1220), .A3(n1219), .ZN(curr_proc_regs[452]) );
  NAND2_X1 U1618 ( .A1(regs[965]), .A2(n20), .ZN(n1224) );
  AOI22_X1 U1619 ( .A1(n29), .A2(regs[1477]), .B1(n28), .B2(regs[453]), .ZN(
        n1223) );
  AOI22_X1 U1620 ( .A1(win[4]), .A2(regs[2501]), .B1(n3), .B2(regs[1989]), 
        .ZN(n1222) );
  NAND3_X1 U1621 ( .A1(n1224), .A2(n1223), .A3(n1222), .ZN(curr_proc_regs[453]) );
  NAND2_X1 U1622 ( .A1(regs[966]), .A2(n14), .ZN(n1227) );
  AOI22_X1 U1623 ( .A1(n29), .A2(regs[1478]), .B1(n25), .B2(regs[454]), .ZN(
        n1226) );
  AOI22_X1 U1624 ( .A1(n37), .A2(regs[2502]), .B1(n35), .B2(regs[1990]), .ZN(
        n1225) );
  NAND3_X1 U1625 ( .A1(n1227), .A2(n1226), .A3(n1225), .ZN(curr_proc_regs[454]) );
  NAND2_X1 U1626 ( .A1(regs[967]), .A2(n20), .ZN(n1230) );
  AOI22_X1 U1627 ( .A1(n29), .A2(regs[1479]), .B1(n5), .B2(regs[455]), .ZN(
        n1229) );
  AOI22_X1 U1628 ( .A1(n38), .A2(regs[2503]), .B1(n9), .B2(regs[1991]), .ZN(
        n1228) );
  NAND3_X1 U1629 ( .A1(n1230), .A2(n1229), .A3(n1228), .ZN(curr_proc_regs[455]) );
  NAND2_X1 U1630 ( .A1(regs[968]), .A2(n20), .ZN(n1233) );
  AOI22_X1 U1631 ( .A1(n29), .A2(regs[1480]), .B1(n5), .B2(regs[456]), .ZN(
        n1232) );
  AOI22_X1 U1632 ( .A1(n37), .A2(regs[2504]), .B1(n9), .B2(regs[1992]), .ZN(
        n1231) );
  NAND3_X1 U1633 ( .A1(n1233), .A2(n1232), .A3(n1231), .ZN(curr_proc_regs[456]) );
  NAND2_X1 U1634 ( .A1(regs[969]), .A2(n14), .ZN(n1236) );
  AOI22_X1 U1635 ( .A1(n29), .A2(regs[1481]), .B1(n5), .B2(regs[457]), .ZN(
        n1235) );
  AOI22_X1 U1636 ( .A1(win[4]), .A2(regs[2505]), .B1(n9), .B2(regs[1993]), 
        .ZN(n1234) );
  NAND3_X1 U1637 ( .A1(n1236), .A2(n1235), .A3(n1234), .ZN(curr_proc_regs[457]) );
  NAND2_X1 U1638 ( .A1(regs[970]), .A2(n14), .ZN(n1239) );
  AOI22_X1 U1639 ( .A1(n29), .A2(regs[1482]), .B1(n1580), .B2(regs[458]), .ZN(
        n1238) );
  AOI22_X1 U1640 ( .A1(n8), .A2(regs[2506]), .B1(n34), .B2(regs[1994]), .ZN(
        n1237) );
  NAND3_X1 U1641 ( .A1(n1239), .A2(n1238), .A3(n1237), .ZN(curr_proc_regs[458]) );
  NAND2_X1 U1642 ( .A1(regs[971]), .A2(n14), .ZN(n1242) );
  AOI22_X1 U1643 ( .A1(n29), .A2(regs[1483]), .B1(n12), .B2(regs[459]), .ZN(
        n1241) );
  AOI22_X1 U1644 ( .A1(n38), .A2(regs[2507]), .B1(n3), .B2(regs[1995]), .ZN(
        n1240) );
  NAND3_X1 U1645 ( .A1(n1242), .A2(n1241), .A3(n1240), .ZN(curr_proc_regs[459]) );
  NAND2_X1 U1646 ( .A1(regs[557]), .A2(n20), .ZN(n1245) );
  AOI22_X1 U1647 ( .A1(n29), .A2(regs[1069]), .B1(n12), .B2(regs[45]), .ZN(
        n1244) );
  AOI22_X1 U1648 ( .A1(n38), .A2(regs[2093]), .B1(n3), .B2(regs[1581]), .ZN(
        n1243) );
  NAND3_X1 U1649 ( .A1(n1245), .A2(n1244), .A3(n1243), .ZN(curr_proc_regs[45])
         );
  NAND2_X1 U1650 ( .A1(regs[972]), .A2(n14), .ZN(n1248) );
  AOI22_X1 U1651 ( .A1(n29), .A2(regs[1484]), .B1(n1580), .B2(regs[460]), .ZN(
        n1247) );
  AOI22_X1 U1652 ( .A1(n38), .A2(regs[2508]), .B1(n34), .B2(regs[1996]), .ZN(
        n1246) );
  NAND3_X1 U1653 ( .A1(n1248), .A2(n1247), .A3(n1246), .ZN(curr_proc_regs[460]) );
  NAND2_X1 U1654 ( .A1(regs[973]), .A2(n20), .ZN(n1251) );
  AOI22_X1 U1655 ( .A1(n29), .A2(regs[1485]), .B1(n24), .B2(regs[461]), .ZN(
        n1250) );
  AOI22_X1 U1656 ( .A1(n38), .A2(regs[2509]), .B1(n35), .B2(regs[1997]), .ZN(
        n1249) );
  NAND3_X1 U1657 ( .A1(n1251), .A2(n1250), .A3(n1249), .ZN(curr_proc_regs[461]) );
  NAND2_X1 U1658 ( .A1(regs[974]), .A2(n14), .ZN(n1254) );
  AOI22_X1 U1659 ( .A1(n29), .A2(regs[1486]), .B1(n12), .B2(regs[462]), .ZN(
        n1253) );
  AOI22_X1 U1660 ( .A1(n38), .A2(regs[2510]), .B1(n3), .B2(regs[1998]), .ZN(
        n1252) );
  NAND3_X1 U1661 ( .A1(n1254), .A2(n1253), .A3(n1252), .ZN(curr_proc_regs[462]) );
  NAND2_X1 U1662 ( .A1(regs[975]), .A2(n20), .ZN(n1257) );
  AOI22_X1 U1663 ( .A1(n29), .A2(regs[1487]), .B1(n12), .B2(regs[463]), .ZN(
        n1256) );
  AOI22_X1 U1664 ( .A1(n38), .A2(regs[2511]), .B1(n3), .B2(regs[1999]), .ZN(
        n1255) );
  NAND3_X1 U1665 ( .A1(n1257), .A2(n1256), .A3(n1255), .ZN(curr_proc_regs[463]) );
  NAND2_X1 U1666 ( .A1(regs[976]), .A2(n14), .ZN(n1260) );
  AOI22_X1 U1667 ( .A1(n29), .A2(regs[1488]), .B1(n5), .B2(regs[464]), .ZN(
        n1259) );
  AOI22_X1 U1668 ( .A1(n38), .A2(regs[2512]), .B1(n9), .B2(regs[2000]), .ZN(
        n1258) );
  NAND3_X1 U1669 ( .A1(n1260), .A2(n1259), .A3(n1258), .ZN(curr_proc_regs[464]) );
  NAND2_X1 U1670 ( .A1(regs[977]), .A2(n20), .ZN(n1263) );
  AOI22_X1 U1671 ( .A1(n29), .A2(regs[1489]), .B1(n24), .B2(regs[465]), .ZN(
        n1262) );
  AOI22_X1 U1672 ( .A1(n38), .A2(regs[2513]), .B1(n9), .B2(regs[2001]), .ZN(
        n1261) );
  NAND3_X1 U1673 ( .A1(n1263), .A2(n1262), .A3(n1261), .ZN(curr_proc_regs[465]) );
  NAND2_X1 U1674 ( .A1(regs[978]), .A2(n14), .ZN(n1266) );
  AOI22_X1 U1675 ( .A1(n29), .A2(regs[1490]), .B1(n12), .B2(regs[466]), .ZN(
        n1265) );
  AOI22_X1 U1676 ( .A1(n38), .A2(regs[2514]), .B1(n34), .B2(regs[2002]), .ZN(
        n1264) );
  NAND3_X1 U1677 ( .A1(n1266), .A2(n1265), .A3(n1264), .ZN(curr_proc_regs[466]) );
  NAND2_X1 U1678 ( .A1(regs[979]), .A2(n11), .ZN(n1269) );
  AOI22_X1 U1679 ( .A1(n29), .A2(regs[1491]), .B1(n28), .B2(regs[467]), .ZN(
        n1268) );
  AOI22_X1 U1680 ( .A1(n38), .A2(regs[2515]), .B1(n3), .B2(regs[2003]), .ZN(
        n1267) );
  NAND3_X1 U1681 ( .A1(n1269), .A2(n1268), .A3(n1267), .ZN(curr_proc_regs[467]) );
  NAND2_X1 U1682 ( .A1(regs[980]), .A2(n17), .ZN(n1272) );
  AOI22_X1 U1683 ( .A1(n29), .A2(regs[1492]), .B1(n26), .B2(regs[468]), .ZN(
        n1271) );
  AOI22_X1 U1684 ( .A1(n38), .A2(regs[2516]), .B1(n3), .B2(regs[2004]), .ZN(
        n1270) );
  NAND3_X1 U1685 ( .A1(n1272), .A2(n1271), .A3(n1270), .ZN(curr_proc_regs[468]) );
  NAND2_X1 U1686 ( .A1(regs[981]), .A2(n1579), .ZN(n1275) );
  AOI22_X1 U1687 ( .A1(n29), .A2(regs[1493]), .B1(n25), .B2(regs[469]), .ZN(
        n1274) );
  AOI22_X1 U1688 ( .A1(n4), .A2(regs[2517]), .B1(n35), .B2(regs[2005]), .ZN(
        n1273) );
  NAND3_X1 U1689 ( .A1(n1275), .A2(n1274), .A3(n1273), .ZN(curr_proc_regs[469]) );
  NAND2_X1 U1690 ( .A1(regs[558]), .A2(n1579), .ZN(n1278) );
  AOI22_X1 U1691 ( .A1(n29), .A2(regs[1070]), .B1(n5), .B2(regs[46]), .ZN(
        n1277) );
  AOI22_X1 U1692 ( .A1(n37), .A2(regs[2094]), .B1(n34), .B2(regs[1582]), .ZN(
        n1276) );
  NAND3_X1 U1693 ( .A1(n1278), .A2(n1277), .A3(n1276), .ZN(curr_proc_regs[46])
         );
  NAND2_X1 U1694 ( .A1(regs[982]), .A2(n7), .ZN(n1281) );
  AOI22_X1 U1695 ( .A1(n29), .A2(regs[1494]), .B1(n26), .B2(regs[470]), .ZN(
        n1280) );
  AOI22_X1 U1696 ( .A1(n39), .A2(regs[2518]), .B1(n9), .B2(regs[2006]), .ZN(
        n1279) );
  NAND3_X1 U1697 ( .A1(n1281), .A2(n1280), .A3(n1279), .ZN(curr_proc_regs[470]) );
  NAND2_X1 U1698 ( .A1(regs[983]), .A2(n11), .ZN(n1284) );
  AOI22_X1 U1699 ( .A1(n29), .A2(regs[1495]), .B1(n26), .B2(regs[471]), .ZN(
        n1283) );
  AOI22_X1 U1700 ( .A1(n8), .A2(regs[2519]), .B1(n9), .B2(regs[2007]), .ZN(
        n1282) );
  NAND3_X1 U1701 ( .A1(n1284), .A2(n1283), .A3(n1282), .ZN(curr_proc_regs[471]) );
  NAND2_X1 U1702 ( .A1(regs[984]), .A2(n1579), .ZN(n1287) );
  AOI22_X1 U1703 ( .A1(n29), .A2(regs[1496]), .B1(n5), .B2(regs[472]), .ZN(
        n1286) );
  AOI22_X1 U1704 ( .A1(n41), .A2(regs[2520]), .B1(n3), .B2(regs[2008]), .ZN(
        n1285) );
  NAND3_X1 U1705 ( .A1(n1287), .A2(n1286), .A3(n1285), .ZN(curr_proc_regs[472]) );
  NAND2_X1 U1706 ( .A1(regs[985]), .A2(n11), .ZN(n1290) );
  AOI22_X1 U1707 ( .A1(n29), .A2(regs[1497]), .B1(n1580), .B2(regs[473]), .ZN(
        n1289) );
  AOI22_X1 U1708 ( .A1(n1), .A2(regs[2521]), .B1(n3), .B2(regs[2009]), .ZN(
        n1288) );
  NAND3_X1 U1709 ( .A1(n1290), .A2(n1289), .A3(n1288), .ZN(curr_proc_regs[473]) );
  NAND2_X1 U1710 ( .A1(regs[986]), .A2(n7), .ZN(n1293) );
  AOI22_X1 U1711 ( .A1(n29), .A2(regs[1498]), .B1(n1580), .B2(regs[474]), .ZN(
        n1292) );
  AOI22_X1 U1712 ( .A1(n10), .A2(regs[2522]), .B1(n35), .B2(regs[2010]), .ZN(
        n1291) );
  NAND3_X1 U1713 ( .A1(n1293), .A2(n1292), .A3(n1291), .ZN(curr_proc_regs[474]) );
  NAND2_X1 U1714 ( .A1(regs[987]), .A2(n11), .ZN(n1296) );
  AOI22_X1 U1715 ( .A1(n29), .A2(regs[1499]), .B1(n1580), .B2(regs[475]), .ZN(
        n1295) );
  AOI22_X1 U1716 ( .A1(n4), .A2(regs[2523]), .B1(n34), .B2(regs[2011]), .ZN(
        n1294) );
  NAND3_X1 U1717 ( .A1(n1296), .A2(n1295), .A3(n1294), .ZN(curr_proc_regs[475]) );
  NAND2_X1 U1718 ( .A1(regs[988]), .A2(n1579), .ZN(n1299) );
  AOI22_X1 U1719 ( .A1(n29), .A2(regs[1500]), .B1(n1580), .B2(regs[476]), .ZN(
        n1298) );
  AOI22_X1 U1720 ( .A1(n37), .A2(regs[2524]), .B1(n9), .B2(regs[2012]), .ZN(
        n1297) );
  NAND3_X1 U1721 ( .A1(n1299), .A2(n1298), .A3(n1297), .ZN(curr_proc_regs[476]) );
  NAND2_X1 U1722 ( .A1(regs[989]), .A2(n19), .ZN(n1302) );
  AOI22_X1 U1723 ( .A1(n29), .A2(regs[1501]), .B1(n12), .B2(regs[477]), .ZN(
        n1301) );
  AOI22_X1 U1724 ( .A1(n39), .A2(regs[2525]), .B1(n3), .B2(regs[2013]), .ZN(
        n1300) );
  NAND3_X1 U1725 ( .A1(n1302), .A2(n1301), .A3(n1300), .ZN(curr_proc_regs[477]) );
  NAND2_X1 U1726 ( .A1(regs[990]), .A2(n7), .ZN(n1305) );
  AOI22_X1 U1727 ( .A1(n29), .A2(regs[1502]), .B1(n12), .B2(regs[478]), .ZN(
        n1304) );
  AOI22_X1 U1728 ( .A1(n8), .A2(regs[2526]), .B1(n33), .B2(regs[2014]), .ZN(
        n1303) );
  NAND3_X1 U1729 ( .A1(n1305), .A2(n1304), .A3(n1303), .ZN(curr_proc_regs[478]) );
  NAND2_X1 U1730 ( .A1(regs[991]), .A2(n19), .ZN(n1308) );
  AOI22_X1 U1731 ( .A1(n29), .A2(regs[1503]), .B1(n12), .B2(regs[479]), .ZN(
        n1307) );
  AOI22_X1 U1732 ( .A1(win[4]), .A2(regs[2527]), .B1(n34), .B2(regs[2015]), 
        .ZN(n1306) );
  NAND3_X1 U1733 ( .A1(n1308), .A2(n1307), .A3(n1306), .ZN(curr_proc_regs[479]) );
  NAND2_X1 U1734 ( .A1(regs[559]), .A2(n7), .ZN(n1311) );
  AOI22_X1 U1735 ( .A1(n29), .A2(regs[1071]), .B1(n12), .B2(regs[47]), .ZN(
        n1310) );
  AOI22_X1 U1736 ( .A1(win[4]), .A2(regs[2095]), .B1(n9), .B2(regs[1583]), 
        .ZN(n1309) );
  NAND3_X1 U1737 ( .A1(n1311), .A2(n1310), .A3(n1309), .ZN(curr_proc_regs[47])
         );
  NAND2_X1 U1738 ( .A1(regs[992]), .A2(n19), .ZN(n1314) );
  AOI22_X1 U1739 ( .A1(n29), .A2(regs[1504]), .B1(n12), .B2(regs[480]), .ZN(
        n1313) );
  AOI22_X1 U1740 ( .A1(win[4]), .A2(regs[2528]), .B1(n9), .B2(regs[2016]), 
        .ZN(n1312) );
  NAND3_X1 U1741 ( .A1(n1314), .A2(n1313), .A3(n1312), .ZN(curr_proc_regs[480]) );
  NAND2_X1 U1742 ( .A1(regs[993]), .A2(n7), .ZN(n1317) );
  AOI22_X1 U1743 ( .A1(n29), .A2(regs[1505]), .B1(n12), .B2(regs[481]), .ZN(
        n1316) );
  AOI22_X1 U1744 ( .A1(win[4]), .A2(regs[2529]), .B1(n35), .B2(regs[2017]), 
        .ZN(n1315) );
  NAND3_X1 U1745 ( .A1(n1317), .A2(n1316), .A3(n1315), .ZN(curr_proc_regs[481]) );
  NAND2_X1 U1746 ( .A1(regs[994]), .A2(n19), .ZN(n1320) );
  AOI22_X1 U1747 ( .A1(n29), .A2(regs[1506]), .B1(n12), .B2(regs[482]), .ZN(
        n1319) );
  AOI22_X1 U1748 ( .A1(win[4]), .A2(regs[2530]), .B1(n3), .B2(regs[2018]), 
        .ZN(n1318) );
  NAND3_X1 U1749 ( .A1(n1320), .A2(n1319), .A3(n1318), .ZN(curr_proc_regs[482]) );
  NAND2_X1 U1750 ( .A1(regs[995]), .A2(n7), .ZN(n1323) );
  AOI22_X1 U1751 ( .A1(n29), .A2(regs[1507]), .B1(n12), .B2(regs[483]), .ZN(
        n1322) );
  AOI22_X1 U1752 ( .A1(win[4]), .A2(regs[2531]), .B1(n3), .B2(regs[2019]), 
        .ZN(n1321) );
  NAND3_X1 U1753 ( .A1(n1323), .A2(n1322), .A3(n1321), .ZN(curr_proc_regs[483]) );
  NAND2_X1 U1754 ( .A1(regs[996]), .A2(n19), .ZN(n1326) );
  AOI22_X1 U1755 ( .A1(n29), .A2(regs[1508]), .B1(n12), .B2(regs[484]), .ZN(
        n1325) );
  AOI22_X1 U1756 ( .A1(win[4]), .A2(regs[2532]), .B1(n34), .B2(regs[2020]), 
        .ZN(n1324) );
  NAND3_X1 U1757 ( .A1(n1326), .A2(n1325), .A3(n1324), .ZN(curr_proc_regs[484]) );
  NAND2_X1 U1758 ( .A1(regs[997]), .A2(n7), .ZN(n1329) );
  AOI22_X1 U1759 ( .A1(n29), .A2(regs[1509]), .B1(n12), .B2(regs[485]), .ZN(
        n1328) );
  AOI22_X1 U1760 ( .A1(win[4]), .A2(regs[2533]), .B1(n2), .B2(regs[2021]), 
        .ZN(n1327) );
  NAND3_X1 U1761 ( .A1(n1329), .A2(n1328), .A3(n1327), .ZN(curr_proc_regs[485]) );
  NAND2_X1 U1762 ( .A1(regs[998]), .A2(n7), .ZN(n1332) );
  AOI22_X1 U1763 ( .A1(n29), .A2(regs[1510]), .B1(n12), .B2(regs[486]), .ZN(
        n1331) );
  AOI22_X1 U1764 ( .A1(win[4]), .A2(regs[2534]), .B1(n9), .B2(regs[2022]), 
        .ZN(n1330) );
  NAND3_X1 U1765 ( .A1(n1332), .A2(n1331), .A3(n1330), .ZN(curr_proc_regs[486]) );
  NAND2_X1 U1766 ( .A1(regs[999]), .A2(n14), .ZN(n1335) );
  AOI22_X1 U1767 ( .A1(n29), .A2(regs[1511]), .B1(n12), .B2(regs[487]), .ZN(
        n1334) );
  AOI22_X1 U1768 ( .A1(win[4]), .A2(regs[2535]), .B1(n34), .B2(regs[2023]), 
        .ZN(n1333) );
  NAND3_X1 U1769 ( .A1(n1335), .A2(n1334), .A3(n1333), .ZN(curr_proc_regs[487]) );
  NAND2_X1 U1770 ( .A1(regs[1000]), .A2(n14), .ZN(n1338) );
  AOI22_X1 U1771 ( .A1(n29), .A2(regs[1512]), .B1(n5), .B2(regs[488]), .ZN(
        n1337) );
  AOI22_X1 U1772 ( .A1(win[4]), .A2(regs[2536]), .B1(n35), .B2(regs[2024]), 
        .ZN(n1336) );
  NAND3_X1 U1773 ( .A1(n1338), .A2(n1337), .A3(n1336), .ZN(curr_proc_regs[488]) );
  NAND2_X1 U1774 ( .A1(regs[1001]), .A2(n14), .ZN(n1341) );
  AOI22_X1 U1775 ( .A1(n29), .A2(regs[1513]), .B1(n26), .B2(regs[489]), .ZN(
        n1340) );
  AOI22_X1 U1776 ( .A1(n4), .A2(regs[2537]), .B1(n3), .B2(regs[2025]), .ZN(
        n1339) );
  NAND3_X1 U1777 ( .A1(n1341), .A2(n1340), .A3(n1339), .ZN(curr_proc_regs[489]) );
  NAND2_X1 U1778 ( .A1(regs[560]), .A2(n14), .ZN(n1344) );
  AOI22_X1 U1779 ( .A1(n29), .A2(regs[1072]), .B1(n25), .B2(regs[48]), .ZN(
        n1343) );
  AOI22_X1 U1780 ( .A1(n4), .A2(regs[2096]), .B1(n35), .B2(regs[1584]), .ZN(
        n1342) );
  NAND3_X1 U1781 ( .A1(n1344), .A2(n1343), .A3(n1342), .ZN(curr_proc_regs[48])
         );
  NAND2_X1 U1782 ( .A1(regs[1002]), .A2(n14), .ZN(n1347) );
  AOI22_X1 U1783 ( .A1(n29), .A2(regs[1514]), .B1(n5), .B2(regs[490]), .ZN(
        n1346) );
  AOI22_X1 U1784 ( .A1(n4), .A2(regs[2538]), .B1(n3), .B2(regs[2026]), .ZN(
        n1345) );
  NAND3_X1 U1785 ( .A1(n1347), .A2(n1346), .A3(n1345), .ZN(curr_proc_regs[490]) );
  NAND2_X1 U1786 ( .A1(regs[1003]), .A2(n14), .ZN(n1350) );
  AOI22_X1 U1787 ( .A1(n29), .A2(regs[1515]), .B1(n1580), .B2(regs[491]), .ZN(
        n1349) );
  AOI22_X1 U1788 ( .A1(n4), .A2(regs[2539]), .B1(n35), .B2(regs[2027]), .ZN(
        n1348) );
  NAND3_X1 U1789 ( .A1(n1350), .A2(n1349), .A3(n1348), .ZN(curr_proc_regs[491]) );
  NAND2_X1 U1790 ( .A1(regs[1004]), .A2(n14), .ZN(n1353) );
  AOI22_X1 U1791 ( .A1(n29), .A2(regs[1516]), .B1(n5), .B2(regs[492]), .ZN(
        n1352) );
  AOI22_X1 U1792 ( .A1(n4), .A2(regs[2540]), .B1(n35), .B2(regs[2028]), .ZN(
        n1351) );
  NAND3_X1 U1793 ( .A1(n1353), .A2(n1352), .A3(n1351), .ZN(curr_proc_regs[492]) );
  NAND2_X1 U1794 ( .A1(regs[1005]), .A2(n14), .ZN(n1356) );
  AOI22_X1 U1795 ( .A1(n29), .A2(regs[1517]), .B1(n1580), .B2(regs[493]), .ZN(
        n1355) );
  AOI22_X1 U1796 ( .A1(n4), .A2(regs[2541]), .B1(n35), .B2(regs[2029]), .ZN(
        n1354) );
  NAND3_X1 U1797 ( .A1(n1356), .A2(n1355), .A3(n1354), .ZN(curr_proc_regs[493]) );
  NAND2_X1 U1798 ( .A1(regs[1006]), .A2(n14), .ZN(n1359) );
  AOI22_X1 U1799 ( .A1(n29), .A2(regs[1518]), .B1(n5), .B2(regs[494]), .ZN(
        n1358) );
  AOI22_X1 U1800 ( .A1(n4), .A2(regs[2542]), .B1(n9), .B2(regs[2030]), .ZN(
        n1357) );
  NAND3_X1 U1801 ( .A1(n1359), .A2(n1358), .A3(n1357), .ZN(curr_proc_regs[494]) );
  NAND2_X1 U1802 ( .A1(regs[1007]), .A2(n14), .ZN(n1362) );
  AOI22_X1 U1803 ( .A1(n29), .A2(regs[1519]), .B1(n1580), .B2(regs[495]), .ZN(
        n1361) );
  AOI22_X1 U1804 ( .A1(n4), .A2(regs[2543]), .B1(n35), .B2(regs[2031]), .ZN(
        n1360) );
  NAND3_X1 U1805 ( .A1(n1362), .A2(n1361), .A3(n1360), .ZN(curr_proc_regs[495]) );
  NAND2_X1 U1806 ( .A1(regs[1008]), .A2(n14), .ZN(n1365) );
  AOI22_X1 U1807 ( .A1(n29), .A2(regs[1520]), .B1(n1580), .B2(regs[496]), .ZN(
        n1364) );
  AOI22_X1 U1808 ( .A1(n4), .A2(regs[2544]), .B1(n35), .B2(regs[2032]), .ZN(
        n1363) );
  NAND3_X1 U1809 ( .A1(n1365), .A2(n1364), .A3(n1363), .ZN(curr_proc_regs[496]) );
  NAND2_X1 U1810 ( .A1(regs[1009]), .A2(n16), .ZN(n1368) );
  AOI22_X1 U1811 ( .A1(n29), .A2(regs[1521]), .B1(n24), .B2(regs[497]), .ZN(
        n1367) );
  AOI22_X1 U1812 ( .A1(n4), .A2(regs[2545]), .B1(n2), .B2(regs[2033]), .ZN(
        n1366) );
  NAND3_X1 U1813 ( .A1(n1368), .A2(n1367), .A3(n1366), .ZN(curr_proc_regs[497]) );
  NAND2_X1 U1814 ( .A1(regs[1010]), .A2(n7), .ZN(n1371) );
  AOI22_X1 U1815 ( .A1(n29), .A2(regs[1522]), .B1(n24), .B2(regs[498]), .ZN(
        n1370) );
  AOI22_X1 U1816 ( .A1(n4), .A2(regs[2546]), .B1(n34), .B2(regs[2034]), .ZN(
        n1369) );
  NAND3_X1 U1817 ( .A1(n1371), .A2(n1370), .A3(n1369), .ZN(curr_proc_regs[498]) );
  NAND2_X1 U1818 ( .A1(regs[1011]), .A2(n1579), .ZN(n1374) );
  AOI22_X1 U1819 ( .A1(n29), .A2(regs[1523]), .B1(n24), .B2(regs[499]), .ZN(
        n1373) );
  AOI22_X1 U1820 ( .A1(n8), .A2(regs[2547]), .B1(n2), .B2(regs[2035]), .ZN(
        n1372) );
  NAND3_X1 U1821 ( .A1(n1374), .A2(n1373), .A3(n1372), .ZN(curr_proc_regs[499]) );
  NAND2_X1 U1822 ( .A1(regs[561]), .A2(n18), .ZN(n1377) );
  AOI22_X1 U1823 ( .A1(n29), .A2(regs[1073]), .B1(n24), .B2(regs[49]), .ZN(
        n1376) );
  AOI22_X1 U1824 ( .A1(n8), .A2(regs[2097]), .B1(n9), .B2(regs[1585]), .ZN(
        n1375) );
  NAND3_X1 U1825 ( .A1(n1377), .A2(n1376), .A3(n1375), .ZN(curr_proc_regs[49])
         );
  NAND2_X1 U1826 ( .A1(regs[516]), .A2(n16), .ZN(n1380) );
  AOI22_X1 U1827 ( .A1(n29), .A2(regs[1028]), .B1(n24), .B2(regs[4]), .ZN(
        n1379) );
  AOI22_X1 U1828 ( .A1(n8), .A2(regs[2052]), .B1(n2), .B2(regs[1540]), .ZN(
        n1378) );
  NAND3_X1 U1829 ( .A1(n1380), .A2(n1379), .A3(n1378), .ZN(curr_proc_regs[4])
         );
  NAND2_X1 U1830 ( .A1(regs[1012]), .A2(n11), .ZN(n1383) );
  AOI22_X1 U1831 ( .A1(n29), .A2(regs[1524]), .B1(n24), .B2(regs[500]), .ZN(
        n1382) );
  AOI22_X1 U1832 ( .A1(n8), .A2(regs[2548]), .B1(n9), .B2(regs[2036]), .ZN(
        n1381) );
  NAND3_X1 U1833 ( .A1(n1383), .A2(n1382), .A3(n1381), .ZN(curr_proc_regs[500]) );
  NAND2_X1 U1834 ( .A1(regs[1013]), .A2(n15), .ZN(n1386) );
  AOI22_X1 U1835 ( .A1(n29), .A2(regs[1525]), .B1(n24), .B2(regs[501]), .ZN(
        n1385) );
  AOI22_X1 U1836 ( .A1(n8), .A2(regs[2549]), .B1(n2), .B2(regs[2037]), .ZN(
        n1384) );
  NAND3_X1 U1837 ( .A1(n1386), .A2(n1385), .A3(n1384), .ZN(curr_proc_regs[501]) );
  NAND2_X1 U1838 ( .A1(regs[1014]), .A2(n16), .ZN(n1389) );
  AOI22_X1 U1839 ( .A1(n29), .A2(regs[1526]), .B1(n24), .B2(regs[502]), .ZN(
        n1388) );
  AOI22_X1 U1840 ( .A1(n8), .A2(regs[2550]), .B1(n35), .B2(regs[2038]), .ZN(
        n1387) );
  NAND3_X1 U1841 ( .A1(n1389), .A2(n1388), .A3(n1387), .ZN(curr_proc_regs[502]) );
  NAND2_X1 U1842 ( .A1(regs[1015]), .A2(n1579), .ZN(n1392) );
  AOI22_X1 U1843 ( .A1(n29), .A2(regs[1527]), .B1(n24), .B2(regs[503]), .ZN(
        n1391) );
  AOI22_X1 U1844 ( .A1(n8), .A2(regs[2551]), .B1(n2), .B2(regs[2039]), .ZN(
        n1390) );
  NAND3_X1 U1845 ( .A1(n1392), .A2(n1391), .A3(n1390), .ZN(curr_proc_regs[503]) );
  NAND2_X1 U1846 ( .A1(regs[1016]), .A2(n16), .ZN(n1395) );
  AOI22_X1 U1847 ( .A1(n29), .A2(regs[1528]), .B1(n24), .B2(regs[504]), .ZN(
        n1394) );
  AOI22_X1 U1848 ( .A1(n8), .A2(regs[2552]), .B1(n3), .B2(regs[2040]), .ZN(
        n1393) );
  NAND3_X1 U1849 ( .A1(n1395), .A2(n1394), .A3(n1393), .ZN(curr_proc_regs[504]) );
  NAND2_X1 U1850 ( .A1(regs[1017]), .A2(n16), .ZN(n1398) );
  AOI22_X1 U1851 ( .A1(n29), .A2(regs[1529]), .B1(n24), .B2(regs[505]), .ZN(
        n1397) );
  AOI22_X1 U1852 ( .A1(n8), .A2(regs[2553]), .B1(n2), .B2(regs[2041]), .ZN(
        n1396) );
  NAND3_X1 U1853 ( .A1(n1398), .A2(n1397), .A3(n1396), .ZN(curr_proc_regs[505]) );
  NAND2_X1 U1854 ( .A1(regs[1018]), .A2(n1579), .ZN(n1401) );
  AOI22_X1 U1855 ( .A1(n29), .A2(regs[1530]), .B1(n24), .B2(regs[506]), .ZN(
        n1400) );
  AOI22_X1 U1856 ( .A1(n8), .A2(regs[2554]), .B1(n34), .B2(regs[2042]), .ZN(
        n1399) );
  NAND3_X1 U1857 ( .A1(n1401), .A2(n1400), .A3(n1399), .ZN(curr_proc_regs[506]) );
  NAND2_X1 U1858 ( .A1(regs[1019]), .A2(n1579), .ZN(n1404) );
  AOI22_X1 U1859 ( .A1(n29), .A2(regs[1531]), .B1(n12), .B2(regs[507]), .ZN(
        n1403) );
  AOI22_X1 U1860 ( .A1(n10), .A2(regs[2555]), .B1(n35), .B2(regs[2043]), .ZN(
        n1402) );
  NAND3_X1 U1861 ( .A1(n1404), .A2(n1403), .A3(n1402), .ZN(curr_proc_regs[507]) );
  NAND2_X1 U1862 ( .A1(regs[1020]), .A2(n1579), .ZN(n1407) );
  AOI22_X1 U1863 ( .A1(n29), .A2(regs[1532]), .B1(n24), .B2(regs[508]), .ZN(
        n1406) );
  AOI22_X1 U1864 ( .A1(win[4]), .A2(regs[2556]), .B1(n9), .B2(regs[2044]), 
        .ZN(n1405) );
  NAND3_X1 U1865 ( .A1(n1407), .A2(n1406), .A3(n1405), .ZN(curr_proc_regs[508]) );
  NAND2_X1 U1866 ( .A1(regs[1021]), .A2(n1579), .ZN(n1410) );
  AOI22_X1 U1867 ( .A1(n29), .A2(regs[1533]), .B1(n12), .B2(regs[509]), .ZN(
        n1409) );
  AOI22_X1 U1868 ( .A1(win[4]), .A2(regs[2557]), .B1(n3), .B2(regs[2045]), 
        .ZN(n1408) );
  NAND3_X1 U1869 ( .A1(n1410), .A2(n1409), .A3(n1408), .ZN(curr_proc_regs[509]) );
  NAND2_X1 U1870 ( .A1(regs[562]), .A2(n1579), .ZN(n1413) );
  AOI22_X1 U1871 ( .A1(n29), .A2(regs[1074]), .B1(n24), .B2(regs[50]), .ZN(
        n1412) );
  AOI22_X1 U1872 ( .A1(n38), .A2(regs[2098]), .B1(n9), .B2(regs[1586]), .ZN(
        n1411) );
  NAND3_X1 U1873 ( .A1(n1413), .A2(n1412), .A3(n1411), .ZN(curr_proc_regs[50])
         );
  NAND2_X1 U1874 ( .A1(regs[1022]), .A2(n1579), .ZN(n1416) );
  AOI22_X1 U1875 ( .A1(n29), .A2(regs[1534]), .B1(n12), .B2(regs[510]), .ZN(
        n1415) );
  AOI22_X1 U1876 ( .A1(win[4]), .A2(regs[2558]), .B1(n3), .B2(regs[2046]), 
        .ZN(n1414) );
  NAND3_X1 U1877 ( .A1(n1416), .A2(n1415), .A3(n1414), .ZN(curr_proc_regs[510]) );
  NAND2_X1 U1878 ( .A1(regs[1023]), .A2(n1579), .ZN(n1419) );
  AOI22_X1 U1879 ( .A1(n29), .A2(regs[1535]), .B1(n24), .B2(regs[511]), .ZN(
        n1418) );
  AOI22_X1 U1880 ( .A1(n41), .A2(regs[2559]), .B1(n35), .B2(regs[2047]), .ZN(
        n1417) );
  NAND3_X1 U1881 ( .A1(n1419), .A2(n1418), .A3(n1417), .ZN(curr_proc_regs[511]) );
  NAND2_X1 U1882 ( .A1(regs[563]), .A2(n1579), .ZN(n1422) );
  AOI22_X1 U1883 ( .A1(n29), .A2(regs[1075]), .B1(n12), .B2(regs[51]), .ZN(
        n1421) );
  AOI22_X1 U1884 ( .A1(win[4]), .A2(regs[2099]), .B1(n9), .B2(regs[1587]), 
        .ZN(n1420) );
  NAND3_X1 U1885 ( .A1(n1422), .A2(n1421), .A3(n1420), .ZN(curr_proc_regs[51])
         );
  NAND2_X1 U1886 ( .A1(regs[564]), .A2(n1579), .ZN(n1425) );
  AOI22_X1 U1887 ( .A1(n29), .A2(regs[1076]), .B1(n24), .B2(regs[52]), .ZN(
        n1424) );
  AOI22_X1 U1888 ( .A1(n37), .A2(regs[2100]), .B1(n3), .B2(regs[1588]), .ZN(
        n1423) );
  NAND3_X1 U1889 ( .A1(n1425), .A2(n1424), .A3(n1423), .ZN(curr_proc_regs[52])
         );
  NAND2_X1 U1890 ( .A1(regs[565]), .A2(n1579), .ZN(n1428) );
  AOI22_X1 U1891 ( .A1(n29), .A2(regs[1077]), .B1(n12), .B2(regs[53]), .ZN(
        n1427) );
  AOI22_X1 U1892 ( .A1(win[4]), .A2(regs[2101]), .B1(n35), .B2(regs[1589]), 
        .ZN(n1426) );
  NAND3_X1 U1893 ( .A1(n1428), .A2(n1427), .A3(n1426), .ZN(curr_proc_regs[53])
         );
  NAND2_X1 U1894 ( .A1(regs[566]), .A2(n1579), .ZN(n1431) );
  AOI22_X1 U1895 ( .A1(n29), .A2(regs[1078]), .B1(n24), .B2(regs[54]), .ZN(
        n1430) );
  AOI22_X1 U1896 ( .A1(n1), .A2(regs[2102]), .B1(n3), .B2(regs[1590]), .ZN(
        n1429) );
  NAND3_X1 U1897 ( .A1(n1431), .A2(n1430), .A3(n1429), .ZN(curr_proc_regs[54])
         );
  NAND2_X1 U1898 ( .A1(regs[567]), .A2(n18), .ZN(n1434) );
  AOI22_X1 U1899 ( .A1(n29), .A2(regs[1079]), .B1(n25), .B2(regs[55]), .ZN(
        n1433) );
  AOI22_X1 U1900 ( .A1(win[4]), .A2(regs[2103]), .B1(n9), .B2(regs[1591]), 
        .ZN(n1432) );
  NAND3_X1 U1901 ( .A1(n1434), .A2(n1433), .A3(n1432), .ZN(curr_proc_regs[55])
         );
  NAND2_X1 U1902 ( .A1(regs[568]), .A2(n11), .ZN(n1437) );
  AOI22_X1 U1903 ( .A1(n29), .A2(regs[1080]), .B1(n25), .B2(regs[56]), .ZN(
        n1436) );
  AOI22_X1 U1904 ( .A1(n37), .A2(regs[2104]), .B1(n35), .B2(regs[1592]), .ZN(
        n1435) );
  NAND3_X1 U1905 ( .A1(n1437), .A2(n1436), .A3(n1435), .ZN(curr_proc_regs[56])
         );
  NAND2_X1 U1906 ( .A1(regs[569]), .A2(n14), .ZN(n1440) );
  AOI22_X1 U1907 ( .A1(n29), .A2(regs[1081]), .B1(n25), .B2(regs[57]), .ZN(
        n1439) );
  AOI22_X1 U1908 ( .A1(n37), .A2(regs[2105]), .B1(n9), .B2(regs[1593]), .ZN(
        n1438) );
  NAND3_X1 U1909 ( .A1(n1440), .A2(n1439), .A3(n1438), .ZN(curr_proc_regs[57])
         );
  NAND2_X1 U1910 ( .A1(regs[570]), .A2(n11), .ZN(n1443) );
  AOI22_X1 U1911 ( .A1(n29), .A2(regs[1082]), .B1(n25), .B2(regs[58]), .ZN(
        n1442) );
  AOI22_X1 U1912 ( .A1(n37), .A2(regs[2106]), .B1(n9), .B2(regs[1594]), .ZN(
        n1441) );
  NAND3_X1 U1913 ( .A1(n1443), .A2(n1442), .A3(n1441), .ZN(curr_proc_regs[58])
         );
  NAND2_X1 U1914 ( .A1(regs[571]), .A2(n7), .ZN(n1446) );
  AOI22_X1 U1915 ( .A1(n29), .A2(regs[1083]), .B1(n25), .B2(regs[59]), .ZN(
        n1445) );
  AOI22_X1 U1916 ( .A1(n37), .A2(regs[2107]), .B1(n3), .B2(regs[1595]), .ZN(
        n1444) );
  NAND3_X1 U1917 ( .A1(n1446), .A2(n1445), .A3(n1444), .ZN(curr_proc_regs[59])
         );
  NAND2_X1 U1918 ( .A1(regs[517]), .A2(n17), .ZN(n1449) );
  AOI22_X1 U1919 ( .A1(n29), .A2(regs[1029]), .B1(n25), .B2(regs[5]), .ZN(
        n1448) );
  AOI22_X1 U1920 ( .A1(n37), .A2(regs[2053]), .B1(n3), .B2(regs[1541]), .ZN(
        n1447) );
  NAND3_X1 U1921 ( .A1(n1449), .A2(n1448), .A3(n1447), .ZN(curr_proc_regs[5])
         );
  NAND2_X1 U1922 ( .A1(regs[572]), .A2(n16), .ZN(n1452) );
  AOI22_X1 U1923 ( .A1(n29), .A2(regs[1084]), .B1(n25), .B2(regs[60]), .ZN(
        n1451) );
  AOI22_X1 U1924 ( .A1(n37), .A2(regs[2108]), .B1(n35), .B2(regs[1596]), .ZN(
        n1450) );
  NAND3_X1 U1925 ( .A1(n1452), .A2(n1451), .A3(n1450), .ZN(curr_proc_regs[60])
         );
  NAND2_X1 U1926 ( .A1(regs[573]), .A2(n13), .ZN(n1455) );
  AOI22_X1 U1927 ( .A1(n29), .A2(regs[1085]), .B1(n25), .B2(regs[61]), .ZN(
        n1454) );
  AOI22_X1 U1928 ( .A1(n37), .A2(regs[2109]), .B1(n34), .B2(regs[1597]), .ZN(
        n1453) );
  NAND3_X1 U1929 ( .A1(n1455), .A2(n1454), .A3(n1453), .ZN(curr_proc_regs[61])
         );
  NAND2_X1 U1930 ( .A1(regs[574]), .A2(n11), .ZN(n1458) );
  AOI22_X1 U1931 ( .A1(n29), .A2(regs[1086]), .B1(n25), .B2(regs[62]), .ZN(
        n1457) );
  AOI22_X1 U1932 ( .A1(n37), .A2(regs[2110]), .B1(n3), .B2(regs[1598]), .ZN(
        n1456) );
  NAND3_X1 U1933 ( .A1(n1458), .A2(n1457), .A3(n1456), .ZN(curr_proc_regs[62])
         );
  NAND2_X1 U1934 ( .A1(regs[575]), .A2(n11), .ZN(n1461) );
  AOI22_X1 U1935 ( .A1(n29), .A2(regs[1087]), .B1(n25), .B2(regs[63]), .ZN(
        n1460) );
  AOI22_X1 U1936 ( .A1(n37), .A2(regs[2111]), .B1(n3), .B2(regs[1599]), .ZN(
        n1459) );
  NAND3_X1 U1937 ( .A1(n1461), .A2(n1460), .A3(n1459), .ZN(curr_proc_regs[63])
         );
  NAND2_X1 U1938 ( .A1(regs[576]), .A2(n13), .ZN(n1464) );
  AOI22_X1 U1939 ( .A1(n29), .A2(regs[1088]), .B1(n25), .B2(regs[64]), .ZN(
        n1463) );
  AOI22_X1 U1940 ( .A1(n37), .A2(regs[2112]), .B1(n34), .B2(regs[1600]), .ZN(
        n1462) );
  NAND3_X1 U1941 ( .A1(n1464), .A2(n1463), .A3(n1462), .ZN(curr_proc_regs[64])
         );
  NAND2_X1 U1942 ( .A1(regs[577]), .A2(n14), .ZN(n1467) );
  AOI22_X1 U1943 ( .A1(n29), .A2(regs[1089]), .B1(n5), .B2(regs[65]), .ZN(
        n1466) );
  AOI22_X1 U1944 ( .A1(n37), .A2(regs[2113]), .B1(n35), .B2(regs[1601]), .ZN(
        n1465) );
  NAND3_X1 U1945 ( .A1(n1467), .A2(n1466), .A3(n1465), .ZN(curr_proc_regs[65])
         );
  NAND2_X1 U1946 ( .A1(regs[578]), .A2(n1579), .ZN(n1470) );
  AOI22_X1 U1947 ( .A1(n29), .A2(regs[1090]), .B1(n5), .B2(regs[66]), .ZN(
        n1469) );
  AOI22_X1 U1948 ( .A1(n36), .A2(regs[2114]), .B1(n35), .B2(regs[1602]), .ZN(
        n1468) );
  NAND3_X1 U1949 ( .A1(n1470), .A2(n1469), .A3(n1468), .ZN(curr_proc_regs[66])
         );
  NAND2_X1 U1950 ( .A1(regs[579]), .A2(n13), .ZN(n1473) );
  AOI22_X1 U1951 ( .A1(n29), .A2(regs[1091]), .B1(n5), .B2(regs[67]), .ZN(
        n1472) );
  AOI22_X1 U1952 ( .A1(n36), .A2(regs[2115]), .B1(n3), .B2(regs[1603]), .ZN(
        n1471) );
  NAND3_X1 U1953 ( .A1(n1473), .A2(n1472), .A3(n1471), .ZN(curr_proc_regs[67])
         );
  NAND2_X1 U1954 ( .A1(regs[580]), .A2(n1579), .ZN(n1476) );
  AOI22_X1 U1955 ( .A1(n29), .A2(regs[1092]), .B1(n5), .B2(regs[68]), .ZN(
        n1475) );
  AOI22_X1 U1956 ( .A1(n36), .A2(regs[2116]), .B1(n3), .B2(regs[1604]), .ZN(
        n1474) );
  NAND3_X1 U1957 ( .A1(n1476), .A2(n1475), .A3(n1474), .ZN(curr_proc_regs[68])
         );
  NAND2_X1 U1958 ( .A1(regs[581]), .A2(n19), .ZN(n1479) );
  AOI22_X1 U1959 ( .A1(n29), .A2(regs[1093]), .B1(n5), .B2(regs[69]), .ZN(
        n1478) );
  AOI22_X1 U1960 ( .A1(n36), .A2(regs[2117]), .B1(n9), .B2(regs[1605]), .ZN(
        n1477) );
  NAND3_X1 U1961 ( .A1(n1479), .A2(n1478), .A3(n1477), .ZN(curr_proc_regs[69])
         );
  NAND2_X1 U1962 ( .A1(regs[518]), .A2(n1579), .ZN(n1482) );
  AOI22_X1 U1963 ( .A1(n29), .A2(regs[1030]), .B1(n5), .B2(regs[6]), .ZN(n1481) );
  AOI22_X1 U1964 ( .A1(n36), .A2(regs[2054]), .B1(n9), .B2(regs[1542]), .ZN(
        n1480) );
  NAND3_X1 U1965 ( .A1(n1482), .A2(n1481), .A3(n1480), .ZN(curr_proc_regs[6])
         );
  NAND2_X1 U1966 ( .A1(regs[582]), .A2(n18), .ZN(n1485) );
  AOI22_X1 U1967 ( .A1(n29), .A2(regs[1094]), .B1(n5), .B2(regs[70]), .ZN(
        n1484) );
  AOI22_X1 U1968 ( .A1(n36), .A2(regs[2118]), .B1(n35), .B2(regs[1606]), .ZN(
        n1483) );
  NAND3_X1 U1969 ( .A1(n1485), .A2(n1484), .A3(n1483), .ZN(curr_proc_regs[70])
         );
  NAND2_X1 U1970 ( .A1(regs[583]), .A2(n1579), .ZN(n1488) );
  AOI22_X1 U1971 ( .A1(n29), .A2(regs[1095]), .B1(n5), .B2(regs[71]), .ZN(
        n1487) );
  AOI22_X1 U1972 ( .A1(n36), .A2(regs[2119]), .B1(n3), .B2(regs[1607]), .ZN(
        n1486) );
  NAND3_X1 U1973 ( .A1(n1488), .A2(n1487), .A3(n1486), .ZN(curr_proc_regs[71])
         );
  NAND2_X1 U1974 ( .A1(regs[584]), .A2(n1579), .ZN(n1491) );
  AOI22_X1 U1975 ( .A1(n29), .A2(regs[1096]), .B1(n5), .B2(regs[72]), .ZN(
        n1490) );
  AOI22_X1 U1976 ( .A1(n36), .A2(regs[2120]), .B1(n9), .B2(regs[1608]), .ZN(
        n1489) );
  NAND3_X1 U1977 ( .A1(n1491), .A2(n1490), .A3(n1489), .ZN(curr_proc_regs[72])
         );
  NAND2_X1 U1978 ( .A1(regs[585]), .A2(n11), .ZN(n1494) );
  AOI22_X1 U1979 ( .A1(n29), .A2(regs[1097]), .B1(n5), .B2(regs[73]), .ZN(
        n1493) );
  AOI22_X1 U1980 ( .A1(n36), .A2(regs[2121]), .B1(n34), .B2(regs[1609]), .ZN(
        n1492) );
  NAND3_X1 U1981 ( .A1(n1494), .A2(n1493), .A3(n1492), .ZN(curr_proc_regs[73])
         );
  NAND2_X1 U1982 ( .A1(regs[586]), .A2(n1579), .ZN(n1497) );
  AOI22_X1 U1983 ( .A1(n29), .A2(regs[1098]), .B1(n5), .B2(regs[74]), .ZN(
        n1496) );
  AOI22_X1 U1984 ( .A1(n36), .A2(regs[2122]), .B1(n9), .B2(regs[1610]), .ZN(
        n1495) );
  NAND3_X1 U1985 ( .A1(n1497), .A2(n1496), .A3(n1495), .ZN(curr_proc_regs[74])
         );
  NAND2_X1 U1986 ( .A1(regs[587]), .A2(n7), .ZN(n1500) );
  AOI22_X1 U1987 ( .A1(n29), .A2(regs[1099]), .B1(n26), .B2(regs[75]), .ZN(
        n1499) );
  AOI22_X1 U1988 ( .A1(n36), .A2(regs[2123]), .B1(n9), .B2(regs[1611]), .ZN(
        n1498) );
  NAND3_X1 U1989 ( .A1(n1500), .A2(n1499), .A3(n1498), .ZN(curr_proc_regs[75])
         );
  NAND2_X1 U1990 ( .A1(regs[588]), .A2(n18), .ZN(n1503) );
  AOI22_X1 U1991 ( .A1(n29), .A2(regs[1100]), .B1(n26), .B2(regs[76]), .ZN(
        n1502) );
  AOI22_X1 U1992 ( .A1(n37), .A2(regs[2124]), .B1(n9), .B2(regs[1612]), .ZN(
        n1501) );
  NAND3_X1 U1993 ( .A1(n1503), .A2(n1502), .A3(n1501), .ZN(curr_proc_regs[76])
         );
  NAND2_X1 U1994 ( .A1(regs[589]), .A2(n11), .ZN(n1506) );
  AOI22_X1 U1995 ( .A1(n29), .A2(regs[1101]), .B1(n26), .B2(regs[77]), .ZN(
        n1505) );
  AOI22_X1 U1996 ( .A1(n38), .A2(regs[2125]), .B1(n35), .B2(regs[1613]), .ZN(
        n1504) );
  NAND3_X1 U1997 ( .A1(n1506), .A2(n1505), .A3(n1504), .ZN(curr_proc_regs[77])
         );
  NAND2_X1 U1998 ( .A1(regs[590]), .A2(n16), .ZN(n1509) );
  AOI22_X1 U1999 ( .A1(n29), .A2(regs[1102]), .B1(n26), .B2(regs[78]), .ZN(
        n1508) );
  AOI22_X1 U2000 ( .A1(n38), .A2(regs[2126]), .B1(n3), .B2(regs[1614]), .ZN(
        n1507) );
  NAND3_X1 U2001 ( .A1(n1509), .A2(n1508), .A3(n1507), .ZN(curr_proc_regs[78])
         );
  NAND2_X1 U2002 ( .A1(regs[591]), .A2(n13), .ZN(n1512) );
  AOI22_X1 U2003 ( .A1(n29), .A2(regs[1103]), .B1(n26), .B2(regs[79]), .ZN(
        n1511) );
  AOI22_X1 U2004 ( .A1(n4), .A2(regs[2127]), .B1(n3), .B2(regs[1615]), .ZN(
        n1510) );
  NAND3_X1 U2005 ( .A1(n1512), .A2(n1511), .A3(n1510), .ZN(curr_proc_regs[79])
         );
  NAND2_X1 U2006 ( .A1(regs[519]), .A2(n11), .ZN(n1515) );
  AOI22_X1 U2007 ( .A1(n29), .A2(regs[1031]), .B1(n26), .B2(regs[7]), .ZN(
        n1514) );
  AOI22_X1 U2008 ( .A1(n1), .A2(regs[2055]), .B1(n34), .B2(regs[1543]), .ZN(
        n1513) );
  NAND3_X1 U2009 ( .A1(n1515), .A2(n1514), .A3(n1513), .ZN(curr_proc_regs[7])
         );
  NAND2_X1 U2010 ( .A1(regs[592]), .A2(n11), .ZN(n1518) );
  AOI22_X1 U2011 ( .A1(n29), .A2(regs[1104]), .B1(n26), .B2(regs[80]), .ZN(
        n1517) );
  AOI22_X1 U2012 ( .A1(n37), .A2(regs[2128]), .B1(n33), .B2(regs[1616]), .ZN(
        n1516) );
  NAND3_X1 U2013 ( .A1(n1518), .A2(n1517), .A3(n1516), .ZN(curr_proc_regs[80])
         );
  NAND2_X1 U2014 ( .A1(regs[593]), .A2(n7), .ZN(n1521) );
  AOI22_X1 U2015 ( .A1(n29), .A2(regs[1105]), .B1(n26), .B2(regs[81]), .ZN(
        n1520) );
  AOI22_X1 U2016 ( .A1(n41), .A2(regs[2129]), .B1(n34), .B2(regs[1617]), .ZN(
        n1519) );
  NAND3_X1 U2017 ( .A1(n1521), .A2(n1520), .A3(n1519), .ZN(curr_proc_regs[81])
         );
  NAND2_X1 U2018 ( .A1(regs[594]), .A2(n15), .ZN(n1524) );
  AOI22_X1 U2019 ( .A1(n29), .A2(regs[1106]), .B1(n26), .B2(regs[82]), .ZN(
        n1523) );
  AOI22_X1 U2020 ( .A1(n39), .A2(regs[2130]), .B1(n9), .B2(regs[1618]), .ZN(
        n1522) );
  NAND3_X1 U2021 ( .A1(n1524), .A2(n1523), .A3(n1522), .ZN(curr_proc_regs[82])
         );
  NAND2_X1 U2022 ( .A1(regs[595]), .A2(n16), .ZN(n1527) );
  AOI22_X1 U2023 ( .A1(n29), .A2(regs[1107]), .B1(n26), .B2(regs[83]), .ZN(
        n1526) );
  AOI22_X1 U2024 ( .A1(n10), .A2(regs[2131]), .B1(n9), .B2(regs[1619]), .ZN(
        n1525) );
  NAND3_X1 U2025 ( .A1(n1527), .A2(n1526), .A3(n1525), .ZN(curr_proc_regs[83])
         );
  NAND2_X1 U2026 ( .A1(regs[596]), .A2(n13), .ZN(n1530) );
  AOI22_X1 U2027 ( .A1(n29), .A2(regs[1108]), .B1(n26), .B2(regs[84]), .ZN(
        n1529) );
  AOI22_X1 U2028 ( .A1(n8), .A2(regs[2132]), .B1(n35), .B2(regs[1620]), .ZN(
        n1528) );
  NAND3_X1 U2029 ( .A1(n1530), .A2(n1529), .A3(n1528), .ZN(curr_proc_regs[84])
         );
  NAND2_X1 U2030 ( .A1(regs[597]), .A2(n1579), .ZN(n1533) );
  AOI22_X1 U2031 ( .A1(n29), .A2(regs[1109]), .B1(n5), .B2(regs[85]), .ZN(
        n1532) );
  AOI22_X1 U2032 ( .A1(win[4]), .A2(regs[2133]), .B1(n35), .B2(regs[1621]), 
        .ZN(n1531) );
  NAND3_X1 U2033 ( .A1(n1533), .A2(n1532), .A3(n1531), .ZN(curr_proc_regs[85])
         );
  NAND2_X1 U2034 ( .A1(regs[598]), .A2(n11), .ZN(n1536) );
  AOI22_X1 U2035 ( .A1(n29), .A2(regs[1110]), .B1(n12), .B2(regs[86]), .ZN(
        n1535) );
  AOI22_X1 U2036 ( .A1(n10), .A2(regs[2134]), .B1(n9), .B2(regs[1622]), .ZN(
        n1534) );
  NAND3_X1 U2037 ( .A1(n1536), .A2(n1535), .A3(n1534), .ZN(curr_proc_regs[86])
         );
  NAND2_X1 U2038 ( .A1(regs[599]), .A2(n1579), .ZN(n1539) );
  AOI22_X1 U2039 ( .A1(n29), .A2(regs[1111]), .B1(n28), .B2(regs[87]), .ZN(
        n1538) );
  AOI22_X1 U2040 ( .A1(n4), .A2(regs[2135]), .B1(n32), .B2(regs[1623]), .ZN(
        n1537) );
  NAND3_X1 U2041 ( .A1(n1539), .A2(n1538), .A3(n1537), .ZN(curr_proc_regs[87])
         );
  NAND2_X1 U2042 ( .A1(regs[600]), .A2(n11), .ZN(n1542) );
  AOI22_X1 U2043 ( .A1(n29), .A2(regs[1112]), .B1(n5), .B2(regs[88]), .ZN(
        n1541) );
  AOI22_X1 U2044 ( .A1(n37), .A2(regs[2136]), .B1(n35), .B2(regs[1624]), .ZN(
        n1540) );
  NAND3_X1 U2045 ( .A1(n1542), .A2(n1541), .A3(n1540), .ZN(curr_proc_regs[88])
         );
  NAND2_X1 U2046 ( .A1(regs[601]), .A2(n1579), .ZN(n1545) );
  AOI22_X1 U2047 ( .A1(n29), .A2(regs[1113]), .B1(n12), .B2(regs[89]), .ZN(
        n1544) );
  AOI22_X1 U2048 ( .A1(n39), .A2(regs[2137]), .B1(n31), .B2(regs[1625]), .ZN(
        n1543) );
  NAND3_X1 U2049 ( .A1(n1545), .A2(n1544), .A3(n1543), .ZN(curr_proc_regs[89])
         );
  NAND2_X1 U2050 ( .A1(regs[520]), .A2(n13), .ZN(n1548) );
  AOI22_X1 U2051 ( .A1(n29), .A2(regs[1032]), .B1(n28), .B2(regs[8]), .ZN(
        n1547) );
  AOI22_X1 U2052 ( .A1(n8), .A2(regs[2056]), .B1(n33), .B2(regs[1544]), .ZN(
        n1546) );
  NAND3_X1 U2053 ( .A1(n1548), .A2(n1547), .A3(n1546), .ZN(curr_proc_regs[8])
         );
  NAND2_X1 U2054 ( .A1(regs[602]), .A2(n1579), .ZN(n1551) );
  AOI22_X1 U2055 ( .A1(n29), .A2(regs[1114]), .B1(n5), .B2(regs[90]), .ZN(
        n1550) );
  AOI22_X1 U2056 ( .A1(n41), .A2(regs[2138]), .B1(n32), .B2(regs[1626]), .ZN(
        n1549) );
  NAND3_X1 U2057 ( .A1(n1551), .A2(n1550), .A3(n1549), .ZN(curr_proc_regs[90])
         );
  NAND2_X1 U2058 ( .A1(regs[603]), .A2(n17), .ZN(n1554) );
  AOI22_X1 U2059 ( .A1(n29), .A2(regs[1115]), .B1(n12), .B2(regs[91]), .ZN(
        n1553) );
  AOI22_X1 U2060 ( .A1(n1), .A2(regs[2139]), .B1(n3), .B2(regs[1627]), .ZN(
        n1552) );
  NAND3_X1 U2061 ( .A1(n1554), .A2(n1553), .A3(n1552), .ZN(curr_proc_regs[91])
         );
  NAND2_X1 U2062 ( .A1(regs[604]), .A2(n14), .ZN(n1557) );
  AOI22_X1 U2063 ( .A1(n29), .A2(regs[1116]), .B1(n28), .B2(regs[92]), .ZN(
        n1556) );
  AOI22_X1 U2064 ( .A1(n10), .A2(regs[2140]), .B1(n3), .B2(regs[1628]), .ZN(
        n1555) );
  NAND3_X1 U2065 ( .A1(n1557), .A2(n1556), .A3(n1555), .ZN(curr_proc_regs[92])
         );
  NAND2_X1 U2066 ( .A1(regs[605]), .A2(n13), .ZN(n1560) );
  AOI22_X1 U2067 ( .A1(n29), .A2(regs[1117]), .B1(n5), .B2(regs[93]), .ZN(
        n1559) );
  AOI22_X1 U2068 ( .A1(n4), .A2(regs[2141]), .B1(n3), .B2(regs[1629]), .ZN(
        n1558) );
  NAND3_X1 U2069 ( .A1(n1560), .A2(n1559), .A3(n1558), .ZN(curr_proc_regs[93])
         );
  NAND2_X1 U2070 ( .A1(regs[606]), .A2(n19), .ZN(n1563) );
  AOI22_X1 U2071 ( .A1(n29), .A2(regs[1118]), .B1(n28), .B2(regs[94]), .ZN(
        n1562) );
  AOI22_X1 U2072 ( .A1(n37), .A2(regs[2142]), .B1(n34), .B2(regs[1630]), .ZN(
        n1561) );
  NAND3_X1 U2073 ( .A1(n1563), .A2(n1562), .A3(n1561), .ZN(curr_proc_regs[94])
         );
  NAND2_X1 U2074 ( .A1(regs[607]), .A2(n20), .ZN(n1566) );
  AOI22_X1 U2075 ( .A1(n29), .A2(regs[1119]), .B1(n5), .B2(regs[95]), .ZN(
        n1565) );
  AOI22_X1 U2076 ( .A1(n39), .A2(regs[2143]), .B1(n3), .B2(regs[1631]), .ZN(
        n1564) );
  NAND3_X1 U2077 ( .A1(n1566), .A2(n1565), .A3(n1564), .ZN(curr_proc_regs[95])
         );
  NAND2_X1 U2078 ( .A1(regs[608]), .A2(n20), .ZN(n1569) );
  AOI22_X1 U2079 ( .A1(n29), .A2(regs[1120]), .B1(n5), .B2(regs[96]), .ZN(
        n1568) );
  AOI22_X1 U2080 ( .A1(n40), .A2(regs[2144]), .B1(n3), .B2(regs[1632]), .ZN(
        n1567) );
  NAND3_X1 U2081 ( .A1(n1569), .A2(n1568), .A3(n1567), .ZN(curr_proc_regs[96])
         );
  NAND2_X1 U2082 ( .A1(regs[609]), .A2(n20), .ZN(n1572) );
  AOI22_X1 U2083 ( .A1(n29), .A2(regs[1121]), .B1(n5), .B2(regs[97]), .ZN(
        n1571) );
  AOI22_X1 U2084 ( .A1(n39), .A2(regs[2145]), .B1(n35), .B2(regs[1633]), .ZN(
        n1570) );
  NAND3_X1 U2085 ( .A1(n1572), .A2(n1571), .A3(n1570), .ZN(curr_proc_regs[97])
         );
  NAND2_X1 U2086 ( .A1(regs[610]), .A2(n20), .ZN(n1575) );
  AOI22_X1 U2087 ( .A1(n29), .A2(regs[1122]), .B1(n5), .B2(regs[98]), .ZN(
        n1574) );
  AOI22_X1 U2088 ( .A1(n8), .A2(regs[2146]), .B1(n34), .B2(regs[1634]), .ZN(
        n1573) );
  NAND3_X1 U2089 ( .A1(n1575), .A2(n1574), .A3(n1573), .ZN(curr_proc_regs[98])
         );
  NAND2_X1 U2090 ( .A1(regs[611]), .A2(n20), .ZN(n1578) );
  AOI22_X1 U2091 ( .A1(n29), .A2(regs[1123]), .B1(n5), .B2(regs[99]), .ZN(
        n1577) );
  AOI22_X1 U2092 ( .A1(n4), .A2(regs[2147]), .B1(n3), .B2(regs[1635]), .ZN(
        n1576) );
  NAND3_X1 U2093 ( .A1(n1578), .A2(n1577), .A3(n1576), .ZN(curr_proc_regs[99])
         );
  NAND2_X1 U2094 ( .A1(regs[521]), .A2(n20), .ZN(n1585) );
  AOI22_X1 U2095 ( .A1(n29), .A2(regs[1033]), .B1(n5), .B2(regs[9]), .ZN(n1584) );
  AOI22_X1 U2096 ( .A1(n41), .A2(regs[2057]), .B1(n3), .B2(regs[1545]), .ZN(
        n1583) );
  NAND3_X1 U2097 ( .A1(n1585), .A2(n1584), .A3(n1583), .ZN(curr_proc_regs[9])
         );
endmodule


module mux_N32_M5_1 ( S, Q, Y );
  input [4:0] S;
  input [1023:0] Q;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688;

  AOI22_X1 U2 ( .A1(n674), .A2(Q[499]), .B1(n673), .B2(Q[563]), .ZN(n1) );
  AOI22_X1 U3 ( .A1(n676), .A2(Q[659]), .B1(n675), .B2(Q[467]), .ZN(n2) );
  AOI22_X1 U4 ( .A1(n678), .A2(Q[371]), .B1(n677), .B2(Q[307]), .ZN(n3) );
  AOI22_X1 U5 ( .A1(n680), .A2(Q[403]), .B1(n679), .B2(Q[275]), .ZN(n4) );
  NAND4_X1 U6 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(n5) );
  AOI22_X1 U7 ( .A1(n682), .A2(Q[339]), .B1(n681), .B2(Q[435]), .ZN(n6) );
  AOI22_X1 U8 ( .A1(n684), .A2(Q[243]), .B1(n683), .B2(Q[147]), .ZN(n7) );
  AOI22_X1 U9 ( .A1(n686), .A2(Q[83]), .B1(n685), .B2(Q[179]), .ZN(n8) );
  AOI22_X1 U10 ( .A1(n688), .A2(Q[211]), .B1(n687), .B2(Q[51]), .ZN(n9) );
  NAND4_X1 U11 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n10) );
  AOI22_X1 U12 ( .A1(n657), .A2(Q[1011]), .B1(n656), .B2(Q[947]), .ZN(n11) );
  AOI22_X1 U13 ( .A1(n659), .A2(Q[979]), .B1(n658), .B2(Q[915]), .ZN(n12) );
  AOI222_X1 U14 ( .A1(n661), .A2(Q[819]), .B1(n662), .B2(Q[115]), .C1(n660), 
        .C2(Q[755]), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n14) );
  AOI22_X1 U16 ( .A1(n664), .A2(Q[851]), .B1(n663), .B2(Q[723]), .ZN(n15) );
  AOI22_X1 U17 ( .A1(n666), .A2(Q[787]), .B1(n665), .B2(Q[883]), .ZN(n16) );
  NAND4_X1 U18 ( .A1(n614), .A2(n615), .A3(n15), .A4(n16), .ZN(n17) );
  OR4_X1 U19 ( .A1(n5), .A2(n10), .A3(n14), .A4(n17), .ZN(Y[19]) );
  AOI22_X1 U20 ( .A1(n674), .A2(Q[509]), .B1(n673), .B2(Q[573]), .ZN(n18) );
  AOI22_X1 U21 ( .A1(n676), .A2(Q[669]), .B1(n675), .B2(Q[477]), .ZN(n19) );
  AOI22_X1 U22 ( .A1(n678), .A2(Q[381]), .B1(n677), .B2(Q[317]), .ZN(n20) );
  AOI22_X1 U23 ( .A1(n680), .A2(Q[413]), .B1(n679), .B2(Q[285]), .ZN(n21) );
  NAND4_X1 U24 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .ZN(n22) );
  AOI22_X1 U25 ( .A1(n682), .A2(Q[349]), .B1(n681), .B2(Q[445]), .ZN(n23) );
  AOI22_X1 U26 ( .A1(n684), .A2(Q[253]), .B1(n683), .B2(Q[157]), .ZN(n24) );
  AOI22_X1 U27 ( .A1(n686), .A2(Q[93]), .B1(n685), .B2(Q[189]), .ZN(n25) );
  AOI22_X1 U28 ( .A1(n688), .A2(Q[221]), .B1(n687), .B2(Q[61]), .ZN(n26) );
  NAND4_X1 U29 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(n27) );
  AOI22_X1 U30 ( .A1(n657), .A2(Q[1021]), .B1(n656), .B2(Q[957]), .ZN(n28) );
  AOI22_X1 U31 ( .A1(n659), .A2(Q[989]), .B1(n658), .B2(Q[925]), .ZN(n29) );
  AOI222_X1 U32 ( .A1(n661), .A2(Q[829]), .B1(n662), .B2(Q[125]), .C1(n660), 
        .C2(Q[765]), .ZN(n30) );
  NAND3_X1 U33 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n31) );
  AOI22_X1 U34 ( .A1(n664), .A2(Q[861]), .B1(n663), .B2(Q[733]), .ZN(n32) );
  AOI22_X1 U35 ( .A1(n666), .A2(Q[797]), .B1(n665), .B2(Q[893]), .ZN(n33) );
  NAND4_X1 U36 ( .A1(n636), .A2(n637), .A3(n32), .A4(n33), .ZN(n34) );
  OR4_X1 U37 ( .A1(n22), .A2(n27), .A3(n31), .A4(n34), .ZN(Y[29]) );
  AOI22_X1 U38 ( .A1(n674), .A2(Q[497]), .B1(n673), .B2(Q[561]), .ZN(n35) );
  AOI22_X1 U39 ( .A1(n676), .A2(Q[657]), .B1(n675), .B2(Q[465]), .ZN(n36) );
  AOI22_X1 U40 ( .A1(n678), .A2(Q[369]), .B1(n677), .B2(Q[305]), .ZN(n37) );
  AOI22_X1 U41 ( .A1(n680), .A2(Q[401]), .B1(n679), .B2(Q[273]), .ZN(n38) );
  NAND4_X1 U42 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(n39) );
  AOI22_X1 U43 ( .A1(n682), .A2(Q[337]), .B1(n681), .B2(Q[433]), .ZN(n40) );
  AOI22_X1 U44 ( .A1(n684), .A2(Q[241]), .B1(n683), .B2(Q[145]), .ZN(n41) );
  AOI22_X1 U45 ( .A1(n686), .A2(Q[81]), .B1(n685), .B2(Q[177]), .ZN(n42) );
  AOI22_X1 U46 ( .A1(n688), .A2(Q[209]), .B1(n687), .B2(Q[49]), .ZN(n43) );
  NAND4_X1 U47 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n44) );
  AOI22_X1 U48 ( .A1(n657), .A2(Q[1009]), .B1(n656), .B2(Q[945]), .ZN(n45) );
  AOI22_X1 U49 ( .A1(n659), .A2(Q[977]), .B1(n658), .B2(Q[913]), .ZN(n46) );
  AOI222_X1 U50 ( .A1(n661), .A2(Q[817]), .B1(n662), .B2(Q[113]), .C1(n660), 
        .C2(Q[753]), .ZN(n47) );
  NAND3_X1 U51 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n48) );
  AOI22_X1 U52 ( .A1(n664), .A2(Q[849]), .B1(n663), .B2(Q[721]), .ZN(n49) );
  AOI22_X1 U53 ( .A1(n666), .A2(Q[785]), .B1(n665), .B2(Q[881]), .ZN(n50) );
  NAND4_X1 U54 ( .A1(n610), .A2(n611), .A3(n49), .A4(n50), .ZN(n51) );
  OR4_X1 U55 ( .A1(n39), .A2(n44), .A3(n48), .A4(n51), .ZN(Y[17]) );
  AOI22_X1 U56 ( .A1(n674), .A2(Q[498]), .B1(n673), .B2(Q[562]), .ZN(n52) );
  AOI22_X1 U57 ( .A1(n676), .A2(Q[658]), .B1(n675), .B2(Q[466]), .ZN(n53) );
  AOI22_X1 U58 ( .A1(n678), .A2(Q[370]), .B1(n677), .B2(Q[306]), .ZN(n54) );
  AOI22_X1 U59 ( .A1(n680), .A2(Q[402]), .B1(n679), .B2(Q[274]), .ZN(n55) );
  NAND4_X1 U60 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .ZN(n56) );
  AOI22_X1 U61 ( .A1(n682), .A2(Q[338]), .B1(n681), .B2(Q[434]), .ZN(n57) );
  AOI22_X1 U62 ( .A1(n684), .A2(Q[242]), .B1(n683), .B2(Q[146]), .ZN(n58) );
  AOI22_X1 U63 ( .A1(n686), .A2(Q[82]), .B1(n685), .B2(Q[178]), .ZN(n59) );
  AOI22_X1 U64 ( .A1(n688), .A2(Q[210]), .B1(n687), .B2(Q[50]), .ZN(n60) );
  NAND4_X1 U65 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(n61) );
  AOI22_X1 U66 ( .A1(n657), .A2(Q[1010]), .B1(n656), .B2(Q[946]), .ZN(n62) );
  AOI22_X1 U67 ( .A1(n659), .A2(Q[978]), .B1(n658), .B2(Q[914]), .ZN(n63) );
  AOI222_X1 U68 ( .A1(n661), .A2(Q[818]), .B1(n662), .B2(Q[114]), .C1(n660), 
        .C2(Q[754]), .ZN(n64) );
  NAND3_X1 U69 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n65) );
  AOI22_X1 U70 ( .A1(n664), .A2(Q[850]), .B1(n663), .B2(Q[722]), .ZN(n66) );
  AOI22_X1 U71 ( .A1(n666), .A2(Q[786]), .B1(n665), .B2(Q[882]), .ZN(n67) );
  NAND4_X1 U72 ( .A1(n612), .A2(n613), .A3(n66), .A4(n67), .ZN(n68) );
  OR4_X1 U73 ( .A1(n56), .A2(n61), .A3(n65), .A4(n68), .ZN(Y[18]) );
  AOI22_X1 U74 ( .A1(n674), .A2(Q[495]), .B1(n673), .B2(Q[559]), .ZN(n69) );
  AOI22_X1 U75 ( .A1(n676), .A2(Q[655]), .B1(n675), .B2(Q[463]), .ZN(n70) );
  AOI22_X1 U76 ( .A1(n678), .A2(Q[367]), .B1(n677), .B2(Q[303]), .ZN(n71) );
  AOI22_X1 U77 ( .A1(n680), .A2(Q[399]), .B1(n679), .B2(Q[271]), .ZN(n72) );
  NAND4_X1 U78 ( .A1(n69), .A2(n70), .A3(n71), .A4(n72), .ZN(n73) );
  AOI22_X1 U79 ( .A1(n682), .A2(Q[335]), .B1(n681), .B2(Q[431]), .ZN(n74) );
  AOI22_X1 U80 ( .A1(n684), .A2(Q[239]), .B1(n683), .B2(Q[143]), .ZN(n75) );
  AOI22_X1 U81 ( .A1(n686), .A2(Q[79]), .B1(n685), .B2(Q[175]), .ZN(n76) );
  AOI22_X1 U82 ( .A1(n688), .A2(Q[207]), .B1(n687), .B2(Q[47]), .ZN(n77) );
  NAND4_X1 U83 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(n78) );
  AOI22_X1 U84 ( .A1(n657), .A2(Q[1007]), .B1(n656), .B2(Q[943]), .ZN(n79) );
  AOI22_X1 U85 ( .A1(n659), .A2(Q[975]), .B1(n658), .B2(Q[911]), .ZN(n80) );
  AOI222_X1 U86 ( .A1(n661), .A2(Q[815]), .B1(n662), .B2(Q[111]), .C1(n660), 
        .C2(Q[751]), .ZN(n81) );
  NAND3_X1 U87 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n82) );
  AOI22_X1 U88 ( .A1(n664), .A2(Q[847]), .B1(n663), .B2(Q[719]), .ZN(n83) );
  AOI22_X1 U89 ( .A1(n666), .A2(Q[783]), .B1(n665), .B2(Q[879]), .ZN(n84) );
  NAND4_X1 U90 ( .A1(n606), .A2(n607), .A3(n83), .A4(n84), .ZN(n85) );
  OR4_X1 U91 ( .A1(n73), .A2(n78), .A3(n82), .A4(n85), .ZN(Y[15]) );
  AOI22_X1 U92 ( .A1(n674), .A2(Q[496]), .B1(n673), .B2(Q[560]), .ZN(n86) );
  AOI22_X1 U93 ( .A1(n676), .A2(Q[656]), .B1(n675), .B2(Q[464]), .ZN(n87) );
  AOI22_X1 U94 ( .A1(n678), .A2(Q[368]), .B1(n677), .B2(Q[304]), .ZN(n88) );
  AOI22_X1 U95 ( .A1(n680), .A2(Q[400]), .B1(n679), .B2(Q[272]), .ZN(n89) );
  NAND4_X1 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(n90) );
  AOI22_X1 U97 ( .A1(n682), .A2(Q[336]), .B1(n681), .B2(Q[432]), .ZN(n91) );
  AOI22_X1 U98 ( .A1(n684), .A2(Q[240]), .B1(n683), .B2(Q[144]), .ZN(n92) );
  AOI22_X1 U99 ( .A1(n686), .A2(Q[80]), .B1(n685), .B2(Q[176]), .ZN(n93) );
  AOI22_X1 U100 ( .A1(n688), .A2(Q[208]), .B1(n687), .B2(Q[48]), .ZN(n94) );
  NAND4_X1 U101 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(n95) );
  AOI22_X1 U102 ( .A1(n657), .A2(Q[1008]), .B1(n656), .B2(Q[944]), .ZN(n96) );
  AOI22_X1 U103 ( .A1(n659), .A2(Q[976]), .B1(n658), .B2(Q[912]), .ZN(n97) );
  AOI222_X1 U104 ( .A1(n661), .A2(Q[816]), .B1(n662), .B2(Q[112]), .C1(n660), 
        .C2(Q[752]), .ZN(n98) );
  NAND3_X1 U105 ( .A1(n96), .A2(n97), .A3(n98), .ZN(n99) );
  AOI22_X1 U106 ( .A1(n664), .A2(Q[848]), .B1(n663), .B2(Q[720]), .ZN(n100) );
  AOI22_X1 U107 ( .A1(n666), .A2(Q[784]), .B1(n665), .B2(Q[880]), .ZN(n101) );
  NAND4_X1 U108 ( .A1(n608), .A2(n609), .A3(n100), .A4(n101), .ZN(n102) );
  OR4_X1 U109 ( .A1(n90), .A2(n95), .A3(n99), .A4(n102), .ZN(Y[16]) );
  AOI22_X1 U110 ( .A1(n674), .A2(Q[493]), .B1(n673), .B2(Q[557]), .ZN(n103) );
  AOI22_X1 U111 ( .A1(n676), .A2(Q[653]), .B1(n675), .B2(Q[461]), .ZN(n104) );
  AOI22_X1 U112 ( .A1(n678), .A2(Q[365]), .B1(n677), .B2(Q[301]), .ZN(n105) );
  AOI22_X1 U113 ( .A1(n680), .A2(Q[397]), .B1(n679), .B2(Q[269]), .ZN(n106) );
  NAND4_X1 U114 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(n107) );
  AOI22_X1 U115 ( .A1(n682), .A2(Q[333]), .B1(n681), .B2(Q[429]), .ZN(n108) );
  AOI22_X1 U116 ( .A1(n684), .A2(Q[237]), .B1(n683), .B2(Q[141]), .ZN(n109) );
  AOI22_X1 U117 ( .A1(n686), .A2(Q[77]), .B1(n685), .B2(Q[173]), .ZN(n110) );
  AOI22_X1 U118 ( .A1(n688), .A2(Q[205]), .B1(n687), .B2(Q[45]), .ZN(n111) );
  NAND4_X1 U119 ( .A1(n108), .A2(n109), .A3(n110), .A4(n111), .ZN(n112) );
  AOI22_X1 U120 ( .A1(n657), .A2(Q[1005]), .B1(n656), .B2(Q[941]), .ZN(n113)
         );
  AOI22_X1 U121 ( .A1(n659), .A2(Q[973]), .B1(n658), .B2(Q[909]), .ZN(n114) );
  AOI222_X1 U122 ( .A1(n661), .A2(Q[813]), .B1(n662), .B2(Q[109]), .C1(n660), 
        .C2(Q[749]), .ZN(n115) );
  NAND3_X1 U123 ( .A1(n113), .A2(n114), .A3(n115), .ZN(n116) );
  AOI22_X1 U124 ( .A1(n664), .A2(Q[845]), .B1(n663), .B2(Q[717]), .ZN(n117) );
  AOI22_X1 U125 ( .A1(n666), .A2(Q[781]), .B1(n665), .B2(Q[877]), .ZN(n118) );
  NAND4_X1 U126 ( .A1(n602), .A2(n603), .A3(n117), .A4(n118), .ZN(n119) );
  OR4_X1 U127 ( .A1(n107), .A2(n112), .A3(n116), .A4(n119), .ZN(Y[13]) );
  AOI22_X1 U128 ( .A1(n674), .A2(Q[494]), .B1(n673), .B2(Q[558]), .ZN(n120) );
  AOI22_X1 U129 ( .A1(n676), .A2(Q[654]), .B1(n675), .B2(Q[462]), .ZN(n121) );
  AOI22_X1 U130 ( .A1(n678), .A2(Q[366]), .B1(n677), .B2(Q[302]), .ZN(n122) );
  AOI22_X1 U131 ( .A1(n680), .A2(Q[398]), .B1(n679), .B2(Q[270]), .ZN(n123) );
  NAND4_X1 U132 ( .A1(n120), .A2(n121), .A3(n122), .A4(n123), .ZN(n124) );
  AOI22_X1 U133 ( .A1(n682), .A2(Q[334]), .B1(n681), .B2(Q[430]), .ZN(n125) );
  AOI22_X1 U134 ( .A1(n684), .A2(Q[238]), .B1(n683), .B2(Q[142]), .ZN(n126) );
  AOI22_X1 U135 ( .A1(n686), .A2(Q[78]), .B1(n685), .B2(Q[174]), .ZN(n127) );
  AOI22_X1 U136 ( .A1(n688), .A2(Q[206]), .B1(n687), .B2(Q[46]), .ZN(n128) );
  NAND4_X1 U137 ( .A1(n125), .A2(n126), .A3(n127), .A4(n128), .ZN(n129) );
  AOI22_X1 U138 ( .A1(n657), .A2(Q[1006]), .B1(n656), .B2(Q[942]), .ZN(n130)
         );
  AOI22_X1 U139 ( .A1(n659), .A2(Q[974]), .B1(n658), .B2(Q[910]), .ZN(n131) );
  AOI222_X1 U140 ( .A1(n661), .A2(Q[814]), .B1(n662), .B2(Q[110]), .C1(n660), 
        .C2(Q[750]), .ZN(n132) );
  NAND3_X1 U141 ( .A1(n130), .A2(n131), .A3(n132), .ZN(n133) );
  AOI22_X1 U142 ( .A1(n664), .A2(Q[846]), .B1(n663), .B2(Q[718]), .ZN(n134) );
  AOI22_X1 U143 ( .A1(n666), .A2(Q[782]), .B1(n665), .B2(Q[878]), .ZN(n135) );
  NAND4_X1 U144 ( .A1(n604), .A2(n605), .A3(n134), .A4(n135), .ZN(n136) );
  OR4_X1 U145 ( .A1(n124), .A2(n129), .A3(n133), .A4(n136), .ZN(Y[14]) );
  AOI22_X1 U146 ( .A1(n562), .A2(Q[510]), .B1(n561), .B2(Q[574]), .ZN(n137) );
  AOI22_X1 U147 ( .A1(n564), .A2(Q[670]), .B1(n563), .B2(Q[478]), .ZN(n138) );
  AOI22_X1 U148 ( .A1(n566), .A2(Q[382]), .B1(n565), .B2(Q[318]), .ZN(n139) );
  AOI22_X1 U149 ( .A1(n568), .A2(Q[414]), .B1(n567), .B2(Q[286]), .ZN(n140) );
  NAND4_X1 U150 ( .A1(n137), .A2(n138), .A3(n139), .A4(n140), .ZN(n141) );
  AOI22_X1 U151 ( .A1(n570), .A2(Q[350]), .B1(n569), .B2(Q[446]), .ZN(n142) );
  AOI22_X1 U152 ( .A1(n572), .A2(Q[254]), .B1(n571), .B2(Q[158]), .ZN(n143) );
  AOI22_X1 U153 ( .A1(n574), .A2(Q[94]), .B1(n573), .B2(Q[190]), .ZN(n144) );
  AOI22_X1 U154 ( .A1(n576), .A2(Q[222]), .B1(n575), .B2(Q[62]), .ZN(n145) );
  NAND4_X1 U155 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(n146) );
  AOI22_X1 U156 ( .A1(n547), .A2(Q[1022]), .B1(n546), .B2(Q[958]), .ZN(n147)
         );
  AOI22_X1 U157 ( .A1(n549), .A2(Q[990]), .B1(n548), .B2(Q[926]), .ZN(n148) );
  AOI222_X1 U158 ( .A1(n551), .A2(Q[830]), .B1(n552), .B2(Q[126]), .C1(n550), 
        .C2(Q[766]), .ZN(n149) );
  NAND3_X1 U159 ( .A1(n147), .A2(n148), .A3(n149), .ZN(n150) );
  AOI22_X1 U160 ( .A1(n554), .A2(Q[862]), .B1(n553), .B2(Q[734]), .ZN(n151) );
  AOI22_X1 U161 ( .A1(n556), .A2(Q[798]), .B1(n555), .B2(Q[894]), .ZN(n152) );
  NAND4_X1 U162 ( .A1(n640), .A2(n641), .A3(n151), .A4(n152), .ZN(n153) );
  OR4_X1 U163 ( .A1(n141), .A2(n146), .A3(n150), .A4(n153), .ZN(Y[30]) );
  AOI22_X1 U164 ( .A1(n562), .A2(Q[508]), .B1(n561), .B2(Q[572]), .ZN(n154) );
  AOI22_X1 U165 ( .A1(n564), .A2(Q[668]), .B1(n563), .B2(Q[476]), .ZN(n155) );
  AOI22_X1 U166 ( .A1(n566), .A2(Q[380]), .B1(n565), .B2(Q[316]), .ZN(n156) );
  AOI22_X1 U167 ( .A1(n568), .A2(Q[412]), .B1(n567), .B2(Q[284]), .ZN(n157) );
  NAND4_X1 U168 ( .A1(n154), .A2(n155), .A3(n156), .A4(n157), .ZN(n158) );
  AOI22_X1 U169 ( .A1(n570), .A2(Q[348]), .B1(n569), .B2(Q[444]), .ZN(n159) );
  AOI22_X1 U170 ( .A1(n572), .A2(Q[252]), .B1(n571), .B2(Q[156]), .ZN(n160) );
  AOI22_X1 U171 ( .A1(n574), .A2(Q[92]), .B1(n573), .B2(Q[188]), .ZN(n161) );
  AOI22_X1 U172 ( .A1(n576), .A2(Q[220]), .B1(n575), .B2(Q[60]), .ZN(n162) );
  NAND4_X1 U173 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(n163) );
  AOI22_X1 U174 ( .A1(n547), .A2(Q[1020]), .B1(n546), .B2(Q[956]), .ZN(n164)
         );
  AOI22_X1 U175 ( .A1(n549), .A2(Q[988]), .B1(n548), .B2(Q[924]), .ZN(n165) );
  AOI222_X1 U176 ( .A1(n551), .A2(Q[828]), .B1(n552), .B2(Q[124]), .C1(n550), 
        .C2(Q[764]), .ZN(n166) );
  NAND3_X1 U177 ( .A1(n164), .A2(n165), .A3(n166), .ZN(n167) );
  AOI22_X1 U178 ( .A1(n554), .A2(Q[860]), .B1(n553), .B2(Q[732]), .ZN(n168) );
  AOI22_X1 U179 ( .A1(n556), .A2(Q[796]), .B1(n555), .B2(Q[892]), .ZN(n169) );
  NAND4_X1 U180 ( .A1(n634), .A2(n635), .A3(n168), .A4(n169), .ZN(n170) );
  OR4_X1 U181 ( .A1(n158), .A2(n163), .A3(n167), .A4(n170), .ZN(Y[28]) );
  AOI22_X1 U182 ( .A1(n562), .A2(Q[507]), .B1(n561), .B2(Q[571]), .ZN(n171) );
  AOI22_X1 U183 ( .A1(n564), .A2(Q[667]), .B1(n563), .B2(Q[475]), .ZN(n172) );
  AOI22_X1 U184 ( .A1(n566), .A2(Q[379]), .B1(n565), .B2(Q[315]), .ZN(n173) );
  AOI22_X1 U185 ( .A1(n568), .A2(Q[411]), .B1(n567), .B2(Q[283]), .ZN(n174) );
  NAND4_X1 U186 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(n175) );
  AOI22_X1 U187 ( .A1(n570), .A2(Q[347]), .B1(n569), .B2(Q[443]), .ZN(n176) );
  AOI22_X1 U188 ( .A1(n572), .A2(Q[251]), .B1(n571), .B2(Q[155]), .ZN(n177) );
  AOI22_X1 U189 ( .A1(n574), .A2(Q[91]), .B1(n573), .B2(Q[187]), .ZN(n178) );
  AOI22_X1 U190 ( .A1(n576), .A2(Q[219]), .B1(n575), .B2(Q[59]), .ZN(n179) );
  NAND4_X1 U191 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(n180) );
  AOI22_X1 U192 ( .A1(n547), .A2(Q[1019]), .B1(n546), .B2(Q[955]), .ZN(n181)
         );
  AOI22_X1 U193 ( .A1(n549), .A2(Q[987]), .B1(n548), .B2(Q[923]), .ZN(n182) );
  AOI222_X1 U194 ( .A1(n551), .A2(Q[827]), .B1(n552), .B2(Q[123]), .C1(n550), 
        .C2(Q[763]), .ZN(n183) );
  NAND3_X1 U195 ( .A1(n181), .A2(n182), .A3(n183), .ZN(n184) );
  AOI22_X1 U196 ( .A1(n554), .A2(Q[859]), .B1(n553), .B2(Q[731]), .ZN(n185) );
  AOI22_X1 U197 ( .A1(n556), .A2(Q[795]), .B1(n555), .B2(Q[891]), .ZN(n186) );
  NAND4_X1 U198 ( .A1(n632), .A2(n633), .A3(n185), .A4(n186), .ZN(n187) );
  OR4_X1 U199 ( .A1(n175), .A2(n180), .A3(n184), .A4(n187), .ZN(Y[27]) );
  AOI22_X1 U200 ( .A1(n562), .A2(Q[506]), .B1(n561), .B2(Q[570]), .ZN(n188) );
  AOI22_X1 U201 ( .A1(n564), .A2(Q[666]), .B1(n563), .B2(Q[474]), .ZN(n189) );
  AOI22_X1 U202 ( .A1(n566), .A2(Q[378]), .B1(n565), .B2(Q[314]), .ZN(n190) );
  AOI22_X1 U203 ( .A1(n568), .A2(Q[410]), .B1(n567), .B2(Q[282]), .ZN(n191) );
  NAND4_X1 U204 ( .A1(n188), .A2(n189), .A3(n190), .A4(n191), .ZN(n192) );
  AOI22_X1 U205 ( .A1(n570), .A2(Q[346]), .B1(n569), .B2(Q[442]), .ZN(n193) );
  AOI22_X1 U206 ( .A1(n572), .A2(Q[250]), .B1(n571), .B2(Q[154]), .ZN(n194) );
  AOI22_X1 U207 ( .A1(n574), .A2(Q[90]), .B1(n573), .B2(Q[186]), .ZN(n195) );
  AOI22_X1 U208 ( .A1(n576), .A2(Q[218]), .B1(n575), .B2(Q[58]), .ZN(n196) );
  NAND4_X1 U209 ( .A1(n193), .A2(n194), .A3(n195), .A4(n196), .ZN(n197) );
  AOI22_X1 U210 ( .A1(n547), .A2(Q[1018]), .B1(n546), .B2(Q[954]), .ZN(n198)
         );
  AOI22_X1 U211 ( .A1(n549), .A2(Q[986]), .B1(n548), .B2(Q[922]), .ZN(n199) );
  AOI222_X1 U212 ( .A1(n551), .A2(Q[826]), .B1(n552), .B2(Q[122]), .C1(n550), 
        .C2(Q[762]), .ZN(n200) );
  NAND3_X1 U213 ( .A1(n198), .A2(n199), .A3(n200), .ZN(n201) );
  AOI22_X1 U214 ( .A1(n554), .A2(Q[858]), .B1(n553), .B2(Q[730]), .ZN(n202) );
  AOI22_X1 U215 ( .A1(n556), .A2(Q[794]), .B1(n555), .B2(Q[890]), .ZN(n203) );
  NAND4_X1 U216 ( .A1(n630), .A2(n631), .A3(n202), .A4(n203), .ZN(n204) );
  OR4_X1 U217 ( .A1(n192), .A2(n197), .A3(n201), .A4(n204), .ZN(Y[26]) );
  AOI22_X1 U218 ( .A1(n562), .A2(Q[505]), .B1(n561), .B2(Q[569]), .ZN(n205) );
  AOI22_X1 U219 ( .A1(n564), .A2(Q[665]), .B1(n563), .B2(Q[473]), .ZN(n206) );
  AOI22_X1 U220 ( .A1(n566), .A2(Q[377]), .B1(n565), .B2(Q[313]), .ZN(n207) );
  AOI22_X1 U221 ( .A1(n568), .A2(Q[409]), .B1(n567), .B2(Q[281]), .ZN(n208) );
  NAND4_X1 U222 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n209) );
  AOI22_X1 U223 ( .A1(n570), .A2(Q[345]), .B1(n569), .B2(Q[441]), .ZN(n210) );
  AOI22_X1 U224 ( .A1(n572), .A2(Q[249]), .B1(n571), .B2(Q[153]), .ZN(n211) );
  AOI22_X1 U225 ( .A1(n574), .A2(Q[89]), .B1(n573), .B2(Q[185]), .ZN(n212) );
  AOI22_X1 U226 ( .A1(n576), .A2(Q[217]), .B1(n575), .B2(Q[57]), .ZN(n213) );
  NAND4_X1 U227 ( .A1(n210), .A2(n211), .A3(n212), .A4(n213), .ZN(n214) );
  AOI22_X1 U228 ( .A1(n547), .A2(Q[1017]), .B1(n546), .B2(Q[953]), .ZN(n215)
         );
  AOI22_X1 U229 ( .A1(n549), .A2(Q[985]), .B1(n548), .B2(Q[921]), .ZN(n216) );
  AOI222_X1 U230 ( .A1(n551), .A2(Q[825]), .B1(n552), .B2(Q[121]), .C1(n550), 
        .C2(Q[761]), .ZN(n217) );
  NAND3_X1 U231 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n218) );
  AOI22_X1 U232 ( .A1(n554), .A2(Q[857]), .B1(n553), .B2(Q[729]), .ZN(n219) );
  AOI22_X1 U233 ( .A1(n556), .A2(Q[793]), .B1(n555), .B2(Q[889]), .ZN(n220) );
  NAND4_X1 U234 ( .A1(n628), .A2(n629), .A3(n219), .A4(n220), .ZN(n221) );
  OR4_X1 U235 ( .A1(n209), .A2(n214), .A3(n218), .A4(n221), .ZN(Y[25]) );
  AOI22_X1 U236 ( .A1(n562), .A2(Q[504]), .B1(n561), .B2(Q[568]), .ZN(n222) );
  AOI22_X1 U237 ( .A1(n564), .A2(Q[664]), .B1(n563), .B2(Q[472]), .ZN(n223) );
  AOI22_X1 U238 ( .A1(n566), .A2(Q[376]), .B1(n565), .B2(Q[312]), .ZN(n224) );
  AOI22_X1 U239 ( .A1(n568), .A2(Q[408]), .B1(n567), .B2(Q[280]), .ZN(n225) );
  NAND4_X1 U240 ( .A1(n222), .A2(n223), .A3(n224), .A4(n225), .ZN(n226) );
  AOI22_X1 U241 ( .A1(n570), .A2(Q[344]), .B1(n569), .B2(Q[440]), .ZN(n227) );
  AOI22_X1 U242 ( .A1(n572), .A2(Q[248]), .B1(n571), .B2(Q[152]), .ZN(n228) );
  AOI22_X1 U243 ( .A1(n574), .A2(Q[88]), .B1(n573), .B2(Q[184]), .ZN(n229) );
  AOI22_X1 U244 ( .A1(n576), .A2(Q[216]), .B1(n575), .B2(Q[56]), .ZN(n230) );
  NAND4_X1 U245 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(n231) );
  AOI22_X1 U246 ( .A1(n547), .A2(Q[1016]), .B1(n546), .B2(Q[952]), .ZN(n232)
         );
  AOI22_X1 U247 ( .A1(n549), .A2(Q[984]), .B1(n548), .B2(Q[920]), .ZN(n233) );
  AOI222_X1 U248 ( .A1(n551), .A2(Q[824]), .B1(n552), .B2(Q[120]), .C1(n550), 
        .C2(Q[760]), .ZN(n234) );
  NAND3_X1 U249 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n235) );
  AOI22_X1 U250 ( .A1(n554), .A2(Q[856]), .B1(n553), .B2(Q[728]), .ZN(n236) );
  AOI22_X1 U251 ( .A1(n556), .A2(Q[792]), .B1(n555), .B2(Q[888]), .ZN(n237) );
  NAND4_X1 U252 ( .A1(n626), .A2(n627), .A3(n236), .A4(n237), .ZN(n238) );
  OR4_X1 U253 ( .A1(n226), .A2(n231), .A3(n235), .A4(n238), .ZN(Y[24]) );
  AOI22_X1 U254 ( .A1(n562), .A2(Q[503]), .B1(n561), .B2(Q[567]), .ZN(n239) );
  AOI22_X1 U255 ( .A1(n564), .A2(Q[663]), .B1(n563), .B2(Q[471]), .ZN(n240) );
  AOI22_X1 U256 ( .A1(n566), .A2(Q[375]), .B1(n565), .B2(Q[311]), .ZN(n241) );
  AOI22_X1 U257 ( .A1(n568), .A2(Q[407]), .B1(n567), .B2(Q[279]), .ZN(n242) );
  NAND4_X1 U258 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(n243) );
  AOI22_X1 U259 ( .A1(n570), .A2(Q[343]), .B1(n569), .B2(Q[439]), .ZN(n244) );
  AOI22_X1 U260 ( .A1(n572), .A2(Q[247]), .B1(n571), .B2(Q[151]), .ZN(n245) );
  AOI22_X1 U261 ( .A1(n574), .A2(Q[87]), .B1(n573), .B2(Q[183]), .ZN(n246) );
  AOI22_X1 U262 ( .A1(n576), .A2(Q[215]), .B1(n575), .B2(Q[55]), .ZN(n247) );
  NAND4_X1 U263 ( .A1(n244), .A2(n245), .A3(n246), .A4(n247), .ZN(n248) );
  AOI22_X1 U264 ( .A1(n547), .A2(Q[1015]), .B1(n546), .B2(Q[951]), .ZN(n249)
         );
  AOI22_X1 U265 ( .A1(n549), .A2(Q[983]), .B1(n548), .B2(Q[919]), .ZN(n250) );
  AOI222_X1 U266 ( .A1(n551), .A2(Q[823]), .B1(n552), .B2(Q[119]), .C1(n550), 
        .C2(Q[759]), .ZN(n251) );
  NAND3_X1 U267 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n252) );
  AOI22_X1 U268 ( .A1(n554), .A2(Q[855]), .B1(n553), .B2(Q[727]), .ZN(n253) );
  AOI22_X1 U269 ( .A1(n556), .A2(Q[791]), .B1(n555), .B2(Q[887]), .ZN(n254) );
  NAND4_X1 U270 ( .A1(n624), .A2(n625), .A3(n253), .A4(n254), .ZN(n255) );
  OR4_X1 U271 ( .A1(n243), .A2(n248), .A3(n252), .A4(n255), .ZN(Y[23]) );
  AOI22_X1 U272 ( .A1(n562), .A2(Q[502]), .B1(n561), .B2(Q[566]), .ZN(n256) );
  AOI22_X1 U273 ( .A1(n564), .A2(Q[662]), .B1(n563), .B2(Q[470]), .ZN(n257) );
  AOI22_X1 U274 ( .A1(n566), .A2(Q[374]), .B1(n565), .B2(Q[310]), .ZN(n258) );
  AOI22_X1 U275 ( .A1(n568), .A2(Q[406]), .B1(n567), .B2(Q[278]), .ZN(n259) );
  NAND4_X1 U276 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(n260) );
  AOI22_X1 U277 ( .A1(n570), .A2(Q[342]), .B1(n569), .B2(Q[438]), .ZN(n261) );
  AOI22_X1 U278 ( .A1(n572), .A2(Q[246]), .B1(n571), .B2(Q[150]), .ZN(n262) );
  AOI22_X1 U279 ( .A1(n574), .A2(Q[86]), .B1(n573), .B2(Q[182]), .ZN(n263) );
  AOI22_X1 U280 ( .A1(n576), .A2(Q[214]), .B1(n575), .B2(Q[54]), .ZN(n264) );
  NAND4_X1 U281 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(n265) );
  AOI22_X1 U282 ( .A1(n547), .A2(Q[1014]), .B1(n546), .B2(Q[950]), .ZN(n266)
         );
  AOI22_X1 U283 ( .A1(n549), .A2(Q[982]), .B1(n548), .B2(Q[918]), .ZN(n267) );
  AOI222_X1 U284 ( .A1(n551), .A2(Q[822]), .B1(n552), .B2(Q[118]), .C1(n550), 
        .C2(Q[758]), .ZN(n268) );
  NAND3_X1 U285 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n269) );
  AOI22_X1 U286 ( .A1(n554), .A2(Q[854]), .B1(n553), .B2(Q[726]), .ZN(n270) );
  AOI22_X1 U287 ( .A1(n556), .A2(Q[790]), .B1(n555), .B2(Q[886]), .ZN(n271) );
  NAND4_X1 U288 ( .A1(n622), .A2(n623), .A3(n270), .A4(n271), .ZN(n272) );
  OR4_X1 U289 ( .A1(n260), .A2(n265), .A3(n269), .A4(n272), .ZN(Y[22]) );
  AOI22_X1 U290 ( .A1(n562), .A2(Q[501]), .B1(n561), .B2(Q[565]), .ZN(n273) );
  AOI22_X1 U291 ( .A1(n564), .A2(Q[661]), .B1(n563), .B2(Q[469]), .ZN(n274) );
  AOI22_X1 U292 ( .A1(n566), .A2(Q[373]), .B1(n565), .B2(Q[309]), .ZN(n275) );
  AOI22_X1 U293 ( .A1(n568), .A2(Q[405]), .B1(n567), .B2(Q[277]), .ZN(n276) );
  NAND4_X1 U294 ( .A1(n273), .A2(n274), .A3(n275), .A4(n276), .ZN(n277) );
  AOI22_X1 U295 ( .A1(n570), .A2(Q[341]), .B1(n569), .B2(Q[437]), .ZN(n278) );
  AOI22_X1 U296 ( .A1(n572), .A2(Q[245]), .B1(n571), .B2(Q[149]), .ZN(n279) );
  AOI22_X1 U297 ( .A1(n574), .A2(Q[85]), .B1(n573), .B2(Q[181]), .ZN(n280) );
  AOI22_X1 U298 ( .A1(n576), .A2(Q[213]), .B1(n575), .B2(Q[53]), .ZN(n281) );
  NAND4_X1 U299 ( .A1(n278), .A2(n279), .A3(n280), .A4(n281), .ZN(n282) );
  AOI22_X1 U300 ( .A1(n547), .A2(Q[1013]), .B1(n546), .B2(Q[949]), .ZN(n283)
         );
  AOI22_X1 U301 ( .A1(n549), .A2(Q[981]), .B1(n548), .B2(Q[917]), .ZN(n284) );
  AOI222_X1 U302 ( .A1(n551), .A2(Q[821]), .B1(n552), .B2(Q[117]), .C1(n550), 
        .C2(Q[757]), .ZN(n285) );
  NAND3_X1 U303 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n286) );
  AOI22_X1 U304 ( .A1(n554), .A2(Q[853]), .B1(n553), .B2(Q[725]), .ZN(n287) );
  AOI22_X1 U305 ( .A1(n556), .A2(Q[789]), .B1(n555), .B2(Q[885]), .ZN(n288) );
  NAND4_X1 U306 ( .A1(n620), .A2(n621), .A3(n287), .A4(n288), .ZN(n289) );
  OR4_X1 U307 ( .A1(n277), .A2(n282), .A3(n286), .A4(n289), .ZN(Y[21]) );
  AOI22_X1 U308 ( .A1(n562), .A2(Q[500]), .B1(n561), .B2(Q[564]), .ZN(n290) );
  AOI22_X1 U309 ( .A1(n564), .A2(Q[660]), .B1(n563), .B2(Q[468]), .ZN(n291) );
  AOI22_X1 U310 ( .A1(n566), .A2(Q[372]), .B1(n565), .B2(Q[308]), .ZN(n292) );
  AOI22_X1 U311 ( .A1(n568), .A2(Q[404]), .B1(n567), .B2(Q[276]), .ZN(n293) );
  NAND4_X1 U312 ( .A1(n290), .A2(n291), .A3(n292), .A4(n293), .ZN(n294) );
  AOI22_X1 U313 ( .A1(n570), .A2(Q[340]), .B1(n569), .B2(Q[436]), .ZN(n295) );
  AOI22_X1 U314 ( .A1(n572), .A2(Q[244]), .B1(n571), .B2(Q[148]), .ZN(n296) );
  AOI22_X1 U315 ( .A1(n574), .A2(Q[84]), .B1(n573), .B2(Q[180]), .ZN(n297) );
  AOI22_X1 U316 ( .A1(n576), .A2(Q[212]), .B1(n575), .B2(Q[52]), .ZN(n298) );
  NAND4_X1 U317 ( .A1(n295), .A2(n296), .A3(n297), .A4(n298), .ZN(n299) );
  AOI22_X1 U318 ( .A1(n547), .A2(Q[1012]), .B1(n546), .B2(Q[948]), .ZN(n300)
         );
  AOI22_X1 U319 ( .A1(n549), .A2(Q[980]), .B1(n548), .B2(Q[916]), .ZN(n301) );
  AOI222_X1 U320 ( .A1(n551), .A2(Q[820]), .B1(n552), .B2(Q[116]), .C1(n550), 
        .C2(Q[756]), .ZN(n302) );
  NAND3_X1 U321 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n303) );
  AOI22_X1 U322 ( .A1(n554), .A2(Q[852]), .B1(n553), .B2(Q[724]), .ZN(n304) );
  AOI22_X1 U323 ( .A1(n556), .A2(Q[788]), .B1(n555), .B2(Q[884]), .ZN(n305) );
  NAND4_X1 U324 ( .A1(n618), .A2(n619), .A3(n304), .A4(n305), .ZN(n306) );
  OR4_X1 U325 ( .A1(n294), .A2(n299), .A3(n303), .A4(n306), .ZN(Y[20]) );
  AOI22_X1 U326 ( .A1(n674), .A2(Q[491]), .B1(n673), .B2(Q[555]), .ZN(n307) );
  AOI22_X1 U327 ( .A1(n676), .A2(Q[651]), .B1(n675), .B2(Q[459]), .ZN(n308) );
  AOI22_X1 U328 ( .A1(n678), .A2(Q[363]), .B1(n677), .B2(Q[299]), .ZN(n309) );
  AOI22_X1 U329 ( .A1(n680), .A2(Q[395]), .B1(n679), .B2(Q[267]), .ZN(n310) );
  NAND4_X1 U330 ( .A1(n307), .A2(n308), .A3(n309), .A4(n310), .ZN(n311) );
  AOI22_X1 U331 ( .A1(n682), .A2(Q[331]), .B1(n681), .B2(Q[427]), .ZN(n312) );
  AOI22_X1 U332 ( .A1(n684), .A2(Q[235]), .B1(n683), .B2(Q[139]), .ZN(n313) );
  AOI22_X1 U333 ( .A1(n686), .A2(Q[75]), .B1(n685), .B2(Q[171]), .ZN(n314) );
  AOI22_X1 U334 ( .A1(n688), .A2(Q[203]), .B1(n687), .B2(Q[43]), .ZN(n315) );
  NAND4_X1 U335 ( .A1(n312), .A2(n313), .A3(n314), .A4(n315), .ZN(n316) );
  AOI22_X1 U336 ( .A1(n657), .A2(Q[1003]), .B1(n656), .B2(Q[939]), .ZN(n317)
         );
  AOI22_X1 U337 ( .A1(n659), .A2(Q[971]), .B1(n658), .B2(Q[907]), .ZN(n318) );
  AOI222_X1 U338 ( .A1(n661), .A2(Q[811]), .B1(n662), .B2(Q[107]), .C1(n660), 
        .C2(Q[747]), .ZN(n319) );
  NAND3_X1 U339 ( .A1(n317), .A2(n318), .A3(n319), .ZN(n320) );
  AOI22_X1 U340 ( .A1(n664), .A2(Q[843]), .B1(n663), .B2(Q[715]), .ZN(n321) );
  AOI22_X1 U341 ( .A1(n666), .A2(Q[779]), .B1(n665), .B2(Q[875]), .ZN(n322) );
  NAND4_X1 U342 ( .A1(n598), .A2(n599), .A3(n321), .A4(n322), .ZN(n323) );
  OR4_X1 U343 ( .A1(n311), .A2(n316), .A3(n320), .A4(n323), .ZN(Y[11]) );
  AOI22_X1 U344 ( .A1(n562), .A2(Q[490]), .B1(n561), .B2(Q[554]), .ZN(n324) );
  AOI22_X1 U345 ( .A1(n564), .A2(Q[650]), .B1(n563), .B2(Q[458]), .ZN(n325) );
  AOI22_X1 U346 ( .A1(n566), .A2(Q[362]), .B1(n565), .B2(Q[298]), .ZN(n326) );
  AOI22_X1 U347 ( .A1(n568), .A2(Q[394]), .B1(n567), .B2(Q[266]), .ZN(n327) );
  NAND4_X1 U348 ( .A1(n324), .A2(n325), .A3(n326), .A4(n327), .ZN(n328) );
  AOI22_X1 U349 ( .A1(n570), .A2(Q[330]), .B1(n569), .B2(Q[426]), .ZN(n329) );
  AOI22_X1 U350 ( .A1(n572), .A2(Q[234]), .B1(n571), .B2(Q[138]), .ZN(n330) );
  AOI22_X1 U351 ( .A1(n574), .A2(Q[74]), .B1(n573), .B2(Q[170]), .ZN(n331) );
  AOI22_X1 U352 ( .A1(n576), .A2(Q[202]), .B1(n575), .B2(Q[42]), .ZN(n332) );
  NAND4_X1 U353 ( .A1(n329), .A2(n330), .A3(n331), .A4(n332), .ZN(n333) );
  AOI22_X1 U354 ( .A1(n547), .A2(Q[1002]), .B1(n546), .B2(Q[938]), .ZN(n334)
         );
  AOI22_X1 U355 ( .A1(n549), .A2(Q[970]), .B1(n548), .B2(Q[906]), .ZN(n335) );
  AOI222_X1 U356 ( .A1(n551), .A2(Q[810]), .B1(n552), .B2(Q[106]), .C1(n550), 
        .C2(Q[746]), .ZN(n336) );
  NAND3_X1 U357 ( .A1(n334), .A2(n335), .A3(n336), .ZN(n337) );
  AOI22_X1 U358 ( .A1(n554), .A2(Q[842]), .B1(n553), .B2(Q[714]), .ZN(n338) );
  AOI22_X1 U359 ( .A1(n556), .A2(Q[778]), .B1(n555), .B2(Q[874]), .ZN(n339) );
  NAND4_X1 U360 ( .A1(n596), .A2(n597), .A3(n338), .A4(n339), .ZN(n340) );
  OR4_X1 U361 ( .A1(n328), .A2(n333), .A3(n337), .A4(n340), .ZN(Y[10]) );
  AOI22_X1 U362 ( .A1(n562), .A2(Q[489]), .B1(n561), .B2(Q[553]), .ZN(n341) );
  AOI22_X1 U363 ( .A1(n564), .A2(Q[649]), .B1(n563), .B2(Q[457]), .ZN(n342) );
  AOI22_X1 U364 ( .A1(n566), .A2(Q[361]), .B1(n565), .B2(Q[297]), .ZN(n343) );
  AOI22_X1 U365 ( .A1(n568), .A2(Q[393]), .B1(n567), .B2(Q[265]), .ZN(n344) );
  NAND4_X1 U366 ( .A1(n341), .A2(n342), .A3(n343), .A4(n344), .ZN(n345) );
  AOI22_X1 U367 ( .A1(n570), .A2(Q[329]), .B1(n569), .B2(Q[425]), .ZN(n346) );
  AOI22_X1 U368 ( .A1(n572), .A2(Q[233]), .B1(n571), .B2(Q[137]), .ZN(n347) );
  AOI22_X1 U369 ( .A1(n574), .A2(Q[73]), .B1(n573), .B2(Q[169]), .ZN(n348) );
  AOI22_X1 U370 ( .A1(n576), .A2(Q[201]), .B1(n575), .B2(Q[41]), .ZN(n349) );
  NAND4_X1 U371 ( .A1(n346), .A2(n347), .A3(n348), .A4(n349), .ZN(n350) );
  AOI22_X1 U372 ( .A1(n547), .A2(Q[1001]), .B1(n546), .B2(Q[937]), .ZN(n351)
         );
  AOI22_X1 U373 ( .A1(n549), .A2(Q[969]), .B1(n548), .B2(Q[905]), .ZN(n352) );
  AOI222_X1 U374 ( .A1(n551), .A2(Q[809]), .B1(n552), .B2(Q[105]), .C1(n550), 
        .C2(Q[745]), .ZN(n353) );
  NAND3_X1 U375 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n354) );
  AOI22_X1 U376 ( .A1(n554), .A2(Q[841]), .B1(n553), .B2(Q[713]), .ZN(n355) );
  AOI22_X1 U377 ( .A1(n556), .A2(Q[777]), .B1(n555), .B2(Q[873]), .ZN(n356) );
  NAND4_X1 U378 ( .A1(n671), .A2(n672), .A3(n355), .A4(n356), .ZN(n357) );
  OR4_X1 U379 ( .A1(n345), .A2(n350), .A3(n354), .A4(n357), .ZN(Y[9]) );
  AOI22_X1 U380 ( .A1(n562), .A2(Q[488]), .B1(n561), .B2(Q[552]), .ZN(n358) );
  AOI22_X1 U381 ( .A1(n564), .A2(Q[648]), .B1(n563), .B2(Q[456]), .ZN(n359) );
  AOI22_X1 U382 ( .A1(n566), .A2(Q[360]), .B1(n565), .B2(Q[296]), .ZN(n360) );
  AOI22_X1 U383 ( .A1(n568), .A2(Q[392]), .B1(n567), .B2(Q[264]), .ZN(n361) );
  NAND4_X1 U384 ( .A1(n358), .A2(n359), .A3(n360), .A4(n361), .ZN(n362) );
  AOI22_X1 U385 ( .A1(n570), .A2(Q[328]), .B1(n569), .B2(Q[424]), .ZN(n363) );
  AOI22_X1 U386 ( .A1(n572), .A2(Q[232]), .B1(n571), .B2(Q[136]), .ZN(n364) );
  AOI22_X1 U387 ( .A1(n574), .A2(Q[72]), .B1(n573), .B2(Q[168]), .ZN(n365) );
  AOI22_X1 U388 ( .A1(n576), .A2(Q[200]), .B1(n575), .B2(Q[40]), .ZN(n366) );
  NAND4_X1 U389 ( .A1(n363), .A2(n364), .A3(n365), .A4(n366), .ZN(n367) );
  AOI22_X1 U390 ( .A1(n547), .A2(Q[1000]), .B1(n546), .B2(Q[936]), .ZN(n368)
         );
  AOI22_X1 U391 ( .A1(n549), .A2(Q[968]), .B1(n548), .B2(Q[904]), .ZN(n369) );
  AOI222_X1 U392 ( .A1(n551), .A2(Q[808]), .B1(n552), .B2(Q[104]), .C1(n550), 
        .C2(Q[744]), .ZN(n370) );
  NAND3_X1 U393 ( .A1(n368), .A2(n369), .A3(n370), .ZN(n371) );
  AOI22_X1 U394 ( .A1(n554), .A2(Q[840]), .B1(n553), .B2(Q[712]), .ZN(n372) );
  AOI22_X1 U395 ( .A1(n556), .A2(Q[776]), .B1(n555), .B2(Q[872]), .ZN(n373) );
  NAND4_X1 U396 ( .A1(n654), .A2(n655), .A3(n372), .A4(n373), .ZN(n374) );
  OR4_X1 U397 ( .A1(n362), .A2(n367), .A3(n371), .A4(n374), .ZN(Y[8]) );
  AOI22_X1 U398 ( .A1(n562), .A2(Q[487]), .B1(n561), .B2(Q[551]), .ZN(n375) );
  AOI22_X1 U399 ( .A1(n564), .A2(Q[647]), .B1(n563), .B2(Q[455]), .ZN(n376) );
  AOI22_X1 U400 ( .A1(n566), .A2(Q[359]), .B1(n565), .B2(Q[295]), .ZN(n377) );
  AOI22_X1 U401 ( .A1(n568), .A2(Q[391]), .B1(n567), .B2(Q[263]), .ZN(n378) );
  NAND4_X1 U402 ( .A1(n375), .A2(n376), .A3(n377), .A4(n378), .ZN(n379) );
  AOI22_X1 U403 ( .A1(n570), .A2(Q[327]), .B1(n569), .B2(Q[423]), .ZN(n380) );
  AOI22_X1 U404 ( .A1(n572), .A2(Q[231]), .B1(n571), .B2(Q[135]), .ZN(n381) );
  AOI22_X1 U405 ( .A1(n574), .A2(Q[71]), .B1(n573), .B2(Q[167]), .ZN(n382) );
  AOI22_X1 U406 ( .A1(n576), .A2(Q[199]), .B1(n575), .B2(Q[39]), .ZN(n383) );
  NAND4_X1 U407 ( .A1(n380), .A2(n381), .A3(n382), .A4(n383), .ZN(n384) );
  AOI22_X1 U408 ( .A1(n547), .A2(Q[999]), .B1(n546), .B2(Q[935]), .ZN(n385) );
  AOI22_X1 U409 ( .A1(n549), .A2(Q[967]), .B1(n548), .B2(Q[903]), .ZN(n386) );
  AOI222_X1 U410 ( .A1(n551), .A2(Q[807]), .B1(n552), .B2(Q[103]), .C1(n550), 
        .C2(Q[743]), .ZN(n387) );
  NAND3_X1 U411 ( .A1(n385), .A2(n386), .A3(n387), .ZN(n388) );
  AOI22_X1 U412 ( .A1(n554), .A2(Q[839]), .B1(n553), .B2(Q[711]), .ZN(n389) );
  AOI22_X1 U413 ( .A1(n556), .A2(Q[775]), .B1(n555), .B2(Q[871]), .ZN(n390) );
  NAND4_X1 U414 ( .A1(n652), .A2(n653), .A3(n389), .A4(n390), .ZN(n391) );
  OR4_X1 U415 ( .A1(n379), .A2(n384), .A3(n388), .A4(n391), .ZN(Y[7]) );
  AOI22_X1 U416 ( .A1(n562), .A2(Q[486]), .B1(n561), .B2(Q[550]), .ZN(n392) );
  AOI22_X1 U417 ( .A1(n564), .A2(Q[646]), .B1(n563), .B2(Q[454]), .ZN(n393) );
  AOI22_X1 U418 ( .A1(n566), .A2(Q[358]), .B1(n565), .B2(Q[294]), .ZN(n394) );
  AOI22_X1 U419 ( .A1(n568), .A2(Q[390]), .B1(n567), .B2(Q[262]), .ZN(n395) );
  NAND4_X1 U420 ( .A1(n392), .A2(n393), .A3(n394), .A4(n395), .ZN(n396) );
  AOI22_X1 U421 ( .A1(n570), .A2(Q[326]), .B1(n569), .B2(Q[422]), .ZN(n397) );
  AOI22_X1 U422 ( .A1(n572), .A2(Q[230]), .B1(n571), .B2(Q[134]), .ZN(n398) );
  AOI22_X1 U423 ( .A1(n574), .A2(Q[70]), .B1(n573), .B2(Q[166]), .ZN(n399) );
  AOI22_X1 U424 ( .A1(n576), .A2(Q[198]), .B1(n575), .B2(Q[38]), .ZN(n400) );
  NAND4_X1 U425 ( .A1(n397), .A2(n398), .A3(n399), .A4(n400), .ZN(n401) );
  AOI22_X1 U426 ( .A1(n547), .A2(Q[998]), .B1(n546), .B2(Q[934]), .ZN(n402) );
  AOI22_X1 U427 ( .A1(n549), .A2(Q[966]), .B1(n548), .B2(Q[902]), .ZN(n403) );
  AOI222_X1 U428 ( .A1(n551), .A2(Q[806]), .B1(n552), .B2(Q[102]), .C1(n550), 
        .C2(Q[742]), .ZN(n404) );
  NAND3_X1 U429 ( .A1(n402), .A2(n403), .A3(n404), .ZN(n405) );
  AOI22_X1 U430 ( .A1(n554), .A2(Q[838]), .B1(n553), .B2(Q[710]), .ZN(n406) );
  AOI22_X1 U431 ( .A1(n556), .A2(Q[774]), .B1(n555), .B2(Q[870]), .ZN(n407) );
  NAND4_X1 U432 ( .A1(n650), .A2(n651), .A3(n406), .A4(n407), .ZN(n408) );
  OR4_X1 U433 ( .A1(n396), .A2(n401), .A3(n405), .A4(n408), .ZN(Y[6]) );
  AOI22_X1 U434 ( .A1(n562), .A2(Q[485]), .B1(n561), .B2(Q[549]), .ZN(n409) );
  AOI22_X1 U435 ( .A1(n564), .A2(Q[645]), .B1(n563), .B2(Q[453]), .ZN(n410) );
  AOI22_X1 U436 ( .A1(n566), .A2(Q[357]), .B1(n565), .B2(Q[293]), .ZN(n411) );
  AOI22_X1 U437 ( .A1(n568), .A2(Q[389]), .B1(n567), .B2(Q[261]), .ZN(n412) );
  NAND4_X1 U438 ( .A1(n409), .A2(n410), .A3(n411), .A4(n412), .ZN(n413) );
  AOI22_X1 U439 ( .A1(n570), .A2(Q[325]), .B1(n569), .B2(Q[421]), .ZN(n414) );
  AOI22_X1 U440 ( .A1(n572), .A2(Q[229]), .B1(n571), .B2(Q[133]), .ZN(n415) );
  AOI22_X1 U441 ( .A1(n574), .A2(Q[69]), .B1(n573), .B2(Q[165]), .ZN(n416) );
  AOI22_X1 U442 ( .A1(n576), .A2(Q[197]), .B1(n575), .B2(Q[37]), .ZN(n417) );
  NAND4_X1 U443 ( .A1(n414), .A2(n415), .A3(n416), .A4(n417), .ZN(n418) );
  AOI22_X1 U444 ( .A1(n547), .A2(Q[997]), .B1(n546), .B2(Q[933]), .ZN(n419) );
  AOI22_X1 U445 ( .A1(n549), .A2(Q[965]), .B1(n548), .B2(Q[901]), .ZN(n420) );
  AOI222_X1 U446 ( .A1(n551), .A2(Q[805]), .B1(n552), .B2(Q[101]), .C1(n550), 
        .C2(Q[741]), .ZN(n421) );
  NAND3_X1 U447 ( .A1(n419), .A2(n420), .A3(n421), .ZN(n422) );
  AOI22_X1 U448 ( .A1(n554), .A2(Q[837]), .B1(n553), .B2(Q[709]), .ZN(n423) );
  AOI22_X1 U449 ( .A1(n556), .A2(Q[773]), .B1(n555), .B2(Q[869]), .ZN(n424) );
  NAND4_X1 U450 ( .A1(n648), .A2(n649), .A3(n423), .A4(n424), .ZN(n425) );
  OR4_X1 U451 ( .A1(n413), .A2(n418), .A3(n422), .A4(n425), .ZN(Y[5]) );
  AOI22_X1 U452 ( .A1(n562), .A2(Q[484]), .B1(n561), .B2(Q[548]), .ZN(n426) );
  AOI22_X1 U453 ( .A1(n564), .A2(Q[644]), .B1(n563), .B2(Q[452]), .ZN(n427) );
  AOI22_X1 U454 ( .A1(n566), .A2(Q[356]), .B1(n565), .B2(Q[292]), .ZN(n428) );
  AOI22_X1 U455 ( .A1(n568), .A2(Q[388]), .B1(n567), .B2(Q[260]), .ZN(n429) );
  NAND4_X1 U456 ( .A1(n426), .A2(n427), .A3(n428), .A4(n429), .ZN(n430) );
  AOI22_X1 U457 ( .A1(n570), .A2(Q[324]), .B1(n569), .B2(Q[420]), .ZN(n431) );
  AOI22_X1 U458 ( .A1(n572), .A2(Q[228]), .B1(n571), .B2(Q[132]), .ZN(n432) );
  AOI22_X1 U459 ( .A1(n574), .A2(Q[68]), .B1(n573), .B2(Q[164]), .ZN(n433) );
  AOI22_X1 U460 ( .A1(n576), .A2(Q[196]), .B1(n575), .B2(Q[36]), .ZN(n434) );
  NAND4_X1 U461 ( .A1(n431), .A2(n432), .A3(n433), .A4(n434), .ZN(n435) );
  AOI22_X1 U462 ( .A1(n547), .A2(Q[996]), .B1(n546), .B2(Q[932]), .ZN(n436) );
  AOI22_X1 U463 ( .A1(n549), .A2(Q[964]), .B1(n548), .B2(Q[900]), .ZN(n437) );
  AOI222_X1 U464 ( .A1(n551), .A2(Q[804]), .B1(n552), .B2(Q[100]), .C1(n550), 
        .C2(Q[740]), .ZN(n438) );
  NAND3_X1 U465 ( .A1(n436), .A2(n437), .A3(n438), .ZN(n439) );
  AOI22_X1 U466 ( .A1(n554), .A2(Q[836]), .B1(n553), .B2(Q[708]), .ZN(n440) );
  AOI22_X1 U467 ( .A1(n556), .A2(Q[772]), .B1(n555), .B2(Q[868]), .ZN(n441) );
  NAND4_X1 U468 ( .A1(n646), .A2(n647), .A3(n440), .A4(n441), .ZN(n442) );
  OR4_X1 U469 ( .A1(n430), .A2(n435), .A3(n439), .A4(n442), .ZN(Y[4]) );
  AOI22_X1 U470 ( .A1(n562), .A2(Q[483]), .B1(n561), .B2(Q[547]), .ZN(n443) );
  AOI22_X1 U471 ( .A1(n564), .A2(Q[643]), .B1(n563), .B2(Q[451]), .ZN(n444) );
  AOI22_X1 U472 ( .A1(n566), .A2(Q[355]), .B1(n565), .B2(Q[291]), .ZN(n445) );
  AOI22_X1 U473 ( .A1(n568), .A2(Q[387]), .B1(n567), .B2(Q[259]), .ZN(n446) );
  NAND4_X1 U474 ( .A1(n443), .A2(n444), .A3(n445), .A4(n446), .ZN(n447) );
  AOI22_X1 U475 ( .A1(n570), .A2(Q[323]), .B1(n569), .B2(Q[419]), .ZN(n448) );
  AOI22_X1 U476 ( .A1(n572), .A2(Q[227]), .B1(n571), .B2(Q[131]), .ZN(n449) );
  AOI22_X1 U477 ( .A1(n574), .A2(Q[67]), .B1(n573), .B2(Q[163]), .ZN(n450) );
  AOI22_X1 U478 ( .A1(n576), .A2(Q[195]), .B1(n575), .B2(Q[35]), .ZN(n451) );
  NAND4_X1 U479 ( .A1(n448), .A2(n449), .A3(n450), .A4(n451), .ZN(n452) );
  AOI22_X1 U480 ( .A1(n547), .A2(Q[995]), .B1(n546), .B2(Q[931]), .ZN(n453) );
  AOI22_X1 U481 ( .A1(n549), .A2(Q[963]), .B1(n548), .B2(Q[899]), .ZN(n454) );
  AOI222_X1 U482 ( .A1(n551), .A2(Q[803]), .B1(n552), .B2(Q[99]), .C1(n550), 
        .C2(Q[739]), .ZN(n455) );
  NAND3_X1 U483 ( .A1(n453), .A2(n454), .A3(n455), .ZN(n456) );
  AOI22_X1 U484 ( .A1(n554), .A2(Q[835]), .B1(n553), .B2(Q[707]), .ZN(n457) );
  AOI22_X1 U485 ( .A1(n556), .A2(Q[771]), .B1(n555), .B2(Q[867]), .ZN(n458) );
  NAND4_X1 U486 ( .A1(n644), .A2(n645), .A3(n457), .A4(n458), .ZN(n459) );
  OR4_X1 U487 ( .A1(n447), .A2(n452), .A3(n456), .A4(n459), .ZN(Y[3]) );
  AOI22_X1 U488 ( .A1(n562), .A2(Q[482]), .B1(n561), .B2(Q[546]), .ZN(n460) );
  AOI22_X1 U489 ( .A1(n564), .A2(Q[642]), .B1(n563), .B2(Q[450]), .ZN(n461) );
  AOI22_X1 U490 ( .A1(n566), .A2(Q[354]), .B1(n565), .B2(Q[290]), .ZN(n462) );
  AOI22_X1 U491 ( .A1(n568), .A2(Q[386]), .B1(n567), .B2(Q[258]), .ZN(n463) );
  NAND4_X1 U492 ( .A1(n460), .A2(n461), .A3(n462), .A4(n463), .ZN(n464) );
  AOI22_X1 U493 ( .A1(n570), .A2(Q[322]), .B1(n569), .B2(Q[418]), .ZN(n465) );
  AOI22_X1 U494 ( .A1(n572), .A2(Q[226]), .B1(n571), .B2(Q[130]), .ZN(n466) );
  AOI22_X1 U495 ( .A1(n574), .A2(Q[66]), .B1(n573), .B2(Q[162]), .ZN(n467) );
  AOI22_X1 U496 ( .A1(n576), .A2(Q[194]), .B1(n575), .B2(Q[34]), .ZN(n468) );
  NAND4_X1 U497 ( .A1(n465), .A2(n466), .A3(n467), .A4(n468), .ZN(n469) );
  AOI22_X1 U498 ( .A1(n547), .A2(Q[994]), .B1(n546), .B2(Q[930]), .ZN(n470) );
  AOI22_X1 U499 ( .A1(n549), .A2(Q[962]), .B1(n548), .B2(Q[898]), .ZN(n471) );
  AOI222_X1 U500 ( .A1(n551), .A2(Q[802]), .B1(n552), .B2(Q[98]), .C1(n550), 
        .C2(Q[738]), .ZN(n472) );
  NAND3_X1 U501 ( .A1(n470), .A2(n471), .A3(n472), .ZN(n473) );
  AOI22_X1 U502 ( .A1(n554), .A2(Q[834]), .B1(n553), .B2(Q[706]), .ZN(n474) );
  AOI22_X1 U503 ( .A1(n556), .A2(Q[770]), .B1(n555), .B2(Q[866]), .ZN(n475) );
  NAND4_X1 U504 ( .A1(n638), .A2(n639), .A3(n474), .A4(n475), .ZN(n476) );
  OR4_X1 U505 ( .A1(n464), .A2(n469), .A3(n473), .A4(n476), .ZN(Y[2]) );
  AOI22_X1 U506 ( .A1(n562), .A2(Q[481]), .B1(n561), .B2(Q[545]), .ZN(n477) );
  AOI22_X1 U507 ( .A1(n564), .A2(Q[641]), .B1(n563), .B2(Q[449]), .ZN(n478) );
  AOI22_X1 U508 ( .A1(n566), .A2(Q[353]), .B1(n565), .B2(Q[289]), .ZN(n479) );
  AOI22_X1 U509 ( .A1(n568), .A2(Q[385]), .B1(n567), .B2(Q[257]), .ZN(n480) );
  NAND4_X1 U510 ( .A1(n477), .A2(n478), .A3(n479), .A4(n480), .ZN(n481) );
  AOI22_X1 U511 ( .A1(n570), .A2(Q[321]), .B1(n569), .B2(Q[417]), .ZN(n482) );
  AOI22_X1 U512 ( .A1(n572), .A2(Q[225]), .B1(n571), .B2(Q[129]), .ZN(n483) );
  AOI22_X1 U513 ( .A1(n574), .A2(Q[65]), .B1(n573), .B2(Q[161]), .ZN(n484) );
  AOI22_X1 U514 ( .A1(n576), .A2(Q[193]), .B1(n575), .B2(Q[33]), .ZN(n485) );
  NAND4_X1 U515 ( .A1(n482), .A2(n483), .A3(n484), .A4(n485), .ZN(n486) );
  AOI22_X1 U516 ( .A1(n547), .A2(Q[993]), .B1(n546), .B2(Q[929]), .ZN(n487) );
  AOI22_X1 U517 ( .A1(n549), .A2(Q[961]), .B1(n548), .B2(Q[897]), .ZN(n488) );
  AOI222_X1 U518 ( .A1(n551), .A2(Q[801]), .B1(n552), .B2(Q[97]), .C1(n550), 
        .C2(Q[737]), .ZN(n489) );
  NAND3_X1 U519 ( .A1(n487), .A2(n488), .A3(n489), .ZN(n490) );
  AOI22_X1 U520 ( .A1(n554), .A2(Q[833]), .B1(n553), .B2(Q[705]), .ZN(n491) );
  AOI22_X1 U521 ( .A1(n556), .A2(Q[769]), .B1(n555), .B2(Q[865]), .ZN(n492) );
  NAND4_X1 U522 ( .A1(n616), .A2(n617), .A3(n491), .A4(n492), .ZN(n493) );
  OR4_X1 U523 ( .A1(n481), .A2(n486), .A3(n490), .A4(n493), .ZN(Y[1]) );
  AOI22_X1 U524 ( .A1(n562), .A2(Q[480]), .B1(n561), .B2(Q[544]), .ZN(n494) );
  AOI22_X1 U525 ( .A1(n564), .A2(Q[640]), .B1(n563), .B2(Q[448]), .ZN(n495) );
  AOI22_X1 U526 ( .A1(n566), .A2(Q[352]), .B1(n565), .B2(Q[288]), .ZN(n496) );
  AOI22_X1 U527 ( .A1(n568), .A2(Q[384]), .B1(n567), .B2(Q[256]), .ZN(n497) );
  NAND4_X1 U528 ( .A1(n494), .A2(n495), .A3(n496), .A4(n497), .ZN(n498) );
  AOI22_X1 U529 ( .A1(n570), .A2(Q[320]), .B1(n569), .B2(Q[416]), .ZN(n499) );
  AOI22_X1 U530 ( .A1(n572), .A2(Q[224]), .B1(n571), .B2(Q[128]), .ZN(n500) );
  AOI22_X1 U531 ( .A1(n574), .A2(Q[64]), .B1(n573), .B2(Q[160]), .ZN(n501) );
  AOI22_X1 U532 ( .A1(n576), .A2(Q[192]), .B1(n575), .B2(Q[32]), .ZN(n502) );
  NAND4_X1 U533 ( .A1(n499), .A2(n500), .A3(n501), .A4(n502), .ZN(n503) );
  AOI22_X1 U534 ( .A1(n547), .A2(Q[992]), .B1(n546), .B2(Q[928]), .ZN(n504) );
  AOI22_X1 U535 ( .A1(n549), .A2(Q[960]), .B1(n548), .B2(Q[896]), .ZN(n505) );
  AOI222_X1 U536 ( .A1(n551), .A2(Q[800]), .B1(n552), .B2(Q[96]), .C1(n550), 
        .C2(Q[736]), .ZN(n506) );
  NAND3_X1 U537 ( .A1(n504), .A2(n505), .A3(n506), .ZN(n507) );
  AOI22_X1 U538 ( .A1(n554), .A2(Q[832]), .B1(n553), .B2(Q[704]), .ZN(n508) );
  AOI22_X1 U539 ( .A1(n556), .A2(Q[768]), .B1(n555), .B2(Q[864]), .ZN(n509) );
  NAND4_X1 U540 ( .A1(n581), .A2(n582), .A3(n508), .A4(n509), .ZN(n510) );
  OR4_X1 U541 ( .A1(n498), .A2(n503), .A3(n507), .A4(n510), .ZN(Y[0]) );
  AOI22_X1 U542 ( .A1(n674), .A2(Q[492]), .B1(n673), .B2(Q[556]), .ZN(n511) );
  AOI22_X1 U543 ( .A1(n676), .A2(Q[652]), .B1(n675), .B2(Q[460]), .ZN(n512) );
  AOI22_X1 U544 ( .A1(n678), .A2(Q[364]), .B1(n677), .B2(Q[300]), .ZN(n513) );
  AOI22_X1 U545 ( .A1(n680), .A2(Q[396]), .B1(n679), .B2(Q[268]), .ZN(n514) );
  NAND4_X1 U546 ( .A1(n511), .A2(n512), .A3(n513), .A4(n514), .ZN(n515) );
  AOI22_X1 U547 ( .A1(n682), .A2(Q[332]), .B1(n681), .B2(Q[428]), .ZN(n516) );
  AOI22_X1 U548 ( .A1(n684), .A2(Q[236]), .B1(n683), .B2(Q[140]), .ZN(n517) );
  AOI22_X1 U549 ( .A1(n686), .A2(Q[76]), .B1(n685), .B2(Q[172]), .ZN(n518) );
  AOI22_X1 U550 ( .A1(n688), .A2(Q[204]), .B1(n687), .B2(Q[44]), .ZN(n519) );
  NAND4_X1 U551 ( .A1(n516), .A2(n517), .A3(n518), .A4(n519), .ZN(n520) );
  AOI22_X1 U552 ( .A1(n657), .A2(Q[1004]), .B1(n656), .B2(Q[940]), .ZN(n521)
         );
  AOI22_X1 U553 ( .A1(n659), .A2(Q[972]), .B1(n658), .B2(Q[908]), .ZN(n522) );
  AOI222_X1 U554 ( .A1(n661), .A2(Q[812]), .B1(n662), .B2(Q[108]), .C1(n660), 
        .C2(Q[748]), .ZN(n523) );
  NAND3_X1 U555 ( .A1(n521), .A2(n522), .A3(n523), .ZN(n524) );
  AOI22_X1 U556 ( .A1(n664), .A2(Q[844]), .B1(n663), .B2(Q[716]), .ZN(n525) );
  AOI22_X1 U557 ( .A1(n666), .A2(Q[780]), .B1(n665), .B2(Q[876]), .ZN(n526) );
  NAND4_X1 U558 ( .A1(n600), .A2(n601), .A3(n525), .A4(n526), .ZN(n527) );
  OR4_X1 U559 ( .A1(n515), .A2(n520), .A3(n524), .A4(n527), .ZN(Y[12]) );
  AOI22_X1 U560 ( .A1(n562), .A2(Q[511]), .B1(n561), .B2(Q[575]), .ZN(n528) );
  AOI22_X1 U561 ( .A1(n564), .A2(Q[671]), .B1(n563), .B2(Q[479]), .ZN(n529) );
  AOI22_X1 U562 ( .A1(n566), .A2(Q[383]), .B1(n565), .B2(Q[319]), .ZN(n530) );
  AOI22_X1 U563 ( .A1(n568), .A2(Q[415]), .B1(n567), .B2(Q[287]), .ZN(n531) );
  NAND4_X1 U564 ( .A1(n528), .A2(n529), .A3(n530), .A4(n531), .ZN(n532) );
  AOI22_X1 U565 ( .A1(n570), .A2(Q[351]), .B1(n569), .B2(Q[447]), .ZN(n533) );
  AOI22_X1 U566 ( .A1(n572), .A2(Q[255]), .B1(n571), .B2(Q[159]), .ZN(n534) );
  AOI22_X1 U567 ( .A1(n574), .A2(Q[95]), .B1(n573), .B2(Q[191]), .ZN(n535) );
  AOI22_X1 U568 ( .A1(n576), .A2(Q[223]), .B1(n575), .B2(Q[63]), .ZN(n536) );
  NAND4_X1 U569 ( .A1(n533), .A2(n534), .A3(n535), .A4(n536), .ZN(n537) );
  AOI22_X1 U570 ( .A1(n547), .A2(Q[1023]), .B1(n546), .B2(Q[959]), .ZN(n538)
         );
  AOI22_X1 U571 ( .A1(n549), .A2(Q[991]), .B1(n548), .B2(Q[927]), .ZN(n539) );
  AOI222_X1 U572 ( .A1(n551), .A2(Q[831]), .B1(n552), .B2(Q[127]), .C1(n550), 
        .C2(Q[767]), .ZN(n540) );
  NAND3_X1 U573 ( .A1(n538), .A2(n539), .A3(n540), .ZN(n541) );
  AOI22_X1 U574 ( .A1(n554), .A2(Q[863]), .B1(n553), .B2(Q[735]), .ZN(n542) );
  AOI22_X1 U575 ( .A1(n556), .A2(Q[799]), .B1(n555), .B2(Q[895]), .ZN(n543) );
  NAND4_X1 U576 ( .A1(n642), .A2(n643), .A3(n542), .A4(n543), .ZN(n544) );
  OR4_X1 U577 ( .A1(n532), .A2(n537), .A3(n541), .A4(n544), .ZN(Y[31]) );
  BUF_X1 U578 ( .A(n687), .Z(n575) );
  BUF_X1 U579 ( .A(n688), .Z(n576) );
  BUF_X1 U580 ( .A(n685), .Z(n573) );
  BUF_X1 U581 ( .A(n686), .Z(n574) );
  BUF_X1 U582 ( .A(n683), .Z(n571) );
  BUF_X1 U583 ( .A(n684), .Z(n572) );
  BUF_X1 U584 ( .A(n681), .Z(n569) );
  BUF_X1 U585 ( .A(n682), .Z(n570) );
  BUF_X1 U586 ( .A(n679), .Z(n567) );
  BUF_X1 U587 ( .A(n680), .Z(n568) );
  BUF_X1 U588 ( .A(n677), .Z(n565) );
  BUF_X1 U589 ( .A(n678), .Z(n566) );
  BUF_X1 U590 ( .A(n675), .Z(n563) );
  BUF_X1 U591 ( .A(n676), .Z(n564) );
  BUF_X1 U592 ( .A(n673), .Z(n561) );
  BUF_X1 U593 ( .A(n674), .Z(n562) );
  BUF_X1 U594 ( .A(n669), .Z(n559) );
  BUF_X1 U595 ( .A(n670), .Z(n560) );
  BUF_X1 U596 ( .A(n667), .Z(n557) );
  BUF_X1 U597 ( .A(n668), .Z(n558) );
  BUF_X1 U598 ( .A(n665), .Z(n555) );
  BUF_X1 U599 ( .A(n666), .Z(n556) );
  BUF_X1 U600 ( .A(n663), .Z(n553) );
  BUF_X1 U601 ( .A(n664), .Z(n554) );
  BUF_X1 U602 ( .A(n662), .Z(n552) );
  BUF_X1 U603 ( .A(n660), .Z(n550) );
  BUF_X1 U604 ( .A(n661), .Z(n551) );
  BUF_X1 U605 ( .A(n658), .Z(n548) );
  BUF_X1 U606 ( .A(n659), .Z(n549) );
  BUF_X1 U607 ( .A(n656), .Z(n546) );
  OR2_X1 U608 ( .A1(n577), .A2(S[1]), .ZN(n591) );
  BUF_X1 U609 ( .A(n657), .Z(n547) );
  NAND2_X1 U610 ( .A1(S[1]), .A2(S[2]), .ZN(n593) );
  NAND3_X1 U611 ( .A1(S[3]), .A2(S[4]), .A3(S[0]), .ZN(n580) );
  NOR2_X1 U612 ( .A1(n593), .A2(n580), .ZN(n657) );
  INV_X1 U613 ( .A(S[2]), .ZN(n577) );
  NOR2_X1 U614 ( .A1(n580), .A2(n591), .ZN(n656) );
  INV_X1 U615 ( .A(S[0]), .ZN(n578) );
  NAND3_X1 U616 ( .A1(S[4]), .A2(S[3]), .A3(n578), .ZN(n579) );
  NOR2_X1 U617 ( .A1(n593), .A2(n579), .ZN(n659) );
  NOR2_X1 U618 ( .A1(n591), .A2(n579), .ZN(n658) );
  OR2_X1 U619 ( .A1(S[1]), .A2(S[2]), .ZN(n594) );
  NOR2_X1 U620 ( .A1(n580), .A2(n594), .ZN(n661) );
  INV_X1 U621 ( .A(S[3]), .ZN(n588) );
  NAND3_X1 U622 ( .A1(S[4]), .A2(S[0]), .A3(n588), .ZN(n584) );
  NOR2_X1 U623 ( .A1(n593), .A2(n584), .ZN(n660) );
  NAND2_X1 U624 ( .A1(S[1]), .A2(n577), .ZN(n590) );
  INV_X1 U625 ( .A(S[4]), .ZN(n583) );
  NAND3_X1 U626 ( .A1(S[0]), .A2(n588), .A3(n583), .ZN(n595) );
  NOR2_X1 U627 ( .A1(n590), .A2(n595), .ZN(n662) );
  NOR2_X1 U628 ( .A1(n590), .A2(n579), .ZN(n664) );
  NAND3_X1 U629 ( .A1(S[4]), .A2(n588), .A3(n578), .ZN(n585) );
  NOR2_X1 U630 ( .A1(n593), .A2(n585), .ZN(n663) );
  NOR2_X1 U631 ( .A1(n579), .A2(n594), .ZN(n666) );
  NOR2_X1 U632 ( .A1(n590), .A2(n580), .ZN(n665) );
  NOR2_X1 U633 ( .A1(n591), .A2(n584), .ZN(n668) );
  NOR2_X1 U634 ( .A1(n590), .A2(n585), .ZN(n667) );
  AOI22_X1 U635 ( .A1(n558), .A2(Q[672]), .B1(n557), .B2(Q[576]), .ZN(n582) );
  NOR2_X1 U636 ( .A1(n594), .A2(n585), .ZN(n670) );
  NOR2_X1 U637 ( .A1(n590), .A2(n584), .ZN(n669) );
  AOI22_X1 U638 ( .A1(n560), .A2(Q[512]), .B1(n559), .B2(Q[608]), .ZN(n581) );
  NAND3_X1 U639 ( .A1(S[3]), .A2(S[0]), .A3(n583), .ZN(n587) );
  NOR2_X1 U640 ( .A1(n593), .A2(n587), .ZN(n674) );
  NOR2_X1 U641 ( .A1(n594), .A2(n584), .ZN(n673) );
  NOR2_X1 U642 ( .A1(n591), .A2(n585), .ZN(n676) );
  NOR2_X1 U643 ( .A1(S[4]), .A2(S[0]), .ZN(n589) );
  NAND2_X1 U644 ( .A1(S[3]), .A2(n589), .ZN(n586) );
  NOR2_X1 U645 ( .A1(n593), .A2(n586), .ZN(n675) );
  NOR2_X1 U646 ( .A1(n590), .A2(n587), .ZN(n678) );
  NOR2_X1 U647 ( .A1(n594), .A2(n587), .ZN(n677) );
  NOR2_X1 U648 ( .A1(n591), .A2(n586), .ZN(n680) );
  NOR2_X1 U649 ( .A1(n594), .A2(n586), .ZN(n679) );
  NOR2_X1 U650 ( .A1(n590), .A2(n586), .ZN(n682) );
  NOR2_X1 U651 ( .A1(n591), .A2(n587), .ZN(n681) );
  NOR2_X1 U652 ( .A1(n595), .A2(n593), .ZN(n684) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n592) );
  NOR2_X1 U654 ( .A1(n591), .A2(n592), .ZN(n683) );
  NOR2_X1 U655 ( .A1(n590), .A2(n592), .ZN(n686) );
  NOR2_X1 U656 ( .A1(n595), .A2(n591), .ZN(n685) );
  NOR2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n688) );
  NOR2_X1 U658 ( .A1(n595), .A2(n594), .ZN(n687) );
  AOI22_X1 U659 ( .A1(n558), .A2(Q[682]), .B1(n557), .B2(Q[586]), .ZN(n597) );
  AOI22_X1 U660 ( .A1(n560), .A2(Q[522]), .B1(n559), .B2(Q[618]), .ZN(n596) );
  AOI22_X1 U661 ( .A1(n668), .A2(Q[683]), .B1(n667), .B2(Q[587]), .ZN(n599) );
  AOI22_X1 U662 ( .A1(n670), .A2(Q[523]), .B1(n669), .B2(Q[619]), .ZN(n598) );
  AOI22_X1 U663 ( .A1(n668), .A2(Q[684]), .B1(n667), .B2(Q[588]), .ZN(n601) );
  AOI22_X1 U664 ( .A1(n670), .A2(Q[524]), .B1(n669), .B2(Q[620]), .ZN(n600) );
  AOI22_X1 U665 ( .A1(n668), .A2(Q[685]), .B1(n667), .B2(Q[589]), .ZN(n603) );
  AOI22_X1 U666 ( .A1(n670), .A2(Q[525]), .B1(n669), .B2(Q[621]), .ZN(n602) );
  AOI22_X1 U667 ( .A1(n668), .A2(Q[686]), .B1(n667), .B2(Q[590]), .ZN(n605) );
  AOI22_X1 U668 ( .A1(n670), .A2(Q[526]), .B1(n669), .B2(Q[622]), .ZN(n604) );
  AOI22_X1 U669 ( .A1(n668), .A2(Q[687]), .B1(n667), .B2(Q[591]), .ZN(n607) );
  AOI22_X1 U670 ( .A1(n670), .A2(Q[527]), .B1(n669), .B2(Q[623]), .ZN(n606) );
  AOI22_X1 U671 ( .A1(n668), .A2(Q[688]), .B1(n667), .B2(Q[592]), .ZN(n609) );
  AOI22_X1 U672 ( .A1(n670), .A2(Q[528]), .B1(n669), .B2(Q[624]), .ZN(n608) );
  AOI22_X1 U673 ( .A1(n668), .A2(Q[689]), .B1(n667), .B2(Q[593]), .ZN(n611) );
  AOI22_X1 U674 ( .A1(n670), .A2(Q[529]), .B1(n669), .B2(Q[625]), .ZN(n610) );
  AOI22_X1 U675 ( .A1(n668), .A2(Q[690]), .B1(n667), .B2(Q[594]), .ZN(n613) );
  AOI22_X1 U676 ( .A1(n670), .A2(Q[530]), .B1(n669), .B2(Q[626]), .ZN(n612) );
  AOI22_X1 U677 ( .A1(n668), .A2(Q[691]), .B1(n667), .B2(Q[595]), .ZN(n615) );
  AOI22_X1 U678 ( .A1(n670), .A2(Q[531]), .B1(n669), .B2(Q[627]), .ZN(n614) );
  AOI22_X1 U679 ( .A1(n558), .A2(Q[673]), .B1(n557), .B2(Q[577]), .ZN(n617) );
  AOI22_X1 U680 ( .A1(n560), .A2(Q[513]), .B1(n559), .B2(Q[609]), .ZN(n616) );
  AOI22_X1 U681 ( .A1(n558), .A2(Q[692]), .B1(n557), .B2(Q[596]), .ZN(n619) );
  AOI22_X1 U682 ( .A1(n560), .A2(Q[532]), .B1(n559), .B2(Q[628]), .ZN(n618) );
  AOI22_X1 U683 ( .A1(n558), .A2(Q[693]), .B1(n557), .B2(Q[597]), .ZN(n621) );
  AOI22_X1 U684 ( .A1(n560), .A2(Q[533]), .B1(n559), .B2(Q[629]), .ZN(n620) );
  AOI22_X1 U685 ( .A1(n558), .A2(Q[694]), .B1(n557), .B2(Q[598]), .ZN(n623) );
  AOI22_X1 U686 ( .A1(n560), .A2(Q[534]), .B1(n559), .B2(Q[630]), .ZN(n622) );
  AOI22_X1 U687 ( .A1(n558), .A2(Q[695]), .B1(n557), .B2(Q[599]), .ZN(n625) );
  AOI22_X1 U688 ( .A1(n560), .A2(Q[535]), .B1(n559), .B2(Q[631]), .ZN(n624) );
  AOI22_X1 U689 ( .A1(n558), .A2(Q[696]), .B1(n557), .B2(Q[600]), .ZN(n627) );
  AOI22_X1 U690 ( .A1(n560), .A2(Q[536]), .B1(n559), .B2(Q[632]), .ZN(n626) );
  AOI22_X1 U691 ( .A1(n558), .A2(Q[697]), .B1(n557), .B2(Q[601]), .ZN(n629) );
  AOI22_X1 U692 ( .A1(n560), .A2(Q[537]), .B1(n559), .B2(Q[633]), .ZN(n628) );
  AOI22_X1 U693 ( .A1(n558), .A2(Q[698]), .B1(n557), .B2(Q[602]), .ZN(n631) );
  AOI22_X1 U694 ( .A1(n560), .A2(Q[538]), .B1(n559), .B2(Q[634]), .ZN(n630) );
  AOI22_X1 U695 ( .A1(n558), .A2(Q[699]), .B1(n557), .B2(Q[603]), .ZN(n633) );
  AOI22_X1 U696 ( .A1(n560), .A2(Q[539]), .B1(n559), .B2(Q[635]), .ZN(n632) );
  AOI22_X1 U697 ( .A1(n558), .A2(Q[700]), .B1(n557), .B2(Q[604]), .ZN(n635) );
  AOI22_X1 U698 ( .A1(n560), .A2(Q[540]), .B1(n559), .B2(Q[636]), .ZN(n634) );
  AOI22_X1 U699 ( .A1(n668), .A2(Q[701]), .B1(n667), .B2(Q[605]), .ZN(n637) );
  AOI22_X1 U700 ( .A1(n670), .A2(Q[541]), .B1(n669), .B2(Q[637]), .ZN(n636) );
  AOI22_X1 U701 ( .A1(n558), .A2(Q[674]), .B1(n557), .B2(Q[578]), .ZN(n639) );
  AOI22_X1 U702 ( .A1(n560), .A2(Q[514]), .B1(n559), .B2(Q[610]), .ZN(n638) );
  AOI22_X1 U703 ( .A1(n558), .A2(Q[702]), .B1(n557), .B2(Q[606]), .ZN(n641) );
  AOI22_X1 U704 ( .A1(n560), .A2(Q[542]), .B1(n559), .B2(Q[638]), .ZN(n640) );
  AOI22_X1 U705 ( .A1(n558), .A2(Q[703]), .B1(n557), .B2(Q[607]), .ZN(n643) );
  AOI22_X1 U706 ( .A1(n560), .A2(Q[543]), .B1(n559), .B2(Q[639]), .ZN(n642) );
  AOI22_X1 U707 ( .A1(n558), .A2(Q[675]), .B1(n557), .B2(Q[579]), .ZN(n645) );
  AOI22_X1 U708 ( .A1(n560), .A2(Q[515]), .B1(n559), .B2(Q[611]), .ZN(n644) );
  AOI22_X1 U709 ( .A1(n558), .A2(Q[676]), .B1(n557), .B2(Q[580]), .ZN(n647) );
  AOI22_X1 U710 ( .A1(n560), .A2(Q[516]), .B1(n559), .B2(Q[612]), .ZN(n646) );
  AOI22_X1 U711 ( .A1(n558), .A2(Q[677]), .B1(n557), .B2(Q[581]), .ZN(n649) );
  AOI22_X1 U712 ( .A1(n560), .A2(Q[517]), .B1(n559), .B2(Q[613]), .ZN(n648) );
  AOI22_X1 U713 ( .A1(n558), .A2(Q[678]), .B1(n557), .B2(Q[582]), .ZN(n651) );
  AOI22_X1 U714 ( .A1(n560), .A2(Q[518]), .B1(n559), .B2(Q[614]), .ZN(n650) );
  AOI22_X1 U715 ( .A1(n558), .A2(Q[679]), .B1(n557), .B2(Q[583]), .ZN(n653) );
  AOI22_X1 U716 ( .A1(n560), .A2(Q[519]), .B1(n559), .B2(Q[615]), .ZN(n652) );
  AOI22_X1 U717 ( .A1(n558), .A2(Q[680]), .B1(n557), .B2(Q[584]), .ZN(n655) );
  AOI22_X1 U718 ( .A1(n560), .A2(Q[520]), .B1(n559), .B2(Q[616]), .ZN(n654) );
  AOI22_X1 U719 ( .A1(n558), .A2(Q[681]), .B1(n557), .B2(Q[585]), .ZN(n672) );
  AOI22_X1 U720 ( .A1(n560), .A2(Q[521]), .B1(n559), .B2(Q[617]), .ZN(n671) );
endmodule


module select_block_NBIT_DATA32_N8_F5 ( regs, win, curr_proc_regs );
  input [2559:0] regs;
  input [4:0] win;
  output [767:0] curr_proc_regs;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221;

  INV_X1 U2 ( .A(n138), .ZN(n7) );
  BUF_X1 U3 ( .A(n102), .Z(n5) );
  CLKBUF_X3 U4 ( .A(n2207), .Z(n65) );
  BUF_X4 U5 ( .A(n77), .Z(n9) );
  BUF_X2 U6 ( .A(n64), .Z(n1) );
  BUF_X2 U7 ( .A(n67), .Z(n77) );
  INV_X2 U8 ( .A(n63), .ZN(n2) );
  INV_X2 U9 ( .A(n2134), .ZN(n3) );
  BUF_X1 U10 ( .A(n101), .Z(n16) );
  NAND2_X2 U11 ( .A1(n141), .A2(win[1]), .ZN(n2207) );
  NAND3_X2 U12 ( .A1(n141), .A2(win[0]), .A3(n140), .ZN(n2134) );
  BUF_X2 U13 ( .A(n2217), .Z(n4) );
  NAND3_X2 U14 ( .A1(n139), .A2(n137), .A3(win[2]), .ZN(n2221) );
  INV_X1 U15 ( .A(n138), .ZN(n20) );
  INV_X2 U16 ( .A(n137), .ZN(n6) );
  INV_X2 U17 ( .A(n63), .ZN(n8) );
  INV_X2 U18 ( .A(n63), .ZN(n10) );
  BUF_X2 U19 ( .A(n2207), .Z(n11) );
  INV_X2 U20 ( .A(n2134), .ZN(n12) );
  INV_X2 U21 ( .A(n63), .ZN(n13) );
  BUF_X2 U22 ( .A(n2134), .Z(n25) );
  BUF_X2 U23 ( .A(n2134), .Z(n24) );
  BUF_X2 U24 ( .A(n4), .Z(n14) );
  BUF_X2 U25 ( .A(n2217), .Z(n73) );
  BUF_X2 U26 ( .A(n2217), .Z(n67) );
  BUF_X2 U27 ( .A(n4), .Z(n15) );
  BUF_X2 U28 ( .A(n2217), .Z(n17) );
  INV_X2 U29 ( .A(n102), .ZN(n18) );
  INV_X2 U30 ( .A(n102), .ZN(n19) );
  INV_X2 U31 ( .A(n137), .ZN(n21) );
  BUF_X4 U32 ( .A(n2217), .Z(n71) );
  INV_X1 U33 ( .A(n63), .ZN(n62) );
  BUF_X1 U34 ( .A(n65), .Z(n63) );
  BUF_X1 U35 ( .A(n2207), .Z(n64) );
  INV_X1 U36 ( .A(n137), .ZN(n103) );
  INV_X1 U37 ( .A(win[4]), .ZN(n137) );
  INV_X1 U38 ( .A(win[4]), .ZN(n138) );
  BUF_X2 U39 ( .A(n4), .Z(n68) );
  BUF_X2 U40 ( .A(n2217), .Z(n72) );
  BUF_X1 U41 ( .A(n102), .Z(n100) );
  BUF_X1 U42 ( .A(n101), .Z(n99) );
  BUF_X1 U43 ( .A(n4), .Z(n66) );
  BUF_X1 U44 ( .A(n14), .Z(n74) );
  BUF_X1 U45 ( .A(n14), .Z(n70) );
  BUF_X1 U46 ( .A(n17), .Z(n76) );
  BUF_X1 U47 ( .A(n17), .Z(n75) );
  BUF_X1 U48 ( .A(n2221), .Z(n101) );
  BUF_X1 U49 ( .A(n2221), .Z(n102) );
  BUF_X1 U50 ( .A(n15), .Z(n69) );
  INV_X1 U51 ( .A(n2134), .ZN(n26) );
  INV_X1 U52 ( .A(n2134), .ZN(n27) );
  INV_X1 U53 ( .A(n24), .ZN(n28) );
  INV_X1 U54 ( .A(n2134), .ZN(n29) );
  INV_X1 U55 ( .A(n2134), .ZN(n30) );
  INV_X1 U56 ( .A(n2134), .ZN(n31) );
  INV_X1 U57 ( .A(n2134), .ZN(n32) );
  INV_X1 U58 ( .A(n2134), .ZN(n33) );
  INV_X1 U59 ( .A(n2134), .ZN(n34) );
  INV_X1 U60 ( .A(n2134), .ZN(n35) );
  INV_X1 U61 ( .A(n2134), .ZN(n36) );
  INV_X1 U62 ( .A(n2134), .ZN(n37) );
  INV_X1 U63 ( .A(n2134), .ZN(n38) );
  INV_X1 U64 ( .A(n2134), .ZN(n39) );
  INV_X1 U65 ( .A(n2134), .ZN(n40) );
  INV_X1 U66 ( .A(n2134), .ZN(n41) );
  INV_X1 U67 ( .A(n2134), .ZN(n42) );
  INV_X1 U68 ( .A(n2134), .ZN(n43) );
  INV_X1 U69 ( .A(n2134), .ZN(n44) );
  INV_X1 U70 ( .A(n2134), .ZN(n45) );
  INV_X1 U71 ( .A(n2134), .ZN(n46) );
  INV_X1 U72 ( .A(n2134), .ZN(n47) );
  INV_X1 U73 ( .A(n2134), .ZN(n48) );
  INV_X1 U74 ( .A(n63), .ZN(n49) );
  INV_X1 U75 ( .A(n2207), .ZN(n50) );
  INV_X1 U76 ( .A(n2207), .ZN(n51) );
  INV_X1 U77 ( .A(n2207), .ZN(n52) );
  INV_X1 U78 ( .A(n2207), .ZN(n53) );
  INV_X1 U79 ( .A(n2207), .ZN(n54) );
  INV_X1 U80 ( .A(n2207), .ZN(n55) );
  INV_X1 U81 ( .A(n63), .ZN(n56) );
  INV_X1 U82 ( .A(n2207), .ZN(n57) );
  INV_X1 U83 ( .A(n2207), .ZN(n58) );
  INV_X1 U84 ( .A(n63), .ZN(n59) );
  INV_X1 U85 ( .A(n63), .ZN(n60) );
  INV_X1 U86 ( .A(n63), .ZN(n61) );
  INV_X1 U87 ( .A(n2221), .ZN(n78) );
  INV_X1 U88 ( .A(n2221), .ZN(n79) );
  INV_X1 U89 ( .A(n2221), .ZN(n80) );
  INV_X1 U90 ( .A(n2221), .ZN(n81) );
  INV_X1 U91 ( .A(n2221), .ZN(n82) );
  INV_X1 U92 ( .A(n2221), .ZN(n83) );
  INV_X1 U93 ( .A(n2221), .ZN(n84) );
  INV_X1 U94 ( .A(n2221), .ZN(n85) );
  INV_X1 U95 ( .A(n2221), .ZN(n86) );
  INV_X1 U96 ( .A(n2221), .ZN(n87) );
  INV_X1 U97 ( .A(n2221), .ZN(n88) );
  INV_X1 U98 ( .A(n102), .ZN(n89) );
  INV_X1 U99 ( .A(n2221), .ZN(n90) );
  INV_X1 U100 ( .A(n102), .ZN(n91) );
  INV_X1 U101 ( .A(n2221), .ZN(n92) );
  INV_X1 U102 ( .A(n2221), .ZN(n93) );
  INV_X1 U103 ( .A(n2221), .ZN(n94) );
  INV_X1 U104 ( .A(n2221), .ZN(n95) );
  INV_X1 U105 ( .A(n2221), .ZN(n96) );
  INV_X1 U106 ( .A(n100), .ZN(n97) );
  INV_X1 U107 ( .A(n2221), .ZN(n98) );
  INV_X1 U108 ( .A(n137), .ZN(n104) );
  INV_X1 U109 ( .A(n137), .ZN(n105) );
  INV_X1 U110 ( .A(n137), .ZN(n106) );
  INV_X1 U111 ( .A(n137), .ZN(n107) );
  INV_X1 U112 ( .A(n137), .ZN(n108) );
  INV_X1 U113 ( .A(n137), .ZN(n109) );
  INV_X1 U114 ( .A(n137), .ZN(n110) );
  INV_X1 U115 ( .A(n137), .ZN(n111) );
  INV_X1 U116 ( .A(n137), .ZN(n112) );
  INV_X1 U117 ( .A(n137), .ZN(n113) );
  INV_X1 U118 ( .A(n137), .ZN(n114) );
  INV_X1 U119 ( .A(n137), .ZN(n115) );
  INV_X1 U120 ( .A(n137), .ZN(n116) );
  INV_X1 U121 ( .A(n137), .ZN(n117) );
  INV_X1 U122 ( .A(n137), .ZN(n118) );
  INV_X1 U123 ( .A(n137), .ZN(n119) );
  INV_X1 U124 ( .A(n137), .ZN(n120) );
  INV_X1 U125 ( .A(n137), .ZN(n121) );
  INV_X1 U126 ( .A(n138), .ZN(n122) );
  INV_X1 U127 ( .A(n138), .ZN(n123) );
  INV_X1 U128 ( .A(n138), .ZN(n124) );
  INV_X1 U129 ( .A(n138), .ZN(n125) );
  INV_X1 U130 ( .A(n138), .ZN(n126) );
  INV_X1 U131 ( .A(n138), .ZN(n127) );
  INV_X1 U132 ( .A(n138), .ZN(n128) );
  INV_X1 U133 ( .A(n138), .ZN(n129) );
  INV_X1 U134 ( .A(n138), .ZN(n130) );
  INV_X1 U135 ( .A(n138), .ZN(n131) );
  INV_X1 U136 ( .A(n138), .ZN(n132) );
  INV_X1 U137 ( .A(n138), .ZN(n133) );
  INV_X1 U138 ( .A(n138), .ZN(n134) );
  INV_X1 U139 ( .A(n138), .ZN(n135) );
  INV_X1 U140 ( .A(n138), .ZN(n136) );
  NOR3_X1 U141 ( .A1(win[3]), .A2(n130), .A3(win[2]), .ZN(n141) );
  INV_X1 U142 ( .A(regs[512]), .ZN(n1316) );
  INV_X1 U143 ( .A(win[3]), .ZN(n139) );
  NOR2_X1 U144 ( .A1(n103), .A2(n139), .ZN(n2217) );
  AOI22_X1 U145 ( .A1(n126), .A2(regs[2048]), .B1(n68), .B2(regs[1536]), .ZN(
        n143) );
  INV_X1 U146 ( .A(win[1]), .ZN(n140) );
  AOI22_X1 U147 ( .A1(n92), .A2(regs[1024]), .B1(n47), .B2(regs[0]), .ZN(n142)
         );
  OAI211_X1 U148 ( .C1(n1), .C2(n1316), .A(n143), .B(n142), .ZN(
        curr_proc_regs[0]) );
  INV_X1 U149 ( .A(regs[1124]), .ZN(n1623) );
  AOI22_X1 U150 ( .A1(n126), .A2(regs[2148]), .B1(n68), .B2(regs[1636]), .ZN(
        n145) );
  AOI22_X1 U151 ( .A1(n59), .A2(regs[612]), .B1(n46), .B2(regs[100]), .ZN(n144) );
  OAI211_X1 U152 ( .C1(n101), .C2(n1623), .A(n145), .B(n144), .ZN(
        curr_proc_regs[100]) );
  INV_X1 U153 ( .A(regs[613]), .ZN(n1626) );
  AOI22_X1 U154 ( .A1(n126), .A2(regs[2149]), .B1(n68), .B2(regs[1637]), .ZN(
        n147) );
  AOI22_X1 U155 ( .A1(n89), .A2(regs[1125]), .B1(n47), .B2(regs[101]), .ZN(
        n146) );
  OAI211_X1 U156 ( .C1(n65), .C2(n1626), .A(n147), .B(n146), .ZN(
        curr_proc_regs[101]) );
  INV_X1 U157 ( .A(regs[614]), .ZN(n1629) );
  AOI22_X1 U158 ( .A1(n126), .A2(regs[2150]), .B1(n68), .B2(regs[1638]), .ZN(
        n149) );
  AOI22_X1 U159 ( .A1(n89), .A2(regs[1126]), .B1(n46), .B2(regs[102]), .ZN(
        n148) );
  OAI211_X1 U160 ( .C1(n1), .C2(n1629), .A(n149), .B(n148), .ZN(
        curr_proc_regs[102]) );
  INV_X1 U161 ( .A(regs[615]), .ZN(n1632) );
  AOI22_X1 U162 ( .A1(n126), .A2(regs[2151]), .B1(n68), .B2(regs[1639]), .ZN(
        n151) );
  AOI22_X1 U163 ( .A1(n18), .A2(regs[1127]), .B1(n46), .B2(regs[103]), .ZN(
        n150) );
  OAI211_X1 U164 ( .C1(n1), .C2(n1632), .A(n151), .B(n150), .ZN(
        curr_proc_regs[103]) );
  INV_X1 U165 ( .A(regs[616]), .ZN(n1635) );
  AOI22_X1 U166 ( .A1(win[4]), .A2(regs[2152]), .B1(n68), .B2(regs[1640]), 
        .ZN(n153) );
  AOI22_X1 U167 ( .A1(n18), .A2(regs[1128]), .B1(n46), .B2(regs[104]), .ZN(
        n152) );
  OAI211_X1 U168 ( .C1(n1), .C2(n1635), .A(n153), .B(n152), .ZN(
        curr_proc_regs[104]) );
  INV_X1 U169 ( .A(regs[617]), .ZN(n1638) );
  AOI22_X1 U170 ( .A1(n130), .A2(regs[2153]), .B1(n68), .B2(regs[1641]), .ZN(
        n155) );
  AOI22_X1 U171 ( .A1(n18), .A2(regs[1129]), .B1(n46), .B2(regs[105]), .ZN(
        n154) );
  OAI211_X1 U172 ( .C1(n2207), .C2(n1638), .A(n155), .B(n154), .ZN(
        curr_proc_regs[105]) );
  INV_X1 U173 ( .A(regs[618]), .ZN(n1641) );
  AOI22_X1 U174 ( .A1(n126), .A2(regs[2154]), .B1(n68), .B2(regs[1642]), .ZN(
        n157) );
  AOI22_X1 U175 ( .A1(n18), .A2(regs[1130]), .B1(n46), .B2(regs[106]), .ZN(
        n156) );
  OAI211_X1 U176 ( .C1(n2207), .C2(n1641), .A(n157), .B(n156), .ZN(
        curr_proc_regs[106]) );
  INV_X1 U177 ( .A(regs[1131]), .ZN(n1644) );
  AOI22_X1 U178 ( .A1(n136), .A2(regs[2155]), .B1(n68), .B2(regs[1643]), .ZN(
        n159) );
  AOI22_X1 U179 ( .A1(n53), .A2(regs[619]), .B1(n46), .B2(regs[107]), .ZN(n158) );
  OAI211_X1 U180 ( .C1(n101), .C2(n1644), .A(n159), .B(n158), .ZN(
        curr_proc_regs[107]) );
  INV_X1 U181 ( .A(regs[620]), .ZN(n1650) );
  AOI22_X1 U182 ( .A1(n135), .A2(regs[2156]), .B1(n68), .B2(regs[1644]), .ZN(
        n161) );
  AOI22_X1 U183 ( .A1(n93), .A2(regs[1132]), .B1(n46), .B2(regs[108]), .ZN(
        n160) );
  OAI211_X1 U184 ( .C1(n1), .C2(n1650), .A(n161), .B(n160), .ZN(
        curr_proc_regs[108]) );
  INV_X1 U185 ( .A(regs[1133]), .ZN(n1653) );
  AOI22_X1 U186 ( .A1(n134), .A2(regs[2157]), .B1(n68), .B2(regs[1645]), .ZN(
        n163) );
  AOI22_X1 U187 ( .A1(n59), .A2(regs[621]), .B1(n46), .B2(regs[109]), .ZN(n162) );
  OAI211_X1 U188 ( .C1(n101), .C2(n1653), .A(n163), .B(n162), .ZN(
        curr_proc_regs[109]) );
  INV_X1 U189 ( .A(regs[522]), .ZN(n1345) );
  AOI22_X1 U190 ( .A1(n133), .A2(regs[2058]), .B1(n67), .B2(regs[1546]), .ZN(
        n165) );
  AOI22_X1 U191 ( .A1(n18), .A2(regs[1034]), .B1(n47), .B2(regs[10]), .ZN(n164) );
  OAI211_X1 U192 ( .C1(n1), .C2(n1345), .A(n165), .B(n164), .ZN(
        curr_proc_regs[10]) );
  INV_X1 U193 ( .A(regs[622]), .ZN(n1656) );
  AOI22_X1 U194 ( .A1(n132), .A2(regs[2158]), .B1(n67), .B2(regs[1646]), .ZN(
        n167) );
  AOI22_X1 U195 ( .A1(n18), .A2(regs[1134]), .B1(n46), .B2(regs[110]), .ZN(
        n166) );
  OAI211_X1 U196 ( .C1(n1), .C2(n1656), .A(n167), .B(n166), .ZN(
        curr_proc_regs[110]) );
  INV_X1 U197 ( .A(regs[623]), .ZN(n1659) );
  AOI22_X1 U198 ( .A1(n127), .A2(regs[2159]), .B1(n67), .B2(regs[1647]), .ZN(
        n169) );
  AOI22_X1 U199 ( .A1(n18), .A2(regs[1135]), .B1(n46), .B2(regs[111]), .ZN(
        n168) );
  OAI211_X1 U200 ( .C1(n2207), .C2(n1659), .A(n169), .B(n168), .ZN(
        curr_proc_regs[111]) );
  INV_X1 U201 ( .A(regs[624]), .ZN(n1662) );
  AOI22_X1 U202 ( .A1(n128), .A2(regs[2160]), .B1(n67), .B2(regs[1648]), .ZN(
        n171) );
  AOI22_X1 U203 ( .A1(n83), .A2(regs[1136]), .B1(n48), .B2(regs[112]), .ZN(
        n170) );
  OAI211_X1 U204 ( .C1(n1), .C2(n1662), .A(n171), .B(n170), .ZN(
        curr_proc_regs[112]) );
  INV_X1 U205 ( .A(regs[625]), .ZN(n1665) );
  AOI22_X1 U206 ( .A1(n129), .A2(regs[2161]), .B1(n67), .B2(regs[1649]), .ZN(
        n173) );
  AOI22_X1 U207 ( .A1(n18), .A2(regs[1137]), .B1(n46), .B2(regs[113]), .ZN(
        n172) );
  OAI211_X1 U208 ( .C1(n1), .C2(n1665), .A(n173), .B(n172), .ZN(
        curr_proc_regs[113]) );
  INV_X1 U209 ( .A(regs[626]), .ZN(n1668) );
  AOI22_X1 U210 ( .A1(n123), .A2(regs[2162]), .B1(n67), .B2(regs[1650]), .ZN(
        n175) );
  AOI22_X1 U211 ( .A1(n18), .A2(regs[1138]), .B1(n48), .B2(regs[114]), .ZN(
        n174) );
  OAI211_X1 U212 ( .C1(n1), .C2(n1668), .A(n175), .B(n174), .ZN(
        curr_proc_regs[114]) );
  INV_X1 U213 ( .A(regs[627]), .ZN(n1671) );
  AOI22_X1 U214 ( .A1(n124), .A2(regs[2163]), .B1(n67), .B2(regs[1651]), .ZN(
        n177) );
  AOI22_X1 U215 ( .A1(n18), .A2(regs[1139]), .B1(n47), .B2(regs[115]), .ZN(
        n176) );
  OAI211_X1 U216 ( .C1(n2207), .C2(n1671), .A(n177), .B(n176), .ZN(
        curr_proc_regs[115]) );
  INV_X1 U217 ( .A(regs[628]), .ZN(n1674) );
  AOI22_X1 U218 ( .A1(n125), .A2(regs[2164]), .B1(n67), .B2(regs[1652]), .ZN(
        n179) );
  AOI22_X1 U219 ( .A1(n90), .A2(regs[1140]), .B1(n47), .B2(regs[116]), .ZN(
        n178) );
  OAI211_X1 U220 ( .C1(n1), .C2(n1674), .A(n179), .B(n178), .ZN(
        curr_proc_regs[116]) );
  INV_X1 U221 ( .A(regs[629]), .ZN(n1677) );
  AOI22_X1 U222 ( .A1(win[4]), .A2(regs[2165]), .B1(n67), .B2(regs[1653]), 
        .ZN(n181) );
  AOI22_X1 U223 ( .A1(n88), .A2(regs[1141]), .B1(n48), .B2(regs[117]), .ZN(
        n180) );
  OAI211_X1 U224 ( .C1(n2207), .C2(n1677), .A(n181), .B(n180), .ZN(
        curr_proc_regs[117]) );
  INV_X1 U225 ( .A(regs[630]), .ZN(n1683) );
  AOI22_X1 U226 ( .A1(n130), .A2(regs[2166]), .B1(n67), .B2(regs[1654]), .ZN(
        n183) );
  AOI22_X1 U227 ( .A1(n87), .A2(regs[1142]), .B1(n46), .B2(regs[118]), .ZN(
        n182) );
  OAI211_X1 U228 ( .C1(n1), .C2(n1683), .A(n183), .B(n182), .ZN(
        curr_proc_regs[118]) );
  INV_X1 U229 ( .A(regs[1143]), .ZN(n1686) );
  AOI22_X1 U230 ( .A1(n126), .A2(regs[2167]), .B1(n67), .B2(regs[1655]), .ZN(
        n185) );
  AOI22_X1 U231 ( .A1(n49), .A2(regs[631]), .B1(n48), .B2(regs[119]), .ZN(n184) );
  OAI211_X1 U232 ( .C1(n101), .C2(n1686), .A(n185), .B(n184), .ZN(
        curr_proc_regs[119]) );
  INV_X1 U233 ( .A(regs[523]), .ZN(n1348) );
  AOI22_X1 U234 ( .A1(n136), .A2(regs[2059]), .B1(n15), .B2(regs[1547]), .ZN(
        n187) );
  AOI22_X1 U235 ( .A1(n92), .A2(regs[1035]), .B1(n47), .B2(regs[11]), .ZN(n186) );
  OAI211_X1 U236 ( .C1(n1), .C2(n1348), .A(n187), .B(n186), .ZN(
        curr_proc_regs[11]) );
  INV_X1 U237 ( .A(regs[1144]), .ZN(n1689) );
  AOI22_X1 U238 ( .A1(n135), .A2(regs[2168]), .B1(n15), .B2(regs[1656]), .ZN(
        n189) );
  AOI22_X1 U239 ( .A1(n50), .A2(regs[632]), .B1(n46), .B2(regs[120]), .ZN(n188) );
  OAI211_X1 U240 ( .C1(n101), .C2(n1689), .A(n189), .B(n188), .ZN(
        curr_proc_regs[120]) );
  INV_X1 U241 ( .A(regs[633]), .ZN(n1692) );
  AOI22_X1 U242 ( .A1(n134), .A2(regs[2169]), .B1(n15), .B2(regs[1657]), .ZN(
        n191) );
  AOI22_X1 U243 ( .A1(n96), .A2(regs[1145]), .B1(n48), .B2(regs[121]), .ZN(
        n190) );
  OAI211_X1 U244 ( .C1(n2207), .C2(n1692), .A(n191), .B(n190), .ZN(
        curr_proc_regs[121]) );
  INV_X1 U245 ( .A(regs[1146]), .ZN(n1695) );
  AOI22_X1 U246 ( .A1(n133), .A2(regs[2170]), .B1(n15), .B2(regs[1658]), .ZN(
        n193) );
  AOI22_X1 U247 ( .A1(n51), .A2(regs[634]), .B1(n47), .B2(regs[122]), .ZN(n192) );
  OAI211_X1 U248 ( .C1(n101), .C2(n1695), .A(n193), .B(n192), .ZN(
        curr_proc_regs[122]) );
  INV_X1 U249 ( .A(regs[635]), .ZN(n1698) );
  AOI22_X1 U250 ( .A1(n132), .A2(regs[2171]), .B1(n15), .B2(regs[1659]), .ZN(
        n195) );
  AOI22_X1 U251 ( .A1(n18), .A2(regs[1147]), .B1(n48), .B2(regs[123]), .ZN(
        n194) );
  OAI211_X1 U252 ( .C1(n1), .C2(n1698), .A(n195), .B(n194), .ZN(
        curr_proc_regs[123]) );
  INV_X1 U253 ( .A(regs[1148]), .ZN(n1701) );
  AOI22_X1 U254 ( .A1(n125), .A2(regs[2172]), .B1(n15), .B2(regs[1660]), .ZN(
        n197) );
  AOI22_X1 U255 ( .A1(n55), .A2(regs[636]), .B1(n46), .B2(regs[124]), .ZN(n196) );
  OAI211_X1 U256 ( .C1(n2221), .C2(n1701), .A(n197), .B(n196), .ZN(
        curr_proc_regs[124]) );
  INV_X1 U257 ( .A(regs[1149]), .ZN(n1704) );
  AOI22_X1 U258 ( .A1(n125), .A2(regs[2173]), .B1(n15), .B2(regs[1661]), .ZN(
        n199) );
  AOI22_X1 U259 ( .A1(n57), .A2(regs[637]), .B1(n48), .B2(regs[125]), .ZN(n198) );
  OAI211_X1 U260 ( .C1(n101), .C2(n1704), .A(n199), .B(n198), .ZN(
        curr_proc_regs[125]) );
  INV_X1 U261 ( .A(regs[1150]), .ZN(n1707) );
  AOI22_X1 U262 ( .A1(n125), .A2(regs[2174]), .B1(n15), .B2(regs[1662]), .ZN(
        n201) );
  AOI22_X1 U263 ( .A1(n57), .A2(regs[638]), .B1(n47), .B2(regs[126]), .ZN(n200) );
  OAI211_X1 U264 ( .C1(n101), .C2(n1707), .A(n201), .B(n200), .ZN(
        curr_proc_regs[126]) );
  INV_X1 U265 ( .A(regs[1151]), .ZN(n1710) );
  AOI22_X1 U266 ( .A1(n125), .A2(regs[2175]), .B1(n15), .B2(regs[1663]), .ZN(
        n203) );
  AOI22_X1 U267 ( .A1(n57), .A2(regs[639]), .B1(n47), .B2(regs[127]), .ZN(n202) );
  OAI211_X1 U268 ( .C1(n101), .C2(n1710), .A(n203), .B(n202), .ZN(
        curr_proc_regs[127]) );
  INV_X1 U269 ( .A(regs[1152]), .ZN(n1716) );
  AOI22_X1 U270 ( .A1(n125), .A2(regs[2176]), .B1(n15), .B2(regs[1664]), .ZN(
        n205) );
  AOI22_X1 U271 ( .A1(n53), .A2(regs[640]), .B1(n46), .B2(regs[128]), .ZN(n204) );
  OAI211_X1 U272 ( .C1(n101), .C2(n1716), .A(n205), .B(n204), .ZN(
        curr_proc_regs[128]) );
  INV_X1 U273 ( .A(regs[641]), .ZN(n1719) );
  AOI22_X1 U274 ( .A1(n125), .A2(regs[2177]), .B1(n15), .B2(regs[1665]), .ZN(
        n207) );
  AOI22_X1 U275 ( .A1(n95), .A2(regs[1153]), .B1(n48), .B2(regs[129]), .ZN(
        n206) );
  OAI211_X1 U276 ( .C1(n2207), .C2(n1719), .A(n207), .B(n206), .ZN(
        curr_proc_regs[129]) );
  INV_X1 U277 ( .A(regs[524]), .ZN(n1351) );
  AOI22_X1 U278 ( .A1(n125), .A2(regs[2060]), .B1(n15), .B2(regs[1548]), .ZN(
        n209) );
  AOI22_X1 U279 ( .A1(n18), .A2(regs[1036]), .B1(n47), .B2(regs[12]), .ZN(n208) );
  OAI211_X1 U280 ( .C1(n2207), .C2(n1351), .A(n209), .B(n208), .ZN(
        curr_proc_regs[12]) );
  INV_X1 U281 ( .A(regs[1154]), .ZN(n1722) );
  AOI22_X1 U282 ( .A1(n125), .A2(regs[2178]), .B1(n15), .B2(regs[1666]), .ZN(
        n211) );
  AOI22_X1 U283 ( .A1(n58), .A2(regs[642]), .B1(n47), .B2(regs[130]), .ZN(n210) );
  OAI211_X1 U284 ( .C1(n101), .C2(n1722), .A(n211), .B(n210), .ZN(
        curr_proc_regs[130]) );
  INV_X1 U285 ( .A(regs[1155]), .ZN(n1725) );
  AOI22_X1 U286 ( .A1(n125), .A2(regs[2179]), .B1(n15), .B2(regs[1667]), .ZN(
        n213) );
  AOI22_X1 U287 ( .A1(n58), .A2(regs[643]), .B1(n47), .B2(regs[131]), .ZN(n212) );
  OAI211_X1 U288 ( .C1(n101), .C2(n1725), .A(n213), .B(n212), .ZN(
        curr_proc_regs[131]) );
  INV_X1 U289 ( .A(regs[1156]), .ZN(n1728) );
  AOI22_X1 U290 ( .A1(n125), .A2(regs[2180]), .B1(n15), .B2(regs[1668]), .ZN(
        n215) );
  AOI22_X1 U291 ( .A1(n55), .A2(regs[644]), .B1(n47), .B2(regs[132]), .ZN(n214) );
  OAI211_X1 U292 ( .C1(n101), .C2(n1728), .A(n215), .B(n214), .ZN(
        curr_proc_regs[132]) );
  INV_X1 U293 ( .A(regs[1157]), .ZN(n1731) );
  AOI22_X1 U294 ( .A1(n125), .A2(regs[2181]), .B1(n15), .B2(regs[1669]), .ZN(
        n217) );
  AOI22_X1 U295 ( .A1(n50), .A2(regs[645]), .B1(n48), .B2(regs[133]), .ZN(n216) );
  OAI211_X1 U296 ( .C1(n2221), .C2(n1731), .A(n217), .B(n216), .ZN(
        curr_proc_regs[133]) );
  INV_X1 U297 ( .A(regs[1158]), .ZN(n1734) );
  AOI22_X1 U298 ( .A1(n124), .A2(regs[2182]), .B1(n15), .B2(regs[1670]), .ZN(
        n219) );
  AOI22_X1 U299 ( .A1(n58), .A2(regs[646]), .B1(n47), .B2(regs[134]), .ZN(n218) );
  OAI211_X1 U300 ( .C1(n101), .C2(n1734), .A(n219), .B(n218), .ZN(
        curr_proc_regs[134]) );
  INV_X1 U301 ( .A(regs[647]), .ZN(n1737) );
  AOI22_X1 U302 ( .A1(n124), .A2(regs[2183]), .B1(n15), .B2(regs[1671]), .ZN(
        n221) );
  AOI22_X1 U303 ( .A1(n18), .A2(regs[1159]), .B1(n46), .B2(regs[135]), .ZN(
        n220) );
  OAI211_X1 U304 ( .C1(n1), .C2(n1737), .A(n221), .B(n220), .ZN(
        curr_proc_regs[135]) );
  INV_X1 U305 ( .A(regs[648]), .ZN(n1740) );
  AOI22_X1 U306 ( .A1(n124), .A2(regs[2184]), .B1(n15), .B2(regs[1672]), .ZN(
        n223) );
  AOI22_X1 U307 ( .A1(n18), .A2(regs[1160]), .B1(n48), .B2(regs[136]), .ZN(
        n222) );
  OAI211_X1 U308 ( .C1(n1), .C2(n1740), .A(n223), .B(n222), .ZN(
        curr_proc_regs[136]) );
  INV_X1 U309 ( .A(regs[1161]), .ZN(n1743) );
  AOI22_X1 U310 ( .A1(n124), .A2(regs[2185]), .B1(n15), .B2(regs[1673]), .ZN(
        n225) );
  AOI22_X1 U311 ( .A1(n60), .A2(regs[649]), .B1(n47), .B2(regs[137]), .ZN(n224) );
  OAI211_X1 U312 ( .C1(n2221), .C2(n1743), .A(n225), .B(n224), .ZN(
        curr_proc_regs[137]) );
  INV_X1 U313 ( .A(regs[650]), .ZN(n1749) );
  AOI22_X1 U314 ( .A1(n124), .A2(regs[2186]), .B1(n15), .B2(regs[1674]), .ZN(
        n227) );
  AOI22_X1 U315 ( .A1(n18), .A2(regs[1162]), .B1(n46), .B2(regs[138]), .ZN(
        n226) );
  OAI211_X1 U316 ( .C1(n2207), .C2(n1749), .A(n227), .B(n226), .ZN(
        curr_proc_regs[138]) );
  INV_X1 U317 ( .A(regs[1163]), .ZN(n1752) );
  AOI22_X1 U318 ( .A1(n124), .A2(regs[2187]), .B1(n15), .B2(regs[1675]), .ZN(
        n229) );
  AOI22_X1 U319 ( .A1(n55), .A2(regs[651]), .B1(n48), .B2(regs[139]), .ZN(n228) );
  OAI211_X1 U320 ( .C1(n101), .C2(n1752), .A(n229), .B(n228), .ZN(
        curr_proc_regs[139]) );
  INV_X1 U321 ( .A(regs[525]), .ZN(n1354) );
  AOI22_X1 U322 ( .A1(n124), .A2(regs[2061]), .B1(n68), .B2(regs[1549]), .ZN(
        n231) );
  AOI22_X1 U323 ( .A1(n18), .A2(regs[1037]), .B1(n48), .B2(regs[13]), .ZN(n230) );
  OAI211_X1 U324 ( .C1(n1), .C2(n1354), .A(n231), .B(n230), .ZN(
        curr_proc_regs[13]) );
  INV_X1 U325 ( .A(regs[652]), .ZN(n1755) );
  AOI22_X1 U326 ( .A1(n124), .A2(regs[2188]), .B1(n66), .B2(regs[1676]), .ZN(
        n233) );
  AOI22_X1 U327 ( .A1(n18), .A2(regs[1164]), .B1(n48), .B2(regs[140]), .ZN(
        n232) );
  OAI211_X1 U328 ( .C1(n2207), .C2(n1755), .A(n233), .B(n232), .ZN(
        curr_proc_regs[140]) );
  INV_X1 U329 ( .A(regs[1165]), .ZN(n1758) );
  AOI22_X1 U330 ( .A1(n124), .A2(regs[2189]), .B1(n15), .B2(regs[1677]), .ZN(
        n235) );
  AOI22_X1 U331 ( .A1(n57), .A2(regs[653]), .B1(n48), .B2(regs[141]), .ZN(n234) );
  OAI211_X1 U332 ( .C1(n2221), .C2(n1758), .A(n235), .B(n234), .ZN(
        curr_proc_regs[141]) );
  INV_X1 U333 ( .A(regs[654]), .ZN(n1761) );
  AOI22_X1 U334 ( .A1(n124), .A2(regs[2190]), .B1(n15), .B2(regs[1678]), .ZN(
        n237) );
  AOI22_X1 U335 ( .A1(n18), .A2(regs[1166]), .B1(n48), .B2(regs[142]), .ZN(
        n236) );
  OAI211_X1 U336 ( .C1(n1), .C2(n1761), .A(n237), .B(n236), .ZN(
        curr_proc_regs[142]) );
  INV_X1 U337 ( .A(regs[1167]), .ZN(n1764) );
  AOI22_X1 U338 ( .A1(n124), .A2(regs[2191]), .B1(n68), .B2(regs[1679]), .ZN(
        n239) );
  AOI22_X1 U339 ( .A1(n55), .A2(regs[655]), .B1(n47), .B2(regs[143]), .ZN(n238) );
  OAI211_X1 U340 ( .C1(n101), .C2(n1764), .A(n239), .B(n238), .ZN(
        curr_proc_regs[143]) );
  INV_X1 U341 ( .A(regs[1168]), .ZN(n1767) );
  AOI22_X1 U342 ( .A1(n123), .A2(regs[2192]), .B1(n4), .B2(regs[1680]), .ZN(
        n241) );
  AOI22_X1 U343 ( .A1(n51), .A2(regs[656]), .B1(n47), .B2(regs[144]), .ZN(n240) );
  OAI211_X1 U344 ( .C1(n102), .C2(n1767), .A(n241), .B(n240), .ZN(
        curr_proc_regs[144]) );
  INV_X1 U345 ( .A(regs[657]), .ZN(n1770) );
  AOI22_X1 U346 ( .A1(n123), .A2(regs[2193]), .B1(n4), .B2(regs[1681]), .ZN(
        n243) );
  AOI22_X1 U347 ( .A1(n93), .A2(regs[1169]), .B1(n47), .B2(regs[145]), .ZN(
        n242) );
  OAI211_X1 U348 ( .C1(n63), .C2(n1770), .A(n243), .B(n242), .ZN(
        curr_proc_regs[145]) );
  INV_X1 U349 ( .A(regs[1170]), .ZN(n1773) );
  AOI22_X1 U350 ( .A1(n123), .A2(regs[2194]), .B1(n66), .B2(regs[1682]), .ZN(
        n245) );
  AOI22_X1 U351 ( .A1(n58), .A2(regs[658]), .B1(n47), .B2(regs[146]), .ZN(n244) );
  OAI211_X1 U352 ( .C1(n100), .C2(n1773), .A(n245), .B(n244), .ZN(
        curr_proc_regs[146]) );
  INV_X1 U353 ( .A(regs[1171]), .ZN(n1776) );
  AOI22_X1 U354 ( .A1(n123), .A2(regs[2195]), .B1(n68), .B2(regs[1683]), .ZN(
        n247) );
  AOI22_X1 U355 ( .A1(n2), .A2(regs[659]), .B1(n47), .B2(regs[147]), .ZN(n246)
         );
  OAI211_X1 U356 ( .C1(n99), .C2(n1776), .A(n247), .B(n246), .ZN(
        curr_proc_regs[147]) );
  INV_X1 U357 ( .A(regs[660]), .ZN(n1782) );
  AOI22_X1 U358 ( .A1(n123), .A2(regs[2196]), .B1(n66), .B2(regs[1684]), .ZN(
        n249) );
  AOI22_X1 U359 ( .A1(n93), .A2(regs[1172]), .B1(n47), .B2(regs[148]), .ZN(
        n248) );
  OAI211_X1 U360 ( .C1(n1), .C2(n1782), .A(n249), .B(n248), .ZN(
        curr_proc_regs[148]) );
  INV_X1 U361 ( .A(regs[1173]), .ZN(n1785) );
  AOI22_X1 U362 ( .A1(n123), .A2(regs[2197]), .B1(n15), .B2(regs[1685]), .ZN(
        n251) );
  AOI22_X1 U363 ( .A1(n55), .A2(regs[661]), .B1(n47), .B2(regs[149]), .ZN(n250) );
  OAI211_X1 U364 ( .C1(n102), .C2(n1785), .A(n251), .B(n250), .ZN(
        curr_proc_regs[149]) );
  INV_X1 U365 ( .A(regs[1038]), .ZN(n1357) );
  AOI22_X1 U366 ( .A1(n123), .A2(regs[2062]), .B1(n15), .B2(regs[1550]), .ZN(
        n253) );
  AOI22_X1 U367 ( .A1(n50), .A2(regs[526]), .B1(n27), .B2(regs[14]), .ZN(n252)
         );
  OAI211_X1 U368 ( .C1(n100), .C2(n1357), .A(n253), .B(n252), .ZN(
        curr_proc_regs[14]) );
  INV_X1 U369 ( .A(regs[1174]), .ZN(n1788) );
  AOI22_X1 U370 ( .A1(n123), .A2(regs[2198]), .B1(n68), .B2(regs[1686]), .ZN(
        n255) );
  AOI22_X1 U371 ( .A1(n51), .A2(regs[662]), .B1(n27), .B2(regs[150]), .ZN(n254) );
  OAI211_X1 U372 ( .C1(n99), .C2(n1788), .A(n255), .B(n254), .ZN(
        curr_proc_regs[150]) );
  INV_X1 U373 ( .A(regs[1175]), .ZN(n1791) );
  AOI22_X1 U374 ( .A1(n123), .A2(regs[2199]), .B1(n68), .B2(regs[1687]), .ZN(
        n257) );
  AOI22_X1 U375 ( .A1(n57), .A2(regs[663]), .B1(n27), .B2(regs[151]), .ZN(n256) );
  OAI211_X1 U376 ( .C1(n102), .C2(n1791), .A(n257), .B(n256), .ZN(
        curr_proc_regs[151]) );
  INV_X1 U377 ( .A(regs[664]), .ZN(n1794) );
  AOI22_X1 U378 ( .A1(n123), .A2(regs[2200]), .B1(n68), .B2(regs[1688]), .ZN(
        n259) );
  AOI22_X1 U379 ( .A1(n93), .A2(regs[1176]), .B1(n26), .B2(regs[152]), .ZN(
        n258) );
  OAI211_X1 U380 ( .C1(n1), .C2(n1794), .A(n259), .B(n258), .ZN(
        curr_proc_regs[152]) );
  INV_X1 U381 ( .A(regs[665]), .ZN(n1797) );
  AOI22_X1 U382 ( .A1(n123), .A2(regs[2201]), .B1(n4), .B2(regs[1689]), .ZN(
        n261) );
  AOI22_X1 U383 ( .A1(n93), .A2(regs[1177]), .B1(n48), .B2(regs[153]), .ZN(
        n260) );
  OAI211_X1 U384 ( .C1(n1), .C2(n1797), .A(n261), .B(n260), .ZN(
        curr_proc_regs[153]) );
  INV_X1 U385 ( .A(regs[666]), .ZN(n1800) );
  AOI22_X1 U386 ( .A1(n122), .A2(regs[2202]), .B1(n66), .B2(regs[1690]), .ZN(
        n263) );
  AOI22_X1 U387 ( .A1(n93), .A2(regs[1178]), .B1(n48), .B2(regs[154]), .ZN(
        n262) );
  OAI211_X1 U388 ( .C1(n64), .C2(n1800), .A(n263), .B(n262), .ZN(
        curr_proc_regs[154]) );
  INV_X1 U389 ( .A(regs[667]), .ZN(n1803) );
  AOI22_X1 U390 ( .A1(n122), .A2(regs[2203]), .B1(n15), .B2(regs[1691]), .ZN(
        n265) );
  AOI22_X1 U391 ( .A1(n93), .A2(regs[1179]), .B1(n48), .B2(regs[155]), .ZN(
        n264) );
  OAI211_X1 U392 ( .C1(n2207), .C2(n1803), .A(n265), .B(n264), .ZN(
        curr_proc_regs[155]) );
  INV_X1 U393 ( .A(regs[668]), .ZN(n1806) );
  AOI22_X1 U394 ( .A1(n122), .A2(regs[2204]), .B1(n15), .B2(regs[1692]), .ZN(
        n267) );
  AOI22_X1 U395 ( .A1(n93), .A2(regs[1180]), .B1(n48), .B2(regs[156]), .ZN(
        n266) );
  OAI211_X1 U396 ( .C1(n65), .C2(n1806), .A(n267), .B(n266), .ZN(
        curr_proc_regs[156]) );
  INV_X1 U397 ( .A(regs[669]), .ZN(n1809) );
  AOI22_X1 U398 ( .A1(n122), .A2(regs[2205]), .B1(n4), .B2(regs[1693]), .ZN(
        n269) );
  AOI22_X1 U399 ( .A1(n93), .A2(regs[1181]), .B1(n48), .B2(regs[157]), .ZN(
        n268) );
  OAI211_X1 U400 ( .C1(n65), .C2(n1809), .A(n269), .B(n268), .ZN(
        curr_proc_regs[157]) );
  INV_X1 U401 ( .A(regs[1182]), .ZN(n1815) );
  AOI22_X1 U402 ( .A1(n122), .A2(regs[2206]), .B1(n68), .B2(regs[1694]), .ZN(
        n271) );
  AOI22_X1 U403 ( .A1(n55), .A2(regs[670]), .B1(n48), .B2(regs[158]), .ZN(n270) );
  OAI211_X1 U404 ( .C1(n2221), .C2(n1815), .A(n271), .B(n270), .ZN(
        curr_proc_regs[158]) );
  INV_X1 U405 ( .A(regs[1183]), .ZN(n1818) );
  AOI22_X1 U406 ( .A1(n122), .A2(regs[2207]), .B1(n68), .B2(regs[1695]), .ZN(
        n273) );
  AOI22_X1 U407 ( .A1(n50), .A2(regs[671]), .B1(n48), .B2(regs[159]), .ZN(n272) );
  OAI211_X1 U408 ( .C1(n2221), .C2(n1818), .A(n273), .B(n272), .ZN(
        curr_proc_regs[159]) );
  INV_X1 U409 ( .A(regs[1039]), .ZN(n1360) );
  AOI22_X1 U410 ( .A1(n122), .A2(regs[2063]), .B1(n66), .B2(regs[1551]), .ZN(
        n275) );
  AOI22_X1 U411 ( .A1(n51), .A2(regs[527]), .B1(n27), .B2(regs[15]), .ZN(n274)
         );
  OAI211_X1 U412 ( .C1(n2221), .C2(n1360), .A(n275), .B(n274), .ZN(
        curr_proc_regs[15]) );
  INV_X1 U413 ( .A(regs[1184]), .ZN(n1821) );
  AOI22_X1 U414 ( .A1(n122), .A2(regs[2208]), .B1(n15), .B2(regs[1696]), .ZN(
        n277) );
  AOI22_X1 U415 ( .A1(n10), .A2(regs[672]), .B1(n47), .B2(regs[160]), .ZN(n276) );
  OAI211_X1 U416 ( .C1(n2221), .C2(n1821), .A(n277), .B(n276), .ZN(
        curr_proc_regs[160]) );
  INV_X1 U417 ( .A(regs[673]), .ZN(n1824) );
  AOI22_X1 U418 ( .A1(n122), .A2(regs[2209]), .B1(n15), .B2(regs[1697]), .ZN(
        n279) );
  AOI22_X1 U419 ( .A1(n93), .A2(regs[1185]), .B1(n26), .B2(regs[161]), .ZN(
        n278) );
  OAI211_X1 U420 ( .C1(n65), .C2(n1824), .A(n279), .B(n278), .ZN(
        curr_proc_regs[161]) );
  INV_X1 U421 ( .A(regs[1186]), .ZN(n1827) );
  AOI22_X1 U422 ( .A1(n122), .A2(regs[2210]), .B1(n68), .B2(regs[1698]), .ZN(
        n281) );
  AOI22_X1 U423 ( .A1(n10), .A2(regs[674]), .B1(n27), .B2(regs[162]), .ZN(n280) );
  OAI211_X1 U424 ( .C1(n2221), .C2(n1827), .A(n281), .B(n280), .ZN(
        curr_proc_regs[162]) );
  INV_X1 U425 ( .A(regs[1187]), .ZN(n1830) );
  AOI22_X1 U426 ( .A1(n122), .A2(regs[2211]), .B1(n4), .B2(regs[1699]), .ZN(
        n283) );
  AOI22_X1 U427 ( .A1(n10), .A2(regs[675]), .B1(n26), .B2(regs[163]), .ZN(n282) );
  OAI211_X1 U428 ( .C1(n2221), .C2(n1830), .A(n283), .B(n282), .ZN(
        curr_proc_regs[163]) );
  INV_X1 U429 ( .A(regs[676]), .ZN(n1833) );
  AOI22_X1 U430 ( .A1(n6), .A2(regs[2212]), .B1(n68), .B2(regs[1700]), .ZN(
        n285) );
  AOI22_X1 U431 ( .A1(n93), .A2(regs[1188]), .B1(n44), .B2(regs[164]), .ZN(
        n284) );
  OAI211_X1 U432 ( .C1(n65), .C2(n1833), .A(n285), .B(n284), .ZN(
        curr_proc_regs[164]) );
  INV_X1 U433 ( .A(regs[1189]), .ZN(n1836) );
  AOI22_X1 U434 ( .A1(n21), .A2(regs[2213]), .B1(n66), .B2(regs[1701]), .ZN(
        n287) );
  AOI22_X1 U435 ( .A1(n51), .A2(regs[677]), .B1(n39), .B2(regs[165]), .ZN(n286) );
  OAI211_X1 U436 ( .C1(n2221), .C2(n1836), .A(n287), .B(n286), .ZN(
        curr_proc_regs[165]) );
  INV_X1 U437 ( .A(regs[678]), .ZN(n1839) );
  AOI22_X1 U438 ( .A1(n21), .A2(regs[2214]), .B1(n15), .B2(regs[1702]), .ZN(
        n289) );
  AOI22_X1 U439 ( .A1(n89), .A2(regs[1190]), .B1(n41), .B2(regs[166]), .ZN(
        n288) );
  OAI211_X1 U440 ( .C1(n65), .C2(n1839), .A(n289), .B(n288), .ZN(
        curr_proc_regs[166]) );
  INV_X1 U441 ( .A(regs[679]), .ZN(n1842) );
  AOI22_X1 U442 ( .A1(n121), .A2(regs[2215]), .B1(n15), .B2(regs[1703]), .ZN(
        n291) );
  AOI22_X1 U443 ( .A1(n18), .A2(regs[1191]), .B1(n45), .B2(regs[167]), .ZN(
        n290) );
  OAI211_X1 U444 ( .C1(n65), .C2(n1842), .A(n291), .B(n290), .ZN(
        curr_proc_regs[167]) );
  INV_X1 U445 ( .A(regs[680]), .ZN(n1848) );
  AOI22_X1 U446 ( .A1(n21), .A2(regs[2216]), .B1(n72), .B2(regs[1704]), .ZN(
        n293) );
  AOI22_X1 U447 ( .A1(n91), .A2(regs[1192]), .B1(n44), .B2(regs[168]), .ZN(
        n292) );
  OAI211_X1 U448 ( .C1(n65), .C2(n1848), .A(n293), .B(n292), .ZN(
        curr_proc_regs[168]) );
  INV_X1 U449 ( .A(regs[1193]), .ZN(n1851) );
  AOI22_X1 U450 ( .A1(n103), .A2(regs[2217]), .B1(n4), .B2(regs[1705]), .ZN(
        n295) );
  AOI22_X1 U451 ( .A1(n51), .A2(regs[681]), .B1(n39), .B2(regs[169]), .ZN(n294) );
  OAI211_X1 U452 ( .C1(n102), .C2(n1851), .A(n295), .B(n294), .ZN(
        curr_proc_regs[169]) );
  INV_X1 U453 ( .A(regs[1040]), .ZN(n1363) );
  AOI22_X1 U454 ( .A1(n103), .A2(regs[2064]), .B1(n66), .B2(regs[1552]), .ZN(
        n297) );
  AOI22_X1 U455 ( .A1(n51), .A2(regs[528]), .B1(n29), .B2(regs[16]), .ZN(n296)
         );
  OAI211_X1 U456 ( .C1(n100), .C2(n1363), .A(n297), .B(n296), .ZN(
        curr_proc_regs[16]) );
  INV_X1 U457 ( .A(regs[1194]), .ZN(n1854) );
  AOI22_X1 U458 ( .A1(n21), .A2(regs[2218]), .B1(n66), .B2(regs[1706]), .ZN(
        n299) );
  AOI22_X1 U459 ( .A1(n51), .A2(regs[682]), .B1(n29), .B2(regs[170]), .ZN(n298) );
  OAI211_X1 U460 ( .C1(n100), .C2(n1854), .A(n299), .B(n298), .ZN(
        curr_proc_regs[170]) );
  INV_X1 U461 ( .A(regs[1195]), .ZN(n1857) );
  AOI22_X1 U462 ( .A1(n103), .A2(regs[2219]), .B1(n66), .B2(regs[1707]), .ZN(
        n301) );
  AOI22_X1 U463 ( .A1(n51), .A2(regs[683]), .B1(n31), .B2(regs[171]), .ZN(n300) );
  OAI211_X1 U464 ( .C1(n99), .C2(n1857), .A(n301), .B(n300), .ZN(
        curr_proc_regs[171]) );
  INV_X1 U465 ( .A(regs[1196]), .ZN(n1860) );
  AOI22_X1 U466 ( .A1(n6), .A2(regs[2220]), .B1(n66), .B2(regs[1708]), .ZN(
        n303) );
  AOI22_X1 U467 ( .A1(n51), .A2(regs[684]), .B1(n30), .B2(regs[172]), .ZN(n302) );
  OAI211_X1 U468 ( .C1(n102), .C2(n1860), .A(n303), .B(n302), .ZN(
        curr_proc_regs[172]) );
  INV_X1 U469 ( .A(regs[1197]), .ZN(n1863) );
  AOI22_X1 U470 ( .A1(n21), .A2(regs[2221]), .B1(n66), .B2(regs[1709]), .ZN(
        n305) );
  AOI22_X1 U471 ( .A1(n51), .A2(regs[685]), .B1(n34), .B2(regs[173]), .ZN(n304) );
  OAI211_X1 U472 ( .C1(n99), .C2(n1863), .A(n305), .B(n304), .ZN(
        curr_proc_regs[173]) );
  INV_X1 U473 ( .A(regs[686]), .ZN(n1866) );
  AOI22_X1 U474 ( .A1(n121), .A2(regs[2222]), .B1(n66), .B2(regs[1710]), .ZN(
        n307) );
  AOI22_X1 U475 ( .A1(n18), .A2(regs[1198]), .B1(n32), .B2(regs[174]), .ZN(
        n306) );
  OAI211_X1 U476 ( .C1(n1), .C2(n1866), .A(n307), .B(n306), .ZN(
        curr_proc_regs[174]) );
  INV_X1 U477 ( .A(regs[687]), .ZN(n1869) );
  AOI22_X1 U478 ( .A1(n121), .A2(regs[2223]), .B1(n66), .B2(regs[1711]), .ZN(
        n309) );
  AOI22_X1 U479 ( .A1(n88), .A2(regs[1199]), .B1(n41), .B2(regs[175]), .ZN(
        n308) );
  OAI211_X1 U480 ( .C1(n1), .C2(n1869), .A(n309), .B(n308), .ZN(
        curr_proc_regs[175]) );
  INV_X1 U481 ( .A(regs[1200]), .ZN(n1872) );
  AOI22_X1 U482 ( .A1(n6), .A2(regs[2224]), .B1(n66), .B2(regs[1712]), .ZN(
        n311) );
  AOI22_X1 U483 ( .A1(n51), .A2(regs[688]), .B1(n43), .B2(regs[176]), .ZN(n310) );
  OAI211_X1 U484 ( .C1(n99), .C2(n1872), .A(n311), .B(n310), .ZN(
        curr_proc_regs[176]) );
  INV_X1 U485 ( .A(regs[689]), .ZN(n1875) );
  AOI22_X1 U486 ( .A1(n6), .A2(regs[2225]), .B1(n66), .B2(regs[1713]), .ZN(
        n313) );
  AOI22_X1 U487 ( .A1(n90), .A2(regs[1201]), .B1(n3), .B2(regs[177]), .ZN(n312) );
  OAI211_X1 U488 ( .C1(n1), .C2(n1875), .A(n313), .B(n312), .ZN(
        curr_proc_regs[177]) );
  INV_X1 U489 ( .A(regs[1202]), .ZN(n1881) );
  AOI22_X1 U490 ( .A1(n103), .A2(regs[2226]), .B1(n66), .B2(regs[1714]), .ZN(
        n315) );
  AOI22_X1 U491 ( .A1(n50), .A2(regs[690]), .B1(n3), .B2(regs[178]), .ZN(n314)
         );
  OAI211_X1 U492 ( .C1(n16), .C2(n1881), .A(n315), .B(n314), .ZN(
        curr_proc_regs[178]) );
  INV_X1 U493 ( .A(regs[691]), .ZN(n1884) );
  AOI22_X1 U494 ( .A1(n6), .A2(regs[2227]), .B1(n66), .B2(regs[1715]), .ZN(
        n317) );
  AOI22_X1 U495 ( .A1(n18), .A2(regs[1203]), .B1(n12), .B2(regs[179]), .ZN(
        n316) );
  OAI211_X1 U496 ( .C1(n1), .C2(n1884), .A(n317), .B(n316), .ZN(
        curr_proc_regs[179]) );
  INV_X1 U497 ( .A(regs[1041]), .ZN(n1366) );
  AOI22_X1 U498 ( .A1(n21), .A2(regs[2065]), .B1(n67), .B2(regs[1553]), .ZN(
        n319) );
  AOI22_X1 U499 ( .A1(n50), .A2(regs[529]), .B1(n32), .B2(regs[17]), .ZN(n318)
         );
  OAI211_X1 U500 ( .C1(n16), .C2(n1366), .A(n319), .B(n318), .ZN(
        curr_proc_regs[17]) );
  INV_X1 U501 ( .A(regs[692]), .ZN(n1887) );
  AOI22_X1 U502 ( .A1(n21), .A2(regs[2228]), .B1(n67), .B2(regs[1716]), .ZN(
        n321) );
  AOI22_X1 U503 ( .A1(n89), .A2(regs[1204]), .B1(n41), .B2(regs[180]), .ZN(
        n320) );
  OAI211_X1 U504 ( .C1(n1), .C2(n1887), .A(n321), .B(n320), .ZN(
        curr_proc_regs[180]) );
  INV_X1 U505 ( .A(regs[693]), .ZN(n1890) );
  AOI22_X1 U506 ( .A1(n121), .A2(regs[2229]), .B1(n67), .B2(regs[1717]), .ZN(
        n323) );
  AOI22_X1 U507 ( .A1(n93), .A2(regs[1205]), .B1(n43), .B2(regs[181]), .ZN(
        n322) );
  OAI211_X1 U508 ( .C1(n1), .C2(n1890), .A(n323), .B(n322), .ZN(
        curr_proc_regs[181]) );
  INV_X1 U509 ( .A(regs[694]), .ZN(n1893) );
  AOI22_X1 U510 ( .A1(n103), .A2(regs[2230]), .B1(n67), .B2(regs[1718]), .ZN(
        n325) );
  AOI22_X1 U511 ( .A1(n18), .A2(regs[1206]), .B1(n3), .B2(regs[182]), .ZN(n324) );
  OAI211_X1 U512 ( .C1(n1), .C2(n1893), .A(n325), .B(n324), .ZN(
        curr_proc_regs[182]) );
  INV_X1 U513 ( .A(regs[695]), .ZN(n1896) );
  AOI22_X1 U514 ( .A1(n21), .A2(regs[2231]), .B1(n67), .B2(regs[1719]), .ZN(
        n327) );
  AOI22_X1 U515 ( .A1(n18), .A2(regs[1207]), .B1(n36), .B2(regs[183]), .ZN(
        n326) );
  OAI211_X1 U516 ( .C1(n1), .C2(n1896), .A(n327), .B(n326), .ZN(
        curr_proc_regs[183]) );
  INV_X1 U517 ( .A(regs[696]), .ZN(n1899) );
  AOI22_X1 U518 ( .A1(n21), .A2(regs[2232]), .B1(n67), .B2(regs[1720]), .ZN(
        n329) );
  AOI22_X1 U519 ( .A1(n93), .A2(regs[1208]), .B1(n33), .B2(regs[184]), .ZN(
        n328) );
  OAI211_X1 U520 ( .C1(n1), .C2(n1899), .A(n329), .B(n328), .ZN(
        curr_proc_regs[184]) );
  INV_X1 U521 ( .A(regs[697]), .ZN(n1902) );
  AOI22_X1 U522 ( .A1(n21), .A2(regs[2233]), .B1(n67), .B2(regs[1721]), .ZN(
        n331) );
  AOI22_X1 U523 ( .A1(n88), .A2(regs[1209]), .B1(n35), .B2(regs[185]), .ZN(
        n330) );
  OAI211_X1 U524 ( .C1(n1), .C2(n1902), .A(n331), .B(n330), .ZN(
        curr_proc_regs[185]) );
  INV_X1 U525 ( .A(regs[1210]), .ZN(n1905) );
  AOI22_X1 U526 ( .A1(n126), .A2(regs[2234]), .B1(n67), .B2(regs[1722]), .ZN(
        n333) );
  AOI22_X1 U527 ( .A1(n50), .A2(regs[698]), .B1(n40), .B2(regs[186]), .ZN(n332) );
  OAI211_X1 U528 ( .C1(n16), .C2(n1905), .A(n333), .B(n332), .ZN(
        curr_proc_regs[186]) );
  INV_X1 U529 ( .A(regs[1211]), .ZN(n1908) );
  AOI22_X1 U530 ( .A1(n6), .A2(regs[2235]), .B1(n67), .B2(regs[1723]), .ZN(
        n335) );
  AOI22_X1 U531 ( .A1(n10), .A2(regs[699]), .B1(n42), .B2(regs[187]), .ZN(n334) );
  OAI211_X1 U532 ( .C1(n16), .C2(n1908), .A(n335), .B(n334), .ZN(
        curr_proc_regs[187]) );
  INV_X1 U533 ( .A(regs[700]), .ZN(n1917) );
  AOI22_X1 U534 ( .A1(n21), .A2(regs[2236]), .B1(n67), .B2(regs[1724]), .ZN(
        n337) );
  AOI22_X1 U535 ( .A1(n90), .A2(regs[1212]), .B1(n31), .B2(regs[188]), .ZN(
        n336) );
  OAI211_X1 U536 ( .C1(n1), .C2(n1917), .A(n337), .B(n336), .ZN(
        curr_proc_regs[188]) );
  INV_X1 U537 ( .A(regs[701]), .ZN(n1920) );
  AOI22_X1 U538 ( .A1(n103), .A2(regs[2237]), .B1(n67), .B2(regs[1725]), .ZN(
        n339) );
  AOI22_X1 U539 ( .A1(n89), .A2(regs[1213]), .B1(n30), .B2(regs[189]), .ZN(
        n338) );
  OAI211_X1 U540 ( .C1(n1), .C2(n1920), .A(n339), .B(n338), .ZN(
        curr_proc_regs[189]) );
  INV_X1 U541 ( .A(regs[1042]), .ZN(n1371) );
  AOI22_X1 U542 ( .A1(n6), .A2(regs[2066]), .B1(n15), .B2(regs[1554]), .ZN(
        n341) );
  AOI22_X1 U543 ( .A1(n10), .A2(regs[530]), .B1(n42), .B2(regs[18]), .ZN(n340)
         );
  OAI211_X1 U544 ( .C1(n16), .C2(n1371), .A(n341), .B(n340), .ZN(
        curr_proc_regs[18]) );
  INV_X1 U545 ( .A(regs[702]), .ZN(n1923) );
  AOI22_X1 U546 ( .A1(n21), .A2(regs[2238]), .B1(n15), .B2(regs[1726]), .ZN(
        n343) );
  AOI22_X1 U547 ( .A1(n88), .A2(regs[1214]), .B1(n31), .B2(regs[190]), .ZN(
        n342) );
  OAI211_X1 U548 ( .C1(n1), .C2(n1923), .A(n343), .B(n342), .ZN(
        curr_proc_regs[190]) );
  INV_X1 U549 ( .A(regs[703]), .ZN(n1926) );
  AOI22_X1 U550 ( .A1(n21), .A2(regs[2239]), .B1(n4), .B2(regs[1727]), .ZN(
        n345) );
  AOI22_X1 U551 ( .A1(n91), .A2(regs[1215]), .B1(n30), .B2(regs[191]), .ZN(
        n344) );
  OAI211_X1 U552 ( .C1(n1), .C2(n1926), .A(n345), .B(n344), .ZN(
        curr_proc_regs[191]) );
  INV_X1 U553 ( .A(regs[1216]), .ZN(n1929) );
  AOI22_X1 U554 ( .A1(n121), .A2(regs[2240]), .B1(n68), .B2(regs[1728]), .ZN(
        n347) );
  AOI22_X1 U555 ( .A1(n10), .A2(regs[704]), .B1(n29), .B2(regs[192]), .ZN(n346) );
  OAI211_X1 U556 ( .C1(n16), .C2(n1929), .A(n347), .B(n346), .ZN(
        curr_proc_regs[192]) );
  INV_X1 U557 ( .A(regs[1217]), .ZN(n1932) );
  AOI22_X1 U558 ( .A1(n21), .A2(regs[2241]), .B1(n66), .B2(regs[1729]), .ZN(
        n349) );
  AOI22_X1 U559 ( .A1(n10), .A2(regs[705]), .B1(n3), .B2(regs[193]), .ZN(n348)
         );
  OAI211_X1 U560 ( .C1(n16), .C2(n1932), .A(n349), .B(n348), .ZN(
        curr_proc_regs[193]) );
  INV_X1 U561 ( .A(regs[1218]), .ZN(n1935) );
  AOI22_X1 U562 ( .A1(n121), .A2(regs[2242]), .B1(n15), .B2(regs[1730]), .ZN(
        n351) );
  AOI22_X1 U563 ( .A1(n10), .A2(regs[706]), .B1(n32), .B2(regs[194]), .ZN(n350) );
  OAI211_X1 U564 ( .C1(n16), .C2(n1935), .A(n351), .B(n350), .ZN(
        curr_proc_regs[194]) );
  INV_X1 U565 ( .A(regs[1219]), .ZN(n1938) );
  AOI22_X1 U566 ( .A1(n21), .A2(regs[2243]), .B1(n9), .B2(regs[1731]), .ZN(
        n353) );
  AOI22_X1 U567 ( .A1(n10), .A2(regs[707]), .B1(n34), .B2(regs[195]), .ZN(n352) );
  OAI211_X1 U568 ( .C1(n16), .C2(n1938), .A(n353), .B(n352), .ZN(
        curr_proc_regs[195]) );
  INV_X1 U569 ( .A(regs[708]), .ZN(n1941) );
  AOI22_X1 U570 ( .A1(n103), .A2(regs[2244]), .B1(n68), .B2(regs[1732]), .ZN(
        n355) );
  AOI22_X1 U571 ( .A1(n18), .A2(regs[1220]), .B1(n34), .B2(regs[196]), .ZN(
        n354) );
  OAI211_X1 U572 ( .C1(n64), .C2(n1941), .A(n355), .B(n354), .ZN(
        curr_proc_regs[196]) );
  INV_X1 U573 ( .A(regs[1221]), .ZN(n1944) );
  AOI22_X1 U574 ( .A1(n6), .A2(regs[2245]), .B1(n9), .B2(regs[1733]), .ZN(n357) );
  AOI22_X1 U575 ( .A1(n10), .A2(regs[709]), .B1(n32), .B2(regs[197]), .ZN(n356) );
  OAI211_X1 U576 ( .C1(n16), .C2(n1944), .A(n357), .B(n356), .ZN(
        curr_proc_regs[197]) );
  INV_X1 U577 ( .A(regs[1222]), .ZN(n1950) );
  AOI22_X1 U578 ( .A1(n21), .A2(regs[2246]), .B1(n68), .B2(regs[1734]), .ZN(
        n359) );
  AOI22_X1 U579 ( .A1(n10), .A2(regs[710]), .B1(n3), .B2(regs[198]), .ZN(n358)
         );
  OAI211_X1 U580 ( .C1(n16), .C2(n1950), .A(n359), .B(n358), .ZN(
        curr_proc_regs[198]) );
  INV_X1 U581 ( .A(regs[711]), .ZN(n1953) );
  AOI22_X1 U582 ( .A1(n21), .A2(regs[2247]), .B1(n15), .B2(regs[1735]), .ZN(
        n361) );
  AOI22_X1 U583 ( .A1(n91), .A2(regs[1223]), .B1(n34), .B2(regs[199]), .ZN(
        n360) );
  OAI211_X1 U584 ( .C1(n11), .C2(n1953), .A(n361), .B(n360), .ZN(
        curr_proc_regs[199]) );
  INV_X1 U585 ( .A(regs[531]), .ZN(n1374) );
  AOI22_X1 U586 ( .A1(n121), .A2(regs[2067]), .B1(n68), .B2(regs[1555]), .ZN(
        n363) );
  AOI22_X1 U587 ( .A1(n92), .A2(regs[1043]), .B1(n44), .B2(regs[19]), .ZN(n362) );
  OAI211_X1 U588 ( .C1(n11), .C2(n1374), .A(n363), .B(n362), .ZN(
        curr_proc_regs[19]) );
  INV_X1 U589 ( .A(regs[513]), .ZN(n1319) );
  AOI22_X1 U590 ( .A1(n121), .A2(regs[2049]), .B1(n66), .B2(regs[1537]), .ZN(
        n365) );
  AOI22_X1 U591 ( .A1(n89), .A2(regs[1025]), .B1(n44), .B2(regs[1]), .ZN(n364)
         );
  OAI211_X1 U592 ( .C1(n2207), .C2(n1319), .A(n365), .B(n364), .ZN(
        curr_proc_regs[1]) );
  INV_X1 U593 ( .A(regs[1224]), .ZN(n1956) );
  AOI22_X1 U594 ( .A1(n103), .A2(regs[2248]), .B1(n15), .B2(regs[1736]), .ZN(
        n367) );
  AOI22_X1 U595 ( .A1(n49), .A2(regs[712]), .B1(n44), .B2(regs[200]), .ZN(n366) );
  OAI211_X1 U596 ( .C1(n16), .C2(n1956), .A(n367), .B(n366), .ZN(
        curr_proc_regs[200]) );
  INV_X1 U597 ( .A(regs[1225]), .ZN(n1959) );
  AOI22_X1 U598 ( .A1(n6), .A2(regs[2249]), .B1(n9), .B2(regs[1737]), .ZN(n369) );
  AOI22_X1 U599 ( .A1(n49), .A2(regs[713]), .B1(n44), .B2(regs[201]), .ZN(n368) );
  OAI211_X1 U600 ( .C1(n16), .C2(n1959), .A(n369), .B(n368), .ZN(
        curr_proc_regs[201]) );
  INV_X1 U601 ( .A(regs[714]), .ZN(n1962) );
  AOI22_X1 U602 ( .A1(n21), .A2(regs[2250]), .B1(n68), .B2(regs[1738]), .ZN(
        n371) );
  AOI22_X1 U603 ( .A1(n91), .A2(regs[1226]), .B1(n29), .B2(regs[202]), .ZN(
        n370) );
  OAI211_X1 U604 ( .C1(n11), .C2(n1962), .A(n371), .B(n370), .ZN(
        curr_proc_regs[202]) );
  INV_X1 U605 ( .A(regs[715]), .ZN(n1965) );
  AOI22_X1 U606 ( .A1(n103), .A2(regs[2251]), .B1(n68), .B2(regs[1739]), .ZN(
        n373) );
  AOI22_X1 U607 ( .A1(n18), .A2(regs[1227]), .B1(n36), .B2(regs[203]), .ZN(
        n372) );
  OAI211_X1 U608 ( .C1(n64), .C2(n1965), .A(n373), .B(n372), .ZN(
        curr_proc_regs[203]) );
  INV_X1 U609 ( .A(regs[1228]), .ZN(n1968) );
  AOI22_X1 U610 ( .A1(n6), .A2(regs[2252]), .B1(n4), .B2(regs[1740]), .ZN(n375) );
  AOI22_X1 U611 ( .A1(n49), .A2(regs[716]), .B1(n30), .B2(regs[204]), .ZN(n374) );
  OAI211_X1 U612 ( .C1(n16), .C2(n1968), .A(n375), .B(n374), .ZN(
        curr_proc_regs[204]) );
  INV_X1 U613 ( .A(regs[1229]), .ZN(n1971) );
  AOI22_X1 U614 ( .A1(n21), .A2(regs[2253]), .B1(n9), .B2(regs[1741]), .ZN(
        n377) );
  AOI22_X1 U615 ( .A1(n50), .A2(regs[717]), .B1(n36), .B2(regs[205]), .ZN(n376) );
  OAI211_X1 U616 ( .C1(n99), .C2(n1971), .A(n377), .B(n376), .ZN(
        curr_proc_regs[205]) );
  INV_X1 U617 ( .A(regs[718]), .ZN(n1974) );
  AOI22_X1 U618 ( .A1(n21), .A2(regs[2254]), .B1(n4), .B2(regs[1742]), .ZN(
        n379) );
  AOI22_X1 U619 ( .A1(n18), .A2(regs[1230]), .B1(n33), .B2(regs[206]), .ZN(
        n378) );
  OAI211_X1 U620 ( .C1(n2207), .C2(n1974), .A(n379), .B(n378), .ZN(
        curr_proc_regs[206]) );
  INV_X1 U621 ( .A(regs[719]), .ZN(n1977) );
  AOI22_X1 U622 ( .A1(n121), .A2(regs[2255]), .B1(n4), .B2(regs[1743]), .ZN(
        n381) );
  AOI22_X1 U623 ( .A1(n92), .A2(regs[1231]), .B1(n35), .B2(regs[207]), .ZN(
        n380) );
  OAI211_X1 U624 ( .C1(n11), .C2(n1977), .A(n381), .B(n380), .ZN(
        curr_proc_regs[207]) );
  INV_X1 U625 ( .A(regs[1232]), .ZN(n1983) );
  AOI22_X1 U626 ( .A1(n103), .A2(regs[2256]), .B1(n66), .B2(regs[1744]), .ZN(
        n383) );
  AOI22_X1 U627 ( .A1(n50), .A2(regs[720]), .B1(n40), .B2(regs[208]), .ZN(n382) );
  OAI211_X1 U628 ( .C1(n99), .C2(n1983), .A(n383), .B(n382), .ZN(
        curr_proc_regs[208]) );
  INV_X1 U629 ( .A(regs[1233]), .ZN(n1986) );
  AOI22_X1 U630 ( .A1(n6), .A2(regs[2257]), .B1(n68), .B2(regs[1745]), .ZN(
        n385) );
  AOI22_X1 U631 ( .A1(n50), .A2(regs[721]), .B1(n32), .B2(regs[209]), .ZN(n384) );
  OAI211_X1 U632 ( .C1(n99), .C2(n1986), .A(n385), .B(n384), .ZN(
        curr_proc_regs[209]) );
  INV_X1 U633 ( .A(regs[1044]), .ZN(n1377) );
  AOI22_X1 U634 ( .A1(n21), .A2(regs[2068]), .B1(n15), .B2(regs[1556]), .ZN(
        n387) );
  AOI22_X1 U635 ( .A1(n50), .A2(regs[532]), .B1(n32), .B2(regs[20]), .ZN(n386)
         );
  OAI211_X1 U636 ( .C1(n99), .C2(n1377), .A(n387), .B(n386), .ZN(
        curr_proc_regs[20]) );
  INV_X1 U637 ( .A(regs[1234]), .ZN(n1989) );
  AOI22_X1 U638 ( .A1(n21), .A2(regs[2258]), .B1(n15), .B2(regs[1746]), .ZN(
        n389) );
  AOI22_X1 U639 ( .A1(n50), .A2(regs[722]), .B1(n41), .B2(regs[210]), .ZN(n388) );
  OAI211_X1 U640 ( .C1(n99), .C2(n1989), .A(n389), .B(n388), .ZN(
        curr_proc_regs[210]) );
  INV_X1 U641 ( .A(regs[1235]), .ZN(n1992) );
  AOI22_X1 U642 ( .A1(n121), .A2(regs[2259]), .B1(n9), .B2(regs[1747]), .ZN(
        n391) );
  AOI22_X1 U643 ( .A1(n50), .A2(regs[723]), .B1(n34), .B2(regs[211]), .ZN(n390) );
  OAI211_X1 U644 ( .C1(n99), .C2(n1992), .A(n391), .B(n390), .ZN(
        curr_proc_regs[211]) );
  INV_X1 U645 ( .A(regs[724]), .ZN(n1995) );
  AOI22_X1 U646 ( .A1(n103), .A2(regs[2260]), .B1(n68), .B2(regs[1748]), .ZN(
        n393) );
  AOI22_X1 U647 ( .A1(n93), .A2(regs[1236]), .B1(n44), .B2(regs[212]), .ZN(
        n392) );
  OAI211_X1 U648 ( .C1(n64), .C2(n1995), .A(n393), .B(n392), .ZN(
        curr_proc_regs[212]) );
  INV_X1 U649 ( .A(regs[1237]), .ZN(n1998) );
  AOI22_X1 U650 ( .A1(n121), .A2(regs[2261]), .B1(n68), .B2(regs[1749]), .ZN(
        n395) );
  AOI22_X1 U651 ( .A1(n50), .A2(regs[725]), .B1(n44), .B2(regs[213]), .ZN(n394) );
  OAI211_X1 U652 ( .C1(n99), .C2(n1998), .A(n395), .B(n394), .ZN(
        curr_proc_regs[213]) );
  INV_X1 U653 ( .A(regs[1238]), .ZN(n2001) );
  AOI22_X1 U654 ( .A1(n121), .A2(regs[2262]), .B1(n4), .B2(regs[1750]), .ZN(
        n397) );
  AOI22_X1 U655 ( .A1(n50), .A2(regs[726]), .B1(n44), .B2(regs[214]), .ZN(n396) );
  OAI211_X1 U656 ( .C1(n16), .C2(n2001), .A(n397), .B(n396), .ZN(
        curr_proc_regs[214]) );
  INV_X1 U657 ( .A(regs[1239]), .ZN(n2004) );
  AOI22_X1 U658 ( .A1(n121), .A2(regs[2263]), .B1(n4), .B2(regs[1751]), .ZN(
        n399) );
  AOI22_X1 U659 ( .A1(n10), .A2(regs[727]), .B1(n44), .B2(regs[215]), .ZN(n398) );
  OAI211_X1 U660 ( .C1(n16), .C2(n2004), .A(n399), .B(n398), .ZN(
        curr_proc_regs[215]) );
  INV_X1 U661 ( .A(regs[1240]), .ZN(n2007) );
  AOI22_X1 U662 ( .A1(n121), .A2(regs[2264]), .B1(n4), .B2(regs[1752]), .ZN(
        n401) );
  AOI22_X1 U663 ( .A1(n10), .A2(regs[728]), .B1(n44), .B2(regs[216]), .ZN(n400) );
  OAI211_X1 U664 ( .C1(n99), .C2(n2007), .A(n401), .B(n400), .ZN(
        curr_proc_regs[216]) );
  INV_X1 U665 ( .A(regs[1241]), .ZN(n2010) );
  AOI22_X1 U666 ( .A1(n121), .A2(regs[2265]), .B1(n4), .B2(regs[1753]), .ZN(
        n403) );
  AOI22_X1 U667 ( .A1(n10), .A2(regs[729]), .B1(n44), .B2(regs[217]), .ZN(n402) );
  OAI211_X1 U668 ( .C1(n100), .C2(n2010), .A(n403), .B(n402), .ZN(
        curr_proc_regs[217]) );
  INV_X1 U669 ( .A(regs[1242]), .ZN(n2016) );
  AOI22_X1 U670 ( .A1(n121), .A2(regs[2266]), .B1(n68), .B2(regs[1754]), .ZN(
        n405) );
  AOI22_X1 U671 ( .A1(n49), .A2(regs[730]), .B1(n44), .B2(regs[218]), .ZN(n404) );
  OAI211_X1 U672 ( .C1(n101), .C2(n2016), .A(n405), .B(n404), .ZN(
        curr_proc_regs[218]) );
  INV_X1 U673 ( .A(regs[731]), .ZN(n2019) );
  AOI22_X1 U674 ( .A1(n121), .A2(regs[2267]), .B1(n9), .B2(regs[1755]), .ZN(
        n407) );
  AOI22_X1 U675 ( .A1(n91), .A2(regs[1243]), .B1(n29), .B2(regs[219]), .ZN(
        n406) );
  OAI211_X1 U676 ( .C1(n2207), .C2(n2019), .A(n407), .B(n406), .ZN(
        curr_proc_regs[219]) );
  INV_X1 U677 ( .A(regs[533]), .ZN(n1380) );
  AOI22_X1 U678 ( .A1(n121), .A2(regs[2069]), .B1(n71), .B2(regs[1557]), .ZN(
        n409) );
  AOI22_X1 U679 ( .A1(n18), .A2(regs[1045]), .B1(n36), .B2(regs[21]), .ZN(n408) );
  OAI211_X1 U680 ( .C1(n2207), .C2(n1380), .A(n409), .B(n408), .ZN(
        curr_proc_regs[21]) );
  INV_X1 U681 ( .A(regs[732]), .ZN(n2022) );
  AOI22_X1 U682 ( .A1(n121), .A2(regs[2268]), .B1(n9), .B2(regs[1756]), .ZN(
        n411) );
  AOI22_X1 U683 ( .A1(n88), .A2(regs[1244]), .B1(n33), .B2(regs[220]), .ZN(
        n410) );
  OAI211_X1 U684 ( .C1(n2207), .C2(n2022), .A(n411), .B(n410), .ZN(
        curr_proc_regs[220]) );
  INV_X1 U685 ( .A(regs[1245]), .ZN(n2025) );
  AOI22_X1 U686 ( .A1(n121), .A2(regs[2269]), .B1(n71), .B2(regs[1757]), .ZN(
        n413) );
  AOI22_X1 U687 ( .A1(n49), .A2(regs[733]), .B1(n36), .B2(regs[221]), .ZN(n412) );
  OAI211_X1 U688 ( .C1(n2221), .C2(n2025), .A(n413), .B(n412), .ZN(
        curr_proc_regs[221]) );
  INV_X1 U689 ( .A(regs[734]), .ZN(n2028) );
  AOI22_X1 U690 ( .A1(n121), .A2(regs[2270]), .B1(n9), .B2(regs[1758]), .ZN(
        n415) );
  AOI22_X1 U691 ( .A1(n90), .A2(regs[1246]), .B1(n12), .B2(regs[222]), .ZN(
        n414) );
  OAI211_X1 U692 ( .C1(n2207), .C2(n2028), .A(n415), .B(n414), .ZN(
        curr_proc_regs[222]) );
  INV_X1 U693 ( .A(regs[735]), .ZN(n2031) );
  AOI22_X1 U694 ( .A1(n119), .A2(regs[2271]), .B1(n9), .B2(regs[1759]), .ZN(
        n417) );
  AOI22_X1 U695 ( .A1(n90), .A2(regs[1247]), .B1(n12), .B2(regs[223]), .ZN(
        n416) );
  OAI211_X1 U696 ( .C1(n2207), .C2(n2031), .A(n417), .B(n416), .ZN(
        curr_proc_regs[223]) );
  INV_X1 U697 ( .A(regs[1248]), .ZN(n2034) );
  AOI22_X1 U698 ( .A1(n118), .A2(regs[2272]), .B1(n9), .B2(regs[1760]), .ZN(
        n419) );
  AOI22_X1 U699 ( .A1(n49), .A2(regs[736]), .B1(n28), .B2(regs[224]), .ZN(n418) );
  OAI211_X1 U700 ( .C1(n5), .C2(n2034), .A(n419), .B(n418), .ZN(
        curr_proc_regs[224]) );
  INV_X1 U701 ( .A(regs[1249]), .ZN(n2037) );
  AOI22_X1 U702 ( .A1(n120), .A2(regs[2273]), .B1(n9), .B2(regs[1761]), .ZN(
        n421) );
  AOI22_X1 U703 ( .A1(n49), .A2(regs[737]), .B1(n32), .B2(regs[225]), .ZN(n420) );
  OAI211_X1 U704 ( .C1(n5), .C2(n2037), .A(n421), .B(n420), .ZN(
        curr_proc_regs[225]) );
  INV_X1 U705 ( .A(regs[738]), .ZN(n2040) );
  AOI22_X1 U706 ( .A1(n120), .A2(regs[2274]), .B1(n9), .B2(regs[1762]), .ZN(
        n423) );
  AOI22_X1 U707 ( .A1(n18), .A2(regs[1250]), .B1(n32), .B2(regs[226]), .ZN(
        n422) );
  OAI211_X1 U708 ( .C1(n11), .C2(n2040), .A(n423), .B(n422), .ZN(
        curr_proc_regs[226]) );
  INV_X1 U709 ( .A(regs[1251]), .ZN(n2043) );
  AOI22_X1 U710 ( .A1(n118), .A2(regs[2275]), .B1(n9), .B2(regs[1763]), .ZN(
        n425) );
  AOI22_X1 U711 ( .A1(n49), .A2(regs[739]), .B1(n12), .B2(regs[227]), .ZN(n424) );
  OAI211_X1 U712 ( .C1(n5), .C2(n2043), .A(n425), .B(n424), .ZN(
        curr_proc_regs[227]) );
  INV_X1 U713 ( .A(regs[1252]), .ZN(n2049) );
  AOI22_X1 U714 ( .A1(n119), .A2(regs[2276]), .B1(n9), .B2(regs[1764]), .ZN(
        n427) );
  AOI22_X1 U715 ( .A1(n49), .A2(regs[740]), .B1(n41), .B2(regs[228]), .ZN(n426) );
  OAI211_X1 U716 ( .C1(n5), .C2(n2049), .A(n427), .B(n426), .ZN(
        curr_proc_regs[228]) );
  INV_X1 U717 ( .A(regs[1253]), .ZN(n2052) );
  AOI22_X1 U718 ( .A1(n118), .A2(regs[2277]), .B1(n15), .B2(regs[1765]), .ZN(
        n429) );
  AOI22_X1 U719 ( .A1(n49), .A2(regs[741]), .B1(n35), .B2(regs[229]), .ZN(n428) );
  OAI211_X1 U720 ( .C1(n5), .C2(n2052), .A(n429), .B(n428), .ZN(
        curr_proc_regs[229]) );
  INV_X1 U721 ( .A(regs[534]), .ZN(n1383) );
  AOI22_X1 U722 ( .A1(n120), .A2(regs[2070]), .B1(n66), .B2(regs[1558]), .ZN(
        n431) );
  AOI22_X1 U723 ( .A1(n92), .A2(regs[1046]), .B1(n40), .B2(regs[22]), .ZN(n430) );
  OAI211_X1 U724 ( .C1(n11), .C2(n1383), .A(n431), .B(n430), .ZN(
        curr_proc_regs[22]) );
  INV_X1 U725 ( .A(regs[1254]), .ZN(n2055) );
  AOI22_X1 U726 ( .A1(n119), .A2(regs[2278]), .B1(n15), .B2(regs[1766]), .ZN(
        n433) );
  AOI22_X1 U727 ( .A1(n56), .A2(regs[742]), .B1(n42), .B2(regs[230]), .ZN(n432) );
  OAI211_X1 U728 ( .C1(n5), .C2(n2055), .A(n433), .B(n432), .ZN(
        curr_proc_regs[230]) );
  INV_X1 U729 ( .A(regs[1255]), .ZN(n2058) );
  AOI22_X1 U730 ( .A1(n120), .A2(regs[2279]), .B1(n15), .B2(regs[1767]), .ZN(
        n435) );
  AOI22_X1 U731 ( .A1(n10), .A2(regs[743]), .B1(n31), .B2(regs[231]), .ZN(n434) );
  OAI211_X1 U732 ( .C1(n5), .C2(n2058), .A(n435), .B(n434), .ZN(
        curr_proc_regs[231]) );
  INV_X1 U733 ( .A(regs[1256]), .ZN(n2061) );
  AOI22_X1 U734 ( .A1(n119), .A2(regs[2280]), .B1(n9), .B2(regs[1768]), .ZN(
        n437) );
  AOI22_X1 U735 ( .A1(n49), .A2(regs[744]), .B1(n36), .B2(regs[232]), .ZN(n436) );
  OAI211_X1 U736 ( .C1(n5), .C2(n2061), .A(n437), .B(n436), .ZN(
        curr_proc_regs[232]) );
  INV_X1 U737 ( .A(regs[1257]), .ZN(n2064) );
  AOI22_X1 U738 ( .A1(n118), .A2(regs[2281]), .B1(n68), .B2(regs[1769]), .ZN(
        n439) );
  AOI22_X1 U739 ( .A1(n10), .A2(regs[745]), .B1(n33), .B2(regs[233]), .ZN(n438) );
  OAI211_X1 U740 ( .C1(n101), .C2(n2064), .A(n439), .B(n438), .ZN(
        curr_proc_regs[233]) );
  INV_X1 U741 ( .A(regs[1258]), .ZN(n2067) );
  AOI22_X1 U742 ( .A1(n119), .A2(regs[2282]), .B1(n9), .B2(regs[1770]), .ZN(
        n441) );
  AOI22_X1 U743 ( .A1(n10), .A2(regs[746]), .B1(n35), .B2(regs[234]), .ZN(n440) );
  OAI211_X1 U744 ( .C1(n102), .C2(n2067), .A(n441), .B(n440), .ZN(
        curr_proc_regs[234]) );
  INV_X1 U745 ( .A(regs[747]), .ZN(n2070) );
  AOI22_X1 U746 ( .A1(n118), .A2(regs[2283]), .B1(n4), .B2(regs[1771]), .ZN(
        n443) );
  AOI22_X1 U747 ( .A1(n92), .A2(regs[1259]), .B1(n40), .B2(regs[235]), .ZN(
        n442) );
  OAI211_X1 U748 ( .C1(n64), .C2(n2070), .A(n443), .B(n442), .ZN(
        curr_proc_regs[235]) );
  INV_X1 U749 ( .A(regs[748]), .ZN(n2073) );
  AOI22_X1 U750 ( .A1(n120), .A2(regs[2284]), .B1(n15), .B2(regs[1772]), .ZN(
        n445) );
  AOI22_X1 U751 ( .A1(n92), .A2(regs[1260]), .B1(n42), .B2(regs[236]), .ZN(
        n444) );
  OAI211_X1 U752 ( .C1(n11), .C2(n2073), .A(n445), .B(n444), .ZN(
        curr_proc_regs[236]) );
  INV_X1 U753 ( .A(regs[1261]), .ZN(n2076) );
  AOI22_X1 U754 ( .A1(n120), .A2(regs[2285]), .B1(n68), .B2(regs[1773]), .ZN(
        n447) );
  AOI22_X1 U755 ( .A1(n10), .A2(regs[749]), .B1(n31), .B2(regs[237]), .ZN(n446) );
  OAI211_X1 U756 ( .C1(n101), .C2(n2076), .A(n447), .B(n446), .ZN(
        curr_proc_regs[237]) );
  INV_X1 U757 ( .A(regs[750]), .ZN(n2082) );
  AOI22_X1 U758 ( .A1(n119), .A2(regs[2286]), .B1(n4), .B2(regs[1774]), .ZN(
        n449) );
  AOI22_X1 U759 ( .A1(n92), .A2(regs[1262]), .B1(n30), .B2(regs[238]), .ZN(
        n448) );
  OAI211_X1 U760 ( .C1(n11), .C2(n2082), .A(n449), .B(n448), .ZN(
        curr_proc_regs[238]) );
  INV_X1 U761 ( .A(regs[751]), .ZN(n2085) );
  AOI22_X1 U762 ( .A1(n118), .A2(regs[2287]), .B1(n68), .B2(regs[1775]), .ZN(
        n451) );
  AOI22_X1 U763 ( .A1(n92), .A2(regs[1263]), .B1(n42), .B2(regs[239]), .ZN(
        n450) );
  OAI211_X1 U764 ( .C1(n64), .C2(n2085), .A(n451), .B(n450), .ZN(
        curr_proc_regs[239]) );
  INV_X1 U765 ( .A(regs[1047]), .ZN(n1386) );
  AOI22_X1 U766 ( .A1(n120), .A2(regs[2071]), .B1(n68), .B2(regs[1559]), .ZN(
        n453) );
  AOI22_X1 U767 ( .A1(n10), .A2(regs[535]), .B1(n36), .B2(regs[23]), .ZN(n452)
         );
  OAI211_X1 U768 ( .C1(n2221), .C2(n1386), .A(n453), .B(n452), .ZN(
        curr_proc_regs[23]) );
  INV_X1 U769 ( .A(regs[1264]), .ZN(n2088) );
  AOI22_X1 U770 ( .A1(n119), .A2(regs[2288]), .B1(n68), .B2(regs[1776]), .ZN(
        n455) );
  AOI22_X1 U771 ( .A1(n10), .A2(regs[752]), .B1(n33), .B2(regs[240]), .ZN(n454) );
  OAI211_X1 U772 ( .C1(n102), .C2(n2088), .A(n455), .B(n454), .ZN(
        curr_proc_regs[240]) );
  INV_X1 U773 ( .A(regs[753]), .ZN(n2091) );
  AOI22_X1 U774 ( .A1(n119), .A2(regs[2289]), .B1(n68), .B2(regs[1777]), .ZN(
        n457) );
  AOI22_X1 U775 ( .A1(n92), .A2(regs[1265]), .B1(n35), .B2(regs[241]), .ZN(
        n456) );
  OAI211_X1 U776 ( .C1(n11), .C2(n2091), .A(n457), .B(n456), .ZN(
        curr_proc_regs[241]) );
  INV_X1 U777 ( .A(regs[1266]), .ZN(n2094) );
  AOI22_X1 U778 ( .A1(n118), .A2(regs[2290]), .B1(n68), .B2(regs[1778]), .ZN(
        n459) );
  AOI22_X1 U779 ( .A1(n10), .A2(regs[754]), .B1(n30), .B2(regs[242]), .ZN(n458) );
  OAI211_X1 U780 ( .C1(n102), .C2(n2094), .A(n459), .B(n458), .ZN(
        curr_proc_regs[242]) );
  INV_X1 U781 ( .A(regs[755]), .ZN(n2097) );
  AOI22_X1 U782 ( .A1(n118), .A2(regs[2291]), .B1(n68), .B2(regs[1779]), .ZN(
        n461) );
  AOI22_X1 U783 ( .A1(n92), .A2(regs[1267]), .B1(n40), .B2(regs[243]), .ZN(
        n460) );
  OAI211_X1 U784 ( .C1(n11), .C2(n2097), .A(n461), .B(n460), .ZN(
        curr_proc_regs[243]) );
  INV_X1 U785 ( .A(regs[756]), .ZN(n2100) );
  AOI22_X1 U786 ( .A1(n120), .A2(regs[2292]), .B1(n68), .B2(regs[1780]), .ZN(
        n463) );
  AOI22_X1 U787 ( .A1(n91), .A2(regs[1268]), .B1(n35), .B2(regs[244]), .ZN(
        n462) );
  OAI211_X1 U788 ( .C1(n2207), .C2(n2100), .A(n463), .B(n462), .ZN(
        curr_proc_regs[244]) );
  INV_X1 U789 ( .A(regs[1269]), .ZN(n2103) );
  AOI22_X1 U790 ( .A1(n119), .A2(regs[2293]), .B1(n68), .B2(regs[1781]), .ZN(
        n465) );
  AOI22_X1 U791 ( .A1(n10), .A2(regs[757]), .B1(n40), .B2(regs[245]), .ZN(n464) );
  OAI211_X1 U792 ( .C1(n2221), .C2(n2103), .A(n465), .B(n464), .ZN(
        curr_proc_regs[245]) );
  INV_X1 U793 ( .A(regs[1270]), .ZN(n2106) );
  AOI22_X1 U794 ( .A1(n118), .A2(regs[2294]), .B1(n68), .B2(regs[1782]), .ZN(
        n467) );
  AOI22_X1 U795 ( .A1(n10), .A2(regs[758]), .B1(n30), .B2(regs[246]), .ZN(n466) );
  OAI211_X1 U796 ( .C1(n5), .C2(n2106), .A(n467), .B(n466), .ZN(
        curr_proc_regs[246]) );
  INV_X1 U797 ( .A(regs[759]), .ZN(n2109) );
  AOI22_X1 U798 ( .A1(n120), .A2(regs[2295]), .B1(n68), .B2(regs[1783]), .ZN(
        n469) );
  AOI22_X1 U799 ( .A1(n91), .A2(regs[1271]), .B1(n36), .B2(regs[247]), .ZN(
        n468) );
  OAI211_X1 U800 ( .C1(n11), .C2(n2109), .A(n469), .B(n468), .ZN(
        curr_proc_regs[247]) );
  INV_X1 U801 ( .A(regs[760]), .ZN(n2115) );
  AOI22_X1 U802 ( .A1(n119), .A2(regs[2296]), .B1(n68), .B2(regs[1784]), .ZN(
        n471) );
  AOI22_X1 U803 ( .A1(n91), .A2(regs[1272]), .B1(n33), .B2(regs[248]), .ZN(
        n470) );
  OAI211_X1 U804 ( .C1(n64), .C2(n2115), .A(n471), .B(n470), .ZN(
        curr_proc_regs[248]) );
  INV_X1 U805 ( .A(regs[761]), .ZN(n2118) );
  AOI22_X1 U806 ( .A1(n118), .A2(regs[2297]), .B1(n68), .B2(regs[1785]), .ZN(
        n473) );
  AOI22_X1 U807 ( .A1(n91), .A2(regs[1273]), .B1(n31), .B2(regs[249]), .ZN(
        n472) );
  OAI211_X1 U808 ( .C1(n11), .C2(n2118), .A(n473), .B(n472), .ZN(
        curr_proc_regs[249]) );
  INV_X1 U809 ( .A(regs[536]), .ZN(n1389) );
  AOI22_X1 U810 ( .A1(n120), .A2(regs[2072]), .B1(n66), .B2(regs[1560]), .ZN(
        n475) );
  AOI22_X1 U811 ( .A1(n91), .A2(regs[1048]), .B1(n42), .B2(regs[24]), .ZN(n474) );
  OAI211_X1 U812 ( .C1(n11), .C2(n1389), .A(n475), .B(n474), .ZN(
        curr_proc_regs[24]) );
  INV_X1 U813 ( .A(regs[762]), .ZN(n2121) );
  AOI22_X1 U814 ( .A1(n119), .A2(regs[2298]), .B1(n15), .B2(regs[1786]), .ZN(
        n477) );
  AOI22_X1 U815 ( .A1(n91), .A2(regs[1274]), .B1(n36), .B2(regs[250]), .ZN(
        n476) );
  OAI211_X1 U816 ( .C1(n11), .C2(n2121), .A(n477), .B(n476), .ZN(
        curr_proc_regs[250]) );
  INV_X1 U817 ( .A(regs[1275]), .ZN(n2124) );
  AOI22_X1 U818 ( .A1(n118), .A2(regs[2299]), .B1(n15), .B2(regs[1787]), .ZN(
        n479) );
  AOI22_X1 U819 ( .A1(n57), .A2(regs[763]), .B1(n33), .B2(regs[251]), .ZN(n478) );
  OAI211_X1 U820 ( .C1(n2221), .C2(n2124), .A(n479), .B(n478), .ZN(
        curr_proc_regs[251]) );
  INV_X1 U821 ( .A(regs[1276]), .ZN(n2127) );
  AOI22_X1 U822 ( .A1(n120), .A2(regs[2300]), .B1(n9), .B2(regs[1788]), .ZN(
        n481) );
  AOI22_X1 U823 ( .A1(n51), .A2(regs[764]), .B1(n29), .B2(regs[252]), .ZN(n480) );
  OAI211_X1 U824 ( .C1(n99), .C2(n2127), .A(n481), .B(n480), .ZN(
        curr_proc_regs[252]) );
  INV_X1 U825 ( .A(regs[765]), .ZN(n2130) );
  AOI22_X1 U826 ( .A1(n120), .A2(regs[2301]), .B1(n68), .B2(regs[1789]), .ZN(
        n483) );
  AOI22_X1 U827 ( .A1(n91), .A2(regs[1277]), .B1(n35), .B2(regs[253]), .ZN(
        n482) );
  OAI211_X1 U828 ( .C1(n11), .C2(n2130), .A(n483), .B(n482), .ZN(
        curr_proc_regs[253]) );
  INV_X1 U829 ( .A(regs[766]), .ZN(n2133) );
  AOI22_X1 U830 ( .A1(n120), .A2(regs[2302]), .B1(n68), .B2(regs[1790]), .ZN(
        n485) );
  AOI22_X1 U831 ( .A1(n91), .A2(regs[1278]), .B1(n36), .B2(regs[254]), .ZN(
        n484) );
  OAI211_X1 U832 ( .C1(n2207), .C2(n2133), .A(n485), .B(n484), .ZN(
        curr_proc_regs[254]) );
  INV_X1 U833 ( .A(regs[1279]), .ZN(n2137) );
  AOI22_X1 U834 ( .A1(n120), .A2(regs[2303]), .B1(n4), .B2(regs[1791]), .ZN(
        n487) );
  AOI22_X1 U835 ( .A1(n52), .A2(regs[767]), .B1(n33), .B2(regs[255]), .ZN(n486) );
  OAI211_X1 U836 ( .C1(n16), .C2(n2137), .A(n487), .B(n486), .ZN(
        curr_proc_regs[255]) );
  NAND2_X1 U837 ( .A1(regs[768]), .A2(n2), .ZN(n490) );
  AOI22_X1 U838 ( .A1(n91), .A2(regs[1280]), .B1(n29), .B2(regs[256]), .ZN(
        n489) );
  AOI22_X1 U839 ( .A1(n120), .A2(regs[2304]), .B1(n2217), .B2(regs[1792]), 
        .ZN(n488) );
  NAND3_X1 U840 ( .A1(n490), .A2(n489), .A3(n488), .ZN(curr_proc_regs[256]) );
  NAND2_X1 U841 ( .A1(regs[1281]), .A2(n19), .ZN(n493) );
  AOI22_X1 U842 ( .A1(n58), .A2(regs[769]), .B1(n42), .B2(regs[257]), .ZN(n492) );
  AOI22_X1 U843 ( .A1(n120), .A2(regs[2305]), .B1(n4), .B2(regs[1793]), .ZN(
        n491) );
  NAND3_X1 U844 ( .A1(n493), .A2(n492), .A3(n491), .ZN(curr_proc_regs[257]) );
  NAND2_X1 U845 ( .A1(regs[1282]), .A2(n18), .ZN(n496) );
  AOI22_X1 U846 ( .A1(n10), .A2(regs[770]), .B1(n40), .B2(regs[258]), .ZN(n495) );
  AOI22_X1 U847 ( .A1(n120), .A2(regs[2306]), .B1(n4), .B2(regs[1794]), .ZN(
        n494) );
  NAND3_X1 U848 ( .A1(n496), .A2(n495), .A3(n494), .ZN(curr_proc_regs[258]) );
  NAND2_X1 U849 ( .A1(regs[1283]), .A2(n18), .ZN(n499) );
  AOI22_X1 U850 ( .A1(n49), .A2(regs[771]), .B1(n30), .B2(regs[259]), .ZN(n498) );
  AOI22_X1 U851 ( .A1(n120), .A2(regs[2307]), .B1(n17), .B2(regs[1795]), .ZN(
        n497) );
  NAND3_X1 U852 ( .A1(n499), .A2(n498), .A3(n497), .ZN(curr_proc_regs[259]) );
  INV_X1 U853 ( .A(regs[1049]), .ZN(n1392) );
  AOI22_X1 U854 ( .A1(n120), .A2(regs[2073]), .B1(n17), .B2(regs[1561]), .ZN(
        n501) );
  AOI22_X1 U855 ( .A1(n10), .A2(regs[537]), .B1(n36), .B2(regs[25]), .ZN(n500)
         );
  OAI211_X1 U856 ( .C1(n100), .C2(n1392), .A(n501), .B(n500), .ZN(
        curr_proc_regs[25]) );
  NAND2_X1 U857 ( .A1(regs[1284]), .A2(n91), .ZN(n504) );
  AOI22_X1 U858 ( .A1(n56), .A2(regs[772]), .B1(n33), .B2(regs[260]), .ZN(n503) );
  AOI22_X1 U859 ( .A1(n120), .A2(regs[2308]), .B1(n17), .B2(regs[1796]), .ZN(
        n502) );
  NAND3_X1 U860 ( .A1(n504), .A2(n503), .A3(n502), .ZN(curr_proc_regs[260]) );
  NAND2_X1 U861 ( .A1(regs[1285]), .A2(n19), .ZN(n507) );
  AOI22_X1 U862 ( .A1(n10), .A2(regs[773]), .B1(n35), .B2(regs[261]), .ZN(n506) );
  AOI22_X1 U863 ( .A1(n120), .A2(regs[2309]), .B1(n17), .B2(regs[1797]), .ZN(
        n505) );
  NAND3_X1 U864 ( .A1(n507), .A2(n506), .A3(n505), .ZN(curr_proc_regs[261]) );
  NAND2_X1 U865 ( .A1(regs[1286]), .A2(n89), .ZN(n510) );
  AOI22_X1 U866 ( .A1(n49), .A2(regs[774]), .B1(n31), .B2(regs[262]), .ZN(n509) );
  AOI22_X1 U867 ( .A1(n120), .A2(regs[2310]), .B1(n17), .B2(regs[1798]), .ZN(
        n508) );
  NAND3_X1 U868 ( .A1(n510), .A2(n509), .A3(n508), .ZN(curr_proc_regs[262]) );
  NAND2_X1 U869 ( .A1(regs[775]), .A2(n62), .ZN(n513) );
  AOI22_X1 U870 ( .A1(n90), .A2(regs[1287]), .B1(n30), .B2(regs[263]), .ZN(
        n512) );
  AOI22_X1 U871 ( .A1(n119), .A2(regs[2311]), .B1(n17), .B2(regs[1799]), .ZN(
        n511) );
  NAND3_X1 U872 ( .A1(n513), .A2(n512), .A3(n511), .ZN(curr_proc_regs[263]) );
  NAND2_X1 U873 ( .A1(regs[1288]), .A2(n18), .ZN(n516) );
  AOI22_X1 U874 ( .A1(n10), .A2(regs[776]), .B1(n29), .B2(regs[264]), .ZN(n515) );
  AOI22_X1 U875 ( .A1(n119), .A2(regs[2312]), .B1(n17), .B2(regs[1800]), .ZN(
        n514) );
  NAND3_X1 U876 ( .A1(n516), .A2(n515), .A3(n514), .ZN(curr_proc_regs[264]) );
  NAND2_X1 U877 ( .A1(regs[1289]), .A2(n78), .ZN(n519) );
  AOI22_X1 U878 ( .A1(n52), .A2(regs[777]), .B1(n40), .B2(regs[265]), .ZN(n518) );
  AOI22_X1 U879 ( .A1(n119), .A2(regs[2313]), .B1(n17), .B2(regs[1801]), .ZN(
        n517) );
  NAND3_X1 U880 ( .A1(n519), .A2(n518), .A3(n517), .ZN(curr_proc_regs[265]) );
  NAND2_X1 U881 ( .A1(regs[778]), .A2(n62), .ZN(n522) );
  AOI22_X1 U882 ( .A1(n90), .A2(regs[1290]), .B1(n33), .B2(regs[266]), .ZN(
        n521) );
  AOI22_X1 U883 ( .A1(n119), .A2(regs[2314]), .B1(n17), .B2(regs[1802]), .ZN(
        n520) );
  NAND3_X1 U884 ( .A1(n522), .A2(n521), .A3(n520), .ZN(curr_proc_regs[266]) );
  NAND2_X1 U885 ( .A1(regs[779]), .A2(n8), .ZN(n525) );
  AOI22_X1 U886 ( .A1(n90), .A2(regs[1291]), .B1(n35), .B2(regs[267]), .ZN(
        n524) );
  AOI22_X1 U887 ( .A1(n119), .A2(regs[2315]), .B1(n17), .B2(regs[1803]), .ZN(
        n523) );
  NAND3_X1 U888 ( .A1(n525), .A2(n524), .A3(n523), .ZN(curr_proc_regs[267]) );
  NAND2_X1 U889 ( .A1(regs[780]), .A2(n8), .ZN(n528) );
  AOI22_X1 U890 ( .A1(n90), .A2(regs[1292]), .B1(n42), .B2(regs[268]), .ZN(
        n527) );
  AOI22_X1 U891 ( .A1(n119), .A2(regs[2316]), .B1(n17), .B2(regs[1804]), .ZN(
        n526) );
  NAND3_X1 U892 ( .A1(n528), .A2(n527), .A3(n526), .ZN(curr_proc_regs[268]) );
  NAND2_X1 U893 ( .A1(regs[781]), .A2(n8), .ZN(n531) );
  AOI22_X1 U894 ( .A1(n90), .A2(regs[1293]), .B1(n35), .B2(regs[269]), .ZN(
        n530) );
  AOI22_X1 U895 ( .A1(n119), .A2(regs[2317]), .B1(n69), .B2(regs[1805]), .ZN(
        n529) );
  NAND3_X1 U896 ( .A1(n531), .A2(n530), .A3(n529), .ZN(curr_proc_regs[269]) );
  INV_X1 U897 ( .A(regs[1050]), .ZN(n1395) );
  AOI22_X1 U898 ( .A1(n119), .A2(regs[2074]), .B1(n69), .B2(regs[1562]), .ZN(
        n533) );
  AOI22_X1 U899 ( .A1(n54), .A2(regs[538]), .B1(n40), .B2(regs[26]), .ZN(n532)
         );
  OAI211_X1 U900 ( .C1(n2221), .C2(n1395), .A(n533), .B(n532), .ZN(
        curr_proc_regs[26]) );
  NAND2_X1 U901 ( .A1(regs[1294]), .A2(n91), .ZN(n536) );
  AOI22_X1 U902 ( .A1(n52), .A2(regs[782]), .B1(n42), .B2(regs[270]), .ZN(n535) );
  AOI22_X1 U903 ( .A1(n119), .A2(regs[2318]), .B1(n69), .B2(regs[1806]), .ZN(
        n534) );
  NAND3_X1 U904 ( .A1(n536), .A2(n535), .A3(n534), .ZN(curr_proc_regs[270]) );
  NAND2_X1 U905 ( .A1(regs[1295]), .A2(n97), .ZN(n539) );
  AOI22_X1 U906 ( .A1(n54), .A2(regs[783]), .B1(n31), .B2(regs[271]), .ZN(n538) );
  AOI22_X1 U907 ( .A1(n119), .A2(regs[2319]), .B1(n69), .B2(regs[1807]), .ZN(
        n537) );
  NAND3_X1 U908 ( .A1(n539), .A2(n538), .A3(n537), .ZN(curr_proc_regs[271]) );
  NAND2_X1 U909 ( .A1(regs[784]), .A2(n62), .ZN(n542) );
  AOI22_X1 U910 ( .A1(n89), .A2(regs[1296]), .B1(n31), .B2(regs[272]), .ZN(
        n541) );
  AOI22_X1 U911 ( .A1(n121), .A2(regs[2320]), .B1(n69), .B2(regs[1808]), .ZN(
        n540) );
  NAND3_X1 U912 ( .A1(n542), .A2(n541), .A3(n540), .ZN(curr_proc_regs[272]) );
  NAND2_X1 U913 ( .A1(regs[785]), .A2(n8), .ZN(n545) );
  AOI22_X1 U914 ( .A1(n89), .A2(regs[1297]), .B1(n30), .B2(regs[273]), .ZN(
        n544) );
  AOI22_X1 U915 ( .A1(n123), .A2(regs[2321]), .B1(n69), .B2(regs[1809]), .ZN(
        n543) );
  NAND3_X1 U916 ( .A1(n545), .A2(n544), .A3(n543), .ZN(curr_proc_regs[273]) );
  NAND2_X1 U917 ( .A1(regs[1298]), .A2(n18), .ZN(n548) );
  AOI22_X1 U918 ( .A1(n53), .A2(regs[786]), .B1(n29), .B2(regs[274]), .ZN(n547) );
  AOI22_X1 U919 ( .A1(n136), .A2(regs[2322]), .B1(n69), .B2(regs[1810]), .ZN(
        n546) );
  NAND3_X1 U920 ( .A1(n548), .A2(n547), .A3(n546), .ZN(curr_proc_regs[274]) );
  NAND2_X1 U921 ( .A1(regs[787]), .A2(n62), .ZN(n551) );
  AOI22_X1 U922 ( .A1(n89), .A2(regs[1299]), .B1(n31), .B2(regs[275]), .ZN(
        n550) );
  AOI22_X1 U923 ( .A1(n135), .A2(regs[2323]), .B1(n69), .B2(regs[1811]), .ZN(
        n549) );
  NAND3_X1 U924 ( .A1(n551), .A2(n550), .A3(n549), .ZN(curr_proc_regs[275]) );
  NAND2_X1 U925 ( .A1(regs[1300]), .A2(n98), .ZN(n554) );
  AOI22_X1 U926 ( .A1(n54), .A2(regs[788]), .B1(n35), .B2(regs[276]), .ZN(n553) );
  AOI22_X1 U927 ( .A1(n131), .A2(regs[2324]), .B1(n69), .B2(regs[1812]), .ZN(
        n552) );
  NAND3_X1 U928 ( .A1(n554), .A2(n553), .A3(n552), .ZN(curr_proc_regs[276]) );
  NAND2_X1 U929 ( .A1(regs[789]), .A2(n8), .ZN(n557) );
  AOI22_X1 U930 ( .A1(n89), .A2(regs[1301]), .B1(n40), .B2(regs[277]), .ZN(
        n556) );
  AOI22_X1 U931 ( .A1(n134), .A2(regs[2325]), .B1(n69), .B2(regs[1813]), .ZN(
        n555) );
  NAND3_X1 U932 ( .A1(n557), .A2(n556), .A3(n555), .ZN(curr_proc_regs[277]) );
  NAND2_X1 U933 ( .A1(regs[1302]), .A2(n19), .ZN(n560) );
  AOI22_X1 U934 ( .A1(n58), .A2(regs[790]), .B1(n40), .B2(regs[278]), .ZN(n559) );
  AOI22_X1 U935 ( .A1(n133), .A2(regs[2326]), .B1(n69), .B2(regs[1814]), .ZN(
        n558) );
  NAND3_X1 U936 ( .A1(n560), .A2(n559), .A3(n558), .ZN(curr_proc_regs[278]) );
  NAND2_X1 U937 ( .A1(regs[791]), .A2(n62), .ZN(n563) );
  AOI22_X1 U938 ( .A1(n88), .A2(regs[1303]), .B1(n41), .B2(regs[279]), .ZN(
        n562) );
  AOI22_X1 U939 ( .A1(n132), .A2(regs[2327]), .B1(n4), .B2(regs[1815]), .ZN(
        n561) );
  NAND3_X1 U940 ( .A1(n563), .A2(n562), .A3(n561), .ZN(curr_proc_regs[279]) );
  INV_X1 U941 ( .A(regs[1051]), .ZN(n1398) );
  AOI22_X1 U942 ( .A1(n126), .A2(regs[2075]), .B1(n4), .B2(regs[1563]), .ZN(
        n565) );
  AOI22_X1 U943 ( .A1(n52), .A2(regs[539]), .B1(n12), .B2(regs[27]), .ZN(n564)
         );
  OAI211_X1 U944 ( .C1(n5), .C2(n1398), .A(n565), .B(n564), .ZN(
        curr_proc_regs[27]) );
  NAND2_X1 U945 ( .A1(regs[792]), .A2(n8), .ZN(n568) );
  AOI22_X1 U946 ( .A1(n88), .A2(regs[1304]), .B1(n43), .B2(regs[280]), .ZN(
        n567) );
  AOI22_X1 U947 ( .A1(n127), .A2(regs[2328]), .B1(n4), .B2(regs[1816]), .ZN(
        n566) );
  NAND3_X1 U948 ( .A1(n568), .A2(n567), .A3(n566), .ZN(curr_proc_regs[280]) );
  NAND2_X1 U949 ( .A1(regs[793]), .A2(n8), .ZN(n571) );
  AOI22_X1 U950 ( .A1(n88), .A2(regs[1305]), .B1(n41), .B2(regs[281]), .ZN(
        n570) );
  AOI22_X1 U951 ( .A1(n128), .A2(regs[2329]), .B1(n4), .B2(regs[1817]), .ZN(
        n569) );
  NAND3_X1 U952 ( .A1(n571), .A2(n570), .A3(n569), .ZN(curr_proc_regs[281]) );
  NAND2_X1 U953 ( .A1(regs[1306]), .A2(n19), .ZN(n574) );
  AOI22_X1 U954 ( .A1(n54), .A2(regs[794]), .B1(n29), .B2(regs[282]), .ZN(n573) );
  AOI22_X1 U955 ( .A1(n129), .A2(regs[2330]), .B1(n4), .B2(regs[1818]), .ZN(
        n572) );
  NAND3_X1 U956 ( .A1(n574), .A2(n573), .A3(n572), .ZN(curr_proc_regs[282]) );
  NAND2_X1 U957 ( .A1(regs[1307]), .A2(n18), .ZN(n577) );
  AOI22_X1 U958 ( .A1(n52), .A2(regs[795]), .B1(n30), .B2(regs[283]), .ZN(n576) );
  AOI22_X1 U959 ( .A1(n134), .A2(regs[2331]), .B1(n4), .B2(regs[1819]), .ZN(
        n575) );
  NAND3_X1 U960 ( .A1(n577), .A2(n576), .A3(n575), .ZN(curr_proc_regs[283]) );
  NAND2_X1 U961 ( .A1(regs[1308]), .A2(n19), .ZN(n580) );
  AOI22_X1 U962 ( .A1(n8), .A2(regs[796]), .B1(n42), .B2(regs[284]), .ZN(n579)
         );
  AOI22_X1 U963 ( .A1(n133), .A2(regs[2332]), .B1(n4), .B2(regs[1820]), .ZN(
        n578) );
  NAND3_X1 U964 ( .A1(n580), .A2(n579), .A3(n578), .ZN(curr_proc_regs[284]) );
  NAND2_X1 U965 ( .A1(regs[797]), .A2(n8), .ZN(n583) );
  AOI22_X1 U966 ( .A1(n88), .A2(regs[1309]), .B1(n42), .B2(regs[285]), .ZN(
        n582) );
  AOI22_X1 U967 ( .A1(n132), .A2(regs[2333]), .B1(n4), .B2(regs[1821]), .ZN(
        n581) );
  NAND3_X1 U968 ( .A1(n583), .A2(n582), .A3(n581), .ZN(curr_proc_regs[285]) );
  NAND2_X1 U969 ( .A1(regs[798]), .A2(n62), .ZN(n586) );
  AOI22_X1 U970 ( .A1(n88), .A2(regs[1310]), .B1(n31), .B2(regs[286]), .ZN(
        n585) );
  AOI22_X1 U971 ( .A1(n127), .A2(regs[2334]), .B1(n4), .B2(regs[1822]), .ZN(
        n584) );
  NAND3_X1 U972 ( .A1(n586), .A2(n585), .A3(n584), .ZN(curr_proc_regs[286]) );
  NAND2_X1 U973 ( .A1(regs[1311]), .A2(n92), .ZN(n589) );
  AOI22_X1 U974 ( .A1(n54), .A2(regs[799]), .B1(n36), .B2(regs[287]), .ZN(n588) );
  AOI22_X1 U975 ( .A1(n128), .A2(regs[2335]), .B1(n4), .B2(regs[1823]), .ZN(
        n587) );
  NAND3_X1 U976 ( .A1(n589), .A2(n588), .A3(n587), .ZN(curr_proc_regs[287]) );
  NAND2_X1 U977 ( .A1(regs[800]), .A2(n8), .ZN(n592) );
  AOI22_X1 U978 ( .A1(n97), .A2(regs[1312]), .B1(n33), .B2(regs[288]), .ZN(
        n591) );
  AOI22_X1 U979 ( .A1(n129), .A2(regs[2336]), .B1(n4), .B2(regs[1824]), .ZN(
        n590) );
  NAND3_X1 U980 ( .A1(n592), .A2(n591), .A3(n590), .ZN(curr_proc_regs[288]) );
  NAND2_X1 U981 ( .A1(regs[801]), .A2(n62), .ZN(n595) );
  AOI22_X1 U982 ( .A1(n89), .A2(regs[1313]), .B1(n43), .B2(regs[289]), .ZN(
        n594) );
  AOI22_X1 U983 ( .A1(n131), .A2(regs[2337]), .B1(n9), .B2(regs[1825]), .ZN(
        n593) );
  NAND3_X1 U984 ( .A1(n595), .A2(n594), .A3(n593), .ZN(curr_proc_regs[289]) );
  INV_X1 U985 ( .A(regs[540]), .ZN(n1403) );
  AOI22_X1 U986 ( .A1(n122), .A2(regs[2076]), .B1(n9), .B2(regs[1564]), .ZN(
        n597) );
  AOI22_X1 U987 ( .A1(n90), .A2(regs[1052]), .B1(n43), .B2(regs[28]), .ZN(n596) );
  OAI211_X1 U988 ( .C1(n64), .C2(n1403), .A(n597), .B(n596), .ZN(
        curr_proc_regs[28]) );
  NAND2_X1 U989 ( .A1(regs[802]), .A2(n8), .ZN(n600) );
  AOI22_X1 U990 ( .A1(n88), .A2(regs[1314]), .B1(n28), .B2(regs[290]), .ZN(
        n599) );
  AOI22_X1 U991 ( .A1(n20), .A2(regs[2338]), .B1(n9), .B2(regs[1826]), .ZN(
        n598) );
  NAND3_X1 U992 ( .A1(n600), .A2(n599), .A3(n598), .ZN(curr_proc_regs[290]) );
  NAND2_X1 U993 ( .A1(regs[803]), .A2(n8), .ZN(n603) );
  AOI22_X1 U994 ( .A1(n88), .A2(regs[1315]), .B1(n3), .B2(regs[291]), .ZN(n602) );
  AOI22_X1 U995 ( .A1(n124), .A2(regs[2339]), .B1(n9), .B2(regs[1827]), .ZN(
        n601) );
  NAND3_X1 U996 ( .A1(n603), .A2(n602), .A3(n601), .ZN(curr_proc_regs[291]) );
  NAND2_X1 U997 ( .A1(regs[804]), .A2(n8), .ZN(n606) );
  AOI22_X1 U998 ( .A1(n88), .A2(regs[1316]), .B1(n43), .B2(regs[292]), .ZN(
        n605) );
  AOI22_X1 U999 ( .A1(n125), .A2(regs[2340]), .B1(n9), .B2(regs[1828]), .ZN(
        n604) );
  NAND3_X1 U1000 ( .A1(n606), .A2(n605), .A3(n604), .ZN(curr_proc_regs[292])
         );
  NAND2_X1 U1001 ( .A1(regs[1317]), .A2(n19), .ZN(n609) );
  AOI22_X1 U1002 ( .A1(n54), .A2(regs[805]), .B1(n3), .B2(regs[293]), .ZN(n608) );
  AOI22_X1 U1003 ( .A1(n20), .A2(regs[2341]), .B1(n9), .B2(regs[1829]), .ZN(
        n607) );
  NAND3_X1 U1004 ( .A1(n609), .A2(n608), .A3(n607), .ZN(curr_proc_regs[293])
         );
  NAND2_X1 U1005 ( .A1(regs[806]), .A2(n8), .ZN(n612) );
  AOI22_X1 U1006 ( .A1(n88), .A2(regs[1318]), .B1(n3), .B2(regs[294]), .ZN(
        n611) );
  AOI22_X1 U1007 ( .A1(n20), .A2(regs[2342]), .B1(n9), .B2(regs[1830]), .ZN(
        n610) );
  NAND3_X1 U1008 ( .A1(n612), .A2(n611), .A3(n610), .ZN(curr_proc_regs[294])
         );
  NAND2_X1 U1009 ( .A1(regs[1319]), .A2(n19), .ZN(n615) );
  AOI22_X1 U1010 ( .A1(n54), .A2(regs[807]), .B1(n12), .B2(regs[295]), .ZN(
        n614) );
  AOI22_X1 U1011 ( .A1(n20), .A2(regs[2343]), .B1(n9), .B2(regs[1831]), .ZN(
        n613) );
  NAND3_X1 U1012 ( .A1(n615), .A2(n614), .A3(n613), .ZN(curr_proc_regs[295])
         );
  NAND2_X1 U1013 ( .A1(regs[808]), .A2(n8), .ZN(n618) );
  AOI22_X1 U1014 ( .A1(n88), .A2(regs[1320]), .B1(n12), .B2(regs[296]), .ZN(
        n617) );
  AOI22_X1 U1015 ( .A1(n20), .A2(regs[2344]), .B1(n9), .B2(regs[1832]), .ZN(
        n616) );
  NAND3_X1 U1016 ( .A1(n618), .A2(n617), .A3(n616), .ZN(curr_proc_regs[296])
         );
  NAND2_X1 U1017 ( .A1(regs[809]), .A2(n8), .ZN(n621) );
  AOI22_X1 U1018 ( .A1(n88), .A2(regs[1321]), .B1(n28), .B2(regs[297]), .ZN(
        n620) );
  AOI22_X1 U1019 ( .A1(n20), .A2(regs[2345]), .B1(n9), .B2(regs[1833]), .ZN(
        n619) );
  NAND3_X1 U1020 ( .A1(n621), .A2(n620), .A3(n619), .ZN(curr_proc_regs[297])
         );
  NAND2_X1 U1021 ( .A1(regs[1322]), .A2(n19), .ZN(n624) );
  AOI22_X1 U1022 ( .A1(n52), .A2(regs[810]), .B1(n41), .B2(regs[298]), .ZN(
        n623) );
  AOI22_X1 U1023 ( .A1(n20), .A2(regs[2346]), .B1(n9), .B2(regs[1834]), .ZN(
        n622) );
  NAND3_X1 U1024 ( .A1(n624), .A2(n623), .A3(n622), .ZN(curr_proc_regs[298])
         );
  NAND2_X1 U1025 ( .A1(regs[811]), .A2(n8), .ZN(n627) );
  AOI22_X1 U1026 ( .A1(n89), .A2(regs[1323]), .B1(n3), .B2(regs[299]), .ZN(
        n626) );
  AOI22_X1 U1027 ( .A1(n20), .A2(regs[2347]), .B1(n71), .B2(regs[1835]), .ZN(
        n625) );
  NAND3_X1 U1028 ( .A1(n627), .A2(n626), .A3(n625), .ZN(curr_proc_regs[299])
         );
  INV_X1 U1029 ( .A(regs[1053]), .ZN(n1406) );
  AOI22_X1 U1030 ( .A1(n20), .A2(regs[2077]), .B1(n71), .B2(regs[1565]), .ZN(
        n629) );
  AOI22_X1 U1031 ( .A1(n54), .A2(regs[541]), .B1(n3), .B2(regs[29]), .ZN(n628)
         );
  OAI211_X1 U1032 ( .C1(n16), .C2(n1406), .A(n629), .B(n628), .ZN(
        curr_proc_regs[29]) );
  INV_X1 U1033 ( .A(regs[514]), .ZN(n1322) );
  AOI22_X1 U1034 ( .A1(n20), .A2(regs[2050]), .B1(n71), .B2(regs[1538]), .ZN(
        n631) );
  AOI22_X1 U1035 ( .A1(n89), .A2(regs[1026]), .B1(n3), .B2(regs[2]), .ZN(n630)
         );
  OAI211_X1 U1036 ( .C1(n11), .C2(n1322), .A(n631), .B(n630), .ZN(
        curr_proc_regs[2]) );
  NAND2_X1 U1037 ( .A1(regs[812]), .A2(n8), .ZN(n634) );
  AOI22_X1 U1038 ( .A1(n89), .A2(regs[1324]), .B1(n34), .B2(regs[300]), .ZN(
        n633) );
  AOI22_X1 U1039 ( .A1(n20), .A2(regs[2348]), .B1(n71), .B2(regs[1836]), .ZN(
        n632) );
  NAND3_X1 U1040 ( .A1(n634), .A2(n633), .A3(n632), .ZN(curr_proc_regs[300])
         );
  NAND2_X1 U1041 ( .A1(regs[813]), .A2(n8), .ZN(n637) );
  AOI22_X1 U1042 ( .A1(n89), .A2(regs[1325]), .B1(n41), .B2(regs[301]), .ZN(
        n636) );
  AOI22_X1 U1043 ( .A1(n20), .A2(regs[2349]), .B1(n71), .B2(regs[1837]), .ZN(
        n635) );
  NAND3_X1 U1044 ( .A1(n637), .A2(n636), .A3(n635), .ZN(curr_proc_regs[301])
         );
  NAND2_X1 U1045 ( .A1(regs[814]), .A2(n8), .ZN(n640) );
  AOI22_X1 U1046 ( .A1(n89), .A2(regs[1326]), .B1(n43), .B2(regs[302]), .ZN(
        n639) );
  AOI22_X1 U1047 ( .A1(n20), .A2(regs[2350]), .B1(n71), .B2(regs[1838]), .ZN(
        n638) );
  NAND3_X1 U1048 ( .A1(n640), .A2(n639), .A3(n638), .ZN(curr_proc_regs[302])
         );
  NAND2_X1 U1049 ( .A1(regs[815]), .A2(n8), .ZN(n643) );
  AOI22_X1 U1050 ( .A1(n89), .A2(regs[1327]), .B1(n3), .B2(regs[303]), .ZN(
        n642) );
  AOI22_X1 U1051 ( .A1(n20), .A2(regs[2351]), .B1(n71), .B2(regs[1839]), .ZN(
        n641) );
  NAND3_X1 U1052 ( .A1(n643), .A2(n642), .A3(n641), .ZN(curr_proc_regs[303])
         );
  NAND2_X1 U1053 ( .A1(regs[1328]), .A2(n19), .ZN(n646) );
  AOI22_X1 U1054 ( .A1(n54), .A2(regs[816]), .B1(n3), .B2(regs[304]), .ZN(n645) );
  AOI22_X1 U1055 ( .A1(n20), .A2(regs[2352]), .B1(n71), .B2(regs[1840]), .ZN(
        n644) );
  NAND3_X1 U1056 ( .A1(n646), .A2(n645), .A3(n644), .ZN(curr_proc_regs[304])
         );
  NAND2_X1 U1057 ( .A1(regs[817]), .A2(n8), .ZN(n649) );
  AOI22_X1 U1058 ( .A1(n89), .A2(regs[1329]), .B1(n12), .B2(regs[305]), .ZN(
        n648) );
  AOI22_X1 U1059 ( .A1(n20), .A2(regs[2353]), .B1(n71), .B2(regs[1841]), .ZN(
        n647) );
  NAND3_X1 U1060 ( .A1(n649), .A2(n648), .A3(n647), .ZN(curr_proc_regs[305])
         );
  NAND2_X1 U1061 ( .A1(regs[1330]), .A2(n19), .ZN(n652) );
  AOI22_X1 U1062 ( .A1(n53), .A2(regs[818]), .B1(n12), .B2(regs[306]), .ZN(
        n651) );
  AOI22_X1 U1063 ( .A1(n20), .A2(regs[2354]), .B1(n71), .B2(regs[1842]), .ZN(
        n650) );
  NAND3_X1 U1064 ( .A1(n652), .A2(n651), .A3(n650), .ZN(curr_proc_regs[306])
         );
  NAND2_X1 U1065 ( .A1(regs[1331]), .A2(n19), .ZN(n655) );
  AOI22_X1 U1066 ( .A1(n52), .A2(regs[819]), .B1(n28), .B2(regs[307]), .ZN(
        n654) );
  AOI22_X1 U1067 ( .A1(n7), .A2(regs[2355]), .B1(n71), .B2(regs[1843]), .ZN(
        n653) );
  NAND3_X1 U1068 ( .A1(n655), .A2(n654), .A3(n653), .ZN(curr_proc_regs[307])
         );
  NAND2_X1 U1069 ( .A1(regs[820]), .A2(n8), .ZN(n658) );
  AOI22_X1 U1070 ( .A1(n90), .A2(regs[1332]), .B1(n45), .B2(regs[308]), .ZN(
        n657) );
  AOI22_X1 U1071 ( .A1(n20), .A2(regs[2356]), .B1(n70), .B2(regs[1844]), .ZN(
        n656) );
  NAND3_X1 U1072 ( .A1(n658), .A2(n657), .A3(n656), .ZN(curr_proc_regs[308])
         );
  NAND2_X1 U1073 ( .A1(regs[821]), .A2(n62), .ZN(n661) );
  AOI22_X1 U1074 ( .A1(n90), .A2(regs[1333]), .B1(n45), .B2(regs[309]), .ZN(
        n660) );
  AOI22_X1 U1075 ( .A1(n20), .A2(regs[2357]), .B1(n70), .B2(regs[1845]), .ZN(
        n659) );
  NAND3_X1 U1076 ( .A1(n661), .A2(n660), .A3(n659), .ZN(curr_proc_regs[309])
         );
  INV_X1 U1077 ( .A(regs[1054]), .ZN(n1409) );
  AOI22_X1 U1078 ( .A1(n20), .A2(regs[2078]), .B1(n70), .B2(regs[1566]), .ZN(
        n663) );
  AOI22_X1 U1079 ( .A1(n54), .A2(regs[542]), .B1(n45), .B2(regs[30]), .ZN(n662) );
  OAI211_X1 U1080 ( .C1(n2221), .C2(n1409), .A(n663), .B(n662), .ZN(
        curr_proc_regs[30]) );
  NAND2_X1 U1081 ( .A1(regs[822]), .A2(n62), .ZN(n666) );
  AOI22_X1 U1082 ( .A1(n90), .A2(regs[1334]), .B1(n45), .B2(regs[310]), .ZN(
        n665) );
  AOI22_X1 U1083 ( .A1(n20), .A2(regs[2358]), .B1(n70), .B2(regs[1846]), .ZN(
        n664) );
  NAND3_X1 U1084 ( .A1(n666), .A2(n665), .A3(n664), .ZN(curr_proc_regs[310])
         );
  NAND2_X1 U1085 ( .A1(regs[823]), .A2(n62), .ZN(n669) );
  AOI22_X1 U1086 ( .A1(n90), .A2(regs[1335]), .B1(n43), .B2(regs[311]), .ZN(
        n668) );
  AOI22_X1 U1087 ( .A1(n20), .A2(regs[2359]), .B1(n70), .B2(regs[1847]), .ZN(
        n667) );
  NAND3_X1 U1088 ( .A1(n669), .A2(n668), .A3(n667), .ZN(curr_proc_regs[311])
         );
  NAND2_X1 U1089 ( .A1(regs[824]), .A2(n62), .ZN(n672) );
  AOI22_X1 U1090 ( .A1(n90), .A2(regs[1336]), .B1(n3), .B2(regs[312]), .ZN(
        n671) );
  AOI22_X1 U1091 ( .A1(n7), .A2(regs[2360]), .B1(n70), .B2(regs[1848]), .ZN(
        n670) );
  NAND3_X1 U1092 ( .A1(n672), .A2(n671), .A3(n670), .ZN(curr_proc_regs[312])
         );
  NAND2_X1 U1093 ( .A1(regs[1337]), .A2(n19), .ZN(n675) );
  AOI22_X1 U1094 ( .A1(n53), .A2(regs[825]), .B1(n3), .B2(regs[313]), .ZN(n674) );
  AOI22_X1 U1095 ( .A1(n7), .A2(regs[2361]), .B1(n70), .B2(regs[1849]), .ZN(
        n673) );
  NAND3_X1 U1096 ( .A1(n675), .A2(n674), .A3(n673), .ZN(curr_proc_regs[313])
         );
  NAND2_X1 U1097 ( .A1(regs[826]), .A2(n62), .ZN(n678) );
  AOI22_X1 U1098 ( .A1(n90), .A2(regs[1338]), .B1(n12), .B2(regs[314]), .ZN(
        n677) );
  AOI22_X1 U1099 ( .A1(n7), .A2(regs[2362]), .B1(n70), .B2(regs[1850]), .ZN(
        n676) );
  NAND3_X1 U1100 ( .A1(n678), .A2(n677), .A3(n676), .ZN(curr_proc_regs[314])
         );
  NAND2_X1 U1101 ( .A1(regs[1339]), .A2(n83), .ZN(n681) );
  AOI22_X1 U1102 ( .A1(n53), .A2(regs[827]), .B1(n12), .B2(regs[315]), .ZN(
        n680) );
  AOI22_X1 U1103 ( .A1(n7), .A2(regs[2363]), .B1(n70), .B2(regs[1851]), .ZN(
        n679) );
  NAND3_X1 U1104 ( .A1(n681), .A2(n680), .A3(n679), .ZN(curr_proc_regs[315])
         );
  NAND2_X1 U1105 ( .A1(regs[1340]), .A2(n84), .ZN(n684) );
  AOI22_X1 U1106 ( .A1(n54), .A2(regs[828]), .B1(n28), .B2(regs[316]), .ZN(
        n683) );
  AOI22_X1 U1107 ( .A1(n7), .A2(regs[2364]), .B1(n70), .B2(regs[1852]), .ZN(
        n682) );
  NAND3_X1 U1108 ( .A1(n684), .A2(n683), .A3(n682), .ZN(curr_proc_regs[316])
         );
  NAND2_X1 U1109 ( .A1(regs[1341]), .A2(n96), .ZN(n687) );
  AOI22_X1 U1110 ( .A1(n53), .A2(regs[829]), .B1(n3), .B2(regs[317]), .ZN(n686) );
  AOI22_X1 U1111 ( .A1(n7), .A2(regs[2365]), .B1(n70), .B2(regs[1853]), .ZN(
        n685) );
  NAND3_X1 U1112 ( .A1(n687), .A2(n686), .A3(n685), .ZN(curr_proc_regs[317])
         );
  NAND2_X1 U1113 ( .A1(regs[1342]), .A2(n81), .ZN(n690) );
  AOI22_X1 U1114 ( .A1(n52), .A2(regs[830]), .B1(n32), .B2(regs[318]), .ZN(
        n689) );
  AOI22_X1 U1115 ( .A1(n7), .A2(regs[2366]), .B1(n67), .B2(regs[1854]), .ZN(
        n688) );
  NAND3_X1 U1116 ( .A1(n690), .A2(n689), .A3(n688), .ZN(curr_proc_regs[318])
         );
  NAND2_X1 U1117 ( .A1(regs[831]), .A2(n8), .ZN(n693) );
  AOI22_X1 U1118 ( .A1(n91), .A2(regs[1343]), .B1(n41), .B2(regs[319]), .ZN(
        n692) );
  AOI22_X1 U1119 ( .A1(n7), .A2(regs[2367]), .B1(n67), .B2(regs[1855]), .ZN(
        n691) );
  NAND3_X1 U1120 ( .A1(n693), .A2(n692), .A3(n691), .ZN(curr_proc_regs[319])
         );
  INV_X1 U1121 ( .A(regs[543]), .ZN(n1412) );
  AOI22_X1 U1122 ( .A1(n7), .A2(regs[2079]), .B1(n67), .B2(regs[1567]), .ZN(
        n695) );
  AOI22_X1 U1123 ( .A1(n91), .A2(regs[1055]), .B1(n43), .B2(regs[31]), .ZN(
        n694) );
  OAI211_X1 U1124 ( .C1(n2207), .C2(n1412), .A(n695), .B(n694), .ZN(
        curr_proc_regs[31]) );
  NAND2_X1 U1125 ( .A1(regs[1344]), .A2(n96), .ZN(n698) );
  AOI22_X1 U1126 ( .A1(n54), .A2(regs[832]), .B1(n3), .B2(regs[320]), .ZN(n697) );
  AOI22_X1 U1127 ( .A1(n7), .A2(regs[2368]), .B1(n67), .B2(regs[1856]), .ZN(
        n696) );
  NAND3_X1 U1128 ( .A1(n698), .A2(n697), .A3(n696), .ZN(curr_proc_regs[320])
         );
  NAND2_X1 U1129 ( .A1(regs[1345]), .A2(n96), .ZN(n701) );
  AOI22_X1 U1130 ( .A1(n54), .A2(regs[833]), .B1(n45), .B2(regs[321]), .ZN(
        n700) );
  AOI22_X1 U1131 ( .A1(n7), .A2(regs[2369]), .B1(n67), .B2(regs[1857]), .ZN(
        n699) );
  NAND3_X1 U1132 ( .A1(n701), .A2(n700), .A3(n699), .ZN(curr_proc_regs[321])
         );
  NAND2_X1 U1133 ( .A1(regs[834]), .A2(n2), .ZN(n704) );
  AOI22_X1 U1134 ( .A1(n92), .A2(regs[1346]), .B1(n45), .B2(regs[322]), .ZN(
        n703) );
  AOI22_X1 U1135 ( .A1(n7), .A2(regs[2370]), .B1(n67), .B2(regs[1858]), .ZN(
        n702) );
  NAND3_X1 U1136 ( .A1(n704), .A2(n703), .A3(n702), .ZN(curr_proc_regs[322])
         );
  NAND2_X1 U1137 ( .A1(regs[835]), .A2(n61), .ZN(n707) );
  AOI22_X1 U1138 ( .A1(n92), .A2(regs[1347]), .B1(n45), .B2(regs[323]), .ZN(
        n706) );
  AOI22_X1 U1139 ( .A1(n7), .A2(regs[2371]), .B1(n67), .B2(regs[1859]), .ZN(
        n705) );
  NAND3_X1 U1140 ( .A1(n707), .A2(n706), .A3(n705), .ZN(curr_proc_regs[323])
         );
  NAND2_X1 U1141 ( .A1(regs[1348]), .A2(n96), .ZN(n710) );
  AOI22_X1 U1142 ( .A1(n54), .A2(regs[836]), .B1(n45), .B2(regs[324]), .ZN(
        n709) );
  AOI22_X1 U1143 ( .A1(n136), .A2(regs[2372]), .B1(n67), .B2(regs[1860]), .ZN(
        n708) );
  NAND3_X1 U1144 ( .A1(n710), .A2(n709), .A3(n708), .ZN(curr_proc_regs[324])
         );
  NAND2_X1 U1145 ( .A1(regs[837]), .A2(n13), .ZN(n713) );
  AOI22_X1 U1146 ( .A1(n92), .A2(regs[1349]), .B1(n45), .B2(regs[325]), .ZN(
        n712) );
  AOI22_X1 U1147 ( .A1(n7), .A2(regs[2373]), .B1(n67), .B2(regs[1861]), .ZN(
        n711) );
  NAND3_X1 U1148 ( .A1(n713), .A2(n712), .A3(n711), .ZN(curr_proc_regs[325])
         );
  NAND2_X1 U1149 ( .A1(regs[838]), .A2(n2), .ZN(n716) );
  AOI22_X1 U1150 ( .A1(n92), .A2(regs[1350]), .B1(n45), .B2(regs[326]), .ZN(
        n715) );
  AOI22_X1 U1151 ( .A1(n7), .A2(regs[2374]), .B1(n67), .B2(regs[1862]), .ZN(
        n714) );
  NAND3_X1 U1152 ( .A1(n716), .A2(n715), .A3(n714), .ZN(curr_proc_regs[326])
         );
  NAND2_X1 U1153 ( .A1(regs[1351]), .A2(n95), .ZN(n719) );
  AOI22_X1 U1154 ( .A1(n54), .A2(regs[839]), .B1(n45), .B2(regs[327]), .ZN(
        n718) );
  AOI22_X1 U1155 ( .A1(n7), .A2(regs[2375]), .B1(n67), .B2(regs[1863]), .ZN(
        n717) );
  NAND3_X1 U1156 ( .A1(n719), .A2(n718), .A3(n717), .ZN(curr_proc_regs[327])
         );
  NAND2_X1 U1157 ( .A1(regs[1352]), .A2(n95), .ZN(n722) );
  AOI22_X1 U1158 ( .A1(n54), .A2(regs[840]), .B1(n12), .B2(regs[328]), .ZN(
        n721) );
  AOI22_X1 U1159 ( .A1(n7), .A2(regs[2376]), .B1(n71), .B2(regs[1864]), .ZN(
        n720) );
  NAND3_X1 U1160 ( .A1(n722), .A2(n721), .A3(n720), .ZN(curr_proc_regs[328])
         );
  NAND2_X1 U1161 ( .A1(regs[841]), .A2(n62), .ZN(n725) );
  AOI22_X1 U1162 ( .A1(n91), .A2(regs[1353]), .B1(n28), .B2(regs[329]), .ZN(
        n724) );
  AOI22_X1 U1163 ( .A1(n7), .A2(regs[2377]), .B1(n71), .B2(regs[1865]), .ZN(
        n723) );
  NAND3_X1 U1164 ( .A1(n725), .A2(n724), .A3(n723), .ZN(curr_proc_regs[329])
         );
  INV_X1 U1165 ( .A(regs[544]), .ZN(n1415) );
  AOI22_X1 U1166 ( .A1(n7), .A2(regs[2080]), .B1(n71), .B2(regs[1568]), .ZN(
        n727) );
  AOI22_X1 U1167 ( .A1(n89), .A2(regs[1056]), .B1(n12), .B2(regs[32]), .ZN(
        n726) );
  OAI211_X1 U1168 ( .C1(n11), .C2(n1415), .A(n727), .B(n726), .ZN(
        curr_proc_regs[32]) );
  NAND2_X1 U1169 ( .A1(regs[1354]), .A2(n95), .ZN(n730) );
  AOI22_X1 U1170 ( .A1(n10), .A2(regs[842]), .B1(n12), .B2(regs[330]), .ZN(
        n729) );
  AOI22_X1 U1171 ( .A1(n7), .A2(regs[2378]), .B1(n71), .B2(regs[1866]), .ZN(
        n728) );
  NAND3_X1 U1172 ( .A1(n730), .A2(n729), .A3(n728), .ZN(curr_proc_regs[330])
         );
  NAND2_X1 U1173 ( .A1(regs[843]), .A2(n2), .ZN(n733) );
  AOI22_X1 U1174 ( .A1(n18), .A2(regs[1355]), .B1(n12), .B2(regs[331]), .ZN(
        n732) );
  AOI22_X1 U1175 ( .A1(n7), .A2(regs[2379]), .B1(n71), .B2(regs[1867]), .ZN(
        n731) );
  NAND3_X1 U1176 ( .A1(n733), .A2(n732), .A3(n731), .ZN(curr_proc_regs[331])
         );
  NAND2_X1 U1177 ( .A1(regs[1356]), .A2(n88), .ZN(n736) );
  AOI22_X1 U1178 ( .A1(n55), .A2(regs[844]), .B1(n12), .B2(regs[332]), .ZN(
        n735) );
  AOI22_X1 U1179 ( .A1(n136), .A2(regs[2380]), .B1(n71), .B2(regs[1868]), .ZN(
        n734) );
  NAND3_X1 U1180 ( .A1(n736), .A2(n735), .A3(n734), .ZN(curr_proc_regs[332])
         );
  NAND2_X1 U1181 ( .A1(regs[845]), .A2(n62), .ZN(n739) );
  AOI22_X1 U1182 ( .A1(n88), .A2(regs[1357]), .B1(n28), .B2(regs[333]), .ZN(
        n738) );
  AOI22_X1 U1183 ( .A1(n136), .A2(regs[2381]), .B1(n71), .B2(regs[1869]), .ZN(
        n737) );
  NAND3_X1 U1184 ( .A1(n739), .A2(n738), .A3(n737), .ZN(curr_proc_regs[333])
         );
  NAND2_X1 U1185 ( .A1(regs[846]), .A2(n60), .ZN(n742) );
  AOI22_X1 U1186 ( .A1(n89), .A2(regs[1358]), .B1(n12), .B2(regs[334]), .ZN(
        n741) );
  AOI22_X1 U1187 ( .A1(n136), .A2(regs[2382]), .B1(n71), .B2(regs[1870]), .ZN(
        n740) );
  NAND3_X1 U1188 ( .A1(n742), .A2(n741), .A3(n740), .ZN(curr_proc_regs[334])
         );
  NAND2_X1 U1189 ( .A1(regs[847]), .A2(n13), .ZN(n745) );
  AOI22_X1 U1190 ( .A1(n18), .A2(regs[1359]), .B1(n3), .B2(regs[335]), .ZN(
        n744) );
  AOI22_X1 U1191 ( .A1(n136), .A2(regs[2383]), .B1(n71), .B2(regs[1871]), .ZN(
        n743) );
  NAND3_X1 U1192 ( .A1(n745), .A2(n744), .A3(n743), .ZN(curr_proc_regs[335])
         );
  NAND2_X1 U1193 ( .A1(regs[1360]), .A2(n94), .ZN(n748) );
  AOI22_X1 U1194 ( .A1(n50), .A2(regs[848]), .B1(n12), .B2(regs[336]), .ZN(
        n747) );
  AOI22_X1 U1195 ( .A1(n136), .A2(regs[2384]), .B1(n71), .B2(regs[1872]), .ZN(
        n746) );
  NAND3_X1 U1196 ( .A1(n748), .A2(n747), .A3(n746), .ZN(curr_proc_regs[336])
         );
  NAND2_X1 U1197 ( .A1(regs[849]), .A2(n62), .ZN(n751) );
  AOI22_X1 U1198 ( .A1(n18), .A2(regs[1361]), .B1(n34), .B2(regs[337]), .ZN(
        n750) );
  AOI22_X1 U1199 ( .A1(n136), .A2(regs[2385]), .B1(n71), .B2(regs[1873]), .ZN(
        n749) );
  NAND3_X1 U1200 ( .A1(n751), .A2(n750), .A3(n749), .ZN(curr_proc_regs[337])
         );
  NAND2_X1 U1201 ( .A1(regs[1362]), .A2(n94), .ZN(n754) );
  AOI22_X1 U1202 ( .A1(n50), .A2(regs[850]), .B1(n46), .B2(regs[338]), .ZN(
        n753) );
  AOI22_X1 U1203 ( .A1(n136), .A2(regs[2386]), .B1(n69), .B2(regs[1874]), .ZN(
        n752) );
  NAND3_X1 U1204 ( .A1(n754), .A2(n753), .A3(n752), .ZN(curr_proc_regs[338])
         );
  NAND2_X1 U1205 ( .A1(regs[1363]), .A2(n95), .ZN(n757) );
  AOI22_X1 U1206 ( .A1(n57), .A2(regs[851]), .B1(n46), .B2(regs[339]), .ZN(
        n756) );
  AOI22_X1 U1207 ( .A1(n136), .A2(regs[2387]), .B1(n9), .B2(regs[1875]), .ZN(
        n755) );
  NAND3_X1 U1208 ( .A1(n757), .A2(n756), .A3(n755), .ZN(curr_proc_regs[339])
         );
  INV_X1 U1209 ( .A(regs[1057]), .ZN(n1418) );
  AOI22_X1 U1210 ( .A1(n136), .A2(regs[2081]), .B1(n73), .B2(regs[1569]), .ZN(
        n759) );
  AOI22_X1 U1211 ( .A1(n55), .A2(regs[545]), .B1(n46), .B2(regs[33]), .ZN(n758) );
  OAI211_X1 U1212 ( .C1(n100), .C2(n1418), .A(n759), .B(n758), .ZN(
        curr_proc_regs[33]) );
  NAND2_X1 U1213 ( .A1(regs[1364]), .A2(n82), .ZN(n762) );
  AOI22_X1 U1214 ( .A1(n49), .A2(regs[852]), .B1(n46), .B2(regs[340]), .ZN(
        n761) );
  AOI22_X1 U1215 ( .A1(n136), .A2(regs[2388]), .B1(n17), .B2(regs[1876]), .ZN(
        n760) );
  NAND3_X1 U1216 ( .A1(n762), .A2(n761), .A3(n760), .ZN(curr_proc_regs[340])
         );
  NAND2_X1 U1217 ( .A1(regs[1365]), .A2(n83), .ZN(n765) );
  AOI22_X1 U1218 ( .A1(n50), .A2(regs[853]), .B1(n34), .B2(regs[341]), .ZN(
        n764) );
  AOI22_X1 U1219 ( .A1(win[4]), .A2(regs[2389]), .B1(n17), .B2(regs[1877]), 
        .ZN(n763) );
  NAND3_X1 U1220 ( .A1(n765), .A2(n764), .A3(n763), .ZN(curr_proc_regs[341])
         );
  NAND2_X1 U1221 ( .A1(regs[1366]), .A2(n85), .ZN(n768) );
  AOI22_X1 U1222 ( .A1(n51), .A2(regs[854]), .B1(n32), .B2(regs[342]), .ZN(
        n767) );
  AOI22_X1 U1223 ( .A1(n135), .A2(regs[2390]), .B1(n69), .B2(regs[1878]), .ZN(
        n766) );
  NAND3_X1 U1224 ( .A1(n768), .A2(n767), .A3(n766), .ZN(curr_proc_regs[342])
         );
  NAND2_X1 U1225 ( .A1(regs[855]), .A2(n62), .ZN(n771) );
  AOI22_X1 U1226 ( .A1(n91), .A2(regs[1367]), .B1(n41), .B2(regs[343]), .ZN(
        n770) );
  AOI22_X1 U1227 ( .A1(n135), .A2(regs[2391]), .B1(n73), .B2(regs[1879]), .ZN(
        n769) );
  NAND3_X1 U1228 ( .A1(n771), .A2(n770), .A3(n769), .ZN(curr_proc_regs[343])
         );
  NAND2_X1 U1229 ( .A1(regs[856]), .A2(n8), .ZN(n774) );
  AOI22_X1 U1230 ( .A1(n92), .A2(regs[1368]), .B1(n43), .B2(regs[344]), .ZN(
        n773) );
  AOI22_X1 U1231 ( .A1(n135), .A2(regs[2392]), .B1(n75), .B2(regs[1880]), .ZN(
        n772) );
  NAND3_X1 U1232 ( .A1(n774), .A2(n773), .A3(n772), .ZN(curr_proc_regs[344])
         );
  NAND2_X1 U1233 ( .A1(regs[1369]), .A2(n98), .ZN(n777) );
  AOI22_X1 U1234 ( .A1(n58), .A2(regs[857]), .B1(n3), .B2(regs[345]), .ZN(n776) );
  AOI22_X1 U1235 ( .A1(n135), .A2(regs[2393]), .B1(n17), .B2(regs[1881]), .ZN(
        n775) );
  NAND3_X1 U1236 ( .A1(n777), .A2(n776), .A3(n775), .ZN(curr_proc_regs[345])
         );
  NAND2_X1 U1237 ( .A1(regs[1370]), .A2(n90), .ZN(n780) );
  AOI22_X1 U1238 ( .A1(n55), .A2(regs[858]), .B1(n3), .B2(regs[346]), .ZN(n779) );
  AOI22_X1 U1239 ( .A1(n135), .A2(regs[2394]), .B1(n69), .B2(regs[1882]), .ZN(
        n778) );
  NAND3_X1 U1240 ( .A1(n780), .A2(n779), .A3(n778), .ZN(curr_proc_regs[346])
         );
  NAND2_X1 U1241 ( .A1(regs[859]), .A2(n8), .ZN(n783) );
  AOI22_X1 U1242 ( .A1(n18), .A2(regs[1371]), .B1(n12), .B2(regs[347]), .ZN(
        n782) );
  AOI22_X1 U1243 ( .A1(n135), .A2(regs[2395]), .B1(n73), .B2(regs[1883]), .ZN(
        n781) );
  NAND3_X1 U1244 ( .A1(n783), .A2(n782), .A3(n781), .ZN(curr_proc_regs[347])
         );
  NAND2_X1 U1245 ( .A1(regs[860]), .A2(n8), .ZN(n786) );
  AOI22_X1 U1246 ( .A1(n18), .A2(regs[1372]), .B1(n37), .B2(regs[348]), .ZN(
        n785) );
  AOI22_X1 U1247 ( .A1(n135), .A2(regs[2396]), .B1(n73), .B2(regs[1884]), .ZN(
        n784) );
  NAND3_X1 U1248 ( .A1(n786), .A2(n785), .A3(n784), .ZN(curr_proc_regs[348])
         );
  NAND2_X1 U1249 ( .A1(regs[861]), .A2(n61), .ZN(n789) );
  AOI22_X1 U1250 ( .A1(n18), .A2(regs[1373]), .B1(n39), .B2(regs[349]), .ZN(
        n788) );
  AOI22_X1 U1251 ( .A1(n135), .A2(regs[2397]), .B1(n15), .B2(regs[1885]), .ZN(
        n787) );
  NAND3_X1 U1252 ( .A1(n789), .A2(n788), .A3(n787), .ZN(curr_proc_regs[349])
         );
  INV_X1 U1253 ( .A(regs[546]), .ZN(n1421) );
  AOI22_X1 U1254 ( .A1(n135), .A2(regs[2082]), .B1(n67), .B2(regs[1570]), .ZN(
        n791) );
  AOI22_X1 U1255 ( .A1(n91), .A2(regs[1058]), .B1(n37), .B2(regs[34]), .ZN(
        n790) );
  OAI211_X1 U1256 ( .C1(n11), .C2(n1421), .A(n791), .B(n790), .ZN(
        curr_proc_regs[34]) );
  NAND2_X1 U1257 ( .A1(regs[862]), .A2(n61), .ZN(n794) );
  AOI22_X1 U1258 ( .A1(n89), .A2(regs[1374]), .B1(n39), .B2(regs[350]), .ZN(
        n793) );
  AOI22_X1 U1259 ( .A1(n135), .A2(regs[2398]), .B1(n17), .B2(regs[1886]), .ZN(
        n792) );
  NAND3_X1 U1260 ( .A1(n794), .A2(n793), .A3(n792), .ZN(curr_proc_regs[350])
         );
  NAND2_X1 U1261 ( .A1(regs[863]), .A2(n59), .ZN(n797) );
  AOI22_X1 U1262 ( .A1(n92), .A2(regs[1375]), .B1(n36), .B2(regs[351]), .ZN(
        n796) );
  AOI22_X1 U1263 ( .A1(n135), .A2(regs[2399]), .B1(n69), .B2(regs[1887]), .ZN(
        n795) );
  NAND3_X1 U1264 ( .A1(n797), .A2(n796), .A3(n795), .ZN(curr_proc_regs[351])
         );
  NAND2_X1 U1265 ( .A1(regs[864]), .A2(n2), .ZN(n800) );
  AOI22_X1 U1266 ( .A1(n90), .A2(regs[1376]), .B1(n36), .B2(regs[352]), .ZN(
        n799) );
  AOI22_X1 U1267 ( .A1(n122), .A2(regs[2400]), .B1(n73), .B2(regs[1888]), .ZN(
        n798) );
  NAND3_X1 U1268 ( .A1(n800), .A2(n799), .A3(n798), .ZN(curr_proc_regs[352])
         );
  NAND2_X1 U1269 ( .A1(regs[1377]), .A2(n81), .ZN(n803) );
  AOI22_X1 U1270 ( .A1(n50), .A2(regs[865]), .B1(n36), .B2(regs[353]), .ZN(
        n802) );
  AOI22_X1 U1271 ( .A1(n123), .A2(regs[2401]), .B1(n73), .B2(regs[1889]), .ZN(
        n801) );
  NAND3_X1 U1272 ( .A1(n803), .A2(n802), .A3(n801), .ZN(curr_proc_regs[353])
         );
  NAND2_X1 U1273 ( .A1(regs[866]), .A2(n2), .ZN(n806) );
  AOI22_X1 U1274 ( .A1(n18), .A2(regs[1378]), .B1(n36), .B2(regs[354]), .ZN(
        n805) );
  AOI22_X1 U1275 ( .A1(n124), .A2(regs[2402]), .B1(n17), .B2(regs[1890]), .ZN(
        n804) );
  NAND3_X1 U1276 ( .A1(n806), .A2(n805), .A3(n804), .ZN(curr_proc_regs[354])
         );
  NAND2_X1 U1277 ( .A1(regs[867]), .A2(n61), .ZN(n809) );
  AOI22_X1 U1278 ( .A1(n91), .A2(regs[1379]), .B1(n36), .B2(regs[355]), .ZN(
        n808) );
  AOI22_X1 U1279 ( .A1(n125), .A2(regs[2403]), .B1(n17), .B2(regs[1891]), .ZN(
        n807) );
  NAND3_X1 U1280 ( .A1(n809), .A2(n808), .A3(n807), .ZN(curr_proc_regs[355])
         );
  NAND2_X1 U1281 ( .A1(regs[868]), .A2(n61), .ZN(n812) );
  AOI22_X1 U1282 ( .A1(n18), .A2(regs[1380]), .B1(n36), .B2(regs[356]), .ZN(
        n811) );
  AOI22_X1 U1283 ( .A1(n122), .A2(regs[2404]), .B1(n69), .B2(regs[1892]), .ZN(
        n810) );
  NAND3_X1 U1284 ( .A1(n812), .A2(n811), .A3(n810), .ZN(curr_proc_regs[356])
         );
  NAND2_X1 U1285 ( .A1(regs[869]), .A2(n61), .ZN(n815) );
  AOI22_X1 U1286 ( .A1(n88), .A2(regs[1381]), .B1(n36), .B2(regs[357]), .ZN(
        n814) );
  AOI22_X1 U1287 ( .A1(n131), .A2(regs[2405]), .B1(n73), .B2(regs[1893]), .ZN(
        n813) );
  NAND3_X1 U1288 ( .A1(n815), .A2(n814), .A3(n813), .ZN(curr_proc_regs[357])
         );
  NAND2_X1 U1289 ( .A1(regs[870]), .A2(n13), .ZN(n818) );
  AOI22_X1 U1290 ( .A1(n93), .A2(regs[1382]), .B1(n37), .B2(regs[358]), .ZN(
        n817) );
  AOI22_X1 U1291 ( .A1(n126), .A2(regs[2406]), .B1(n72), .B2(regs[1894]), .ZN(
        n816) );
  NAND3_X1 U1292 ( .A1(n818), .A2(n817), .A3(n816), .ZN(curr_proc_regs[358])
         );
  NAND2_X1 U1293 ( .A1(regs[871]), .A2(n13), .ZN(n821) );
  AOI22_X1 U1294 ( .A1(n93), .A2(regs[1383]), .B1(n39), .B2(regs[359]), .ZN(
        n820) );
  AOI22_X1 U1295 ( .A1(n136), .A2(regs[2407]), .B1(n72), .B2(regs[1895]), .ZN(
        n819) );
  NAND3_X1 U1296 ( .A1(n821), .A2(n820), .A3(n819), .ZN(curr_proc_regs[359])
         );
  INV_X1 U1297 ( .A(regs[1059]), .ZN(n1424) );
  AOI22_X1 U1298 ( .A1(n135), .A2(regs[2083]), .B1(n72), .B2(regs[1571]), .ZN(
        n823) );
  AOI22_X1 U1299 ( .A1(n8), .A2(regs[547]), .B1(n39), .B2(regs[35]), .ZN(n822)
         );
  OAI211_X1 U1300 ( .C1(n5), .C2(n1424), .A(n823), .B(n822), .ZN(
        curr_proc_regs[35]) );
  NAND2_X1 U1301 ( .A1(regs[872]), .A2(n13), .ZN(n826) );
  AOI22_X1 U1302 ( .A1(n18), .A2(regs[1384]), .B1(n38), .B2(regs[360]), .ZN(
        n825) );
  AOI22_X1 U1303 ( .A1(n134), .A2(regs[2408]), .B1(n72), .B2(regs[1896]), .ZN(
        n824) );
  NAND3_X1 U1304 ( .A1(n826), .A2(n825), .A3(n824), .ZN(curr_proc_regs[360])
         );
  NAND2_X1 U1305 ( .A1(regs[1385]), .A2(n98), .ZN(n829) );
  AOI22_X1 U1306 ( .A1(n51), .A2(regs[873]), .B1(n39), .B2(regs[361]), .ZN(
        n828) );
  AOI22_X1 U1307 ( .A1(n134), .A2(regs[2409]), .B1(n72), .B2(regs[1897]), .ZN(
        n827) );
  NAND3_X1 U1308 ( .A1(n829), .A2(n828), .A3(n827), .ZN(curr_proc_regs[361])
         );
  NAND2_X1 U1309 ( .A1(regs[1386]), .A2(n84), .ZN(n832) );
  AOI22_X1 U1310 ( .A1(n51), .A2(regs[874]), .B1(n38), .B2(regs[362]), .ZN(
        n831) );
  AOI22_X1 U1311 ( .A1(n134), .A2(regs[2410]), .B1(n72), .B2(regs[1898]), .ZN(
        n830) );
  NAND3_X1 U1312 ( .A1(n832), .A2(n831), .A3(n830), .ZN(curr_proc_regs[362])
         );
  NAND2_X1 U1313 ( .A1(regs[875]), .A2(n60), .ZN(n835) );
  AOI22_X1 U1314 ( .A1(n18), .A2(regs[1387]), .B1(n37), .B2(regs[363]), .ZN(
        n834) );
  AOI22_X1 U1315 ( .A1(n134), .A2(regs[2411]), .B1(n72), .B2(regs[1899]), .ZN(
        n833) );
  NAND3_X1 U1316 ( .A1(n835), .A2(n834), .A3(n833), .ZN(curr_proc_regs[363])
         );
  NAND2_X1 U1317 ( .A1(regs[876]), .A2(n13), .ZN(n838) );
  AOI22_X1 U1318 ( .A1(n80), .A2(regs[1388]), .B1(n37), .B2(regs[364]), .ZN(
        n837) );
  AOI22_X1 U1319 ( .A1(n134), .A2(regs[2412]), .B1(n72), .B2(regs[1900]), .ZN(
        n836) );
  NAND3_X1 U1320 ( .A1(n838), .A2(n837), .A3(n836), .ZN(curr_proc_regs[364])
         );
  NAND2_X1 U1321 ( .A1(regs[877]), .A2(n2), .ZN(n841) );
  AOI22_X1 U1322 ( .A1(n94), .A2(regs[1389]), .B1(n38), .B2(regs[365]), .ZN(
        n840) );
  AOI22_X1 U1323 ( .A1(n134), .A2(regs[2413]), .B1(n72), .B2(regs[1901]), .ZN(
        n839) );
  NAND3_X1 U1324 ( .A1(n841), .A2(n840), .A3(n839), .ZN(curr_proc_regs[365])
         );
  NAND2_X1 U1325 ( .A1(regs[1390]), .A2(n86), .ZN(n844) );
  AOI22_X1 U1326 ( .A1(n57), .A2(regs[878]), .B1(n39), .B2(regs[366]), .ZN(
        n843) );
  AOI22_X1 U1327 ( .A1(n134), .A2(regs[2414]), .B1(n72), .B2(regs[1902]), .ZN(
        n842) );
  NAND3_X1 U1328 ( .A1(n844), .A2(n843), .A3(n842), .ZN(curr_proc_regs[366])
         );
  NAND2_X1 U1329 ( .A1(regs[1391]), .A2(n98), .ZN(n847) );
  AOI22_X1 U1330 ( .A1(n55), .A2(regs[879]), .B1(n38), .B2(regs[367]), .ZN(
        n846) );
  AOI22_X1 U1331 ( .A1(n134), .A2(regs[2415]), .B1(n72), .B2(regs[1903]), .ZN(
        n845) );
  NAND3_X1 U1332 ( .A1(n847), .A2(n846), .A3(n845), .ZN(curr_proc_regs[367])
         );
  NAND2_X1 U1333 ( .A1(regs[1392]), .A2(n19), .ZN(n850) );
  AOI22_X1 U1334 ( .A1(n54), .A2(regs[880]), .B1(n37), .B2(regs[368]), .ZN(
        n849) );
  AOI22_X1 U1335 ( .A1(n134), .A2(regs[2416]), .B1(n73), .B2(regs[1904]), .ZN(
        n848) );
  NAND3_X1 U1336 ( .A1(n850), .A2(n849), .A3(n848), .ZN(curr_proc_regs[368])
         );
  NAND2_X1 U1337 ( .A1(regs[1393]), .A2(n19), .ZN(n853) );
  AOI22_X1 U1338 ( .A1(n50), .A2(regs[881]), .B1(n39), .B2(regs[369]), .ZN(
        n852) );
  AOI22_X1 U1339 ( .A1(n134), .A2(regs[2417]), .B1(n74), .B2(regs[1905]), .ZN(
        n851) );
  NAND3_X1 U1340 ( .A1(n853), .A2(n852), .A3(n851), .ZN(curr_proc_regs[369])
         );
  INV_X1 U1341 ( .A(regs[1060]), .ZN(n1427) );
  AOI22_X1 U1342 ( .A1(n134), .A2(regs[2084]), .B1(n70), .B2(regs[1572]), .ZN(
        n855) );
  AOI22_X1 U1343 ( .A1(n57), .A2(regs[548]), .B1(n38), .B2(regs[36]), .ZN(n854) );
  OAI211_X1 U1344 ( .C1(n99), .C2(n1427), .A(n855), .B(n854), .ZN(
        curr_proc_regs[36]) );
  NAND2_X1 U1345 ( .A1(regs[1394]), .A2(n19), .ZN(n858) );
  AOI22_X1 U1346 ( .A1(n58), .A2(regs[882]), .B1(n37), .B2(regs[370]), .ZN(
        n857) );
  AOI22_X1 U1347 ( .A1(n133), .A2(regs[2418]), .B1(n69), .B2(regs[1906]), .ZN(
        n856) );
  NAND3_X1 U1348 ( .A1(n858), .A2(n857), .A3(n856), .ZN(curr_proc_regs[370])
         );
  NAND2_X1 U1349 ( .A1(regs[883]), .A2(n2), .ZN(n861) );
  AOI22_X1 U1350 ( .A1(n18), .A2(regs[1395]), .B1(n38), .B2(regs[371]), .ZN(
        n860) );
  AOI22_X1 U1351 ( .A1(n133), .A2(regs[2419]), .B1(n17), .B2(regs[1907]), .ZN(
        n859) );
  NAND3_X1 U1352 ( .A1(n861), .A2(n860), .A3(n859), .ZN(curr_proc_regs[371])
         );
  NAND2_X1 U1353 ( .A1(regs[1396]), .A2(n19), .ZN(n864) );
  AOI22_X1 U1354 ( .A1(n57), .A2(regs[884]), .B1(n39), .B2(regs[372]), .ZN(
        n863) );
  AOI22_X1 U1355 ( .A1(n133), .A2(regs[2420]), .B1(n73), .B2(regs[1908]), .ZN(
        n862) );
  NAND3_X1 U1356 ( .A1(n864), .A2(n863), .A3(n862), .ZN(curr_proc_regs[372])
         );
  NAND2_X1 U1357 ( .A1(regs[885]), .A2(n13), .ZN(n867) );
  AOI22_X1 U1358 ( .A1(n18), .A2(regs[1397]), .B1(n38), .B2(regs[373]), .ZN(
        n866) );
  AOI22_X1 U1359 ( .A1(n133), .A2(regs[2421]), .B1(n72), .B2(regs[1909]), .ZN(
        n865) );
  NAND3_X1 U1360 ( .A1(n867), .A2(n866), .A3(n865), .ZN(curr_proc_regs[373])
         );
  NAND2_X1 U1361 ( .A1(regs[886]), .A2(n13), .ZN(n870) );
  AOI22_X1 U1362 ( .A1(n18), .A2(regs[1398]), .B1(n37), .B2(regs[374]), .ZN(
        n869) );
  AOI22_X1 U1363 ( .A1(n133), .A2(regs[2422]), .B1(n73), .B2(regs[1910]), .ZN(
        n868) );
  NAND3_X1 U1364 ( .A1(n870), .A2(n869), .A3(n868), .ZN(curr_proc_regs[374])
         );
  NAND2_X1 U1365 ( .A1(regs[887]), .A2(n2), .ZN(n873) );
  AOI22_X1 U1366 ( .A1(n93), .A2(regs[1399]), .B1(n37), .B2(regs[375]), .ZN(
        n872) );
  AOI22_X1 U1367 ( .A1(n133), .A2(regs[2423]), .B1(n66), .B2(regs[1911]), .ZN(
        n871) );
  NAND3_X1 U1368 ( .A1(n873), .A2(n872), .A3(n871), .ZN(curr_proc_regs[375])
         );
  NAND2_X1 U1369 ( .A1(regs[1400]), .A2(n19), .ZN(n876) );
  AOI22_X1 U1370 ( .A1(n50), .A2(regs[888]), .B1(n39), .B2(regs[376]), .ZN(
        n875) );
  AOI22_X1 U1371 ( .A1(n133), .A2(regs[2424]), .B1(n17), .B2(regs[1912]), .ZN(
        n874) );
  NAND3_X1 U1372 ( .A1(n876), .A2(n875), .A3(n874), .ZN(curr_proc_regs[376])
         );
  NAND2_X1 U1373 ( .A1(regs[889]), .A2(n2), .ZN(n879) );
  AOI22_X1 U1374 ( .A1(n18), .A2(regs[1401]), .B1(n38), .B2(regs[377]), .ZN(
        n878) );
  AOI22_X1 U1375 ( .A1(n133), .A2(regs[2425]), .B1(n15), .B2(regs[1913]), .ZN(
        n877) );
  NAND3_X1 U1376 ( .A1(n879), .A2(n878), .A3(n877), .ZN(curr_proc_regs[377])
         );
  NAND2_X1 U1377 ( .A1(regs[890]), .A2(n13), .ZN(n882) );
  AOI22_X1 U1378 ( .A1(n89), .A2(regs[1402]), .B1(n37), .B2(regs[378]), .ZN(
        n881) );
  AOI22_X1 U1379 ( .A1(n133), .A2(regs[2426]), .B1(n73), .B2(regs[1914]), .ZN(
        n880) );
  NAND3_X1 U1380 ( .A1(n882), .A2(n881), .A3(n880), .ZN(curr_proc_regs[378])
         );
  NAND2_X1 U1381 ( .A1(regs[1403]), .A2(n19), .ZN(n885) );
  AOI22_X1 U1382 ( .A1(n58), .A2(regs[891]), .B1(n37), .B2(regs[379]), .ZN(
        n884) );
  AOI22_X1 U1383 ( .A1(n133), .A2(regs[2427]), .B1(n73), .B2(regs[1915]), .ZN(
        n883) );
  NAND3_X1 U1384 ( .A1(n885), .A2(n884), .A3(n883), .ZN(curr_proc_regs[379])
         );
  INV_X1 U1385 ( .A(regs[549]), .ZN(n1430) );
  AOI22_X1 U1386 ( .A1(n133), .A2(regs[2085]), .B1(n73), .B2(regs[1573]), .ZN(
        n887) );
  AOI22_X1 U1387 ( .A1(n91), .A2(regs[1061]), .B1(n37), .B2(regs[37]), .ZN(
        n886) );
  OAI211_X1 U1388 ( .C1(n11), .C2(n1430), .A(n887), .B(n886), .ZN(
        curr_proc_regs[37]) );
  NAND2_X1 U1389 ( .A1(regs[1404]), .A2(n19), .ZN(n890) );
  AOI22_X1 U1390 ( .A1(n58), .A2(regs[892]), .B1(n37), .B2(regs[380]), .ZN(
        n889) );
  AOI22_X1 U1391 ( .A1(n132), .A2(regs[2428]), .B1(n73), .B2(regs[1916]), .ZN(
        n888) );
  NAND3_X1 U1392 ( .A1(n890), .A2(n889), .A3(n888), .ZN(curr_proc_regs[380])
         );
  NAND2_X1 U1393 ( .A1(regs[893]), .A2(n2), .ZN(n893) );
  AOI22_X1 U1394 ( .A1(n93), .A2(regs[1405]), .B1(n38), .B2(regs[381]), .ZN(
        n892) );
  AOI22_X1 U1395 ( .A1(n132), .A2(regs[2429]), .B1(n73), .B2(regs[1917]), .ZN(
        n891) );
  NAND3_X1 U1396 ( .A1(n893), .A2(n892), .A3(n891), .ZN(curr_proc_regs[381])
         );
  NAND2_X1 U1397 ( .A1(regs[1406]), .A2(n90), .ZN(n896) );
  AOI22_X1 U1398 ( .A1(n13), .A2(regs[894]), .B1(n37), .B2(regs[382]), .ZN(
        n895) );
  AOI22_X1 U1399 ( .A1(n132), .A2(regs[2430]), .B1(n73), .B2(regs[1918]), .ZN(
        n894) );
  NAND3_X1 U1400 ( .A1(n896), .A2(n895), .A3(n894), .ZN(curr_proc_regs[382])
         );
  NAND2_X1 U1401 ( .A1(regs[895]), .A2(n2), .ZN(n899) );
  AOI22_X1 U1402 ( .A1(n81), .A2(regs[1407]), .B1(n39), .B2(regs[383]), .ZN(
        n898) );
  AOI22_X1 U1403 ( .A1(n132), .A2(regs[2431]), .B1(n73), .B2(regs[1919]), .ZN(
        n897) );
  NAND3_X1 U1404 ( .A1(n899), .A2(n898), .A3(n897), .ZN(curr_proc_regs[383])
         );
  NAND2_X1 U1405 ( .A1(regs[1408]), .A2(n95), .ZN(n902) );
  AOI22_X1 U1406 ( .A1(n56), .A2(regs[896]), .B1(n38), .B2(regs[384]), .ZN(
        n901) );
  AOI22_X1 U1407 ( .A1(n132), .A2(regs[2432]), .B1(n73), .B2(regs[1920]), .ZN(
        n900) );
  NAND3_X1 U1408 ( .A1(n902), .A2(n901), .A3(n900), .ZN(curr_proc_regs[384])
         );
  NAND2_X1 U1409 ( .A1(regs[897]), .A2(n2), .ZN(n905) );
  AOI22_X1 U1410 ( .A1(n81), .A2(regs[1409]), .B1(n37), .B2(regs[385]), .ZN(
        n904) );
  AOI22_X1 U1411 ( .A1(n132), .A2(regs[2433]), .B1(n73), .B2(regs[1921]), .ZN(
        n903) );
  NAND3_X1 U1412 ( .A1(n905), .A2(n904), .A3(n903), .ZN(curr_proc_regs[385])
         );
  NAND2_X1 U1413 ( .A1(regs[898]), .A2(n8), .ZN(n908) );
  AOI22_X1 U1414 ( .A1(n81), .A2(regs[1410]), .B1(n39), .B2(regs[386]), .ZN(
        n907) );
  AOI22_X1 U1415 ( .A1(n132), .A2(regs[2434]), .B1(n73), .B2(regs[1922]), .ZN(
        n906) );
  NAND3_X1 U1416 ( .A1(n908), .A2(n907), .A3(n906), .ZN(curr_proc_regs[386])
         );
  NAND2_X1 U1417 ( .A1(regs[899]), .A2(n8), .ZN(n911) );
  AOI22_X1 U1418 ( .A1(n81), .A2(regs[1411]), .B1(n38), .B2(regs[387]), .ZN(
        n910) );
  AOI22_X1 U1419 ( .A1(n132), .A2(regs[2435]), .B1(n73), .B2(regs[1923]), .ZN(
        n909) );
  NAND3_X1 U1420 ( .A1(n911), .A2(n910), .A3(n909), .ZN(curr_proc_regs[387])
         );
  NAND2_X1 U1421 ( .A1(regs[1412]), .A2(n19), .ZN(n914) );
  AOI22_X1 U1422 ( .A1(n55), .A2(regs[900]), .B1(n38), .B2(regs[388]), .ZN(
        n913) );
  AOI22_X1 U1423 ( .A1(n132), .A2(regs[2436]), .B1(n69), .B2(regs[1924]), .ZN(
        n912) );
  NAND3_X1 U1424 ( .A1(n914), .A2(n913), .A3(n912), .ZN(curr_proc_regs[388])
         );
  NAND2_X1 U1425 ( .A1(regs[1413]), .A2(n19), .ZN(n917) );
  AOI22_X1 U1426 ( .A1(n51), .A2(regs[901]), .B1(n38), .B2(regs[389]), .ZN(
        n916) );
  AOI22_X1 U1427 ( .A1(n132), .A2(regs[2437]), .B1(n17), .B2(regs[1925]), .ZN(
        n915) );
  NAND3_X1 U1428 ( .A1(n917), .A2(n916), .A3(n915), .ZN(curr_proc_regs[389])
         );
  INV_X1 U1429 ( .A(regs[550]), .ZN(n1435) );
  AOI22_X1 U1430 ( .A1(n132), .A2(regs[2086]), .B1(n69), .B2(regs[1574]), .ZN(
        n919) );
  AOI22_X1 U1431 ( .A1(n81), .A2(regs[1062]), .B1(n38), .B2(regs[38]), .ZN(
        n918) );
  OAI211_X1 U1432 ( .C1(n11), .C2(n1435), .A(n919), .B(n918), .ZN(
        curr_proc_regs[38]) );
  NAND2_X1 U1433 ( .A1(regs[1414]), .A2(n97), .ZN(n922) );
  AOI22_X1 U1434 ( .A1(n50), .A2(regs[902]), .B1(n38), .B2(regs[390]), .ZN(
        n921) );
  AOI22_X1 U1435 ( .A1(n131), .A2(regs[2438]), .B1(n14), .B2(regs[1926]), .ZN(
        n920) );
  NAND3_X1 U1436 ( .A1(n922), .A2(n921), .A3(n920), .ZN(curr_proc_regs[390])
         );
  NAND2_X1 U1437 ( .A1(regs[903]), .A2(n8), .ZN(n925) );
  AOI22_X1 U1438 ( .A1(n81), .A2(regs[1415]), .B1(n37), .B2(regs[391]), .ZN(
        n924) );
  AOI22_X1 U1439 ( .A1(n131), .A2(regs[2439]), .B1(n69), .B2(regs[1927]), .ZN(
        n923) );
  NAND3_X1 U1440 ( .A1(n925), .A2(n924), .A3(n923), .ZN(curr_proc_regs[391])
         );
  NAND2_X1 U1441 ( .A1(regs[904]), .A2(n2), .ZN(n928) );
  AOI22_X1 U1442 ( .A1(n81), .A2(regs[1416]), .B1(n37), .B2(regs[392]), .ZN(
        n927) );
  AOI22_X1 U1443 ( .A1(n131), .A2(regs[2440]), .B1(n4), .B2(regs[1928]), .ZN(
        n926) );
  NAND3_X1 U1444 ( .A1(n928), .A2(n927), .A3(n926), .ZN(curr_proc_regs[392])
         );
  NAND2_X1 U1445 ( .A1(regs[905]), .A2(n8), .ZN(n931) );
  AOI22_X1 U1446 ( .A1(n81), .A2(regs[1417]), .B1(n37), .B2(regs[393]), .ZN(
        n930) );
  AOI22_X1 U1447 ( .A1(n131), .A2(regs[2441]), .B1(n69), .B2(regs[1929]), .ZN(
        n929) );
  NAND3_X1 U1448 ( .A1(n931), .A2(n930), .A3(n929), .ZN(curr_proc_regs[393])
         );
  NAND2_X1 U1449 ( .A1(regs[1418]), .A2(n19), .ZN(n934) );
  AOI22_X1 U1450 ( .A1(n62), .A2(regs[906]), .B1(n37), .B2(regs[394]), .ZN(
        n933) );
  AOI22_X1 U1451 ( .A1(n131), .A2(regs[2442]), .B1(n4), .B2(regs[1930]), .ZN(
        n932) );
  NAND3_X1 U1452 ( .A1(n934), .A2(n933), .A3(n932), .ZN(curr_proc_regs[394])
         );
  NAND2_X1 U1453 ( .A1(regs[907]), .A2(n60), .ZN(n937) );
  AOI22_X1 U1454 ( .A1(n81), .A2(regs[1419]), .B1(n37), .B2(regs[395]), .ZN(
        n936) );
  AOI22_X1 U1455 ( .A1(n131), .A2(regs[2443]), .B1(n76), .B2(regs[1931]), .ZN(
        n935) );
  NAND3_X1 U1456 ( .A1(n937), .A2(n936), .A3(n935), .ZN(curr_proc_regs[395])
         );
  NAND2_X1 U1457 ( .A1(regs[908]), .A2(n61), .ZN(n940) );
  AOI22_X1 U1458 ( .A1(n81), .A2(regs[1420]), .B1(n37), .B2(regs[396]), .ZN(
        n939) );
  AOI22_X1 U1459 ( .A1(n131), .A2(regs[2444]), .B1(n69), .B2(regs[1932]), .ZN(
        n938) );
  NAND3_X1 U1460 ( .A1(n940), .A2(n939), .A3(n938), .ZN(curr_proc_regs[396])
         );
  NAND2_X1 U1461 ( .A1(regs[909]), .A2(n8), .ZN(n943) );
  AOI22_X1 U1462 ( .A1(n98), .A2(regs[1421]), .B1(n37), .B2(regs[397]), .ZN(
        n942) );
  AOI22_X1 U1463 ( .A1(n131), .A2(regs[2445]), .B1(n75), .B2(regs[1933]), .ZN(
        n941) );
  NAND3_X1 U1464 ( .A1(n943), .A2(n942), .A3(n941), .ZN(curr_proc_regs[397])
         );
  NAND2_X1 U1465 ( .A1(regs[910]), .A2(n2), .ZN(n946) );
  AOI22_X1 U1466 ( .A1(n96), .A2(regs[1422]), .B1(n39), .B2(regs[398]), .ZN(
        n945) );
  AOI22_X1 U1467 ( .A1(n131), .A2(regs[2446]), .B1(n73), .B2(regs[1934]), .ZN(
        n944) );
  NAND3_X1 U1468 ( .A1(n946), .A2(n945), .A3(n944), .ZN(curr_proc_regs[398])
         );
  NAND2_X1 U1469 ( .A1(regs[1423]), .A2(n19), .ZN(n949) );
  AOI22_X1 U1470 ( .A1(n60), .A2(regs[911]), .B1(n39), .B2(regs[399]), .ZN(
        n948) );
  AOI22_X1 U1471 ( .A1(n131), .A2(regs[2447]), .B1(n73), .B2(regs[1935]), .ZN(
        n947) );
  NAND3_X1 U1472 ( .A1(n949), .A2(n948), .A3(n947), .ZN(curr_proc_regs[399])
         );
  INV_X1 U1473 ( .A(regs[551]), .ZN(n1438) );
  AOI22_X1 U1474 ( .A1(n131), .A2(regs[2087]), .B1(n73), .B2(regs[1575]), .ZN(
        n951) );
  AOI22_X1 U1475 ( .A1(n94), .A2(regs[1063]), .B1(n39), .B2(regs[39]), .ZN(
        n950) );
  OAI211_X1 U1476 ( .C1(n11), .C2(n1438), .A(n951), .B(n950), .ZN(
        curr_proc_regs[39]) );
  INV_X1 U1477 ( .A(regs[515]), .ZN(n1325) );
  AOI22_X1 U1478 ( .A1(n130), .A2(regs[2051]), .B1(n73), .B2(regs[1539]), .ZN(
        n953) );
  AOI22_X1 U1479 ( .A1(n96), .A2(regs[1027]), .B1(n39), .B2(regs[3]), .ZN(n952) );
  OAI211_X1 U1480 ( .C1(n2207), .C2(n1325), .A(n953), .B(n952), .ZN(
        curr_proc_regs[3]) );
  NAND2_X1 U1481 ( .A1(regs[912]), .A2(n8), .ZN(n956) );
  AOI22_X1 U1482 ( .A1(n96), .A2(regs[1424]), .B1(n38), .B2(regs[400]), .ZN(
        n955) );
  AOI22_X1 U1483 ( .A1(n130), .A2(regs[2448]), .B1(n73), .B2(regs[1936]), .ZN(
        n954) );
  NAND3_X1 U1484 ( .A1(n956), .A2(n955), .A3(n954), .ZN(curr_proc_regs[400])
         );
  NAND2_X1 U1485 ( .A1(regs[913]), .A2(n2), .ZN(n959) );
  AOI22_X1 U1486 ( .A1(n95), .A2(regs[1425]), .B1(n38), .B2(regs[401]), .ZN(
        n958) );
  AOI22_X1 U1487 ( .A1(n130), .A2(regs[2449]), .B1(n73), .B2(regs[1937]), .ZN(
        n957) );
  NAND3_X1 U1488 ( .A1(n959), .A2(n958), .A3(n957), .ZN(curr_proc_regs[401])
         );
  NAND2_X1 U1489 ( .A1(regs[1426]), .A2(n19), .ZN(n962) );
  AOI22_X1 U1490 ( .A1(n50), .A2(regs[914]), .B1(n38), .B2(regs[402]), .ZN(
        n961) );
  AOI22_X1 U1491 ( .A1(n130), .A2(regs[2450]), .B1(n73), .B2(regs[1938]), .ZN(
        n960) );
  NAND3_X1 U1492 ( .A1(n962), .A2(n961), .A3(n960), .ZN(curr_proc_regs[402])
         );
  NAND2_X1 U1493 ( .A1(regs[1427]), .A2(n85), .ZN(n965) );
  AOI22_X1 U1494 ( .A1(n60), .A2(regs[915]), .B1(n38), .B2(regs[403]), .ZN(
        n964) );
  AOI22_X1 U1495 ( .A1(n130), .A2(regs[2451]), .B1(n73), .B2(regs[1939]), .ZN(
        n963) );
  NAND3_X1 U1496 ( .A1(n965), .A2(n964), .A3(n963), .ZN(curr_proc_regs[403])
         );
  NAND2_X1 U1497 ( .A1(regs[1428]), .A2(n19), .ZN(n968) );
  AOI22_X1 U1498 ( .A1(n51), .A2(regs[916]), .B1(n38), .B2(regs[404]), .ZN(
        n967) );
  AOI22_X1 U1499 ( .A1(n130), .A2(regs[2452]), .B1(n73), .B2(regs[1940]), .ZN(
        n966) );
  NAND3_X1 U1500 ( .A1(n968), .A2(n967), .A3(n966), .ZN(curr_proc_regs[404])
         );
  NAND2_X1 U1501 ( .A1(regs[917]), .A2(n8), .ZN(n971) );
  AOI22_X1 U1502 ( .A1(n94), .A2(regs[1429]), .B1(n38), .B2(regs[405]), .ZN(
        n970) );
  AOI22_X1 U1503 ( .A1(n130), .A2(regs[2453]), .B1(n73), .B2(regs[1941]), .ZN(
        n969) );
  NAND3_X1 U1504 ( .A1(n971), .A2(n970), .A3(n969), .ZN(curr_proc_regs[405])
         );
  NAND2_X1 U1505 ( .A1(regs[1430]), .A2(n19), .ZN(n974) );
  AOI22_X1 U1506 ( .A1(n60), .A2(regs[918]), .B1(n38), .B2(regs[406]), .ZN(
        n973) );
  AOI22_X1 U1507 ( .A1(n130), .A2(regs[2454]), .B1(n73), .B2(regs[1942]), .ZN(
        n972) );
  NAND3_X1 U1508 ( .A1(n974), .A2(n973), .A3(n972), .ZN(curr_proc_regs[406])
         );
  NAND2_X1 U1509 ( .A1(regs[919]), .A2(n2), .ZN(n977) );
  AOI22_X1 U1510 ( .A1(n80), .A2(regs[1431]), .B1(n39), .B2(regs[407]), .ZN(
        n976) );
  AOI22_X1 U1511 ( .A1(n130), .A2(regs[2455]), .B1(n68), .B2(regs[1943]), .ZN(
        n975) );
  NAND3_X1 U1512 ( .A1(n977), .A2(n976), .A3(n975), .ZN(curr_proc_regs[407])
         );
  NAND2_X1 U1513 ( .A1(regs[1432]), .A2(n98), .ZN(n980) );
  AOI22_X1 U1514 ( .A1(n61), .A2(regs[920]), .B1(n38), .B2(regs[408]), .ZN(
        n979) );
  AOI22_X1 U1515 ( .A1(n130), .A2(regs[2456]), .B1(n72), .B2(regs[1944]), .ZN(
        n978) );
  NAND3_X1 U1516 ( .A1(n980), .A2(n979), .A3(n978), .ZN(curr_proc_regs[408])
         );
  NAND2_X1 U1517 ( .A1(regs[921]), .A2(n13), .ZN(n983) );
  AOI22_X1 U1518 ( .A1(n80), .A2(regs[1433]), .B1(n37), .B2(regs[409]), .ZN(
        n982) );
  AOI22_X1 U1519 ( .A1(n130), .A2(regs[2457]), .B1(n68), .B2(regs[1945]), .ZN(
        n981) );
  NAND3_X1 U1520 ( .A1(n983), .A2(n982), .A3(n981), .ZN(curr_proc_regs[409])
         );
  INV_X1 U1521 ( .A(regs[552]), .ZN(n1441) );
  AOI22_X1 U1522 ( .A1(n129), .A2(regs[2088]), .B1(n72), .B2(regs[1576]), .ZN(
        n985) );
  AOI22_X1 U1523 ( .A1(n81), .A2(regs[1064]), .B1(n27), .B2(regs[40]), .ZN(
        n984) );
  OAI211_X1 U1524 ( .C1(n11), .C2(n1441), .A(n985), .B(n984), .ZN(
        curr_proc_regs[40]) );
  NAND2_X1 U1525 ( .A1(regs[1434]), .A2(n78), .ZN(n988) );
  AOI22_X1 U1526 ( .A1(n52), .A2(regs[922]), .B1(n39), .B2(regs[410]), .ZN(
        n987) );
  AOI22_X1 U1527 ( .A1(n129), .A2(regs[2458]), .B1(n72), .B2(regs[1946]), .ZN(
        n986) );
  NAND3_X1 U1528 ( .A1(n988), .A2(n987), .A3(n986), .ZN(curr_proc_regs[410])
         );
  NAND2_X1 U1529 ( .A1(regs[1435]), .A2(n83), .ZN(n991) );
  AOI22_X1 U1530 ( .A1(n53), .A2(regs[923]), .B1(n39), .B2(regs[411]), .ZN(
        n990) );
  AOI22_X1 U1531 ( .A1(n129), .A2(regs[2459]), .B1(n72), .B2(regs[1947]), .ZN(
        n989) );
  NAND3_X1 U1532 ( .A1(n991), .A2(n990), .A3(n989), .ZN(curr_proc_regs[411])
         );
  NAND2_X1 U1533 ( .A1(regs[924]), .A2(n13), .ZN(n994) );
  AOI22_X1 U1534 ( .A1(n82), .A2(regs[1436]), .B1(n39), .B2(regs[412]), .ZN(
        n993) );
  AOI22_X1 U1535 ( .A1(n129), .A2(regs[2460]), .B1(n72), .B2(regs[1948]), .ZN(
        n992) );
  NAND3_X1 U1536 ( .A1(n994), .A2(n993), .A3(n992), .ZN(curr_proc_regs[412])
         );
  NAND2_X1 U1537 ( .A1(regs[1437]), .A2(n86), .ZN(n997) );
  AOI22_X1 U1538 ( .A1(n10), .A2(regs[925]), .B1(n39), .B2(regs[413]), .ZN(
        n996) );
  AOI22_X1 U1539 ( .A1(n129), .A2(regs[2461]), .B1(n72), .B2(regs[1949]), .ZN(
        n995) );
  NAND3_X1 U1540 ( .A1(n997), .A2(n996), .A3(n995), .ZN(curr_proc_regs[413])
         );
  NAND2_X1 U1541 ( .A1(regs[1438]), .A2(n79), .ZN(n1000) );
  AOI22_X1 U1542 ( .A1(n58), .A2(regs[926]), .B1(n39), .B2(regs[414]), .ZN(
        n999) );
  AOI22_X1 U1543 ( .A1(n129), .A2(regs[2462]), .B1(n72), .B2(regs[1950]), .ZN(
        n998) );
  NAND3_X1 U1544 ( .A1(n1000), .A2(n999), .A3(n998), .ZN(curr_proc_regs[414])
         );
  NAND2_X1 U1545 ( .A1(regs[927]), .A2(n2), .ZN(n1003) );
  AOI22_X1 U1546 ( .A1(n83), .A2(regs[1439]), .B1(n39), .B2(regs[415]), .ZN(
        n1002) );
  AOI22_X1 U1547 ( .A1(n129), .A2(regs[2463]), .B1(n72), .B2(regs[1951]), .ZN(
        n1001) );
  NAND3_X1 U1548 ( .A1(n1003), .A2(n1002), .A3(n1001), .ZN(curr_proc_regs[415]) );
  NAND2_X1 U1549 ( .A1(regs[1440]), .A2(n94), .ZN(n1006) );
  AOI22_X1 U1550 ( .A1(n57), .A2(regs[928]), .B1(n39), .B2(regs[416]), .ZN(
        n1005) );
  AOI22_X1 U1551 ( .A1(n129), .A2(regs[2464]), .B1(n72), .B2(regs[1952]), .ZN(
        n1004) );
  NAND3_X1 U1552 ( .A1(n1006), .A2(n1005), .A3(n1004), .ZN(curr_proc_regs[416]) );
  NAND2_X1 U1553 ( .A1(regs[929]), .A2(n2), .ZN(n1009) );
  AOI22_X1 U1554 ( .A1(n84), .A2(regs[1441]), .B1(n41), .B2(regs[417]), .ZN(
        n1008) );
  AOI22_X1 U1555 ( .A1(n129), .A2(regs[2465]), .B1(n77), .B2(regs[1953]), .ZN(
        n1007) );
  NAND3_X1 U1556 ( .A1(n1009), .A2(n1008), .A3(n1007), .ZN(curr_proc_regs[417]) );
  NAND2_X1 U1557 ( .A1(regs[1442]), .A2(n96), .ZN(n1012) );
  AOI22_X1 U1558 ( .A1(n2), .A2(regs[930]), .B1(n43), .B2(regs[418]), .ZN(
        n1011) );
  AOI22_X1 U1559 ( .A1(n129), .A2(regs[2466]), .B1(n76), .B2(regs[1954]), .ZN(
        n1010) );
  NAND3_X1 U1560 ( .A1(n1012), .A2(n1011), .A3(n1010), .ZN(curr_proc_regs[418]) );
  NAND2_X1 U1561 ( .A1(regs[1443]), .A2(n96), .ZN(n1015) );
  AOI22_X1 U1562 ( .A1(n51), .A2(regs[931]), .B1(n48), .B2(regs[419]), .ZN(
        n1014) );
  AOI22_X1 U1563 ( .A1(n129), .A2(regs[2467]), .B1(n75), .B2(regs[1955]), .ZN(
        n1013) );
  NAND3_X1 U1564 ( .A1(n1015), .A2(n1014), .A3(n1013), .ZN(curr_proc_regs[419]) );
  INV_X1 U1565 ( .A(regs[1065]), .ZN(n1444) );
  AOI22_X1 U1566 ( .A1(n128), .A2(regs[2089]), .B1(n69), .B2(regs[1577]), .ZN(
        n1017) );
  AOI22_X1 U1567 ( .A1(n2), .A2(regs[553]), .B1(n47), .B2(regs[41]), .ZN(n1016) );
  OAI211_X1 U1568 ( .C1(n16), .C2(n1444), .A(n1017), .B(n1016), .ZN(
        curr_proc_regs[41]) );
  NAND2_X1 U1569 ( .A1(regs[1444]), .A2(n96), .ZN(n1020) );
  AOI22_X1 U1570 ( .A1(n60), .A2(regs[932]), .B1(n43), .B2(regs[420]), .ZN(
        n1019) );
  AOI22_X1 U1571 ( .A1(n128), .A2(regs[2468]), .B1(n77), .B2(regs[1956]), .ZN(
        n1018) );
  NAND3_X1 U1572 ( .A1(n1020), .A2(n1019), .A3(n1018), .ZN(curr_proc_regs[420]) );
  NAND2_X1 U1573 ( .A1(regs[933]), .A2(n13), .ZN(n1023) );
  AOI22_X1 U1574 ( .A1(n85), .A2(regs[1445]), .B1(n48), .B2(regs[421]), .ZN(
        n1022) );
  AOI22_X1 U1575 ( .A1(n128), .A2(regs[2469]), .B1(n9), .B2(regs[1957]), .ZN(
        n1021) );
  NAND3_X1 U1576 ( .A1(n1023), .A2(n1022), .A3(n1021), .ZN(curr_proc_regs[421]) );
  NAND2_X1 U1577 ( .A1(regs[1446]), .A2(n95), .ZN(n1026) );
  AOI22_X1 U1578 ( .A1(n2), .A2(regs[934]), .B1(n47), .B2(regs[422]), .ZN(
        n1025) );
  AOI22_X1 U1579 ( .A1(n128), .A2(regs[2470]), .B1(n73), .B2(regs[1958]), .ZN(
        n1024) );
  NAND3_X1 U1580 ( .A1(n1026), .A2(n1025), .A3(n1024), .ZN(curr_proc_regs[422]) );
  NAND2_X1 U1581 ( .A1(regs[1447]), .A2(n95), .ZN(n1029) );
  AOI22_X1 U1582 ( .A1(n55), .A2(regs[935]), .B1(n46), .B2(regs[423]), .ZN(
        n1028) );
  AOI22_X1 U1583 ( .A1(n128), .A2(regs[2471]), .B1(n17), .B2(regs[1959]), .ZN(
        n1027) );
  NAND3_X1 U1584 ( .A1(n1029), .A2(n1028), .A3(n1027), .ZN(curr_proc_regs[423]) );
  NAND2_X1 U1585 ( .A1(regs[1448]), .A2(n95), .ZN(n1032) );
  AOI22_X1 U1586 ( .A1(n10), .A2(regs[936]), .B1(n30), .B2(regs[424]), .ZN(
        n1031) );
  AOI22_X1 U1587 ( .A1(n128), .A2(regs[2472]), .B1(n72), .B2(regs[1960]), .ZN(
        n1030) );
  NAND3_X1 U1588 ( .A1(n1032), .A2(n1031), .A3(n1030), .ZN(curr_proc_regs[424]) );
  NAND2_X1 U1589 ( .A1(regs[1449]), .A2(n95), .ZN(n1035) );
  AOI22_X1 U1590 ( .A1(n10), .A2(regs[937]), .B1(n29), .B2(regs[425]), .ZN(
        n1034) );
  AOI22_X1 U1591 ( .A1(n128), .A2(regs[2473]), .B1(n72), .B2(regs[1961]), .ZN(
        n1033) );
  NAND3_X1 U1592 ( .A1(n1035), .A2(n1034), .A3(n1033), .ZN(curr_proc_regs[425]) );
  NAND2_X1 U1593 ( .A1(regs[938]), .A2(n13), .ZN(n1038) );
  AOI22_X1 U1594 ( .A1(n86), .A2(regs[1450]), .B1(n28), .B2(regs[426]), .ZN(
        n1037) );
  AOI22_X1 U1595 ( .A1(n128), .A2(regs[2474]), .B1(n74), .B2(regs[1962]), .ZN(
        n1036) );
  NAND3_X1 U1596 ( .A1(n1038), .A2(n1037), .A3(n1036), .ZN(curr_proc_regs[426]) );
  NAND2_X1 U1597 ( .A1(regs[1451]), .A2(n94), .ZN(n1041) );
  AOI22_X1 U1598 ( .A1(n56), .A2(regs[939]), .B1(n31), .B2(regs[427]), .ZN(
        n1040) );
  AOI22_X1 U1599 ( .A1(n128), .A2(regs[2475]), .B1(n73), .B2(regs[1963]), .ZN(
        n1039) );
  NAND3_X1 U1600 ( .A1(n1041), .A2(n1040), .A3(n1039), .ZN(curr_proc_regs[427]) );
  NAND2_X1 U1601 ( .A1(regs[1452]), .A2(n94), .ZN(n1044) );
  AOI22_X1 U1602 ( .A1(n10), .A2(regs[940]), .B1(n30), .B2(regs[428]), .ZN(
        n1043) );
  AOI22_X1 U1603 ( .A1(n128), .A2(regs[2476]), .B1(n70), .B2(regs[1964]), .ZN(
        n1042) );
  NAND3_X1 U1604 ( .A1(n1044), .A2(n1043), .A3(n1042), .ZN(curr_proc_regs[428]) );
  NAND2_X1 U1605 ( .A1(regs[941]), .A2(n2), .ZN(n1047) );
  AOI22_X1 U1606 ( .A1(n87), .A2(regs[1453]), .B1(n29), .B2(regs[429]), .ZN(
        n1046) );
  AOI22_X1 U1607 ( .A1(n128), .A2(regs[2477]), .B1(n17), .B2(regs[1965]), .ZN(
        n1045) );
  NAND3_X1 U1608 ( .A1(n1047), .A2(n1046), .A3(n1045), .ZN(curr_proc_regs[429]) );
  INV_X1 U1609 ( .A(regs[1066]), .ZN(n1447) );
  AOI22_X1 U1610 ( .A1(n127), .A2(regs[2090]), .B1(n17), .B2(regs[1578]), .ZN(
        n1049) );
  AOI22_X1 U1611 ( .A1(n49), .A2(regs[554]), .B1(n35), .B2(regs[42]), .ZN(
        n1048) );
  OAI211_X1 U1612 ( .C1(n100), .C2(n1447), .A(n1049), .B(n1048), .ZN(
        curr_proc_regs[42]) );
  NAND2_X1 U1613 ( .A1(regs[942]), .A2(n13), .ZN(n1052) );
  AOI22_X1 U1614 ( .A1(n94), .A2(regs[1454]), .B1(n38), .B2(regs[430]), .ZN(
        n1051) );
  AOI22_X1 U1615 ( .A1(n127), .A2(regs[2478]), .B1(n17), .B2(regs[1966]), .ZN(
        n1050) );
  NAND3_X1 U1616 ( .A1(n1052), .A2(n1051), .A3(n1050), .ZN(curr_proc_regs[430]) );
  NAND2_X1 U1617 ( .A1(regs[1455]), .A2(n94), .ZN(n1055) );
  AOI22_X1 U1618 ( .A1(n10), .A2(regs[943]), .B1(n37), .B2(regs[431]), .ZN(
        n1054) );
  AOI22_X1 U1619 ( .A1(n127), .A2(regs[2479]), .B1(n73), .B2(regs[1967]), .ZN(
        n1053) );
  NAND3_X1 U1620 ( .A1(n1055), .A2(n1054), .A3(n1053), .ZN(curr_proc_regs[431]) );
  NAND2_X1 U1621 ( .A1(regs[1456]), .A2(n94), .ZN(n1058) );
  AOI22_X1 U1622 ( .A1(n56), .A2(regs[944]), .B1(n27), .B2(regs[432]), .ZN(
        n1057) );
  AOI22_X1 U1623 ( .A1(n127), .A2(regs[2480]), .B1(n72), .B2(regs[1968]), .ZN(
        n1056) );
  NAND3_X1 U1624 ( .A1(n1058), .A2(n1057), .A3(n1056), .ZN(curr_proc_regs[432]) );
  NAND2_X1 U1625 ( .A1(regs[945]), .A2(n13), .ZN(n1061) );
  AOI22_X1 U1626 ( .A1(n96), .A2(regs[1457]), .B1(n26), .B2(regs[433]), .ZN(
        n1060) );
  AOI22_X1 U1627 ( .A1(n127), .A2(regs[2481]), .B1(n72), .B2(regs[1969]), .ZN(
        n1059) );
  NAND3_X1 U1628 ( .A1(n1061), .A2(n1060), .A3(n1059), .ZN(curr_proc_regs[433]) );
  NAND2_X1 U1629 ( .A1(regs[1458]), .A2(n94), .ZN(n1064) );
  AOI22_X1 U1630 ( .A1(n56), .A2(regs[946]), .B1(n28), .B2(regs[434]), .ZN(
        n1063) );
  AOI22_X1 U1631 ( .A1(n127), .A2(regs[2482]), .B1(n69), .B2(regs[1970]), .ZN(
        n1062) );
  NAND3_X1 U1632 ( .A1(n1064), .A2(n1063), .A3(n1062), .ZN(curr_proc_regs[434]) );
  NAND2_X1 U1633 ( .A1(regs[947]), .A2(n2), .ZN(n1067) );
  AOI22_X1 U1634 ( .A1(n96), .A2(regs[1459]), .B1(n45), .B2(regs[435]), .ZN(
        n1066) );
  AOI22_X1 U1635 ( .A1(n127), .A2(regs[2483]), .B1(n17), .B2(regs[1971]), .ZN(
        n1065) );
  NAND3_X1 U1636 ( .A1(n1067), .A2(n1066), .A3(n1065), .ZN(curr_proc_regs[435]) );
  NAND2_X1 U1637 ( .A1(regs[948]), .A2(n2), .ZN(n1070) );
  AOI22_X1 U1638 ( .A1(n96), .A2(regs[1460]), .B1(n44), .B2(regs[436]), .ZN(
        n1069) );
  AOI22_X1 U1639 ( .A1(n127), .A2(regs[2484]), .B1(n73), .B2(regs[1972]), .ZN(
        n1068) );
  NAND3_X1 U1640 ( .A1(n1070), .A2(n1069), .A3(n1068), .ZN(curr_proc_regs[436]) );
  NAND2_X1 U1641 ( .A1(regs[1461]), .A2(n84), .ZN(n1073) );
  AOI22_X1 U1642 ( .A1(n10), .A2(regs[949]), .B1(n26), .B2(regs[437]), .ZN(
        n1072) );
  AOI22_X1 U1643 ( .A1(n127), .A2(regs[2485]), .B1(n77), .B2(regs[1973]), .ZN(
        n1071) );
  NAND3_X1 U1644 ( .A1(n1073), .A2(n1072), .A3(n1071), .ZN(curr_proc_regs[437]) );
  NAND2_X1 U1645 ( .A1(regs[1462]), .A2(n92), .ZN(n1076) );
  AOI22_X1 U1646 ( .A1(n49), .A2(regs[950]), .B1(n26), .B2(regs[438]), .ZN(
        n1075) );
  AOI22_X1 U1647 ( .A1(n127), .A2(regs[2486]), .B1(n67), .B2(regs[1974]), .ZN(
        n1074) );
  NAND3_X1 U1648 ( .A1(n1076), .A2(n1075), .A3(n1074), .ZN(curr_proc_regs[438]) );
  NAND2_X1 U1649 ( .A1(regs[951]), .A2(n13), .ZN(n1079) );
  AOI22_X1 U1650 ( .A1(n82), .A2(regs[1463]), .B1(n37), .B2(regs[439]), .ZN(
        n1078) );
  AOI22_X1 U1651 ( .A1(n127), .A2(regs[2487]), .B1(n77), .B2(regs[1975]), .ZN(
        n1077) );
  NAND3_X1 U1652 ( .A1(n1079), .A2(n1078), .A3(n1077), .ZN(curr_proc_regs[439]) );
  INV_X1 U1653 ( .A(regs[1067]), .ZN(n1450) );
  AOI22_X1 U1654 ( .A1(n126), .A2(regs[2091]), .B1(n9), .B2(regs[1579]), .ZN(
        n1081) );
  AOI22_X1 U1655 ( .A1(n54), .A2(regs[555]), .B1(n45), .B2(regs[43]), .ZN(
        n1080) );
  OAI211_X1 U1656 ( .C1(n5), .C2(n1450), .A(n1081), .B(n1080), .ZN(
        curr_proc_regs[43]) );
  NAND2_X1 U1657 ( .A1(regs[952]), .A2(n13), .ZN(n1084) );
  AOI22_X1 U1658 ( .A1(n98), .A2(regs[1464]), .B1(n29), .B2(regs[440]), .ZN(
        n1083) );
  AOI22_X1 U1659 ( .A1(n126), .A2(regs[2488]), .B1(n77), .B2(regs[1976]), .ZN(
        n1082) );
  NAND3_X1 U1660 ( .A1(n1084), .A2(n1083), .A3(n1082), .ZN(curr_proc_regs[440]) );
  NAND2_X1 U1661 ( .A1(regs[1465]), .A2(n93), .ZN(n1087) );
  AOI22_X1 U1662 ( .A1(n55), .A2(regs[953]), .B1(n33), .B2(regs[441]), .ZN(
        n1086) );
  AOI22_X1 U1663 ( .A1(n126), .A2(regs[2489]), .B1(n67), .B2(regs[1977]), .ZN(
        n1085) );
  NAND3_X1 U1664 ( .A1(n1087), .A2(n1086), .A3(n1085), .ZN(curr_proc_regs[441]) );
  NAND2_X1 U1665 ( .A1(regs[954]), .A2(n13), .ZN(n1090) );
  AOI22_X1 U1666 ( .A1(n80), .A2(regs[1466]), .B1(n36), .B2(regs[442]), .ZN(
        n1089) );
  AOI22_X1 U1667 ( .A1(n126), .A2(regs[2490]), .B1(n77), .B2(regs[1978]), .ZN(
        n1088) );
  NAND3_X1 U1668 ( .A1(n1090), .A2(n1089), .A3(n1088), .ZN(curr_proc_regs[442]) );
  NAND2_X1 U1669 ( .A1(regs[955]), .A2(n13), .ZN(n1093) );
  AOI22_X1 U1670 ( .A1(n80), .A2(regs[1467]), .B1(n33), .B2(regs[443]), .ZN(
        n1092) );
  AOI22_X1 U1671 ( .A1(n126), .A2(regs[2491]), .B1(n9), .B2(regs[1979]), .ZN(
        n1091) );
  NAND3_X1 U1672 ( .A1(n1093), .A2(n1092), .A3(n1091), .ZN(curr_proc_regs[443]) );
  NAND2_X1 U1673 ( .A1(regs[956]), .A2(n13), .ZN(n1096) );
  AOI22_X1 U1674 ( .A1(n80), .A2(regs[1468]), .B1(n35), .B2(regs[444]), .ZN(
        n1095) );
  AOI22_X1 U1675 ( .A1(n130), .A2(regs[2492]), .B1(n77), .B2(regs[1980]), .ZN(
        n1094) );
  NAND3_X1 U1676 ( .A1(n1096), .A2(n1095), .A3(n1094), .ZN(curr_proc_regs[444]) );
  NAND2_X1 U1677 ( .A1(regs[957]), .A2(n13), .ZN(n1099) );
  AOI22_X1 U1678 ( .A1(n80), .A2(regs[1469]), .B1(n40), .B2(regs[445]), .ZN(
        n1098) );
  AOI22_X1 U1679 ( .A1(n111), .A2(regs[2493]), .B1(n67), .B2(regs[1981]), .ZN(
        n1097) );
  NAND3_X1 U1680 ( .A1(n1099), .A2(n1098), .A3(n1097), .ZN(curr_proc_regs[445]) );
  NAND2_X1 U1681 ( .A1(regs[1470]), .A2(n88), .ZN(n1102) );
  AOI22_X1 U1682 ( .A1(n55), .A2(regs[958]), .B1(n42), .B2(regs[446]), .ZN(
        n1101) );
  AOI22_X1 U1683 ( .A1(n111), .A2(regs[2494]), .B1(n77), .B2(regs[1982]), .ZN(
        n1100) );
  NAND3_X1 U1684 ( .A1(n1102), .A2(n1101), .A3(n1100), .ZN(curr_proc_regs[446]) );
  NAND2_X1 U1685 ( .A1(regs[959]), .A2(n13), .ZN(n1105) );
  AOI22_X1 U1686 ( .A1(n80), .A2(regs[1471]), .B1(n35), .B2(regs[447]), .ZN(
        n1104) );
  AOI22_X1 U1687 ( .A1(n111), .A2(regs[2495]), .B1(n67), .B2(regs[1983]), .ZN(
        n1103) );
  NAND3_X1 U1688 ( .A1(n1105), .A2(n1104), .A3(n1103), .ZN(curr_proc_regs[447]) );
  NAND2_X1 U1689 ( .A1(regs[960]), .A2(n13), .ZN(n1108) );
  AOI22_X1 U1690 ( .A1(n80), .A2(regs[1472]), .B1(n40), .B2(regs[448]), .ZN(
        n1107) );
  AOI22_X1 U1691 ( .A1(n111), .A2(regs[2496]), .B1(n77), .B2(regs[1984]), .ZN(
        n1106) );
  NAND3_X1 U1692 ( .A1(n1108), .A2(n1107), .A3(n1106), .ZN(curr_proc_regs[448]) );
  NAND2_X1 U1693 ( .A1(regs[961]), .A2(n61), .ZN(n1111) );
  AOI22_X1 U1694 ( .A1(n80), .A2(regs[1473]), .B1(n42), .B2(regs[449]), .ZN(
        n1110) );
  AOI22_X1 U1695 ( .A1(n111), .A2(regs[2497]), .B1(n9), .B2(regs[1985]), .ZN(
        n1109) );
  NAND3_X1 U1696 ( .A1(n1111), .A2(n1110), .A3(n1109), .ZN(curr_proc_regs[449]) );
  INV_X1 U1697 ( .A(regs[556]), .ZN(n1453) );
  AOI22_X1 U1698 ( .A1(n111), .A2(regs[2092]), .B1(n9), .B2(regs[1580]), .ZN(
        n1113) );
  AOI22_X1 U1699 ( .A1(n80), .A2(regs[1068]), .B1(n31), .B2(regs[44]), .ZN(
        n1112) );
  OAI211_X1 U1700 ( .C1(n11), .C2(n1453), .A(n1113), .B(n1112), .ZN(
        curr_proc_regs[44]) );
  NAND2_X1 U1701 ( .A1(regs[962]), .A2(n13), .ZN(n1116) );
  AOI22_X1 U1702 ( .A1(n80), .A2(regs[1474]), .B1(n27), .B2(regs[450]), .ZN(
        n1115) );
  AOI22_X1 U1703 ( .A1(n111), .A2(regs[2498]), .B1(n77), .B2(regs[1986]), .ZN(
        n1114) );
  NAND3_X1 U1704 ( .A1(n1116), .A2(n1115), .A3(n1114), .ZN(curr_proc_regs[450]) );
  NAND2_X1 U1705 ( .A1(regs[1475]), .A2(n93), .ZN(n1119) );
  AOI22_X1 U1706 ( .A1(n55), .A2(regs[963]), .B1(n26), .B2(regs[451]), .ZN(
        n1118) );
  AOI22_X1 U1707 ( .A1(n110), .A2(regs[2499]), .B1(n67), .B2(regs[1987]), .ZN(
        n1117) );
  NAND3_X1 U1708 ( .A1(n1119), .A2(n1118), .A3(n1117), .ZN(curr_proc_regs[451]) );
  NAND2_X1 U1709 ( .A1(regs[1476]), .A2(n92), .ZN(n1122) );
  AOI22_X1 U1710 ( .A1(n55), .A2(regs[964]), .B1(n27), .B2(regs[452]), .ZN(
        n1121) );
  AOI22_X1 U1711 ( .A1(n110), .A2(regs[2500]), .B1(n77), .B2(regs[1988]), .ZN(
        n1120) );
  NAND3_X1 U1712 ( .A1(n1122), .A2(n1121), .A3(n1120), .ZN(curr_proc_regs[452]) );
  NAND2_X1 U1713 ( .A1(regs[1477]), .A2(n92), .ZN(n1125) );
  AOI22_X1 U1714 ( .A1(n55), .A2(regs[965]), .B1(n38), .B2(regs[453]), .ZN(
        n1124) );
  AOI22_X1 U1715 ( .A1(n110), .A2(regs[2501]), .B1(n77), .B2(regs[1989]), .ZN(
        n1123) );
  NAND3_X1 U1716 ( .A1(n1125), .A2(n1124), .A3(n1123), .ZN(curr_proc_regs[453]) );
  NAND2_X1 U1717 ( .A1(regs[1478]), .A2(n93), .ZN(n1128) );
  AOI22_X1 U1718 ( .A1(n55), .A2(regs[966]), .B1(n45), .B2(regs[454]), .ZN(
        n1127) );
  AOI22_X1 U1719 ( .A1(n110), .A2(regs[2502]), .B1(n9), .B2(regs[1990]), .ZN(
        n1126) );
  NAND3_X1 U1720 ( .A1(n1128), .A2(n1127), .A3(n1126), .ZN(curr_proc_regs[454]) );
  NAND2_X1 U1721 ( .A1(regs[967]), .A2(n13), .ZN(n1131) );
  AOI22_X1 U1722 ( .A1(n80), .A2(regs[1479]), .B1(n44), .B2(regs[455]), .ZN(
        n1130) );
  AOI22_X1 U1723 ( .A1(n110), .A2(regs[2503]), .B1(n77), .B2(regs[1991]), .ZN(
        n1129) );
  NAND3_X1 U1724 ( .A1(n1131), .A2(n1130), .A3(n1129), .ZN(curr_proc_regs[455]) );
  NAND2_X1 U1725 ( .A1(regs[968]), .A2(n59), .ZN(n1134) );
  AOI22_X1 U1726 ( .A1(n80), .A2(regs[1480]), .B1(n27), .B2(regs[456]), .ZN(
        n1133) );
  AOI22_X1 U1727 ( .A1(n110), .A2(regs[2504]), .B1(n67), .B2(regs[1992]), .ZN(
        n1132) );
  NAND3_X1 U1728 ( .A1(n1134), .A2(n1133), .A3(n1132), .ZN(curr_proc_regs[456]) );
  NAND2_X1 U1729 ( .A1(regs[1481]), .A2(n80), .ZN(n1137) );
  AOI22_X1 U1730 ( .A1(n55), .A2(regs[969]), .B1(n3), .B2(regs[457]), .ZN(
        n1136) );
  AOI22_X1 U1731 ( .A1(n110), .A2(regs[2505]), .B1(n77), .B2(regs[1993]), .ZN(
        n1135) );
  NAND3_X1 U1732 ( .A1(n1137), .A2(n1136), .A3(n1135), .ZN(curr_proc_regs[457]) );
  NAND2_X1 U1733 ( .A1(regs[1482]), .A2(n79), .ZN(n1140) );
  AOI22_X1 U1734 ( .A1(n55), .A2(regs[970]), .B1(n12), .B2(regs[458]), .ZN(
        n1139) );
  AOI22_X1 U1735 ( .A1(n110), .A2(regs[2506]), .B1(n77), .B2(regs[1994]), .ZN(
        n1138) );
  NAND3_X1 U1736 ( .A1(n1140), .A2(n1139), .A3(n1138), .ZN(curr_proc_regs[458]) );
  NAND2_X1 U1737 ( .A1(regs[1483]), .A2(n78), .ZN(n1143) );
  AOI22_X1 U1738 ( .A1(n55), .A2(regs[971]), .B1(n12), .B2(regs[459]), .ZN(
        n1142) );
  AOI22_X1 U1739 ( .A1(n110), .A2(regs[2507]), .B1(n77), .B2(regs[1995]), .ZN(
        n1141) );
  NAND3_X1 U1740 ( .A1(n1143), .A2(n1142), .A3(n1141), .ZN(curr_proc_regs[459]) );
  INV_X1 U1741 ( .A(regs[557]), .ZN(n1456) );
  AOI22_X1 U1742 ( .A1(n110), .A2(regs[2093]), .B1(n77), .B2(regs[1581]), .ZN(
        n1145) );
  AOI22_X1 U1743 ( .A1(n79), .A2(regs[1069]), .B1(n28), .B2(regs[45]), .ZN(
        n1144) );
  OAI211_X1 U1744 ( .C1(n11), .C2(n1456), .A(n1145), .B(n1144), .ZN(
        curr_proc_regs[45]) );
  NAND2_X1 U1745 ( .A1(regs[1484]), .A2(n83), .ZN(n1148) );
  AOI22_X1 U1746 ( .A1(n55), .A2(regs[972]), .B1(n40), .B2(regs[460]), .ZN(
        n1147) );
  AOI22_X1 U1747 ( .A1(n110), .A2(regs[2508]), .B1(n77), .B2(regs[1996]), .ZN(
        n1146) );
  NAND3_X1 U1748 ( .A1(n1148), .A2(n1147), .A3(n1146), .ZN(curr_proc_regs[460]) );
  NAND2_X1 U1749 ( .A1(regs[973]), .A2(n13), .ZN(n1151) );
  AOI22_X1 U1750 ( .A1(n79), .A2(regs[1485]), .B1(n42), .B2(regs[461]), .ZN(
        n1150) );
  AOI22_X1 U1751 ( .A1(n107), .A2(regs[2509]), .B1(n77), .B2(regs[1997]), .ZN(
        n1149) );
  NAND3_X1 U1752 ( .A1(n1151), .A2(n1150), .A3(n1149), .ZN(curr_proc_regs[461]) );
  NAND2_X1 U1753 ( .A1(regs[974]), .A2(n61), .ZN(n1154) );
  AOI22_X1 U1754 ( .A1(n79), .A2(regs[1486]), .B1(n31), .B2(regs[462]), .ZN(
        n1153) );
  AOI22_X1 U1755 ( .A1(n108), .A2(regs[2510]), .B1(n77), .B2(regs[1998]), .ZN(
        n1152) );
  NAND3_X1 U1756 ( .A1(n1154), .A2(n1153), .A3(n1152), .ZN(curr_proc_regs[462]) );
  NAND2_X1 U1757 ( .A1(regs[975]), .A2(n61), .ZN(n1157) );
  AOI22_X1 U1758 ( .A1(n79), .A2(regs[1487]), .B1(n30), .B2(regs[463]), .ZN(
        n1156) );
  AOI22_X1 U1759 ( .A1(n109), .A2(regs[2511]), .B1(n77), .B2(regs[1999]), .ZN(
        n1155) );
  NAND3_X1 U1760 ( .A1(n1157), .A2(n1156), .A3(n1155), .ZN(curr_proc_regs[463]) );
  NAND2_X1 U1761 ( .A1(regs[1488]), .A2(n94), .ZN(n1160) );
  AOI22_X1 U1762 ( .A1(n49), .A2(regs[976]), .B1(n29), .B2(regs[464]), .ZN(
        n1159) );
  AOI22_X1 U1763 ( .A1(n109), .A2(regs[2512]), .B1(n77), .B2(regs[2000]), .ZN(
        n1158) );
  NAND3_X1 U1764 ( .A1(n1160), .A2(n1159), .A3(n1158), .ZN(curr_proc_regs[464]) );
  NAND2_X1 U1765 ( .A1(regs[977]), .A2(n61), .ZN(n1163) );
  AOI22_X1 U1766 ( .A1(n79), .A2(regs[1489]), .B1(n36), .B2(regs[465]), .ZN(
        n1162) );
  AOI22_X1 U1767 ( .A1(n108), .A2(regs[2513]), .B1(n77), .B2(regs[2001]), .ZN(
        n1161) );
  NAND3_X1 U1768 ( .A1(n1163), .A2(n1162), .A3(n1161), .ZN(curr_proc_regs[465]) );
  NAND2_X1 U1769 ( .A1(regs[1490]), .A2(n94), .ZN(n1166) );
  AOI22_X1 U1770 ( .A1(n56), .A2(regs[978]), .B1(n33), .B2(regs[466]), .ZN(
        n1165) );
  AOI22_X1 U1771 ( .A1(n107), .A2(regs[2514]), .B1(n77), .B2(regs[2002]), .ZN(
        n1164) );
  NAND3_X1 U1772 ( .A1(n1166), .A2(n1165), .A3(n1164), .ZN(curr_proc_regs[466]) );
  NAND2_X1 U1773 ( .A1(regs[979]), .A2(n61), .ZN(n1169) );
  AOI22_X1 U1774 ( .A1(n79), .A2(regs[1491]), .B1(n40), .B2(regs[467]), .ZN(
        n1168) );
  AOI22_X1 U1775 ( .A1(n108), .A2(regs[2515]), .B1(n77), .B2(regs[2003]), .ZN(
        n1167) );
  NAND3_X1 U1776 ( .A1(n1169), .A2(n1168), .A3(n1167), .ZN(curr_proc_regs[467]) );
  NAND2_X1 U1777 ( .A1(regs[1492]), .A2(n94), .ZN(n1172) );
  AOI22_X1 U1778 ( .A1(n10), .A2(regs[980]), .B1(n40), .B2(regs[468]), .ZN(
        n1171) );
  AOI22_X1 U1779 ( .A1(n109), .A2(regs[2516]), .B1(n77), .B2(regs[2004]), .ZN(
        n1170) );
  NAND3_X1 U1780 ( .A1(n1172), .A2(n1171), .A3(n1170), .ZN(curr_proc_regs[468]) );
  NAND2_X1 U1781 ( .A1(regs[981]), .A2(n2), .ZN(n1175) );
  AOI22_X1 U1782 ( .A1(n79), .A2(regs[1493]), .B1(n40), .B2(regs[469]), .ZN(
        n1174) );
  AOI22_X1 U1783 ( .A1(n107), .A2(regs[2517]), .B1(n67), .B2(regs[2005]), .ZN(
        n1173) );
  NAND3_X1 U1784 ( .A1(n1175), .A2(n1174), .A3(n1173), .ZN(curr_proc_regs[469]) );
  INV_X1 U1785 ( .A(regs[558]), .ZN(n1459) );
  AOI22_X1 U1786 ( .A1(n109), .A2(regs[2094]), .B1(n77), .B2(regs[1582]), .ZN(
        n1177) );
  AOI22_X1 U1787 ( .A1(n79), .A2(regs[1070]), .B1(n40), .B2(regs[46]), .ZN(
        n1176) );
  OAI211_X1 U1788 ( .C1(n65), .C2(n1459), .A(n1177), .B(n1176), .ZN(
        curr_proc_regs[46]) );
  NAND2_X1 U1789 ( .A1(regs[982]), .A2(n59), .ZN(n1180) );
  AOI22_X1 U1790 ( .A1(n79), .A2(regs[1494]), .B1(n28), .B2(regs[470]), .ZN(
        n1179) );
  AOI22_X1 U1791 ( .A1(n107), .A2(regs[2518]), .B1(n67), .B2(regs[2006]), .ZN(
        n1178) );
  NAND3_X1 U1792 ( .A1(n1180), .A2(n1179), .A3(n1178), .ZN(curr_proc_regs[470]) );
  NAND2_X1 U1793 ( .A1(regs[1495]), .A2(n94), .ZN(n1183) );
  AOI22_X1 U1794 ( .A1(n49), .A2(regs[983]), .B1(n28), .B2(regs[471]), .ZN(
        n1182) );
  AOI22_X1 U1795 ( .A1(n108), .A2(regs[2519]), .B1(n9), .B2(regs[2007]), .ZN(
        n1181) );
  NAND3_X1 U1796 ( .A1(n1183), .A2(n1182), .A3(n1181), .ZN(curr_proc_regs[471]) );
  NAND2_X1 U1797 ( .A1(regs[1496]), .A2(n94), .ZN(n1186) );
  AOI22_X1 U1798 ( .A1(n10), .A2(regs[984]), .B1(n34), .B2(regs[472]), .ZN(
        n1185) );
  AOI22_X1 U1799 ( .A1(n107), .A2(regs[2520]), .B1(n77), .B2(regs[2008]), .ZN(
        n1184) );
  NAND3_X1 U1800 ( .A1(n1186), .A2(n1185), .A3(n1184), .ZN(curr_proc_regs[472]) );
  NAND2_X1 U1801 ( .A1(regs[985]), .A2(n13), .ZN(n1189) );
  AOI22_X1 U1802 ( .A1(n79), .A2(regs[1497]), .B1(n32), .B2(regs[473]), .ZN(
        n1188) );
  AOI22_X1 U1803 ( .A1(n108), .A2(regs[2521]), .B1(n77), .B2(regs[2009]), .ZN(
        n1187) );
  NAND3_X1 U1804 ( .A1(n1189), .A2(n1188), .A3(n1187), .ZN(curr_proc_regs[473]) );
  NAND2_X1 U1805 ( .A1(regs[986]), .A2(n13), .ZN(n1192) );
  AOI22_X1 U1806 ( .A1(n79), .A2(regs[1498]), .B1(n41), .B2(regs[474]), .ZN(
        n1191) );
  AOI22_X1 U1807 ( .A1(n109), .A2(regs[2522]), .B1(n67), .B2(regs[2010]), .ZN(
        n1190) );
  NAND3_X1 U1808 ( .A1(n1192), .A2(n1191), .A3(n1190), .ZN(curr_proc_regs[474]) );
  NAND2_X1 U1809 ( .A1(regs[1499]), .A2(n95), .ZN(n1195) );
  AOI22_X1 U1810 ( .A1(n49), .A2(regs[987]), .B1(n43), .B2(regs[475]), .ZN(
        n1194) );
  AOI22_X1 U1811 ( .A1(n109), .A2(regs[2523]), .B1(n77), .B2(regs[2011]), .ZN(
        n1193) );
  NAND3_X1 U1812 ( .A1(n1195), .A2(n1194), .A3(n1193), .ZN(curr_proc_regs[475]) );
  NAND2_X1 U1813 ( .A1(regs[1500]), .A2(n95), .ZN(n1198) );
  AOI22_X1 U1814 ( .A1(n10), .A2(regs[988]), .B1(n3), .B2(regs[476]), .ZN(
        n1197) );
  AOI22_X1 U1815 ( .A1(n107), .A2(regs[2524]), .B1(n9), .B2(regs[2012]), .ZN(
        n1196) );
  NAND3_X1 U1816 ( .A1(n1198), .A2(n1197), .A3(n1196), .ZN(curr_proc_regs[476]) );
  NAND2_X1 U1817 ( .A1(regs[989]), .A2(n60), .ZN(n1201) );
  AOI22_X1 U1818 ( .A1(n79), .A2(regs[1501]), .B1(n41), .B2(regs[477]), .ZN(
        n1200) );
  AOI22_X1 U1819 ( .A1(n108), .A2(regs[2525]), .B1(n9), .B2(regs[2013]), .ZN(
        n1199) );
  NAND3_X1 U1820 ( .A1(n1201), .A2(n1200), .A3(n1199), .ZN(curr_proc_regs[477]) );
  NAND2_X1 U1821 ( .A1(regs[990]), .A2(n61), .ZN(n1204) );
  AOI22_X1 U1822 ( .A1(n80), .A2(regs[1502]), .B1(n41), .B2(regs[478]), .ZN(
        n1203) );
  AOI22_X1 U1823 ( .A1(n109), .A2(regs[2526]), .B1(n77), .B2(regs[2014]), .ZN(
        n1202) );
  NAND3_X1 U1824 ( .A1(n1204), .A2(n1203), .A3(n1202), .ZN(curr_proc_regs[478]) );
  NAND2_X1 U1825 ( .A1(regs[991]), .A2(n2), .ZN(n1207) );
  AOI22_X1 U1826 ( .A1(n87), .A2(regs[1503]), .B1(n41), .B2(regs[479]), .ZN(
        n1206) );
  AOI22_X1 U1827 ( .A1(n107), .A2(regs[2527]), .B1(n67), .B2(regs[2015]), .ZN(
        n1205) );
  NAND3_X1 U1828 ( .A1(n1207), .A2(n1206), .A3(n1205), .ZN(curr_proc_regs[479]) );
  INV_X1 U1829 ( .A(regs[559]), .ZN(n1462) );
  AOI22_X1 U1830 ( .A1(n107), .A2(regs[2095]), .B1(n77), .B2(regs[1583]), .ZN(
        n1209) );
  AOI22_X1 U1831 ( .A1(n87), .A2(regs[1071]), .B1(n41), .B2(regs[47]), .ZN(
        n1208) );
  OAI211_X1 U1832 ( .C1(n65), .C2(n1462), .A(n1209), .B(n1208), .ZN(
        curr_proc_regs[47]) );
  NAND2_X1 U1833 ( .A1(regs[992]), .A2(n61), .ZN(n1212) );
  AOI22_X1 U1834 ( .A1(n85), .A2(regs[1504]), .B1(n40), .B2(regs[480]), .ZN(
        n1211) );
  AOI22_X1 U1835 ( .A1(n108), .A2(regs[2528]), .B1(n77), .B2(regs[2016]), .ZN(
        n1210) );
  NAND3_X1 U1836 ( .A1(n1212), .A2(n1211), .A3(n1210), .ZN(curr_proc_regs[480]) );
  NAND2_X1 U1837 ( .A1(regs[1505]), .A2(n95), .ZN(n1215) );
  AOI22_X1 U1838 ( .A1(n56), .A2(regs[993]), .B1(n40), .B2(regs[481]), .ZN(
        n1214) );
  AOI22_X1 U1839 ( .A1(n108), .A2(regs[2529]), .B1(n9), .B2(regs[2017]), .ZN(
        n1213) );
  NAND3_X1 U1840 ( .A1(n1215), .A2(n1214), .A3(n1213), .ZN(curr_proc_regs[481]) );
  NAND2_X1 U1841 ( .A1(regs[1506]), .A2(n95), .ZN(n1218) );
  AOI22_X1 U1842 ( .A1(n10), .A2(regs[994]), .B1(n40), .B2(regs[482]), .ZN(
        n1217) );
  AOI22_X1 U1843 ( .A1(n109), .A2(regs[2530]), .B1(n77), .B2(regs[2018]), .ZN(
        n1216) );
  NAND3_X1 U1844 ( .A1(n1218), .A2(n1217), .A3(n1216), .ZN(curr_proc_regs[482]) );
  NAND2_X1 U1845 ( .A1(regs[995]), .A2(n62), .ZN(n1221) );
  AOI22_X1 U1846 ( .A1(n94), .A2(regs[1507]), .B1(n40), .B2(regs[483]), .ZN(
        n1220) );
  AOI22_X1 U1847 ( .A1(n107), .A2(regs[2531]), .B1(n9), .B2(regs[2019]), .ZN(
        n1219) );
  NAND3_X1 U1848 ( .A1(n1221), .A2(n1220), .A3(n1219), .ZN(curr_proc_regs[483]) );
  NAND2_X1 U1849 ( .A1(regs[996]), .A2(n8), .ZN(n1224) );
  AOI22_X1 U1850 ( .A1(n98), .A2(regs[1508]), .B1(n40), .B2(regs[484]), .ZN(
        n1223) );
  AOI22_X1 U1851 ( .A1(n108), .A2(regs[2532]), .B1(n77), .B2(regs[2020]), .ZN(
        n1222) );
  NAND3_X1 U1852 ( .A1(n1224), .A2(n1223), .A3(n1222), .ZN(curr_proc_regs[484]) );
  NAND2_X1 U1853 ( .A1(regs[997]), .A2(n8), .ZN(n1227) );
  AOI22_X1 U1854 ( .A1(n95), .A2(regs[1509]), .B1(n40), .B2(regs[485]), .ZN(
        n1226) );
  AOI22_X1 U1855 ( .A1(n109), .A2(regs[2533]), .B1(n77), .B2(regs[2021]), .ZN(
        n1225) );
  NAND3_X1 U1856 ( .A1(n1227), .A2(n1226), .A3(n1225), .ZN(curr_proc_regs[485]) );
  NAND2_X1 U1857 ( .A1(regs[998]), .A2(n8), .ZN(n1230) );
  AOI22_X1 U1858 ( .A1(n78), .A2(regs[1510]), .B1(n40), .B2(regs[486]), .ZN(
        n1229) );
  AOI22_X1 U1859 ( .A1(n107), .A2(regs[2534]), .B1(n77), .B2(regs[2022]), .ZN(
        n1228) );
  NAND3_X1 U1860 ( .A1(n1230), .A2(n1229), .A3(n1228), .ZN(curr_proc_regs[486]) );
  NAND2_X1 U1861 ( .A1(regs[1511]), .A2(n96), .ZN(n1233) );
  AOI22_X1 U1862 ( .A1(n49), .A2(regs[999]), .B1(n27), .B2(regs[487]), .ZN(
        n1232) );
  AOI22_X1 U1863 ( .A1(n108), .A2(regs[2535]), .B1(n67), .B2(regs[2023]), .ZN(
        n1231) );
  NAND3_X1 U1864 ( .A1(n1233), .A2(n1232), .A3(n1231), .ZN(curr_proc_regs[487]) );
  NAND2_X1 U1865 ( .A1(regs[1000]), .A2(n8), .ZN(n1236) );
  AOI22_X1 U1866 ( .A1(n86), .A2(regs[1512]), .B1(n45), .B2(regs[488]), .ZN(
        n1235) );
  AOI22_X1 U1867 ( .A1(n109), .A2(regs[2536]), .B1(n77), .B2(regs[2024]), .ZN(
        n1234) );
  NAND3_X1 U1868 ( .A1(n1236), .A2(n1235), .A3(n1234), .ZN(curr_proc_regs[488]) );
  NAND2_X1 U1869 ( .A1(regs[1513]), .A2(n96), .ZN(n1239) );
  AOI22_X1 U1870 ( .A1(n10), .A2(regs[1001]), .B1(n45), .B2(regs[489]), .ZN(
        n1238) );
  AOI22_X1 U1871 ( .A1(n107), .A2(regs[2537]), .B1(n77), .B2(regs[2025]), .ZN(
        n1237) );
  NAND3_X1 U1872 ( .A1(n1239), .A2(n1238), .A3(n1237), .ZN(curr_proc_regs[489]) );
  INV_X1 U1873 ( .A(regs[560]), .ZN(n1467) );
  AOI22_X1 U1874 ( .A1(n108), .A2(regs[2096]), .B1(n77), .B2(regs[1584]), .ZN(
        n1241) );
  AOI22_X1 U1875 ( .A1(n78), .A2(regs[1072]), .B1(n45), .B2(regs[48]), .ZN(
        n1240) );
  OAI211_X1 U1876 ( .C1(n65), .C2(n1467), .A(n1241), .B(n1240), .ZN(
        curr_proc_regs[48]) );
  NAND2_X1 U1877 ( .A1(regs[1002]), .A2(n8), .ZN(n1244) );
  AOI22_X1 U1878 ( .A1(n78), .A2(regs[1514]), .B1(n41), .B2(regs[490]), .ZN(
        n1243) );
  AOI22_X1 U1879 ( .A1(n109), .A2(regs[2538]), .B1(n77), .B2(regs[2026]), .ZN(
        n1242) );
  NAND3_X1 U1880 ( .A1(n1244), .A2(n1243), .A3(n1242), .ZN(curr_proc_regs[490]) );
  NAND2_X1 U1881 ( .A1(regs[1003]), .A2(n8), .ZN(n1247) );
  AOI22_X1 U1882 ( .A1(n78), .A2(regs[1515]), .B1(n41), .B2(regs[491]), .ZN(
        n1246) );
  AOI22_X1 U1883 ( .A1(n109), .A2(regs[2539]), .B1(n77), .B2(regs[2027]), .ZN(
        n1245) );
  NAND3_X1 U1884 ( .A1(n1247), .A2(n1246), .A3(n1245), .ZN(curr_proc_regs[491]) );
  NAND2_X1 U1885 ( .A1(regs[1516]), .A2(n96), .ZN(n1250) );
  AOI22_X1 U1886 ( .A1(n55), .A2(regs[1004]), .B1(n41), .B2(regs[492]), .ZN(
        n1249) );
  AOI22_X1 U1887 ( .A1(n109), .A2(regs[2540]), .B1(n9), .B2(regs[2028]), .ZN(
        n1248) );
  NAND3_X1 U1888 ( .A1(n1250), .A2(n1249), .A3(n1248), .ZN(curr_proc_regs[492]) );
  NAND2_X1 U1889 ( .A1(regs[1517]), .A2(n96), .ZN(n1253) );
  AOI22_X1 U1890 ( .A1(n2), .A2(regs[1005]), .B1(n41), .B2(regs[493]), .ZN(
        n1252) );
  AOI22_X1 U1891 ( .A1(n109), .A2(regs[2541]), .B1(n77), .B2(regs[2029]), .ZN(
        n1251) );
  NAND3_X1 U1892 ( .A1(n1253), .A2(n1252), .A3(n1251), .ZN(curr_proc_regs[493]) );
  NAND2_X1 U1893 ( .A1(regs[1518]), .A2(n96), .ZN(n1256) );
  AOI22_X1 U1894 ( .A1(n61), .A2(regs[1006]), .B1(n41), .B2(regs[494]), .ZN(
        n1255) );
  AOI22_X1 U1895 ( .A1(n109), .A2(regs[2542]), .B1(n77), .B2(regs[2030]), .ZN(
        n1254) );
  NAND3_X1 U1896 ( .A1(n1256), .A2(n1255), .A3(n1254), .ZN(curr_proc_regs[494]) );
  NAND2_X1 U1897 ( .A1(regs[1519]), .A2(n82), .ZN(n1259) );
  AOI22_X1 U1898 ( .A1(n2), .A2(regs[1007]), .B1(n41), .B2(regs[495]), .ZN(
        n1258) );
  AOI22_X1 U1899 ( .A1(n109), .A2(regs[2543]), .B1(n77), .B2(regs[2031]), .ZN(
        n1257) );
  NAND3_X1 U1900 ( .A1(n1259), .A2(n1258), .A3(n1257), .ZN(curr_proc_regs[495]) );
  NAND2_X1 U1901 ( .A1(regs[1008]), .A2(n8), .ZN(n1262) );
  AOI22_X1 U1902 ( .A1(n78), .A2(regs[1520]), .B1(n41), .B2(regs[496]), .ZN(
        n1261) );
  AOI22_X1 U1903 ( .A1(n109), .A2(regs[2544]), .B1(n77), .B2(regs[2032]), .ZN(
        n1260) );
  NAND3_X1 U1904 ( .A1(n1262), .A2(n1261), .A3(n1260), .ZN(curr_proc_regs[496]) );
  NAND2_X1 U1905 ( .A1(regs[1009]), .A2(n8), .ZN(n1265) );
  AOI22_X1 U1906 ( .A1(n78), .A2(regs[1521]), .B1(n42), .B2(regs[497]), .ZN(
        n1264) );
  AOI22_X1 U1907 ( .A1(n109), .A2(regs[2545]), .B1(n71), .B2(regs[2033]), .ZN(
        n1263) );
  NAND3_X1 U1908 ( .A1(n1265), .A2(n1264), .A3(n1263), .ZN(curr_proc_regs[497]) );
  NAND2_X1 U1909 ( .A1(regs[1010]), .A2(n62), .ZN(n1268) );
  AOI22_X1 U1910 ( .A1(n78), .A2(regs[1522]), .B1(n42), .B2(regs[498]), .ZN(
        n1267) );
  AOI22_X1 U1911 ( .A1(n109), .A2(regs[2546]), .B1(n71), .B2(regs[2034]), .ZN(
        n1266) );
  NAND3_X1 U1912 ( .A1(n1268), .A2(n1267), .A3(n1266), .ZN(curr_proc_regs[498]) );
  NAND2_X1 U1913 ( .A1(regs[1523]), .A2(n95), .ZN(n1271) );
  AOI22_X1 U1914 ( .A1(n59), .A2(regs[1011]), .B1(n42), .B2(regs[499]), .ZN(
        n1270) );
  AOI22_X1 U1915 ( .A1(n109), .A2(regs[2547]), .B1(n71), .B2(regs[2035]), .ZN(
        n1269) );
  NAND3_X1 U1916 ( .A1(n1271), .A2(n1270), .A3(n1269), .ZN(curr_proc_regs[499]) );
  INV_X1 U1917 ( .A(regs[1073]), .ZN(n1470) );
  AOI22_X1 U1918 ( .A1(n109), .A2(regs[2097]), .B1(n71), .B2(regs[1585]), .ZN(
        n1273) );
  AOI22_X1 U1919 ( .A1(n60), .A2(regs[561]), .B1(n42), .B2(regs[49]), .ZN(
        n1272) );
  OAI211_X1 U1920 ( .C1(n2221), .C2(n1470), .A(n1273), .B(n1272), .ZN(
        curr_proc_regs[49]) );
  INV_X1 U1921 ( .A(regs[1028]), .ZN(n1328) );
  AOI22_X1 U1922 ( .A1(n109), .A2(regs[2052]), .B1(n71), .B2(regs[1540]), .ZN(
        n1275) );
  AOI22_X1 U1923 ( .A1(n61), .A2(regs[516]), .B1(n44), .B2(regs[4]), .ZN(n1274) );
  OAI211_X1 U1924 ( .C1(n99), .C2(n1328), .A(n1275), .B(n1274), .ZN(
        curr_proc_regs[4]) );
  NAND2_X1 U1925 ( .A1(regs[1012]), .A2(n8), .ZN(n1278) );
  AOI22_X1 U1926 ( .A1(n78), .A2(regs[1524]), .B1(n46), .B2(regs[500]), .ZN(
        n1277) );
  AOI22_X1 U1927 ( .A1(n108), .A2(regs[2548]), .B1(n71), .B2(regs[2036]), .ZN(
        n1276) );
  NAND3_X1 U1928 ( .A1(n1278), .A2(n1277), .A3(n1276), .ZN(curr_proc_regs[500]) );
  NAND2_X1 U1929 ( .A1(regs[1525]), .A2(n85), .ZN(n1281) );
  AOI22_X1 U1930 ( .A1(n2), .A2(regs[1013]), .B1(n26), .B2(regs[501]), .ZN(
        n1280) );
  AOI22_X1 U1931 ( .A1(n108), .A2(regs[2549]), .B1(n71), .B2(regs[2037]), .ZN(
        n1279) );
  NAND3_X1 U1932 ( .A1(n1281), .A2(n1280), .A3(n1279), .ZN(curr_proc_regs[501]) );
  NAND2_X1 U1933 ( .A1(regs[1526]), .A2(n80), .ZN(n1284) );
  AOI22_X1 U1934 ( .A1(n51), .A2(regs[1014]), .B1(n45), .B2(regs[502]), .ZN(
        n1283) );
  AOI22_X1 U1935 ( .A1(n108), .A2(regs[2550]), .B1(n71), .B2(regs[2038]), .ZN(
        n1282) );
  NAND3_X1 U1936 ( .A1(n1284), .A2(n1283), .A3(n1282), .ZN(curr_proc_regs[502]) );
  NAND2_X1 U1937 ( .A1(regs[1527]), .A2(n87), .ZN(n1287) );
  AOI22_X1 U1938 ( .A1(n51), .A2(regs[1015]), .B1(n44), .B2(regs[503]), .ZN(
        n1286) );
  AOI22_X1 U1939 ( .A1(n108), .A2(regs[2551]), .B1(n71), .B2(regs[2039]), .ZN(
        n1285) );
  NAND3_X1 U1940 ( .A1(n1287), .A2(n1286), .A3(n1285), .ZN(curr_proc_regs[503]) );
  NAND2_X1 U1941 ( .A1(regs[1528]), .A2(n19), .ZN(n1290) );
  AOI22_X1 U1942 ( .A1(n57), .A2(regs[1016]), .B1(n27), .B2(regs[504]), .ZN(
        n1289) );
  AOI22_X1 U1943 ( .A1(n108), .A2(regs[2552]), .B1(n71), .B2(regs[2040]), .ZN(
        n1288) );
  NAND3_X1 U1944 ( .A1(n1290), .A2(n1289), .A3(n1288), .ZN(curr_proc_regs[504]) );
  NAND2_X1 U1945 ( .A1(regs[1017]), .A2(n62), .ZN(n1293) );
  AOI22_X1 U1946 ( .A1(n78), .A2(regs[1529]), .B1(n26), .B2(regs[505]), .ZN(
        n1292) );
  AOI22_X1 U1947 ( .A1(n108), .A2(regs[2553]), .B1(n71), .B2(regs[2041]), .ZN(
        n1291) );
  NAND3_X1 U1948 ( .A1(n1293), .A2(n1292), .A3(n1291), .ZN(curr_proc_regs[505]) );
  NAND2_X1 U1949 ( .A1(regs[1018]), .A2(n62), .ZN(n1296) );
  AOI22_X1 U1950 ( .A1(n78), .A2(regs[1530]), .B1(n43), .B2(regs[506]), .ZN(
        n1295) );
  AOI22_X1 U1951 ( .A1(n108), .A2(regs[2554]), .B1(n71), .B2(regs[2042]), .ZN(
        n1294) );
  NAND3_X1 U1952 ( .A1(n1296), .A2(n1295), .A3(n1294), .ZN(curr_proc_regs[506]) );
  NAND2_X1 U1953 ( .A1(regs[1531]), .A2(n19), .ZN(n1299) );
  AOI22_X1 U1954 ( .A1(n13), .A2(regs[1019]), .B1(n43), .B2(regs[507]), .ZN(
        n1298) );
  AOI22_X1 U1955 ( .A1(n108), .A2(regs[2555]), .B1(n71), .B2(regs[2043]), .ZN(
        n1297) );
  NAND3_X1 U1956 ( .A1(n1299), .A2(n1298), .A3(n1297), .ZN(curr_proc_regs[507]) );
  NAND2_X1 U1957 ( .A1(regs[1020]), .A2(n62), .ZN(n1302) );
  AOI22_X1 U1958 ( .A1(n78), .A2(regs[1532]), .B1(n43), .B2(regs[508]), .ZN(
        n1301) );
  AOI22_X1 U1959 ( .A1(n108), .A2(regs[2556]), .B1(n71), .B2(regs[2044]), .ZN(
        n1300) );
  NAND3_X1 U1960 ( .A1(n1302), .A2(n1301), .A3(n1300), .ZN(curr_proc_regs[508]) );
  NAND2_X1 U1961 ( .A1(regs[1021]), .A2(n8), .ZN(n1305) );
  AOI22_X1 U1962 ( .A1(n78), .A2(regs[1533]), .B1(n43), .B2(regs[509]), .ZN(
        n1304) );
  AOI22_X1 U1963 ( .A1(n108), .A2(regs[2557]), .B1(n71), .B2(regs[2045]), .ZN(
        n1303) );
  NAND3_X1 U1964 ( .A1(n1305), .A2(n1304), .A3(n1303), .ZN(curr_proc_regs[509]) );
  INV_X1 U1965 ( .A(regs[562]), .ZN(n1473) );
  AOI22_X1 U1966 ( .A1(n108), .A2(regs[2098]), .B1(n71), .B2(regs[1586]), .ZN(
        n1307) );
  AOI22_X1 U1967 ( .A1(n94), .A2(regs[1074]), .B1(n42), .B2(regs[50]), .ZN(
        n1306) );
  OAI211_X1 U1968 ( .C1(n65), .C2(n1473), .A(n1307), .B(n1306), .ZN(
        curr_proc_regs[50]) );
  NAND2_X1 U1969 ( .A1(regs[1022]), .A2(n2), .ZN(n1310) );
  AOI22_X1 U1970 ( .A1(n96), .A2(regs[1534]), .B1(n42), .B2(regs[510]), .ZN(
        n1309) );
  AOI22_X1 U1971 ( .A1(n107), .A2(regs[2558]), .B1(n71), .B2(regs[2046]), .ZN(
        n1308) );
  NAND3_X1 U1972 ( .A1(n1310), .A2(n1309), .A3(n1308), .ZN(curr_proc_regs[510]) );
  NAND2_X1 U1973 ( .A1(regs[1535]), .A2(n19), .ZN(n1313) );
  AOI22_X1 U1974 ( .A1(n2), .A2(regs[1023]), .B1(n42), .B2(regs[511]), .ZN(
        n1312) );
  AOI22_X1 U1975 ( .A1(n107), .A2(regs[2559]), .B1(n71), .B2(regs[2047]), .ZN(
        n1311) );
  NAND3_X1 U1976 ( .A1(n1313), .A2(n1312), .A3(n1311), .ZN(curr_proc_regs[511]) );
  AOI22_X1 U1977 ( .A1(n107), .A2(regs[0]), .B1(n71), .B2(regs[2048]), .ZN(
        n1315) );
  AOI22_X1 U1978 ( .A1(n59), .A2(regs[1024]), .B1(n98), .B2(regs[1536]), .ZN(
        n1314) );
  OAI211_X1 U1979 ( .C1(n1316), .C2(n24), .A(n1315), .B(n1314), .ZN(
        curr_proc_regs[512]) );
  AOI22_X1 U1980 ( .A1(n107), .A2(regs[1]), .B1(n71), .B2(regs[2049]), .ZN(
        n1318) );
  AOI22_X1 U1981 ( .A1(n60), .A2(regs[1025]), .B1(n98), .B2(regs[1537]), .ZN(
        n1317) );
  OAI211_X1 U1982 ( .C1(n24), .C2(n1319), .A(n1318), .B(n1317), .ZN(
        curr_proc_regs[513]) );
  AOI22_X1 U1983 ( .A1(n107), .A2(regs[2]), .B1(n71), .B2(regs[2050]), .ZN(
        n1321) );
  AOI22_X1 U1984 ( .A1(n13), .A2(regs[1026]), .B1(n98), .B2(regs[1538]), .ZN(
        n1320) );
  OAI211_X1 U1985 ( .C1(n24), .C2(n1322), .A(n1321), .B(n1320), .ZN(
        curr_proc_regs[514]) );
  AOI22_X1 U1986 ( .A1(n107), .A2(regs[3]), .B1(n71), .B2(regs[2051]), .ZN(
        n1324) );
  AOI22_X1 U1987 ( .A1(n2), .A2(regs[1027]), .B1(n98), .B2(regs[1539]), .ZN(
        n1323) );
  OAI211_X1 U1988 ( .C1(n24), .C2(n1325), .A(n1324), .B(n1323), .ZN(
        curr_proc_regs[515]) );
  AOI22_X1 U1989 ( .A1(n107), .A2(regs[4]), .B1(n71), .B2(regs[2052]), .ZN(
        n1327) );
  AOI22_X1 U1990 ( .A1(n95), .A2(regs[1540]), .B1(n42), .B2(regs[516]), .ZN(
        n1326) );
  OAI211_X1 U1991 ( .C1(n65), .C2(n1328), .A(n1327), .B(n1326), .ZN(
        curr_proc_regs[516]) );
  INV_X1 U1992 ( .A(regs[1541]), .ZN(n1331) );
  AOI22_X1 U1993 ( .A1(n107), .A2(regs[5]), .B1(n71), .B2(regs[2053]), .ZN(
        n1330) );
  AOI22_X1 U1994 ( .A1(n13), .A2(regs[1029]), .B1(n42), .B2(regs[517]), .ZN(
        n1329) );
  OAI211_X1 U1995 ( .C1(n16), .C2(n1331), .A(n1330), .B(n1329), .ZN(
        curr_proc_regs[517]) );
  INV_X1 U1996 ( .A(regs[1030]), .ZN(n1914) );
  AOI22_X1 U1997 ( .A1(n107), .A2(regs[6]), .B1(n71), .B2(regs[2054]), .ZN(
        n1333) );
  AOI22_X1 U1998 ( .A1(n94), .A2(regs[1542]), .B1(n42), .B2(regs[518]), .ZN(
        n1332) );
  OAI211_X1 U1999 ( .C1(n63), .C2(n1914), .A(n1333), .B(n1332), .ZN(
        curr_proc_regs[518]) );
  INV_X1 U2000 ( .A(regs[1031]), .ZN(n2152) );
  AOI22_X1 U2001 ( .A1(n107), .A2(regs[7]), .B1(n71), .B2(regs[2055]), .ZN(
        n1335) );
  AOI22_X1 U2002 ( .A1(n78), .A2(regs[1543]), .B1(n42), .B2(regs[519]), .ZN(
        n1334) );
  OAI211_X1 U2003 ( .C1(n65), .C2(n2152), .A(n1335), .B(n1334), .ZN(
        curr_proc_regs[519]) );
  INV_X1 U2004 ( .A(regs[563]), .ZN(n1476) );
  AOI22_X1 U2005 ( .A1(n107), .A2(regs[2099]), .B1(n71), .B2(regs[1587]), .ZN(
        n1337) );
  AOI22_X1 U2006 ( .A1(n95), .A2(regs[1075]), .B1(n12), .B2(regs[51]), .ZN(
        n1336) );
  OAI211_X1 U2007 ( .C1(n65), .C2(n1476), .A(n1337), .B(n1336), .ZN(
        curr_proc_regs[51]) );
  INV_X1 U2008 ( .A(regs[1032]), .ZN(n2185) );
  AOI22_X1 U2009 ( .A1(n106), .A2(regs[8]), .B1(n71), .B2(regs[2056]), .ZN(
        n1339) );
  AOI22_X1 U2010 ( .A1(n81), .A2(regs[1544]), .B1(n28), .B2(regs[520]), .ZN(
        n1338) );
  OAI211_X1 U2011 ( .C1(n63), .C2(n2185), .A(n1339), .B(n1338), .ZN(
        curr_proc_regs[520]) );
  INV_X1 U2012 ( .A(regs[1545]), .ZN(n1342) );
  AOI22_X1 U2013 ( .A1(n104), .A2(regs[9]), .B1(n71), .B2(regs[2057]), .ZN(
        n1341) );
  AOI22_X1 U2014 ( .A1(n2), .A2(regs[1033]), .B1(n34), .B2(regs[521]), .ZN(
        n1340) );
  OAI211_X1 U2015 ( .C1(n100), .C2(n1342), .A(n1341), .B(n1340), .ZN(
        curr_proc_regs[521]) );
  AOI22_X1 U2016 ( .A1(n105), .A2(regs[10]), .B1(n71), .B2(regs[2058]), .ZN(
        n1344) );
  AOI22_X1 U2017 ( .A1(n13), .A2(regs[1034]), .B1(n98), .B2(regs[1546]), .ZN(
        n1343) );
  OAI211_X1 U2018 ( .C1(n24), .C2(n1345), .A(n1344), .B(n1343), .ZN(
        curr_proc_regs[522]) );
  AOI22_X1 U2019 ( .A1(n105), .A2(regs[11]), .B1(n71), .B2(regs[2059]), .ZN(
        n1347) );
  AOI22_X1 U2020 ( .A1(n13), .A2(regs[1035]), .B1(n98), .B2(regs[1547]), .ZN(
        n1346) );
  OAI211_X1 U2021 ( .C1(n24), .C2(n1348), .A(n1347), .B(n1346), .ZN(
        curr_proc_regs[523]) );
  AOI22_X1 U2022 ( .A1(n104), .A2(regs[12]), .B1(n71), .B2(regs[2060]), .ZN(
        n1350) );
  AOI22_X1 U2023 ( .A1(n61), .A2(regs[1036]), .B1(n98), .B2(regs[1548]), .ZN(
        n1349) );
  OAI211_X1 U2024 ( .C1(n24), .C2(n1351), .A(n1350), .B(n1349), .ZN(
        curr_proc_regs[524]) );
  AOI22_X1 U2025 ( .A1(n106), .A2(regs[13]), .B1(n71), .B2(regs[2061]), .ZN(
        n1353) );
  AOI22_X1 U2026 ( .A1(n57), .A2(regs[1037]), .B1(n98), .B2(regs[1549]), .ZN(
        n1352) );
  OAI211_X1 U2027 ( .C1(n24), .C2(n1354), .A(n1353), .B(n1352), .ZN(
        curr_proc_regs[525]) );
  AOI22_X1 U2028 ( .A1(n104), .A2(regs[14]), .B1(n71), .B2(regs[2062]), .ZN(
        n1356) );
  AOI22_X1 U2029 ( .A1(n96), .A2(regs[1550]), .B1(n34), .B2(regs[526]), .ZN(
        n1355) );
  OAI211_X1 U2030 ( .C1(n65), .C2(n1357), .A(n1356), .B(n1355), .ZN(
        curr_proc_regs[526]) );
  AOI22_X1 U2031 ( .A1(n105), .A2(regs[15]), .B1(n71), .B2(regs[2063]), .ZN(
        n1359) );
  AOI22_X1 U2032 ( .A1(n78), .A2(regs[1551]), .B1(n43), .B2(regs[527]), .ZN(
        n1358) );
  OAI211_X1 U2033 ( .C1(n63), .C2(n1360), .A(n1359), .B(n1358), .ZN(
        curr_proc_regs[527]) );
  AOI22_X1 U2034 ( .A1(n106), .A2(regs[16]), .B1(n71), .B2(regs[2064]), .ZN(
        n1362) );
  AOI22_X1 U2035 ( .A1(n81), .A2(regs[1552]), .B1(n43), .B2(regs[528]), .ZN(
        n1361) );
  OAI211_X1 U2036 ( .C1(n65), .C2(n1363), .A(n1362), .B(n1361), .ZN(
        curr_proc_regs[528]) );
  AOI22_X1 U2037 ( .A1(n105), .A2(regs[17]), .B1(n71), .B2(regs[2065]), .ZN(
        n1365) );
  AOI22_X1 U2038 ( .A1(n82), .A2(regs[1553]), .B1(n43), .B2(regs[529]), .ZN(
        n1364) );
  OAI211_X1 U2039 ( .C1(n63), .C2(n1366), .A(n1365), .B(n1364), .ZN(
        curr_proc_regs[529]) );
  INV_X1 U2040 ( .A(regs[1076]), .ZN(n1479) );
  AOI22_X1 U2041 ( .A1(n106), .A2(regs[2100]), .B1(n71), .B2(regs[1588]), .ZN(
        n1368) );
  AOI22_X1 U2042 ( .A1(n57), .A2(regs[564]), .B1(n43), .B2(regs[52]), .ZN(
        n1367) );
  OAI211_X1 U2043 ( .C1(n5), .C2(n1479), .A(n1368), .B(n1367), .ZN(
        curr_proc_regs[52]) );
  AOI22_X1 U2044 ( .A1(n106), .A2(regs[18]), .B1(n71), .B2(regs[2066]), .ZN(
        n1370) );
  AOI22_X1 U2045 ( .A1(n79), .A2(regs[1554]), .B1(n43), .B2(regs[530]), .ZN(
        n1369) );
  OAI211_X1 U2046 ( .C1(n65), .C2(n1371), .A(n1370), .B(n1369), .ZN(
        curr_proc_regs[530]) );
  AOI22_X1 U2047 ( .A1(n106), .A2(regs[19]), .B1(n71), .B2(regs[2067]), .ZN(
        n1373) );
  AOI22_X1 U2048 ( .A1(n57), .A2(regs[1043]), .B1(n82), .B2(regs[1555]), .ZN(
        n1372) );
  OAI211_X1 U2049 ( .C1(n24), .C2(n1374), .A(n1373), .B(n1372), .ZN(
        curr_proc_regs[531]) );
  AOI22_X1 U2050 ( .A1(n106), .A2(regs[20]), .B1(n71), .B2(regs[2068]), .ZN(
        n1376) );
  AOI22_X1 U2051 ( .A1(n80), .A2(regs[1556]), .B1(n43), .B2(regs[532]), .ZN(
        n1375) );
  OAI211_X1 U2052 ( .C1(n65), .C2(n1377), .A(n1376), .B(n1375), .ZN(
        curr_proc_regs[532]) );
  AOI22_X1 U2053 ( .A1(n106), .A2(regs[21]), .B1(n71), .B2(regs[2069]), .ZN(
        n1379) );
  AOI22_X1 U2054 ( .A1(n57), .A2(regs[1045]), .B1(n81), .B2(regs[1557]), .ZN(
        n1378) );
  OAI211_X1 U2055 ( .C1(n24), .C2(n1380), .A(n1379), .B(n1378), .ZN(
        curr_proc_regs[533]) );
  AOI22_X1 U2056 ( .A1(n106), .A2(regs[22]), .B1(n71), .B2(regs[2070]), .ZN(
        n1382) );
  AOI22_X1 U2057 ( .A1(n57), .A2(regs[1046]), .B1(n85), .B2(regs[1558]), .ZN(
        n1381) );
  OAI211_X1 U2058 ( .C1(n24), .C2(n1383), .A(n1382), .B(n1381), .ZN(
        curr_proc_regs[534]) );
  AOI22_X1 U2059 ( .A1(n106), .A2(regs[23]), .B1(n71), .B2(regs[2071]), .ZN(
        n1385) );
  AOI22_X1 U2060 ( .A1(n83), .A2(regs[1559]), .B1(n43), .B2(regs[535]), .ZN(
        n1384) );
  OAI211_X1 U2061 ( .C1(n65), .C2(n1386), .A(n1385), .B(n1384), .ZN(
        curr_proc_regs[535]) );
  AOI22_X1 U2062 ( .A1(n106), .A2(regs[24]), .B1(n71), .B2(regs[2072]), .ZN(
        n1388) );
  AOI22_X1 U2063 ( .A1(n57), .A2(regs[1048]), .B1(n84), .B2(regs[1560]), .ZN(
        n1387) );
  OAI211_X1 U2064 ( .C1(n24), .C2(n1389), .A(n1388), .B(n1387), .ZN(
        curr_proc_regs[536]) );
  AOI22_X1 U2065 ( .A1(n106), .A2(regs[25]), .B1(n71), .B2(regs[2073]), .ZN(
        n1391) );
  AOI22_X1 U2066 ( .A1(n84), .A2(regs[1561]), .B1(n26), .B2(regs[537]), .ZN(
        n1390) );
  OAI211_X1 U2067 ( .C1(n65), .C2(n1392), .A(n1391), .B(n1390), .ZN(
        curr_proc_regs[537]) );
  AOI22_X1 U2068 ( .A1(n106), .A2(regs[26]), .B1(n71), .B2(regs[2074]), .ZN(
        n1394) );
  AOI22_X1 U2069 ( .A1(n85), .A2(regs[1562]), .B1(n26), .B2(regs[538]), .ZN(
        n1393) );
  OAI211_X1 U2070 ( .C1(n65), .C2(n1395), .A(n1394), .B(n1393), .ZN(
        curr_proc_regs[538]) );
  AOI22_X1 U2071 ( .A1(n106), .A2(regs[27]), .B1(n71), .B2(regs[2075]), .ZN(
        n1397) );
  AOI22_X1 U2072 ( .A1(n86), .A2(regs[1563]), .B1(n26), .B2(regs[539]), .ZN(
        n1396) );
  OAI211_X1 U2073 ( .C1(n65), .C2(n1398), .A(n1397), .B(n1396), .ZN(
        curr_proc_regs[539]) );
  INV_X1 U2074 ( .A(regs[565]), .ZN(n1482) );
  AOI22_X1 U2075 ( .A1(n104), .A2(regs[2101]), .B1(n71), .B2(regs[1589]), .ZN(
        n1400) );
  AOI22_X1 U2076 ( .A1(n87), .A2(regs[1077]), .B1(n26), .B2(regs[53]), .ZN(
        n1399) );
  OAI211_X1 U2077 ( .C1(n65), .C2(n1482), .A(n1400), .B(n1399), .ZN(
        curr_proc_regs[53]) );
  AOI22_X1 U2078 ( .A1(n106), .A2(regs[28]), .B1(n71), .B2(regs[2076]), .ZN(
        n1402) );
  AOI22_X1 U2079 ( .A1(n61), .A2(regs[1052]), .B1(n86), .B2(regs[1564]), .ZN(
        n1401) );
  OAI211_X1 U2080 ( .C1(n24), .C2(n1403), .A(n1402), .B(n1401), .ZN(
        curr_proc_regs[540]) );
  AOI22_X1 U2081 ( .A1(n104), .A2(regs[29]), .B1(n71), .B2(regs[2077]), .ZN(
        n1405) );
  AOI22_X1 U2082 ( .A1(n98), .A2(regs[1565]), .B1(n26), .B2(regs[541]), .ZN(
        n1404) );
  OAI211_X1 U2083 ( .C1(n65), .C2(n1406), .A(n1405), .B(n1404), .ZN(
        curr_proc_regs[541]) );
  AOI22_X1 U2084 ( .A1(n105), .A2(regs[30]), .B1(n71), .B2(regs[2078]), .ZN(
        n1408) );
  AOI22_X1 U2085 ( .A1(n84), .A2(regs[1566]), .B1(n26), .B2(regs[542]), .ZN(
        n1407) );
  OAI211_X1 U2086 ( .C1(n63), .C2(n1409), .A(n1408), .B(n1407), .ZN(
        curr_proc_regs[542]) );
  AOI22_X1 U2087 ( .A1(n105), .A2(regs[31]), .B1(n71), .B2(regs[2079]), .ZN(
        n1411) );
  AOI22_X1 U2088 ( .A1(n2), .A2(regs[1055]), .B1(n95), .B2(regs[1567]), .ZN(
        n1410) );
  OAI211_X1 U2089 ( .C1(n24), .C2(n1412), .A(n1411), .B(n1410), .ZN(
        curr_proc_regs[543]) );
  AOI22_X1 U2090 ( .A1(n106), .A2(regs[32]), .B1(n71), .B2(regs[2080]), .ZN(
        n1414) );
  AOI22_X1 U2091 ( .A1(n13), .A2(regs[1056]), .B1(n98), .B2(regs[1568]), .ZN(
        n1413) );
  OAI211_X1 U2092 ( .C1(n24), .C2(n1415), .A(n1414), .B(n1413), .ZN(
        curr_proc_regs[544]) );
  AOI22_X1 U2093 ( .A1(n104), .A2(regs[33]), .B1(n71), .B2(regs[2081]), .ZN(
        n1417) );
  AOI22_X1 U2094 ( .A1(n95), .A2(regs[1569]), .B1(n26), .B2(regs[545]), .ZN(
        n1416) );
  OAI211_X1 U2095 ( .C1(n2207), .C2(n1418), .A(n1417), .B(n1416), .ZN(
        curr_proc_regs[545]) );
  AOI22_X1 U2096 ( .A1(n105), .A2(regs[34]), .B1(n71), .B2(regs[2082]), .ZN(
        n1420) );
  AOI22_X1 U2097 ( .A1(n13), .A2(regs[1058]), .B1(n79), .B2(regs[1570]), .ZN(
        n1419) );
  OAI211_X1 U2098 ( .C1(n25), .C2(n1421), .A(n1420), .B(n1419), .ZN(
        curr_proc_regs[546]) );
  AOI22_X1 U2099 ( .A1(n106), .A2(regs[35]), .B1(n71), .B2(regs[2083]), .ZN(
        n1423) );
  AOI22_X1 U2100 ( .A1(n94), .A2(regs[1571]), .B1(n26), .B2(regs[547]), .ZN(
        n1422) );
  OAI211_X1 U2101 ( .C1(n64), .C2(n1424), .A(n1423), .B(n1422), .ZN(
        curr_proc_regs[547]) );
  AOI22_X1 U2102 ( .A1(n106), .A2(regs[36]), .B1(n71), .B2(regs[2084]), .ZN(
        n1426) );
  AOI22_X1 U2103 ( .A1(n88), .A2(regs[1572]), .B1(n26), .B2(regs[548]), .ZN(
        n1425) );
  OAI211_X1 U2104 ( .C1(n2207), .C2(n1427), .A(n1426), .B(n1425), .ZN(
        curr_proc_regs[548]) );
  AOI22_X1 U2105 ( .A1(n104), .A2(regs[37]), .B1(n71), .B2(regs[2085]), .ZN(
        n1429) );
  AOI22_X1 U2106 ( .A1(n13), .A2(regs[1061]), .B1(n87), .B2(regs[1573]), .ZN(
        n1428) );
  OAI211_X1 U2107 ( .C1(n2134), .C2(n1430), .A(n1429), .B(n1428), .ZN(
        curr_proc_regs[549]) );
  INV_X1 U2108 ( .A(regs[1078]), .ZN(n1485) );
  AOI22_X1 U2109 ( .A1(n104), .A2(regs[2102]), .B1(n71), .B2(regs[1590]), .ZN(
        n1432) );
  AOI22_X1 U2110 ( .A1(n58), .A2(regs[566]), .B1(n26), .B2(regs[54]), .ZN(
        n1431) );
  OAI211_X1 U2111 ( .C1(n99), .C2(n1485), .A(n1432), .B(n1431), .ZN(
        curr_proc_regs[54]) );
  AOI22_X1 U2112 ( .A1(n105), .A2(regs[38]), .B1(n71), .B2(regs[2086]), .ZN(
        n1434) );
  AOI22_X1 U2113 ( .A1(n58), .A2(regs[1062]), .B1(n85), .B2(regs[1574]), .ZN(
        n1433) );
  OAI211_X1 U2114 ( .C1(n2134), .C2(n1435), .A(n1434), .B(n1433), .ZN(
        curr_proc_regs[550]) );
  AOI22_X1 U2115 ( .A1(n106), .A2(regs[39]), .B1(n71), .B2(regs[2087]), .ZN(
        n1437) );
  AOI22_X1 U2116 ( .A1(n58), .A2(regs[1063]), .B1(n84), .B2(regs[1575]), .ZN(
        n1436) );
  OAI211_X1 U2117 ( .C1(n2134), .C2(n1438), .A(n1437), .B(n1436), .ZN(
        curr_proc_regs[551]) );
  AOI22_X1 U2118 ( .A1(n104), .A2(regs[40]), .B1(n71), .B2(regs[2088]), .ZN(
        n1440) );
  AOI22_X1 U2119 ( .A1(n58), .A2(regs[1064]), .B1(n97), .B2(regs[1576]), .ZN(
        n1439) );
  OAI211_X1 U2120 ( .C1(n2134), .C2(n1441), .A(n1440), .B(n1439), .ZN(
        curr_proc_regs[552]) );
  AOI22_X1 U2121 ( .A1(n105), .A2(regs[41]), .B1(n71), .B2(regs[2089]), .ZN(
        n1443) );
  AOI22_X1 U2122 ( .A1(n90), .A2(regs[1577]), .B1(n26), .B2(regs[553]), .ZN(
        n1442) );
  OAI211_X1 U2123 ( .C1(n2207), .C2(n1444), .A(n1443), .B(n1442), .ZN(
        curr_proc_regs[553]) );
  AOI22_X1 U2124 ( .A1(n106), .A2(regs[42]), .B1(n71), .B2(regs[2090]), .ZN(
        n1446) );
  AOI22_X1 U2125 ( .A1(n92), .A2(regs[1578]), .B1(n27), .B2(regs[554]), .ZN(
        n1445) );
  OAI211_X1 U2126 ( .C1(n2207), .C2(n1447), .A(n1446), .B(n1445), .ZN(
        curr_proc_regs[554]) );
  AOI22_X1 U2127 ( .A1(n104), .A2(regs[43]), .B1(n71), .B2(regs[2091]), .ZN(
        n1449) );
  AOI22_X1 U2128 ( .A1(n93), .A2(regs[1579]), .B1(n27), .B2(regs[555]), .ZN(
        n1448) );
  OAI211_X1 U2129 ( .C1(n63), .C2(n1450), .A(n1449), .B(n1448), .ZN(
        curr_proc_regs[555]) );
  AOI22_X1 U2130 ( .A1(n105), .A2(regs[44]), .B1(n74), .B2(regs[2092]), .ZN(
        n1452) );
  AOI22_X1 U2131 ( .A1(n58), .A2(regs[1068]), .B1(n81), .B2(regs[1580]), .ZN(
        n1451) );
  OAI211_X1 U2132 ( .C1(n2134), .C2(n1453), .A(n1452), .B(n1451), .ZN(
        curr_proc_regs[556]) );
  AOI22_X1 U2133 ( .A1(n106), .A2(regs[45]), .B1(n4), .B2(regs[2093]), .ZN(
        n1455) );
  AOI22_X1 U2134 ( .A1(n58), .A2(regs[1069]), .B1(n82), .B2(regs[1581]), .ZN(
        n1454) );
  OAI211_X1 U2135 ( .C1(n24), .C2(n1456), .A(n1455), .B(n1454), .ZN(
        curr_proc_regs[557]) );
  AOI22_X1 U2136 ( .A1(n104), .A2(regs[46]), .B1(n14), .B2(regs[2094]), .ZN(
        n1458) );
  AOI22_X1 U2137 ( .A1(n57), .A2(regs[1070]), .B1(n78), .B2(regs[1582]), .ZN(
        n1457) );
  OAI211_X1 U2138 ( .C1(n24), .C2(n1459), .A(n1458), .B(n1457), .ZN(
        curr_proc_regs[558]) );
  AOI22_X1 U2139 ( .A1(n105), .A2(regs[47]), .B1(n70), .B2(regs[2095]), .ZN(
        n1461) );
  AOI22_X1 U2140 ( .A1(n57), .A2(regs[1071]), .B1(n79), .B2(regs[1583]), .ZN(
        n1460) );
  OAI211_X1 U2141 ( .C1(n24), .C2(n1462), .A(n1461), .B(n1460), .ZN(
        curr_proc_regs[559]) );
  INV_X1 U2142 ( .A(regs[1079]), .ZN(n1488) );
  AOI22_X1 U2143 ( .A1(n105), .A2(regs[2103]), .B1(n74), .B2(regs[1591]), .ZN(
        n1464) );
  AOI22_X1 U2144 ( .A1(n57), .A2(regs[567]), .B1(n27), .B2(regs[55]), .ZN(
        n1463) );
  OAI211_X1 U2145 ( .C1(n5), .C2(n1488), .A(n1464), .B(n1463), .ZN(
        curr_proc_regs[55]) );
  AOI22_X1 U2146 ( .A1(n105), .A2(regs[48]), .B1(n4), .B2(regs[2096]), .ZN(
        n1466) );
  AOI22_X1 U2147 ( .A1(n57), .A2(regs[1072]), .B1(n80), .B2(regs[1584]), .ZN(
        n1465) );
  OAI211_X1 U2148 ( .C1(n24), .C2(n1467), .A(n1466), .B(n1465), .ZN(
        curr_proc_regs[560]) );
  AOI22_X1 U2149 ( .A1(n105), .A2(regs[49]), .B1(n14), .B2(regs[2097]), .ZN(
        n1469) );
  AOI22_X1 U2150 ( .A1(n88), .A2(regs[1585]), .B1(n27), .B2(regs[561]), .ZN(
        n1468) );
  OAI211_X1 U2151 ( .C1(n2207), .C2(n1470), .A(n1469), .B(n1468), .ZN(
        curr_proc_regs[561]) );
  AOI22_X1 U2152 ( .A1(n105), .A2(regs[50]), .B1(n70), .B2(regs[2098]), .ZN(
        n1472) );
  AOI22_X1 U2153 ( .A1(n57), .A2(regs[1074]), .B1(n82), .B2(regs[1586]), .ZN(
        n1471) );
  OAI211_X1 U2154 ( .C1(n24), .C2(n1473), .A(n1472), .B(n1471), .ZN(
        curr_proc_regs[562]) );
  AOI22_X1 U2155 ( .A1(n105), .A2(regs[51]), .B1(n74), .B2(regs[2099]), .ZN(
        n1475) );
  AOI22_X1 U2156 ( .A1(n59), .A2(regs[1075]), .B1(n78), .B2(regs[1587]), .ZN(
        n1474) );
  OAI211_X1 U2157 ( .C1(n24), .C2(n1476), .A(n1475), .B(n1474), .ZN(
        curr_proc_regs[563]) );
  AOI22_X1 U2158 ( .A1(n105), .A2(regs[52]), .B1(n4), .B2(regs[2100]), .ZN(
        n1478) );
  AOI22_X1 U2159 ( .A1(n90), .A2(regs[1588]), .B1(n27), .B2(regs[564]), .ZN(
        n1477) );
  OAI211_X1 U2160 ( .C1(n63), .C2(n1479), .A(n1478), .B(n1477), .ZN(
        curr_proc_regs[564]) );
  AOI22_X1 U2161 ( .A1(n105), .A2(regs[53]), .B1(n14), .B2(regs[2101]), .ZN(
        n1481) );
  AOI22_X1 U2162 ( .A1(n59), .A2(regs[1077]), .B1(n80), .B2(regs[1589]), .ZN(
        n1480) );
  OAI211_X1 U2163 ( .C1(n24), .C2(n1482), .A(n1481), .B(n1480), .ZN(
        curr_proc_regs[565]) );
  AOI22_X1 U2164 ( .A1(n105), .A2(regs[54]), .B1(n4), .B2(regs[2102]), .ZN(
        n1484) );
  AOI22_X1 U2165 ( .A1(n92), .A2(regs[1590]), .B1(n27), .B2(regs[566]), .ZN(
        n1483) );
  OAI211_X1 U2166 ( .C1(n64), .C2(n1485), .A(n1484), .B(n1483), .ZN(
        curr_proc_regs[566]) );
  AOI22_X1 U2167 ( .A1(n105), .A2(regs[55]), .B1(n14), .B2(regs[2103]), .ZN(
        n1487) );
  AOI22_X1 U2168 ( .A1(n93), .A2(regs[1591]), .B1(n27), .B2(regs[567]), .ZN(
        n1486) );
  OAI211_X1 U2169 ( .C1(n63), .C2(n1488), .A(n1487), .B(n1486), .ZN(
        curr_proc_regs[567]) );
  INV_X1 U2170 ( .A(regs[1592]), .ZN(n1491) );
  AOI22_X1 U2171 ( .A1(n105), .A2(regs[56]), .B1(n70), .B2(regs[2104]), .ZN(
        n1490) );
  AOI22_X1 U2172 ( .A1(n59), .A2(regs[1080]), .B1(n27), .B2(regs[568]), .ZN(
        n1489) );
  OAI211_X1 U2173 ( .C1(n5), .C2(n1491), .A(n1490), .B(n1489), .ZN(
        curr_proc_regs[568]) );
  INV_X1 U2174 ( .A(regs[1593]), .ZN(n1494) );
  AOI22_X1 U2175 ( .A1(n105), .A2(regs[57]), .B1(n70), .B2(regs[2105]), .ZN(
        n1493) );
  AOI22_X1 U2176 ( .A1(n59), .A2(regs[1081]), .B1(n27), .B2(regs[569]), .ZN(
        n1492) );
  OAI211_X1 U2177 ( .C1(n5), .C2(n1494), .A(n1493), .B(n1492), .ZN(
        curr_proc_regs[569]) );
  INV_X1 U2178 ( .A(regs[1080]), .ZN(n1497) );
  AOI22_X1 U2179 ( .A1(n104), .A2(regs[2104]), .B1(n74), .B2(regs[1592]), .ZN(
        n1496) );
  AOI22_X1 U2180 ( .A1(n59), .A2(regs[568]), .B1(n27), .B2(regs[56]), .ZN(
        n1495) );
  OAI211_X1 U2181 ( .C1(n5), .C2(n1497), .A(n1496), .B(n1495), .ZN(
        curr_proc_regs[56]) );
  INV_X1 U2182 ( .A(regs[1594]), .ZN(n1500) );
  AOI22_X1 U2183 ( .A1(n104), .A2(regs[58]), .B1(n4), .B2(regs[2106]), .ZN(
        n1499) );
  AOI22_X1 U2184 ( .A1(n59), .A2(regs[1082]), .B1(n27), .B2(regs[570]), .ZN(
        n1498) );
  OAI211_X1 U2185 ( .C1(n5), .C2(n1500), .A(n1499), .B(n1498), .ZN(
        curr_proc_regs[570]) );
  INV_X1 U2186 ( .A(regs[1595]), .ZN(n1503) );
  AOI22_X1 U2187 ( .A1(n104), .A2(regs[59]), .B1(n14), .B2(regs[2107]), .ZN(
        n1502) );
  AOI22_X1 U2188 ( .A1(n58), .A2(regs[1083]), .B1(n34), .B2(regs[571]), .ZN(
        n1501) );
  OAI211_X1 U2189 ( .C1(n5), .C2(n1503), .A(n1502), .B(n1501), .ZN(
        curr_proc_regs[571]) );
  INV_X1 U2190 ( .A(regs[1084]), .ZN(n1615) );
  AOI22_X1 U2191 ( .A1(n104), .A2(regs[60]), .B1(n74), .B2(regs[2108]), .ZN(
        n1505) );
  AOI22_X1 U2192 ( .A1(n88), .A2(regs[1596]), .B1(n32), .B2(regs[572]), .ZN(
        n1504) );
  OAI211_X1 U2193 ( .C1(n2207), .C2(n1615), .A(n1505), .B(n1504), .ZN(
        curr_proc_regs[572]) );
  INV_X1 U2194 ( .A(regs[1597]), .ZN(n1508) );
  AOI22_X1 U2195 ( .A1(n104), .A2(regs[61]), .B1(n70), .B2(regs[2109]), .ZN(
        n1507) );
  AOI22_X1 U2196 ( .A1(n58), .A2(regs[1085]), .B1(n41), .B2(regs[573]), .ZN(
        n1506) );
  OAI211_X1 U2197 ( .C1(n5), .C2(n1508), .A(n1507), .B(n1506), .ZN(
        curr_proc_regs[573]) );
  INV_X1 U2198 ( .A(regs[1598]), .ZN(n1511) );
  AOI22_X1 U2199 ( .A1(n104), .A2(regs[62]), .B1(n74), .B2(regs[2110]), .ZN(
        n1510) );
  AOI22_X1 U2200 ( .A1(n58), .A2(regs[1086]), .B1(n43), .B2(regs[574]), .ZN(
        n1509) );
  OAI211_X1 U2201 ( .C1(n100), .C2(n1511), .A(n1510), .B(n1509), .ZN(
        curr_proc_regs[574]) );
  INV_X1 U2202 ( .A(regs[1599]), .ZN(n1514) );
  AOI22_X1 U2203 ( .A1(n104), .A2(regs[63]), .B1(n4), .B2(regs[2111]), .ZN(
        n1513) );
  AOI22_X1 U2204 ( .A1(n58), .A2(regs[1087]), .B1(n3), .B2(regs[575]), .ZN(
        n1512) );
  OAI211_X1 U2205 ( .C1(n5), .C2(n1514), .A(n1513), .B(n1512), .ZN(
        curr_proc_regs[575]) );
  INV_X1 U2206 ( .A(regs[1088]), .ZN(n1746) );
  AOI22_X1 U2207 ( .A1(n104), .A2(regs[64]), .B1(n74), .B2(regs[2112]), .ZN(
        n1516) );
  AOI22_X1 U2208 ( .A1(n90), .A2(regs[1600]), .B1(n3), .B2(regs[576]), .ZN(
        n1515) );
  OAI211_X1 U2209 ( .C1(n64), .C2(n1746), .A(n1516), .B(n1515), .ZN(
        curr_proc_regs[576]) );
  INV_X1 U2210 ( .A(regs[1601]), .ZN(n1519) );
  AOI22_X1 U2211 ( .A1(n104), .A2(regs[65]), .B1(n74), .B2(regs[2113]), .ZN(
        n1518) );
  AOI22_X1 U2212 ( .A1(n58), .A2(regs[1089]), .B1(n12), .B2(regs[577]), .ZN(
        n1517) );
  OAI211_X1 U2213 ( .C1(n16), .C2(n1519), .A(n1518), .B(n1517), .ZN(
        curr_proc_regs[577]) );
  INV_X1 U2214 ( .A(regs[1090]), .ZN(n1812) );
  AOI22_X1 U2215 ( .A1(n104), .A2(regs[66]), .B1(n74), .B2(regs[2114]), .ZN(
        n1521) );
  AOI22_X1 U2216 ( .A1(n78), .A2(regs[1602]), .B1(n12), .B2(regs[578]), .ZN(
        n1520) );
  OAI211_X1 U2217 ( .C1(n63), .C2(n1812), .A(n1521), .B(n1520), .ZN(
        curr_proc_regs[578]) );
  INV_X1 U2218 ( .A(regs[1603]), .ZN(n1524) );
  AOI22_X1 U2219 ( .A1(n104), .A2(regs[67]), .B1(n74), .B2(regs[2115]), .ZN(
        n1523) );
  AOI22_X1 U2220 ( .A1(n50), .A2(regs[1091]), .B1(n28), .B2(regs[579]), .ZN(
        n1522) );
  OAI211_X1 U2221 ( .C1(n99), .C2(n1524), .A(n1523), .B(n1522), .ZN(
        curr_proc_regs[579]) );
  INV_X1 U2222 ( .A(regs[569]), .ZN(n1527) );
  AOI22_X1 U2223 ( .A1(n21), .A2(regs[2105]), .B1(n74), .B2(regs[1593]), .ZN(
        n1526) );
  AOI22_X1 U2224 ( .A1(n92), .A2(regs[1081]), .B1(n34), .B2(regs[57]), .ZN(
        n1525) );
  OAI211_X1 U2225 ( .C1(n2207), .C2(n1527), .A(n1526), .B(n1525), .ZN(
        curr_proc_regs[57]) );
  INV_X1 U2226 ( .A(regs[1604]), .ZN(n1530) );
  AOI22_X1 U2227 ( .A1(n21), .A2(regs[68]), .B1(n74), .B2(regs[2116]), .ZN(
        n1529) );
  AOI22_X1 U2228 ( .A1(n57), .A2(regs[1092]), .B1(n32), .B2(regs[580]), .ZN(
        n1528) );
  OAI211_X1 U2229 ( .C1(n100), .C2(n1530), .A(n1529), .B(n1528), .ZN(
        curr_proc_regs[580]) );
  INV_X1 U2230 ( .A(regs[1605]), .ZN(n1533) );
  AOI22_X1 U2231 ( .A1(n21), .A2(regs[69]), .B1(n74), .B2(regs[2117]), .ZN(
        n1532) );
  AOI22_X1 U2232 ( .A1(n52), .A2(regs[1093]), .B1(n28), .B2(regs[581]), .ZN(
        n1531) );
  OAI211_X1 U2233 ( .C1(n102), .C2(n1533), .A(n1532), .B(n1531), .ZN(
        curr_proc_regs[581]) );
  INV_X1 U2234 ( .A(regs[1094]), .ZN(n1947) );
  AOI22_X1 U2235 ( .A1(n21), .A2(regs[70]), .B1(n74), .B2(regs[2118]), .ZN(
        n1535) );
  AOI22_X1 U2236 ( .A1(n93), .A2(regs[1606]), .B1(n28), .B2(regs[582]), .ZN(
        n1534) );
  OAI211_X1 U2237 ( .C1(n2207), .C2(n1947), .A(n1535), .B(n1534), .ZN(
        curr_proc_regs[582]) );
  INV_X1 U2238 ( .A(regs[1607]), .ZN(n1538) );
  AOI22_X1 U2239 ( .A1(n21), .A2(regs[71]), .B1(n74), .B2(regs[2119]), .ZN(
        n1537) );
  AOI22_X1 U2240 ( .A1(n62), .A2(regs[1095]), .B1(n28), .B2(regs[583]), .ZN(
        n1536) );
  OAI211_X1 U2241 ( .C1(n5), .C2(n1538), .A(n1537), .B(n1536), .ZN(
        curr_proc_regs[583]) );
  INV_X1 U2242 ( .A(regs[1096]), .ZN(n2013) );
  AOI22_X1 U2243 ( .A1(n21), .A2(regs[72]), .B1(n74), .B2(regs[2120]), .ZN(
        n1540) );
  AOI22_X1 U2244 ( .A1(n88), .A2(regs[1608]), .B1(n28), .B2(regs[584]), .ZN(
        n1539) );
  OAI211_X1 U2245 ( .C1(n63), .C2(n2013), .A(n1540), .B(n1539), .ZN(
        curr_proc_regs[584]) );
  INV_X1 U2246 ( .A(regs[1097]), .ZN(n2046) );
  AOI22_X1 U2247 ( .A1(n21), .A2(regs[73]), .B1(n74), .B2(regs[2121]), .ZN(
        n1542) );
  AOI22_X1 U2248 ( .A1(n90), .A2(regs[1609]), .B1(n28), .B2(regs[585]), .ZN(
        n1541) );
  OAI211_X1 U2249 ( .C1(n64), .C2(n2046), .A(n1542), .B(n1541), .ZN(
        curr_proc_regs[585]) );
  INV_X1 U2250 ( .A(regs[1098]), .ZN(n2079) );
  AOI22_X1 U2251 ( .A1(n21), .A2(regs[74]), .B1(n74), .B2(regs[2122]), .ZN(
        n1544) );
  AOI22_X1 U2252 ( .A1(n89), .A2(regs[1610]), .B1(n28), .B2(regs[586]), .ZN(
        n1543) );
  OAI211_X1 U2253 ( .C1(n2207), .C2(n2079), .A(n1544), .B(n1543), .ZN(
        curr_proc_regs[586]) );
  INV_X1 U2254 ( .A(regs[1611]), .ZN(n1547) );
  AOI22_X1 U2255 ( .A1(n21), .A2(regs[75]), .B1(n14), .B2(regs[2123]), .ZN(
        n1546) );
  AOI22_X1 U2256 ( .A1(n59), .A2(regs[1099]), .B1(n28), .B2(regs[587]), .ZN(
        n1545) );
  OAI211_X1 U2257 ( .C1(n99), .C2(n1547), .A(n1546), .B(n1545), .ZN(
        curr_proc_regs[587]) );
  INV_X1 U2258 ( .A(regs[1100]), .ZN(n2140) );
  AOI22_X1 U2259 ( .A1(n21), .A2(regs[76]), .B1(n4), .B2(regs[2124]), .ZN(
        n1549) );
  AOI22_X1 U2260 ( .A1(n91), .A2(regs[1612]), .B1(n28), .B2(regs[588]), .ZN(
        n1548) );
  OAI211_X1 U2261 ( .C1(n1), .C2(n2140), .A(n1549), .B(n1548), .ZN(
        curr_proc_regs[588]) );
  INV_X1 U2262 ( .A(regs[1613]), .ZN(n1552) );
  AOI22_X1 U2263 ( .A1(n21), .A2(regs[77]), .B1(n14), .B2(regs[2125]), .ZN(
        n1551) );
  AOI22_X1 U2264 ( .A1(n54), .A2(regs[1101]), .B1(n28), .B2(regs[589]), .ZN(
        n1550) );
  OAI211_X1 U2265 ( .C1(n2221), .C2(n1552), .A(n1551), .B(n1550), .ZN(
        curr_proc_regs[589]) );
  INV_X1 U2266 ( .A(regs[570]), .ZN(n1555) );
  AOI22_X1 U2267 ( .A1(n21), .A2(regs[2106]), .B1(n4), .B2(regs[1594]), .ZN(
        n1554) );
  AOI22_X1 U2268 ( .A1(n97), .A2(regs[1082]), .B1(n28), .B2(regs[58]), .ZN(
        n1553) );
  OAI211_X1 U2269 ( .C1(n63), .C2(n1555), .A(n1554), .B(n1553), .ZN(
        curr_proc_regs[58]) );
  INV_X1 U2270 ( .A(regs[1102]), .ZN(n2146) );
  AOI22_X1 U2271 ( .A1(n21), .A2(regs[78]), .B1(n70), .B2(regs[2126]), .ZN(
        n1557) );
  AOI22_X1 U2272 ( .A1(n86), .A2(regs[1614]), .B1(n28), .B2(regs[590]), .ZN(
        n1556) );
  OAI211_X1 U2273 ( .C1(n11), .C2(n2146), .A(n1557), .B(n1556), .ZN(
        curr_proc_regs[590]) );
  INV_X1 U2274 ( .A(regs[1103]), .ZN(n2149) );
  AOI22_X1 U2275 ( .A1(n21), .A2(regs[79]), .B1(n74), .B2(regs[2127]), .ZN(
        n1559) );
  AOI22_X1 U2276 ( .A1(n81), .A2(regs[1615]), .B1(n29), .B2(regs[591]), .ZN(
        n1558) );
  OAI211_X1 U2277 ( .C1(n11), .C2(n2149), .A(n1559), .B(n1558), .ZN(
        curr_proc_regs[591]) );
  INV_X1 U2278 ( .A(regs[1104]), .ZN(n2155) );
  AOI22_X1 U2279 ( .A1(n21), .A2(regs[80]), .B1(n14), .B2(regs[2128]), .ZN(
        n1561) );
  AOI22_X1 U2280 ( .A1(n82), .A2(regs[1616]), .B1(n29), .B2(regs[592]), .ZN(
        n1560) );
  OAI211_X1 U2281 ( .C1(n11), .C2(n2155), .A(n1561), .B(n1560), .ZN(
        curr_proc_regs[592]) );
  INV_X1 U2282 ( .A(regs[1105]), .ZN(n2158) );
  AOI22_X1 U2283 ( .A1(n21), .A2(regs[81]), .B1(n4), .B2(regs[2129]), .ZN(
        n1563) );
  AOI22_X1 U2284 ( .A1(n86), .A2(regs[1617]), .B1(n29), .B2(regs[593]), .ZN(
        n1562) );
  OAI211_X1 U2285 ( .C1(n11), .C2(n2158), .A(n1563), .B(n1562), .ZN(
        curr_proc_regs[593]) );
  INV_X1 U2286 ( .A(regs[1618]), .ZN(n1566) );
  AOI22_X1 U2287 ( .A1(n21), .A2(regs[82]), .B1(n14), .B2(regs[2130]), .ZN(
        n1565) );
  AOI22_X1 U2288 ( .A1(n53), .A2(regs[1106]), .B1(n29), .B2(regs[594]), .ZN(
        n1564) );
  OAI211_X1 U2289 ( .C1(n100), .C2(n1566), .A(n1565), .B(n1564), .ZN(
        curr_proc_regs[594]) );
  INV_X1 U2290 ( .A(regs[1619]), .ZN(n1569) );
  AOI22_X1 U2291 ( .A1(n21), .A2(regs[83]), .B1(n70), .B2(regs[2131]), .ZN(
        n1568) );
  AOI22_X1 U2292 ( .A1(n59), .A2(regs[1107]), .B1(n29), .B2(regs[595]), .ZN(
        n1567) );
  OAI211_X1 U2293 ( .C1(n99), .C2(n1569), .A(n1568), .B(n1567), .ZN(
        curr_proc_regs[595]) );
  INV_X1 U2294 ( .A(regs[1620]), .ZN(n1572) );
  AOI22_X1 U2295 ( .A1(n21), .A2(regs[84]), .B1(n70), .B2(regs[2132]), .ZN(
        n1571) );
  AOI22_X1 U2296 ( .A1(n59), .A2(regs[1108]), .B1(n29), .B2(regs[596]), .ZN(
        n1570) );
  OAI211_X1 U2297 ( .C1(n100), .C2(n1572), .A(n1571), .B(n1570), .ZN(
        curr_proc_regs[596]) );
  INV_X1 U2298 ( .A(regs[1621]), .ZN(n1575) );
  AOI22_X1 U2299 ( .A1(n21), .A2(regs[85]), .B1(n74), .B2(regs[2133]), .ZN(
        n1574) );
  AOI22_X1 U2300 ( .A1(n59), .A2(regs[1109]), .B1(n29), .B2(regs[597]), .ZN(
        n1573) );
  OAI211_X1 U2301 ( .C1(n16), .C2(n1575), .A(n1574), .B(n1573), .ZN(
        curr_proc_regs[597]) );
  INV_X1 U2302 ( .A(regs[1110]), .ZN(n2173) );
  AOI22_X1 U2303 ( .A1(n21), .A2(regs[86]), .B1(n4), .B2(regs[2134]), .ZN(
        n1577) );
  AOI22_X1 U2304 ( .A1(n78), .A2(regs[1622]), .B1(n29), .B2(regs[598]), .ZN(
        n1576) );
  OAI211_X1 U2305 ( .C1(n11), .C2(n2173), .A(n1577), .B(n1576), .ZN(
        curr_proc_regs[598]) );
  INV_X1 U2306 ( .A(regs[1111]), .ZN(n2176) );
  AOI22_X1 U2307 ( .A1(n21), .A2(regs[87]), .B1(n14), .B2(regs[2135]), .ZN(
        n1579) );
  AOI22_X1 U2308 ( .A1(n79), .A2(regs[1623]), .B1(n29), .B2(regs[599]), .ZN(
        n1578) );
  OAI211_X1 U2309 ( .C1(n11), .C2(n2176), .A(n1579), .B(n1578), .ZN(
        curr_proc_regs[599]) );
  INV_X1 U2310 ( .A(regs[571]), .ZN(n1582) );
  AOI22_X1 U2311 ( .A1(n6), .A2(regs[2107]), .B1(n14), .B2(regs[1595]), .ZN(
        n1581) );
  AOI22_X1 U2312 ( .A1(n80), .A2(regs[1083]), .B1(n29), .B2(regs[59]), .ZN(
        n1580) );
  OAI211_X1 U2313 ( .C1(n11), .C2(n1582), .A(n1581), .B(n1580), .ZN(
        curr_proc_regs[59]) );
  INV_X1 U2314 ( .A(regs[517]), .ZN(n1585) );
  AOI22_X1 U2315 ( .A1(n6), .A2(regs[2053]), .B1(n70), .B2(regs[1541]), .ZN(
        n1584) );
  AOI22_X1 U2316 ( .A1(n87), .A2(regs[1029]), .B1(n29), .B2(regs[5]), .ZN(
        n1583) );
  OAI211_X1 U2317 ( .C1(n64), .C2(n1585), .A(n1584), .B(n1583), .ZN(
        curr_proc_regs[5]) );
  INV_X1 U2318 ( .A(regs[1112]), .ZN(n2179) );
  AOI22_X1 U2319 ( .A1(n6), .A2(regs[88]), .B1(n74), .B2(regs[2136]), .ZN(
        n1587) );
  AOI22_X1 U2320 ( .A1(n95), .A2(regs[1624]), .B1(n30), .B2(regs[600]), .ZN(
        n1586) );
  OAI211_X1 U2321 ( .C1(n64), .C2(n2179), .A(n1587), .B(n1586), .ZN(
        curr_proc_regs[600]) );
  INV_X1 U2322 ( .A(regs[1625]), .ZN(n1590) );
  AOI22_X1 U2323 ( .A1(n6), .A2(regs[89]), .B1(n70), .B2(regs[2137]), .ZN(
        n1589) );
  AOI22_X1 U2324 ( .A1(n49), .A2(regs[1113]), .B1(n30), .B2(regs[601]), .ZN(
        n1588) );
  OAI211_X1 U2325 ( .C1(n99), .C2(n1590), .A(n1589), .B(n1588), .ZN(
        curr_proc_regs[601]) );
  INV_X1 U2326 ( .A(regs[1626]), .ZN(n1593) );
  AOI22_X1 U2327 ( .A1(n6), .A2(regs[90]), .B1(n74), .B2(regs[2138]), .ZN(
        n1592) );
  AOI22_X1 U2328 ( .A1(n54), .A2(regs[1114]), .B1(n30), .B2(regs[602]), .ZN(
        n1591) );
  OAI211_X1 U2329 ( .C1(n102), .C2(n1593), .A(n1592), .B(n1591), .ZN(
        curr_proc_regs[602]) );
  INV_X1 U2330 ( .A(regs[1627]), .ZN(n1596) );
  AOI22_X1 U2331 ( .A1(n6), .A2(regs[91]), .B1(n14), .B2(regs[2139]), .ZN(
        n1595) );
  AOI22_X1 U2332 ( .A1(n54), .A2(regs[1115]), .B1(n30), .B2(regs[603]), .ZN(
        n1594) );
  OAI211_X1 U2333 ( .C1(n5), .C2(n1596), .A(n1595), .B(n1594), .ZN(
        curr_proc_regs[603]) );
  INV_X1 U2334 ( .A(regs[1116]), .ZN(n2194) );
  AOI22_X1 U2335 ( .A1(n6), .A2(regs[92]), .B1(n14), .B2(regs[2140]), .ZN(
        n1598) );
  AOI22_X1 U2336 ( .A1(n94), .A2(regs[1628]), .B1(n30), .B2(regs[604]), .ZN(
        n1597) );
  OAI211_X1 U2337 ( .C1(n64), .C2(n2194), .A(n1598), .B(n1597), .ZN(
        curr_proc_regs[604]) );
  INV_X1 U2338 ( .A(regs[1629]), .ZN(n1601) );
  AOI22_X1 U2339 ( .A1(n6), .A2(regs[93]), .B1(n4), .B2(regs[2141]), .ZN(n1600) );
  AOI22_X1 U2340 ( .A1(n53), .A2(regs[1117]), .B1(n30), .B2(regs[605]), .ZN(
        n1599) );
  OAI211_X1 U2341 ( .C1(n101), .C2(n1601), .A(n1600), .B(n1599), .ZN(
        curr_proc_regs[605]) );
  INV_X1 U2342 ( .A(regs[1630]), .ZN(n1604) );
  AOI22_X1 U2343 ( .A1(n6), .A2(regs[94]), .B1(n14), .B2(regs[2142]), .ZN(
        n1603) );
  AOI22_X1 U2344 ( .A1(n53), .A2(regs[1118]), .B1(n30), .B2(regs[606]), .ZN(
        n1602) );
  OAI211_X1 U2345 ( .C1(n102), .C2(n1604), .A(n1603), .B(n1602), .ZN(
        curr_proc_regs[606]) );
  INV_X1 U2346 ( .A(regs[1119]), .ZN(n2203) );
  AOI22_X1 U2347 ( .A1(n6), .A2(regs[95]), .B1(n14), .B2(regs[2143]), .ZN(
        n1606) );
  AOI22_X1 U2348 ( .A1(n83), .A2(regs[1631]), .B1(n30), .B2(regs[607]), .ZN(
        n1605) );
  OAI211_X1 U2349 ( .C1(n64), .C2(n2203), .A(n1606), .B(n1605), .ZN(
        curr_proc_regs[607]) );
  INV_X1 U2350 ( .A(regs[1632]), .ZN(n1609) );
  AOI22_X1 U2351 ( .A1(n6), .A2(regs[96]), .B1(n14), .B2(regs[2144]), .ZN(
        n1608) );
  AOI22_X1 U2352 ( .A1(n53), .A2(regs[1120]), .B1(n30), .B2(regs[608]), .ZN(
        n1607) );
  OAI211_X1 U2353 ( .C1(n102), .C2(n1609), .A(n1608), .B(n1607), .ZN(
        curr_proc_regs[608]) );
  INV_X1 U2354 ( .A(regs[1633]), .ZN(n1612) );
  AOI22_X1 U2355 ( .A1(n103), .A2(regs[97]), .B1(n14), .B2(regs[2145]), .ZN(
        n1611) );
  AOI22_X1 U2356 ( .A1(n53), .A2(regs[1121]), .B1(n30), .B2(regs[609]), .ZN(
        n1610) );
  OAI211_X1 U2357 ( .C1(n99), .C2(n1612), .A(n1611), .B(n1610), .ZN(
        curr_proc_regs[609]) );
  AOI22_X1 U2358 ( .A1(n103), .A2(regs[2108]), .B1(n14), .B2(regs[1596]), .ZN(
        n1614) );
  AOI22_X1 U2359 ( .A1(n52), .A2(regs[572]), .B1(n30), .B2(regs[60]), .ZN(
        n1613) );
  OAI211_X1 U2360 ( .C1(n100), .C2(n1615), .A(n1614), .B(n1613), .ZN(
        curr_proc_regs[60]) );
  INV_X1 U2361 ( .A(regs[1634]), .ZN(n1618) );
  AOI22_X1 U2362 ( .A1(n103), .A2(regs[98]), .B1(n70), .B2(regs[2146]), .ZN(
        n1617) );
  AOI22_X1 U2363 ( .A1(n54), .A2(regs[1122]), .B1(n31), .B2(regs[610]), .ZN(
        n1616) );
  OAI211_X1 U2364 ( .C1(n100), .C2(n1618), .A(n1617), .B(n1616), .ZN(
        curr_proc_regs[610]) );
  INV_X1 U2365 ( .A(regs[1123]), .ZN(n2216) );
  AOI22_X1 U2366 ( .A1(n103), .A2(regs[99]), .B1(n74), .B2(regs[2147]), .ZN(
        n1620) );
  AOI22_X1 U2367 ( .A1(n96), .A2(regs[1635]), .B1(n31), .B2(regs[611]), .ZN(
        n1619) );
  OAI211_X1 U2368 ( .C1(n64), .C2(n2216), .A(n1620), .B(n1619), .ZN(
        curr_proc_regs[611]) );
  AOI22_X1 U2369 ( .A1(n103), .A2(regs[100]), .B1(n14), .B2(regs[2148]), .ZN(
        n1622) );
  AOI22_X1 U2370 ( .A1(n87), .A2(regs[1636]), .B1(n31), .B2(regs[612]), .ZN(
        n1621) );
  OAI211_X1 U2371 ( .C1(n64), .C2(n1623), .A(n1622), .B(n1621), .ZN(
        curr_proc_regs[612]) );
  AOI22_X1 U2372 ( .A1(n103), .A2(regs[101]), .B1(n14), .B2(regs[2149]), .ZN(
        n1625) );
  AOI22_X1 U2373 ( .A1(n53), .A2(regs[1125]), .B1(n98), .B2(regs[1637]), .ZN(
        n1624) );
  OAI211_X1 U2374 ( .C1(n24), .C2(n1626), .A(n1625), .B(n1624), .ZN(
        curr_proc_regs[613]) );
  AOI22_X1 U2375 ( .A1(n103), .A2(regs[102]), .B1(n14), .B2(regs[2150]), .ZN(
        n1628) );
  AOI22_X1 U2376 ( .A1(n52), .A2(regs[1126]), .B1(n98), .B2(regs[1638]), .ZN(
        n1627) );
  OAI211_X1 U2377 ( .C1(n24), .C2(n1629), .A(n1628), .B(n1627), .ZN(
        curr_proc_regs[614]) );
  AOI22_X1 U2378 ( .A1(n103), .A2(regs[103]), .B1(n75), .B2(regs[2151]), .ZN(
        n1631) );
  AOI22_X1 U2379 ( .A1(n54), .A2(regs[1127]), .B1(n98), .B2(regs[1639]), .ZN(
        n1630) );
  OAI211_X1 U2380 ( .C1(n24), .C2(n1632), .A(n1631), .B(n1630), .ZN(
        curr_proc_regs[615]) );
  AOI22_X1 U2381 ( .A1(n103), .A2(regs[104]), .B1(n75), .B2(regs[2152]), .ZN(
        n1634) );
  AOI22_X1 U2382 ( .A1(n53), .A2(regs[1128]), .B1(n84), .B2(regs[1640]), .ZN(
        n1633) );
  OAI211_X1 U2383 ( .C1(n24), .C2(n1635), .A(n1634), .B(n1633), .ZN(
        curr_proc_regs[616]) );
  AOI22_X1 U2384 ( .A1(n106), .A2(regs[105]), .B1(n75), .B2(regs[2153]), .ZN(
        n1637) );
  AOI22_X1 U2385 ( .A1(n52), .A2(regs[1129]), .B1(n83), .B2(regs[1641]), .ZN(
        n1636) );
  OAI211_X1 U2386 ( .C1(n2134), .C2(n1638), .A(n1637), .B(n1636), .ZN(
        curr_proc_regs[617]) );
  AOI22_X1 U2387 ( .A1(n118), .A2(regs[106]), .B1(n75), .B2(regs[2154]), .ZN(
        n1640) );
  AOI22_X1 U2388 ( .A1(n52), .A2(regs[1130]), .B1(n84), .B2(regs[1642]), .ZN(
        n1639) );
  OAI211_X1 U2389 ( .C1(n24), .C2(n1641), .A(n1640), .B(n1639), .ZN(
        curr_proc_regs[618]) );
  AOI22_X1 U2390 ( .A1(n118), .A2(regs[107]), .B1(n75), .B2(regs[2155]), .ZN(
        n1643) );
  AOI22_X1 U2391 ( .A1(n87), .A2(regs[1643]), .B1(n31), .B2(regs[619]), .ZN(
        n1642) );
  OAI211_X1 U2392 ( .C1(n64), .C2(n1644), .A(n1643), .B(n1642), .ZN(
        curr_proc_regs[619]) );
  INV_X1 U2393 ( .A(regs[1085]), .ZN(n1647) );
  AOI22_X1 U2394 ( .A1(n118), .A2(regs[2109]), .B1(n75), .B2(regs[1597]), .ZN(
        n1646) );
  AOI22_X1 U2395 ( .A1(n52), .A2(regs[573]), .B1(n31), .B2(regs[61]), .ZN(
        n1645) );
  OAI211_X1 U2396 ( .C1(n100), .C2(n1647), .A(n1646), .B(n1645), .ZN(
        curr_proc_regs[61]) );
  AOI22_X1 U2397 ( .A1(n118), .A2(regs[108]), .B1(n75), .B2(regs[2156]), .ZN(
        n1649) );
  AOI22_X1 U2398 ( .A1(n52), .A2(regs[1132]), .B1(n85), .B2(regs[1644]), .ZN(
        n1648) );
  OAI211_X1 U2399 ( .C1(n24), .C2(n1650), .A(n1649), .B(n1648), .ZN(
        curr_proc_regs[620]) );
  AOI22_X1 U2400 ( .A1(n118), .A2(regs[109]), .B1(n75), .B2(regs[2157]), .ZN(
        n1652) );
  AOI22_X1 U2401 ( .A1(n87), .A2(regs[1645]), .B1(n31), .B2(regs[621]), .ZN(
        n1651) );
  OAI211_X1 U2402 ( .C1(n11), .C2(n1653), .A(n1652), .B(n1651), .ZN(
        curr_proc_regs[621]) );
  AOI22_X1 U2403 ( .A1(n118), .A2(regs[110]), .B1(n75), .B2(regs[2158]), .ZN(
        n1655) );
  AOI22_X1 U2404 ( .A1(n53), .A2(regs[1134]), .B1(n81), .B2(regs[1646]), .ZN(
        n1654) );
  OAI211_X1 U2405 ( .C1(n24), .C2(n1656), .A(n1655), .B(n1654), .ZN(
        curr_proc_regs[622]) );
  AOI22_X1 U2406 ( .A1(n118), .A2(regs[111]), .B1(n75), .B2(regs[2159]), .ZN(
        n1658) );
  AOI22_X1 U2407 ( .A1(n53), .A2(regs[1135]), .B1(n82), .B2(regs[1647]), .ZN(
        n1657) );
  OAI211_X1 U2408 ( .C1(n24), .C2(n1659), .A(n1658), .B(n1657), .ZN(
        curr_proc_regs[623]) );
  AOI22_X1 U2409 ( .A1(n118), .A2(regs[112]), .B1(n75), .B2(regs[2160]), .ZN(
        n1661) );
  AOI22_X1 U2410 ( .A1(n53), .A2(regs[1136]), .B1(n97), .B2(regs[1648]), .ZN(
        n1660) );
  OAI211_X1 U2411 ( .C1(n24), .C2(n1662), .A(n1661), .B(n1660), .ZN(
        curr_proc_regs[624]) );
  AOI22_X1 U2412 ( .A1(n118), .A2(regs[113]), .B1(n76), .B2(regs[2161]), .ZN(
        n1664) );
  AOI22_X1 U2413 ( .A1(n53), .A2(regs[1137]), .B1(n78), .B2(regs[1649]), .ZN(
        n1663) );
  OAI211_X1 U2414 ( .C1(n24), .C2(n1665), .A(n1664), .B(n1663), .ZN(
        curr_proc_regs[625]) );
  AOI22_X1 U2415 ( .A1(n118), .A2(regs[114]), .B1(n17), .B2(regs[2162]), .ZN(
        n1667) );
  AOI22_X1 U2416 ( .A1(n53), .A2(regs[1138]), .B1(n98), .B2(regs[1650]), .ZN(
        n1666) );
  OAI211_X1 U2417 ( .C1(n24), .C2(n1668), .A(n1667), .B(n1666), .ZN(
        curr_proc_regs[626]) );
  AOI22_X1 U2418 ( .A1(n118), .A2(regs[115]), .B1(n75), .B2(regs[2163]), .ZN(
        n1670) );
  AOI22_X1 U2419 ( .A1(n53), .A2(regs[1139]), .B1(n81), .B2(regs[1651]), .ZN(
        n1669) );
  OAI211_X1 U2420 ( .C1(n24), .C2(n1671), .A(n1670), .B(n1669), .ZN(
        curr_proc_regs[627]) );
  AOI22_X1 U2421 ( .A1(n115), .A2(regs[116]), .B1(n76), .B2(regs[2164]), .ZN(
        n1673) );
  AOI22_X1 U2422 ( .A1(n53), .A2(regs[1140]), .B1(n85), .B2(regs[1652]), .ZN(
        n1672) );
  OAI211_X1 U2423 ( .C1(n24), .C2(n1674), .A(n1673), .B(n1672), .ZN(
        curr_proc_regs[628]) );
  AOI22_X1 U2424 ( .A1(n116), .A2(regs[117]), .B1(n17), .B2(regs[2165]), .ZN(
        n1676) );
  AOI22_X1 U2425 ( .A1(n53), .A2(regs[1141]), .B1(n86), .B2(regs[1653]), .ZN(
        n1675) );
  OAI211_X1 U2426 ( .C1(n24), .C2(n1677), .A(n1676), .B(n1675), .ZN(
        curr_proc_regs[629]) );
  INV_X1 U2427 ( .A(regs[1086]), .ZN(n1680) );
  AOI22_X1 U2428 ( .A1(n117), .A2(regs[2110]), .B1(n75), .B2(regs[1598]), .ZN(
        n1679) );
  AOI22_X1 U2429 ( .A1(n51), .A2(regs[574]), .B1(n31), .B2(regs[62]), .ZN(
        n1678) );
  OAI211_X1 U2430 ( .C1(n100), .C2(n1680), .A(n1679), .B(n1678), .ZN(
        curr_proc_regs[62]) );
  AOI22_X1 U2431 ( .A1(n117), .A2(regs[118]), .B1(n76), .B2(regs[2166]), .ZN(
        n1682) );
  AOI22_X1 U2432 ( .A1(n51), .A2(regs[1142]), .B1(n80), .B2(regs[1654]), .ZN(
        n1681) );
  OAI211_X1 U2433 ( .C1(n24), .C2(n1683), .A(n1682), .B(n1681), .ZN(
        curr_proc_regs[630]) );
  AOI22_X1 U2434 ( .A1(n116), .A2(regs[119]), .B1(n17), .B2(regs[2167]), .ZN(
        n1685) );
  AOI22_X1 U2435 ( .A1(n87), .A2(regs[1655]), .B1(n31), .B2(regs[631]), .ZN(
        n1684) );
  OAI211_X1 U2436 ( .C1(n2207), .C2(n1686), .A(n1685), .B(n1684), .ZN(
        curr_proc_regs[631]) );
  AOI22_X1 U2437 ( .A1(n115), .A2(regs[120]), .B1(n75), .B2(regs[2168]), .ZN(
        n1688) );
  AOI22_X1 U2438 ( .A1(n87), .A2(regs[1656]), .B1(n31), .B2(regs[632]), .ZN(
        n1687) );
  OAI211_X1 U2439 ( .C1(n11), .C2(n1689), .A(n1688), .B(n1687), .ZN(
        curr_proc_regs[632]) );
  AOI22_X1 U2440 ( .A1(n116), .A2(regs[121]), .B1(n76), .B2(regs[2169]), .ZN(
        n1691) );
  AOI22_X1 U2441 ( .A1(n51), .A2(regs[1145]), .B1(n86), .B2(regs[1657]), .ZN(
        n1690) );
  OAI211_X1 U2442 ( .C1(n24), .C2(n1692), .A(n1691), .B(n1690), .ZN(
        curr_proc_regs[633]) );
  AOI22_X1 U2443 ( .A1(n117), .A2(regs[122]), .B1(n17), .B2(regs[2170]), .ZN(
        n1694) );
  AOI22_X1 U2444 ( .A1(n87), .A2(regs[1658]), .B1(n31), .B2(regs[634]), .ZN(
        n1693) );
  OAI211_X1 U2445 ( .C1(n2207), .C2(n1695), .A(n1694), .B(n1693), .ZN(
        curr_proc_regs[634]) );
  AOI22_X1 U2446 ( .A1(n115), .A2(regs[123]), .B1(n76), .B2(regs[2171]), .ZN(
        n1697) );
  AOI22_X1 U2447 ( .A1(n52), .A2(regs[1147]), .B1(n87), .B2(regs[1659]), .ZN(
        n1696) );
  OAI211_X1 U2448 ( .C1(n24), .C2(n1698), .A(n1697), .B(n1696), .ZN(
        curr_proc_regs[635]) );
  AOI22_X1 U2449 ( .A1(n117), .A2(regs[124]), .B1(n76), .B2(regs[2172]), .ZN(
        n1700) );
  AOI22_X1 U2450 ( .A1(n87), .A2(regs[1660]), .B1(n31), .B2(regs[636]), .ZN(
        n1699) );
  OAI211_X1 U2451 ( .C1(n11), .C2(n1701), .A(n1700), .B(n1699), .ZN(
        curr_proc_regs[636]) );
  AOI22_X1 U2452 ( .A1(n115), .A2(regs[125]), .B1(n76), .B2(regs[2173]), .ZN(
        n1703) );
  AOI22_X1 U2453 ( .A1(n87), .A2(regs[1661]), .B1(n12), .B2(regs[637]), .ZN(
        n1702) );
  OAI211_X1 U2454 ( .C1(n2207), .C2(n1704), .A(n1703), .B(n1702), .ZN(
        curr_proc_regs[637]) );
  AOI22_X1 U2455 ( .A1(n116), .A2(regs[126]), .B1(n76), .B2(regs[2174]), .ZN(
        n1706) );
  AOI22_X1 U2456 ( .A1(n87), .A2(regs[1662]), .B1(n12), .B2(regs[638]), .ZN(
        n1705) );
  OAI211_X1 U2457 ( .C1(n11), .C2(n1707), .A(n1706), .B(n1705), .ZN(
        curr_proc_regs[638]) );
  AOI22_X1 U2458 ( .A1(n115), .A2(regs[127]), .B1(n76), .B2(regs[2175]), .ZN(
        n1709) );
  AOI22_X1 U2459 ( .A1(n87), .A2(regs[1663]), .B1(n12), .B2(regs[639]), .ZN(
        n1708) );
  OAI211_X1 U2460 ( .C1(n11), .C2(n1710), .A(n1709), .B(n1708), .ZN(
        curr_proc_regs[639]) );
  INV_X1 U2461 ( .A(regs[1087]), .ZN(n1713) );
  AOI22_X1 U2462 ( .A1(n116), .A2(regs[2111]), .B1(n76), .B2(regs[1599]), .ZN(
        n1712) );
  AOI22_X1 U2463 ( .A1(n52), .A2(regs[575]), .B1(n12), .B2(regs[63]), .ZN(
        n1711) );
  OAI211_X1 U2464 ( .C1(n100), .C2(n1713), .A(n1712), .B(n1711), .ZN(
        curr_proc_regs[63]) );
  AOI22_X1 U2465 ( .A1(n117), .A2(regs[128]), .B1(n76), .B2(regs[2176]), .ZN(
        n1715) );
  AOI22_X1 U2466 ( .A1(n87), .A2(regs[1664]), .B1(n12), .B2(regs[640]), .ZN(
        n1714) );
  OAI211_X1 U2467 ( .C1(n11), .C2(n1716), .A(n1715), .B(n1714), .ZN(
        curr_proc_regs[640]) );
  AOI22_X1 U2468 ( .A1(n117), .A2(regs[129]), .B1(n76), .B2(regs[2177]), .ZN(
        n1718) );
  AOI22_X1 U2469 ( .A1(n52), .A2(regs[1153]), .B1(n81), .B2(regs[1665]), .ZN(
        n1717) );
  OAI211_X1 U2470 ( .C1(n24), .C2(n1719), .A(n1718), .B(n1717), .ZN(
        curr_proc_regs[641]) );
  AOI22_X1 U2471 ( .A1(n115), .A2(regs[130]), .B1(n76), .B2(regs[2178]), .ZN(
        n1721) );
  AOI22_X1 U2472 ( .A1(n86), .A2(regs[1666]), .B1(n12), .B2(regs[642]), .ZN(
        n1720) );
  OAI211_X1 U2473 ( .C1(n11), .C2(n1722), .A(n1721), .B(n1720), .ZN(
        curr_proc_regs[642]) );
  AOI22_X1 U2474 ( .A1(n116), .A2(regs[131]), .B1(n76), .B2(regs[2179]), .ZN(
        n1724) );
  AOI22_X1 U2475 ( .A1(n86), .A2(regs[1667]), .B1(n12), .B2(regs[643]), .ZN(
        n1723) );
  OAI211_X1 U2476 ( .C1(n11), .C2(n1725), .A(n1724), .B(n1723), .ZN(
        curr_proc_regs[643]) );
  AOI22_X1 U2477 ( .A1(n117), .A2(regs[132]), .B1(n76), .B2(regs[2180]), .ZN(
        n1727) );
  AOI22_X1 U2478 ( .A1(n86), .A2(regs[1668]), .B1(n12), .B2(regs[644]), .ZN(
        n1726) );
  OAI211_X1 U2479 ( .C1(n11), .C2(n1728), .A(n1727), .B(n1726), .ZN(
        curr_proc_regs[644]) );
  AOI22_X1 U2480 ( .A1(n115), .A2(regs[133]), .B1(n17), .B2(regs[2181]), .ZN(
        n1730) );
  AOI22_X1 U2481 ( .A1(n86), .A2(regs[1669]), .B1(n12), .B2(regs[645]), .ZN(
        n1729) );
  OAI211_X1 U2482 ( .C1(n11), .C2(n1731), .A(n1730), .B(n1729), .ZN(
        curr_proc_regs[645]) );
  AOI22_X1 U2483 ( .A1(n115), .A2(regs[134]), .B1(n75), .B2(regs[2182]), .ZN(
        n1733) );
  AOI22_X1 U2484 ( .A1(n86), .A2(regs[1670]), .B1(n12), .B2(regs[646]), .ZN(
        n1732) );
  OAI211_X1 U2485 ( .C1(n11), .C2(n1734), .A(n1733), .B(n1732), .ZN(
        curr_proc_regs[646]) );
  AOI22_X1 U2486 ( .A1(n116), .A2(regs[135]), .B1(n75), .B2(regs[2183]), .ZN(
        n1736) );
  AOI22_X1 U2487 ( .A1(n52), .A2(regs[1159]), .B1(n83), .B2(regs[1671]), .ZN(
        n1735) );
  OAI211_X1 U2488 ( .C1(n24), .C2(n1737), .A(n1736), .B(n1735), .ZN(
        curr_proc_regs[647]) );
  AOI22_X1 U2489 ( .A1(n116), .A2(regs[136]), .B1(n76), .B2(regs[2184]), .ZN(
        n1739) );
  AOI22_X1 U2490 ( .A1(n52), .A2(regs[1160]), .B1(n84), .B2(regs[1672]), .ZN(
        n1738) );
  OAI211_X1 U2491 ( .C1(n24), .C2(n1740), .A(n1739), .B(n1738), .ZN(
        curr_proc_regs[648]) );
  AOI22_X1 U2492 ( .A1(n117), .A2(regs[137]), .B1(n17), .B2(regs[2185]), .ZN(
        n1742) );
  AOI22_X1 U2493 ( .A1(n86), .A2(regs[1673]), .B1(n12), .B2(regs[649]), .ZN(
        n1741) );
  OAI211_X1 U2494 ( .C1(n64), .C2(n1743), .A(n1742), .B(n1741), .ZN(
        curr_proc_regs[649]) );
  AOI22_X1 U2495 ( .A1(n115), .A2(regs[2112]), .B1(n76), .B2(regs[1600]), .ZN(
        n1745) );
  AOI22_X1 U2496 ( .A1(n52), .A2(regs[576]), .B1(n12), .B2(regs[64]), .ZN(
        n1744) );
  OAI211_X1 U2497 ( .C1(n100), .C2(n1746), .A(n1745), .B(n1744), .ZN(
        curr_proc_regs[64]) );
  AOI22_X1 U2498 ( .A1(n116), .A2(regs[138]), .B1(n75), .B2(regs[2186]), .ZN(
        n1748) );
  AOI22_X1 U2499 ( .A1(n52), .A2(regs[1162]), .B1(n81), .B2(regs[1674]), .ZN(
        n1747) );
  OAI211_X1 U2500 ( .C1(n25), .C2(n1749), .A(n1748), .B(n1747), .ZN(
        curr_proc_regs[650]) );
  AOI22_X1 U2501 ( .A1(n117), .A2(regs[139]), .B1(n76), .B2(regs[2187]), .ZN(
        n1751) );
  AOI22_X1 U2502 ( .A1(n86), .A2(regs[1675]), .B1(n12), .B2(regs[651]), .ZN(
        n1750) );
  OAI211_X1 U2503 ( .C1(n2207), .C2(n1752), .A(n1751), .B(n1750), .ZN(
        curr_proc_regs[651]) );
  AOI22_X1 U2504 ( .A1(n115), .A2(regs[140]), .B1(n17), .B2(regs[2188]), .ZN(
        n1754) );
  AOI22_X1 U2505 ( .A1(n52), .A2(regs[1164]), .B1(n82), .B2(regs[1676]), .ZN(
        n1753) );
  OAI211_X1 U2506 ( .C1(n25), .C2(n1755), .A(n1754), .B(n1753), .ZN(
        curr_proc_regs[652]) );
  AOI22_X1 U2507 ( .A1(n116), .A2(regs[141]), .B1(n17), .B2(regs[2189]), .ZN(
        n1757) );
  AOI22_X1 U2508 ( .A1(n86), .A2(regs[1677]), .B1(n12), .B2(regs[653]), .ZN(
        n1756) );
  OAI211_X1 U2509 ( .C1(n64), .C2(n1758), .A(n1757), .B(n1756), .ZN(
        curr_proc_regs[653]) );
  AOI22_X1 U2510 ( .A1(n117), .A2(regs[142]), .B1(n75), .B2(regs[2190]), .ZN(
        n1760) );
  AOI22_X1 U2511 ( .A1(n8), .A2(regs[1166]), .B1(n87), .B2(regs[1678]), .ZN(
        n1759) );
  OAI211_X1 U2512 ( .C1(n25), .C2(n1761), .A(n1760), .B(n1759), .ZN(
        curr_proc_regs[654]) );
  AOI22_X1 U2513 ( .A1(n115), .A2(regs[143]), .B1(n76), .B2(regs[2191]), .ZN(
        n1763) );
  AOI22_X1 U2514 ( .A1(n86), .A2(regs[1679]), .B1(n12), .B2(regs[655]), .ZN(
        n1762) );
  OAI211_X1 U2515 ( .C1(n2207), .C2(n1764), .A(n1763), .B(n1762), .ZN(
        curr_proc_regs[655]) );
  AOI22_X1 U2516 ( .A1(n116), .A2(regs[144]), .B1(n75), .B2(regs[2192]), .ZN(
        n1766) );
  AOI22_X1 U2517 ( .A1(n86), .A2(regs[1680]), .B1(n12), .B2(regs[656]), .ZN(
        n1765) );
  OAI211_X1 U2518 ( .C1(n64), .C2(n1767), .A(n1766), .B(n1765), .ZN(
        curr_proc_regs[656]) );
  AOI22_X1 U2519 ( .A1(n117), .A2(regs[145]), .B1(n75), .B2(regs[2193]), .ZN(
        n1769) );
  AOI22_X1 U2520 ( .A1(n13), .A2(regs[1169]), .B1(n98), .B2(regs[1681]), .ZN(
        n1768) );
  OAI211_X1 U2521 ( .C1(n25), .C2(n1770), .A(n1769), .B(n1768), .ZN(
        curr_proc_regs[657]) );
  AOI22_X1 U2522 ( .A1(n117), .A2(regs[146]), .B1(n76), .B2(regs[2194]), .ZN(
        n1772) );
  AOI22_X1 U2523 ( .A1(n86), .A2(regs[1682]), .B1(n12), .B2(regs[658]), .ZN(
        n1771) );
  OAI211_X1 U2524 ( .C1(n64), .C2(n1773), .A(n1772), .B(n1771), .ZN(
        curr_proc_regs[658]) );
  AOI22_X1 U2525 ( .A1(n117), .A2(regs[147]), .B1(n17), .B2(regs[2195]), .ZN(
        n1775) );
  AOI22_X1 U2526 ( .A1(n85), .A2(regs[1683]), .B1(n12), .B2(regs[659]), .ZN(
        n1774) );
  OAI211_X1 U2527 ( .C1(n64), .C2(n1776), .A(n1775), .B(n1774), .ZN(
        curr_proc_regs[659]) );
  INV_X1 U2528 ( .A(regs[577]), .ZN(n1779) );
  AOI22_X1 U2529 ( .A1(n117), .A2(regs[2113]), .B1(n17), .B2(regs[1601]), .ZN(
        n1778) );
  AOI22_X1 U2530 ( .A1(n85), .A2(regs[1089]), .B1(n12), .B2(regs[65]), .ZN(
        n1777) );
  OAI211_X1 U2531 ( .C1(n11), .C2(n1779), .A(n1778), .B(n1777), .ZN(
        curr_proc_regs[65]) );
  AOI22_X1 U2532 ( .A1(n117), .A2(regs[148]), .B1(n76), .B2(regs[2196]), .ZN(
        n1781) );
  AOI22_X1 U2533 ( .A1(n2), .A2(regs[1172]), .B1(n85), .B2(regs[1684]), .ZN(
        n1780) );
  OAI211_X1 U2534 ( .C1(n25), .C2(n1782), .A(n1781), .B(n1780), .ZN(
        curr_proc_regs[660]) );
  AOI22_X1 U2535 ( .A1(n117), .A2(regs[149]), .B1(n75), .B2(regs[2197]), .ZN(
        n1784) );
  AOI22_X1 U2536 ( .A1(n85), .A2(regs[1685]), .B1(n12), .B2(regs[661]), .ZN(
        n1783) );
  OAI211_X1 U2537 ( .C1(n11), .C2(n1785), .A(n1784), .B(n1783), .ZN(
        curr_proc_regs[661]) );
  AOI22_X1 U2538 ( .A1(n117), .A2(regs[150]), .B1(n17), .B2(regs[2198]), .ZN(
        n1787) );
  AOI22_X1 U2539 ( .A1(n85), .A2(regs[1686]), .B1(n12), .B2(regs[662]), .ZN(
        n1786) );
  OAI211_X1 U2540 ( .C1(n11), .C2(n1788), .A(n1787), .B(n1786), .ZN(
        curr_proc_regs[662]) );
  AOI22_X1 U2541 ( .A1(n117), .A2(regs[151]), .B1(n17), .B2(regs[2199]), .ZN(
        n1790) );
  AOI22_X1 U2542 ( .A1(n85), .A2(regs[1687]), .B1(n12), .B2(regs[663]), .ZN(
        n1789) );
  OAI211_X1 U2543 ( .C1(n11), .C2(n1791), .A(n1790), .B(n1789), .ZN(
        curr_proc_regs[663]) );
  AOI22_X1 U2544 ( .A1(n117), .A2(regs[152]), .B1(n17), .B2(regs[2200]), .ZN(
        n1793) );
  AOI22_X1 U2545 ( .A1(n10), .A2(regs[1176]), .B1(n85), .B2(regs[1688]), .ZN(
        n1792) );
  OAI211_X1 U2546 ( .C1(n25), .C2(n1794), .A(n1793), .B(n1792), .ZN(
        curr_proc_regs[664]) );
  AOI22_X1 U2547 ( .A1(n117), .A2(regs[153]), .B1(n76), .B2(regs[2201]), .ZN(
        n1796) );
  AOI22_X1 U2548 ( .A1(n8), .A2(regs[1177]), .B1(n78), .B2(regs[1689]), .ZN(
        n1795) );
  OAI211_X1 U2549 ( .C1(n2134), .C2(n1797), .A(n1796), .B(n1795), .ZN(
        curr_proc_regs[665]) );
  AOI22_X1 U2550 ( .A1(n117), .A2(regs[154]), .B1(n17), .B2(regs[2202]), .ZN(
        n1799) );
  AOI22_X1 U2551 ( .A1(n13), .A2(regs[1178]), .B1(n79), .B2(regs[1690]), .ZN(
        n1798) );
  OAI211_X1 U2552 ( .C1(n25), .C2(n1800), .A(n1799), .B(n1798), .ZN(
        curr_proc_regs[666]) );
  AOI22_X1 U2553 ( .A1(n117), .A2(regs[155]), .B1(n17), .B2(regs[2203]), .ZN(
        n1802) );
  AOI22_X1 U2554 ( .A1(n2), .A2(regs[1179]), .B1(n80), .B2(regs[1691]), .ZN(
        n1801) );
  OAI211_X1 U2555 ( .C1(n24), .C2(n1803), .A(n1802), .B(n1801), .ZN(
        curr_proc_regs[667]) );
  AOI22_X1 U2556 ( .A1(n116), .A2(regs[156]), .B1(n17), .B2(regs[2204]), .ZN(
        n1805) );
  AOI22_X1 U2557 ( .A1(n10), .A2(regs[1180]), .B1(n86), .B2(regs[1692]), .ZN(
        n1804) );
  OAI211_X1 U2558 ( .C1(n2134), .C2(n1806), .A(n1805), .B(n1804), .ZN(
        curr_proc_regs[668]) );
  AOI22_X1 U2559 ( .A1(n116), .A2(regs[157]), .B1(n17), .B2(regs[2205]), .ZN(
        n1808) );
  AOI22_X1 U2560 ( .A1(n8), .A2(regs[1181]), .B1(n87), .B2(regs[1693]), .ZN(
        n1807) );
  OAI211_X1 U2561 ( .C1(n25), .C2(n1809), .A(n1808), .B(n1807), .ZN(
        curr_proc_regs[669]) );
  AOI22_X1 U2562 ( .A1(n116), .A2(regs[2114]), .B1(n75), .B2(regs[1602]), .ZN(
        n1811) );
  AOI22_X1 U2563 ( .A1(n13), .A2(regs[578]), .B1(n26), .B2(regs[66]), .ZN(
        n1810) );
  OAI211_X1 U2564 ( .C1(n100), .C2(n1812), .A(n1811), .B(n1810), .ZN(
        curr_proc_regs[66]) );
  AOI22_X1 U2565 ( .A1(n116), .A2(regs[158]), .B1(n76), .B2(regs[2206]), .ZN(
        n1814) );
  AOI22_X1 U2566 ( .A1(n85), .A2(regs[1694]), .B1(n26), .B2(regs[670]), .ZN(
        n1813) );
  OAI211_X1 U2567 ( .C1(n11), .C2(n1815), .A(n1814), .B(n1813), .ZN(
        curr_proc_regs[670]) );
  AOI22_X1 U2568 ( .A1(n116), .A2(regs[159]), .B1(n17), .B2(regs[2207]), .ZN(
        n1817) );
  AOI22_X1 U2569 ( .A1(n85), .A2(regs[1695]), .B1(n44), .B2(regs[671]), .ZN(
        n1816) );
  OAI211_X1 U2570 ( .C1(n11), .C2(n1818), .A(n1817), .B(n1816), .ZN(
        curr_proc_regs[671]) );
  AOI22_X1 U2571 ( .A1(n116), .A2(regs[160]), .B1(n17), .B2(regs[2208]), .ZN(
        n1820) );
  AOI22_X1 U2572 ( .A1(n85), .A2(regs[1696]), .B1(n44), .B2(regs[672]), .ZN(
        n1819) );
  OAI211_X1 U2573 ( .C1(n11), .C2(n1821), .A(n1820), .B(n1819), .ZN(
        curr_proc_regs[672]) );
  AOI22_X1 U2574 ( .A1(n116), .A2(regs[161]), .B1(n17), .B2(regs[2209]), .ZN(
        n1823) );
  AOI22_X1 U2575 ( .A1(n56), .A2(regs[1185]), .B1(n82), .B2(regs[1697]), .ZN(
        n1822) );
  OAI211_X1 U2576 ( .C1(n24), .C2(n1824), .A(n1823), .B(n1822), .ZN(
        curr_proc_regs[673]) );
  AOI22_X1 U2577 ( .A1(n116), .A2(regs[162]), .B1(n17), .B2(regs[2210]), .ZN(
        n1826) );
  AOI22_X1 U2578 ( .A1(n85), .A2(regs[1698]), .B1(n45), .B2(regs[674]), .ZN(
        n1825) );
  OAI211_X1 U2579 ( .C1(n65), .C2(n1827), .A(n1826), .B(n1825), .ZN(
        curr_proc_regs[674]) );
  AOI22_X1 U2580 ( .A1(n116), .A2(regs[163]), .B1(n72), .B2(regs[2211]), .ZN(
        n1829) );
  AOI22_X1 U2581 ( .A1(n85), .A2(regs[1699]), .B1(n44), .B2(regs[675]), .ZN(
        n1828) );
  OAI211_X1 U2582 ( .C1(n65), .C2(n1830), .A(n1829), .B(n1828), .ZN(
        curr_proc_regs[675]) );
  AOI22_X1 U2583 ( .A1(n116), .A2(regs[164]), .B1(n73), .B2(regs[2212]), .ZN(
        n1832) );
  AOI22_X1 U2584 ( .A1(n56), .A2(regs[1188]), .B1(n86), .B2(regs[1700]), .ZN(
        n1831) );
  OAI211_X1 U2585 ( .C1(n2134), .C2(n1833), .A(n1832), .B(n1831), .ZN(
        curr_proc_regs[676]) );
  AOI22_X1 U2586 ( .A1(n116), .A2(regs[165]), .B1(n2217), .B2(regs[2213]), 
        .ZN(n1835) );
  AOI22_X1 U2587 ( .A1(n85), .A2(regs[1701]), .B1(n45), .B2(regs[677]), .ZN(
        n1834) );
  OAI211_X1 U2588 ( .C1(n65), .C2(n1836), .A(n1835), .B(n1834), .ZN(
        curr_proc_regs[677]) );
  AOI22_X1 U2589 ( .A1(n115), .A2(regs[166]), .B1(n2217), .B2(regs[2214]), 
        .ZN(n1838) );
  AOI22_X1 U2590 ( .A1(n10), .A2(regs[1190]), .B1(n79), .B2(regs[1702]), .ZN(
        n1837) );
  OAI211_X1 U2591 ( .C1(n25), .C2(n1839), .A(n1838), .B(n1837), .ZN(
        curr_proc_regs[678]) );
  AOI22_X1 U2592 ( .A1(n115), .A2(regs[167]), .B1(n72), .B2(regs[2215]), .ZN(
        n1841) );
  AOI22_X1 U2593 ( .A1(n49), .A2(regs[1191]), .B1(n98), .B2(regs[1703]), .ZN(
        n1840) );
  OAI211_X1 U2594 ( .C1(n25), .C2(n1842), .A(n1841), .B(n1840), .ZN(
        curr_proc_regs[679]) );
  INV_X1 U2595 ( .A(regs[579]), .ZN(n1845) );
  AOI22_X1 U2596 ( .A1(n115), .A2(regs[2115]), .B1(n73), .B2(regs[1603]), .ZN(
        n1844) );
  AOI22_X1 U2597 ( .A1(n84), .A2(regs[1091]), .B1(n27), .B2(regs[67]), .ZN(
        n1843) );
  OAI211_X1 U2598 ( .C1(n65), .C2(n1845), .A(n1844), .B(n1843), .ZN(
        curr_proc_regs[67]) );
  AOI22_X1 U2599 ( .A1(n115), .A2(regs[168]), .B1(n9), .B2(regs[2216]), .ZN(
        n1847) );
  AOI22_X1 U2600 ( .A1(n10), .A2(regs[1192]), .B1(n84), .B2(regs[1704]), .ZN(
        n1846) );
  OAI211_X1 U2601 ( .C1(n25), .C2(n1848), .A(n1847), .B(n1846), .ZN(
        curr_proc_regs[680]) );
  AOI22_X1 U2602 ( .A1(n115), .A2(regs[169]), .B1(n9), .B2(regs[2217]), .ZN(
        n1850) );
  AOI22_X1 U2603 ( .A1(n84), .A2(regs[1705]), .B1(n26), .B2(regs[681]), .ZN(
        n1849) );
  OAI211_X1 U2604 ( .C1(n65), .C2(n1851), .A(n1850), .B(n1849), .ZN(
        curr_proc_regs[681]) );
  AOI22_X1 U2605 ( .A1(n115), .A2(regs[170]), .B1(n9), .B2(regs[2218]), .ZN(
        n1853) );
  AOI22_X1 U2606 ( .A1(n84), .A2(regs[1706]), .B1(n44), .B2(regs[682]), .ZN(
        n1852) );
  OAI211_X1 U2607 ( .C1(n65), .C2(n1854), .A(n1853), .B(n1852), .ZN(
        curr_proc_regs[682]) );
  AOI22_X1 U2608 ( .A1(n115), .A2(regs[171]), .B1(n9), .B2(regs[2219]), .ZN(
        n1856) );
  AOI22_X1 U2609 ( .A1(n84), .A2(regs[1707]), .B1(n48), .B2(regs[683]), .ZN(
        n1855) );
  OAI211_X1 U2610 ( .C1(n65), .C2(n1857), .A(n1856), .B(n1855), .ZN(
        curr_proc_regs[683]) );
  AOI22_X1 U2611 ( .A1(n115), .A2(regs[172]), .B1(n9), .B2(regs[2220]), .ZN(
        n1859) );
  AOI22_X1 U2612 ( .A1(n84), .A2(regs[1708]), .B1(n3), .B2(regs[684]), .ZN(
        n1858) );
  OAI211_X1 U2613 ( .C1(n65), .C2(n1860), .A(n1859), .B(n1858), .ZN(
        curr_proc_regs[684]) );
  AOI22_X1 U2614 ( .A1(n115), .A2(regs[173]), .B1(n9), .B2(regs[2221]), .ZN(
        n1862) );
  AOI22_X1 U2615 ( .A1(n84), .A2(regs[1709]), .B1(n3), .B2(regs[685]), .ZN(
        n1861) );
  OAI211_X1 U2616 ( .C1(n65), .C2(n1863), .A(n1862), .B(n1861), .ZN(
        curr_proc_regs[685]) );
  AOI22_X1 U2617 ( .A1(n115), .A2(regs[174]), .B1(n9), .B2(regs[2222]), .ZN(
        n1865) );
  AOI22_X1 U2618 ( .A1(n10), .A2(regs[1198]), .B1(n97), .B2(regs[1710]), .ZN(
        n1864) );
  OAI211_X1 U2619 ( .C1(n25), .C2(n1866), .A(n1865), .B(n1864), .ZN(
        curr_proc_regs[686]) );
  AOI22_X1 U2620 ( .A1(n115), .A2(regs[175]), .B1(n4), .B2(regs[2223]), .ZN(
        n1868) );
  AOI22_X1 U2621 ( .A1(n56), .A2(regs[1199]), .B1(n19), .B2(regs[1711]), .ZN(
        n1867) );
  OAI211_X1 U2622 ( .C1(n25), .C2(n1869), .A(n1868), .B(n1867), .ZN(
        curr_proc_regs[687]) );
  AOI22_X1 U2623 ( .A1(n6), .A2(regs[176]), .B1(n9), .B2(regs[2224]), .ZN(
        n1871) );
  AOI22_X1 U2624 ( .A1(n84), .A2(regs[1712]), .B1(n3), .B2(regs[688]), .ZN(
        n1870) );
  OAI211_X1 U2625 ( .C1(n1), .C2(n1872), .A(n1871), .B(n1870), .ZN(
        curr_proc_regs[688]) );
  AOI22_X1 U2626 ( .A1(n113), .A2(regs[177]), .B1(n9), .B2(regs[2225]), .ZN(
        n1874) );
  AOI22_X1 U2627 ( .A1(n10), .A2(regs[1201]), .B1(n19), .B2(regs[1713]), .ZN(
        n1873) );
  OAI211_X1 U2628 ( .C1(n25), .C2(n1875), .A(n1874), .B(n1873), .ZN(
        curr_proc_regs[689]) );
  INV_X1 U2629 ( .A(regs[580]), .ZN(n1878) );
  AOI22_X1 U2630 ( .A1(n114), .A2(regs[2116]), .B1(n67), .B2(regs[1604]), .ZN(
        n1877) );
  AOI22_X1 U2631 ( .A1(n84), .A2(regs[1092]), .B1(n3), .B2(regs[68]), .ZN(
        n1876) );
  OAI211_X1 U2632 ( .C1(n1), .C2(n1878), .A(n1877), .B(n1876), .ZN(
        curr_proc_regs[68]) );
  AOI22_X1 U2633 ( .A1(n114), .A2(regs[178]), .B1(n9), .B2(regs[2226]), .ZN(
        n1880) );
  AOI22_X1 U2634 ( .A1(n84), .A2(regs[1714]), .B1(n3), .B2(regs[690]), .ZN(
        n1879) );
  OAI211_X1 U2635 ( .C1(n65), .C2(n1881), .A(n1880), .B(n1879), .ZN(
        curr_proc_regs[690]) );
  AOI22_X1 U2636 ( .A1(n113), .A2(regs[179]), .B1(n9), .B2(regs[2227]), .ZN(
        n1883) );
  AOI22_X1 U2637 ( .A1(n56), .A2(regs[1203]), .B1(n19), .B2(regs[1715]), .ZN(
        n1882) );
  OAI211_X1 U2638 ( .C1(n25), .C2(n1884), .A(n1883), .B(n1882), .ZN(
        curr_proc_regs[691]) );
  AOI22_X1 U2639 ( .A1(n6), .A2(regs[180]), .B1(n73), .B2(regs[2228]), .ZN(
        n1886) );
  AOI22_X1 U2640 ( .A1(n49), .A2(regs[1204]), .B1(n19), .B2(regs[1716]), .ZN(
        n1885) );
  OAI211_X1 U2641 ( .C1(n25), .C2(n1887), .A(n1886), .B(n1885), .ZN(
        curr_proc_regs[692]) );
  AOI22_X1 U2642 ( .A1(n113), .A2(regs[181]), .B1(n9), .B2(regs[2229]), .ZN(
        n1889) );
  AOI22_X1 U2643 ( .A1(n10), .A2(regs[1205]), .B1(n97), .B2(regs[1717]), .ZN(
        n1888) );
  OAI211_X1 U2644 ( .C1(n25), .C2(n1890), .A(n1889), .B(n1888), .ZN(
        curr_proc_regs[693]) );
  AOI22_X1 U2645 ( .A1(n114), .A2(regs[182]), .B1(n9), .B2(regs[2230]), .ZN(
        n1892) );
  AOI22_X1 U2646 ( .A1(n10), .A2(regs[1206]), .B1(n19), .B2(regs[1718]), .ZN(
        n1891) );
  OAI211_X1 U2647 ( .C1(n25), .C2(n1893), .A(n1892), .B(n1891), .ZN(
        curr_proc_regs[694]) );
  AOI22_X1 U2648 ( .A1(n6), .A2(regs[183]), .B1(n9), .B2(regs[2231]), .ZN(
        n1895) );
  AOI22_X1 U2649 ( .A1(n56), .A2(regs[1207]), .B1(n97), .B2(regs[1719]), .ZN(
        n1894) );
  OAI211_X1 U2650 ( .C1(n25), .C2(n1896), .A(n1895), .B(n1894), .ZN(
        curr_proc_regs[695]) );
  AOI22_X1 U2651 ( .A1(n114), .A2(regs[184]), .B1(n9), .B2(regs[2232]), .ZN(
        n1898) );
  AOI22_X1 U2652 ( .A1(n56), .A2(regs[1208]), .B1(n19), .B2(regs[1720]), .ZN(
        n1897) );
  OAI211_X1 U2653 ( .C1(n25), .C2(n1899), .A(n1898), .B(n1897), .ZN(
        curr_proc_regs[696]) );
  AOI22_X1 U2654 ( .A1(n6), .A2(regs[185]), .B1(n9), .B2(regs[2233]), .ZN(
        n1901) );
  AOI22_X1 U2655 ( .A1(n56), .A2(regs[1209]), .B1(n19), .B2(regs[1721]), .ZN(
        n1900) );
  OAI211_X1 U2656 ( .C1(n25), .C2(n1902), .A(n1901), .B(n1900), .ZN(
        curr_proc_regs[697]) );
  AOI22_X1 U2657 ( .A1(n6), .A2(regs[186]), .B1(n9), .B2(regs[2234]), .ZN(
        n1904) );
  AOI22_X1 U2658 ( .A1(n84), .A2(regs[1722]), .B1(n3), .B2(regs[698]), .ZN(
        n1903) );
  OAI211_X1 U2659 ( .C1(n65), .C2(n1905), .A(n1904), .B(n1903), .ZN(
        curr_proc_regs[698]) );
  AOI22_X1 U2660 ( .A1(n6), .A2(regs[187]), .B1(n9), .B2(regs[2235]), .ZN(
        n1907) );
  AOI22_X1 U2661 ( .A1(n79), .A2(regs[1723]), .B1(n3), .B2(regs[699]), .ZN(
        n1906) );
  OAI211_X1 U2662 ( .C1(n1), .C2(n1908), .A(n1907), .B(n1906), .ZN(
        curr_proc_regs[699]) );
  INV_X1 U2663 ( .A(regs[581]), .ZN(n1911) );
  AOI22_X1 U2664 ( .A1(n6), .A2(regs[2117]), .B1(n9), .B2(regs[1605]), .ZN(
        n1910) );
  AOI22_X1 U2665 ( .A1(n83), .A2(regs[1093]), .B1(n3), .B2(regs[69]), .ZN(
        n1909) );
  OAI211_X1 U2666 ( .C1(n65), .C2(n1911), .A(n1910), .B(n1909), .ZN(
        curr_proc_regs[69]) );
  AOI22_X1 U2667 ( .A1(n6), .A2(regs[2054]), .B1(n9), .B2(regs[1542]), .ZN(
        n1913) );
  AOI22_X1 U2668 ( .A1(n56), .A2(regs[518]), .B1(n3), .B2(regs[6]), .ZN(n1912)
         );
  OAI211_X1 U2669 ( .C1(n100), .C2(n1914), .A(n1913), .B(n1912), .ZN(
        curr_proc_regs[6]) );
  AOI22_X1 U2670 ( .A1(n6), .A2(regs[188]), .B1(n9), .B2(regs[2236]), .ZN(
        n1916) );
  AOI22_X1 U2671 ( .A1(n56), .A2(regs[1212]), .B1(n97), .B2(regs[1724]), .ZN(
        n1915) );
  OAI211_X1 U2672 ( .C1(n25), .C2(n1917), .A(n1916), .B(n1915), .ZN(
        curr_proc_regs[700]) );
  AOI22_X1 U2673 ( .A1(n6), .A2(regs[189]), .B1(n9), .B2(regs[2237]), .ZN(
        n1919) );
  AOI22_X1 U2674 ( .A1(n56), .A2(regs[1213]), .B1(n97), .B2(regs[1725]), .ZN(
        n1918) );
  OAI211_X1 U2675 ( .C1(n25), .C2(n1920), .A(n1919), .B(n1918), .ZN(
        curr_proc_regs[701]) );
  AOI22_X1 U2676 ( .A1(n6), .A2(regs[190]), .B1(n9), .B2(regs[2238]), .ZN(
        n1922) );
  AOI22_X1 U2677 ( .A1(n56), .A2(regs[1214]), .B1(n97), .B2(regs[1726]), .ZN(
        n1921) );
  OAI211_X1 U2678 ( .C1(n25), .C2(n1923), .A(n1922), .B(n1921), .ZN(
        curr_proc_regs[702]) );
  AOI22_X1 U2679 ( .A1(n6), .A2(regs[191]), .B1(n9), .B2(regs[2239]), .ZN(
        n1925) );
  AOI22_X1 U2680 ( .A1(n56), .A2(regs[1215]), .B1(n97), .B2(regs[1727]), .ZN(
        n1924) );
  OAI211_X1 U2681 ( .C1(n25), .C2(n1926), .A(n1925), .B(n1924), .ZN(
        curr_proc_regs[703]) );
  AOI22_X1 U2682 ( .A1(n6), .A2(regs[192]), .B1(n9), .B2(regs[2240]), .ZN(
        n1928) );
  AOI22_X1 U2683 ( .A1(n83), .A2(regs[1728]), .B1(n3), .B2(regs[704]), .ZN(
        n1927) );
  OAI211_X1 U2684 ( .C1(n65), .C2(n1929), .A(n1928), .B(n1927), .ZN(
        curr_proc_regs[704]) );
  AOI22_X1 U2685 ( .A1(n6), .A2(regs[193]), .B1(n73), .B2(regs[2241]), .ZN(
        n1931) );
  AOI22_X1 U2686 ( .A1(n83), .A2(regs[1729]), .B1(n3), .B2(regs[705]), .ZN(
        n1930) );
  OAI211_X1 U2687 ( .C1(n65), .C2(n1932), .A(n1931), .B(n1930), .ZN(
        curr_proc_regs[705]) );
  AOI22_X1 U2688 ( .A1(n113), .A2(regs[194]), .B1(n17), .B2(regs[2242]), .ZN(
        n1934) );
  AOI22_X1 U2689 ( .A1(n83), .A2(regs[1730]), .B1(n3), .B2(regs[706]), .ZN(
        n1933) );
  OAI211_X1 U2690 ( .C1(n65), .C2(n1935), .A(n1934), .B(n1933), .ZN(
        curr_proc_regs[706]) );
  AOI22_X1 U2691 ( .A1(n6), .A2(regs[195]), .B1(n9), .B2(regs[2243]), .ZN(
        n1937) );
  AOI22_X1 U2692 ( .A1(n83), .A2(regs[1731]), .B1(n3), .B2(regs[707]), .ZN(
        n1936) );
  OAI211_X1 U2693 ( .C1(n65), .C2(n1938), .A(n1937), .B(n1936), .ZN(
        curr_proc_regs[707]) );
  AOI22_X1 U2694 ( .A1(n113), .A2(regs[196]), .B1(n9), .B2(regs[2244]), .ZN(
        n1940) );
  AOI22_X1 U2695 ( .A1(n56), .A2(regs[1220]), .B1(n97), .B2(regs[1732]), .ZN(
        n1939) );
  OAI211_X1 U2696 ( .C1(n25), .C2(n1941), .A(n1940), .B(n1939), .ZN(
        curr_proc_regs[708]) );
  AOI22_X1 U2697 ( .A1(n114), .A2(regs[197]), .B1(n9), .B2(regs[2245]), .ZN(
        n1943) );
  AOI22_X1 U2698 ( .A1(n83), .A2(regs[1733]), .B1(n3), .B2(regs[709]), .ZN(
        n1942) );
  OAI211_X1 U2699 ( .C1(n65), .C2(n1944), .A(n1943), .B(n1942), .ZN(
        curr_proc_regs[709]) );
  AOI22_X1 U2700 ( .A1(n114), .A2(regs[2118]), .B1(n72), .B2(regs[1606]), .ZN(
        n1946) );
  AOI22_X1 U2701 ( .A1(n56), .A2(regs[582]), .B1(n3), .B2(regs[70]), .ZN(n1945) );
  OAI211_X1 U2702 ( .C1(n101), .C2(n1947), .A(n1946), .B(n1945), .ZN(
        curr_proc_regs[70]) );
  AOI22_X1 U2703 ( .A1(n6), .A2(regs[198]), .B1(n9), .B2(regs[2246]), .ZN(
        n1949) );
  AOI22_X1 U2704 ( .A1(n83), .A2(regs[1734]), .B1(n3), .B2(regs[710]), .ZN(
        n1948) );
  OAI211_X1 U2705 ( .C1(n65), .C2(n1950), .A(n1949), .B(n1948), .ZN(
        curr_proc_regs[710]) );
  AOI22_X1 U2706 ( .A1(n113), .A2(regs[199]), .B1(n9), .B2(regs[2247]), .ZN(
        n1952) );
  AOI22_X1 U2707 ( .A1(n60), .A2(regs[1223]), .B1(n19), .B2(regs[1735]), .ZN(
        n1951) );
  OAI211_X1 U2708 ( .C1(n25), .C2(n1953), .A(n1952), .B(n1951), .ZN(
        curr_proc_regs[711]) );
  AOI22_X1 U2709 ( .A1(n114), .A2(regs[200]), .B1(n9), .B2(regs[2248]), .ZN(
        n1955) );
  AOI22_X1 U2710 ( .A1(n83), .A2(regs[1736]), .B1(n3), .B2(regs[712]), .ZN(
        n1954) );
  OAI211_X1 U2711 ( .C1(n1), .C2(n1956), .A(n1955), .B(n1954), .ZN(
        curr_proc_regs[712]) );
  AOI22_X1 U2712 ( .A1(n6), .A2(regs[201]), .B1(n72), .B2(regs[2249]), .ZN(
        n1958) );
  AOI22_X1 U2713 ( .A1(n83), .A2(regs[1737]), .B1(n3), .B2(regs[713]), .ZN(
        n1957) );
  OAI211_X1 U2714 ( .C1(n65), .C2(n1959), .A(n1958), .B(n1957), .ZN(
        curr_proc_regs[713]) );
  AOI22_X1 U2715 ( .A1(n6), .A2(regs[202]), .B1(n9), .B2(regs[2250]), .ZN(
        n1961) );
  AOI22_X1 U2716 ( .A1(n2), .A2(regs[1226]), .B1(n97), .B2(regs[1738]), .ZN(
        n1960) );
  OAI211_X1 U2717 ( .C1(n25), .C2(n1962), .A(n1961), .B(n1960), .ZN(
        curr_proc_regs[714]) );
  AOI22_X1 U2718 ( .A1(n113), .A2(regs[203]), .B1(n73), .B2(regs[2251]), .ZN(
        n1964) );
  AOI22_X1 U2719 ( .A1(n13), .A2(regs[1227]), .B1(n97), .B2(regs[1739]), .ZN(
        n1963) );
  OAI211_X1 U2720 ( .C1(n25), .C2(n1965), .A(n1964), .B(n1963), .ZN(
        curr_proc_regs[715]) );
  AOI22_X1 U2721 ( .A1(n113), .A2(regs[204]), .B1(n72), .B2(regs[2252]), .ZN(
        n1967) );
  AOI22_X1 U2722 ( .A1(n83), .A2(regs[1740]), .B1(n3), .B2(regs[716]), .ZN(
        n1966) );
  OAI211_X1 U2723 ( .C1(n1), .C2(n1968), .A(n1967), .B(n1966), .ZN(
        curr_proc_regs[716]) );
  AOI22_X1 U2724 ( .A1(n114), .A2(regs[205]), .B1(n9), .B2(regs[2253]), .ZN(
        n1970) );
  AOI22_X1 U2725 ( .A1(n98), .A2(regs[1741]), .B1(n3), .B2(regs[717]), .ZN(
        n1969) );
  OAI211_X1 U2726 ( .C1(n65), .C2(n1971), .A(n1970), .B(n1969), .ZN(
        curr_proc_regs[717]) );
  AOI22_X1 U2727 ( .A1(n6), .A2(regs[206]), .B1(n9), .B2(regs[2254]), .ZN(
        n1973) );
  AOI22_X1 U2728 ( .A1(n13), .A2(regs[1230]), .B1(n97), .B2(regs[1742]), .ZN(
        n1972) );
  OAI211_X1 U2729 ( .C1(n25), .C2(n1974), .A(n1973), .B(n1972), .ZN(
        curr_proc_regs[718]) );
  AOI22_X1 U2730 ( .A1(n113), .A2(regs[207]), .B1(n9), .B2(regs[2255]), .ZN(
        n1976) );
  AOI22_X1 U2731 ( .A1(n13), .A2(regs[1231]), .B1(n19), .B2(regs[1743]), .ZN(
        n1975) );
  OAI211_X1 U2732 ( .C1(n25), .C2(n1977), .A(n1976), .B(n1975), .ZN(
        curr_proc_regs[719]) );
  INV_X1 U2733 ( .A(regs[583]), .ZN(n1980) );
  AOI22_X1 U2734 ( .A1(n114), .A2(regs[2119]), .B1(n9), .B2(regs[1607]), .ZN(
        n1979) );
  AOI22_X1 U2735 ( .A1(n83), .A2(regs[1095]), .B1(n3), .B2(regs[71]), .ZN(
        n1978) );
  OAI211_X1 U2736 ( .C1(n1), .C2(n1980), .A(n1979), .B(n1978), .ZN(
        curr_proc_regs[71]) );
  AOI22_X1 U2737 ( .A1(n6), .A2(regs[208]), .B1(n72), .B2(regs[2256]), .ZN(
        n1982) );
  AOI22_X1 U2738 ( .A1(n79), .A2(regs[1744]), .B1(n3), .B2(regs[720]), .ZN(
        n1981) );
  OAI211_X1 U2739 ( .C1(n65), .C2(n1983), .A(n1982), .B(n1981), .ZN(
        curr_proc_regs[720]) );
  AOI22_X1 U2740 ( .A1(n113), .A2(regs[209]), .B1(n9), .B2(regs[2257]), .ZN(
        n1985) );
  AOI22_X1 U2741 ( .A1(n87), .A2(regs[1745]), .B1(n32), .B2(regs[721]), .ZN(
        n1984) );
  OAI211_X1 U2742 ( .C1(n65), .C2(n1986), .A(n1985), .B(n1984), .ZN(
        curr_proc_regs[721]) );
  AOI22_X1 U2743 ( .A1(n114), .A2(regs[210]), .B1(n9), .B2(regs[2258]), .ZN(
        n1988) );
  AOI22_X1 U2744 ( .A1(n96), .A2(regs[1746]), .B1(n45), .B2(regs[722]), .ZN(
        n1987) );
  OAI211_X1 U2745 ( .C1(n65), .C2(n1989), .A(n1988), .B(n1987), .ZN(
        curr_proc_regs[722]) );
  AOI22_X1 U2746 ( .A1(n6), .A2(regs[211]), .B1(n9), .B2(regs[2259]), .ZN(
        n1991) );
  AOI22_X1 U2747 ( .A1(n95), .A2(regs[1747]), .B1(n44), .B2(regs[723]), .ZN(
        n1990) );
  OAI211_X1 U2748 ( .C1(n65), .C2(n1992), .A(n1991), .B(n1990), .ZN(
        curr_proc_regs[723]) );
  AOI22_X1 U2749 ( .A1(n113), .A2(regs[212]), .B1(n9), .B2(regs[2260]), .ZN(
        n1994) );
  AOI22_X1 U2750 ( .A1(n59), .A2(regs[1236]), .B1(n97), .B2(regs[1748]), .ZN(
        n1993) );
  OAI211_X1 U2751 ( .C1(n25), .C2(n1995), .A(n1994), .B(n1993), .ZN(
        curr_proc_regs[724]) );
  AOI22_X1 U2752 ( .A1(n114), .A2(regs[213]), .B1(n9), .B2(regs[2261]), .ZN(
        n1997) );
  AOI22_X1 U2753 ( .A1(n94), .A2(regs[1749]), .B1(n44), .B2(regs[725]), .ZN(
        n1996) );
  OAI211_X1 U2754 ( .C1(n65), .C2(n1998), .A(n1997), .B(n1996), .ZN(
        curr_proc_regs[725]) );
  AOI22_X1 U2755 ( .A1(n114), .A2(regs[214]), .B1(n9), .B2(regs[2262]), .ZN(
        n2000) );
  AOI22_X1 U2756 ( .A1(n96), .A2(regs[1750]), .B1(n44), .B2(regs[726]), .ZN(
        n1999) );
  OAI211_X1 U2757 ( .C1(n65), .C2(n2001), .A(n2000), .B(n1999), .ZN(
        curr_proc_regs[726]) );
  AOI22_X1 U2758 ( .A1(n114), .A2(regs[215]), .B1(n9), .B2(regs[2263]), .ZN(
        n2003) );
  AOI22_X1 U2759 ( .A1(n79), .A2(regs[1751]), .B1(n27), .B2(regs[727]), .ZN(
        n2002) );
  OAI211_X1 U2760 ( .C1(n1), .C2(n2004), .A(n2003), .B(n2002), .ZN(
        curr_proc_regs[727]) );
  AOI22_X1 U2761 ( .A1(n114), .A2(regs[216]), .B1(n9), .B2(regs[2264]), .ZN(
        n2006) );
  AOI22_X1 U2762 ( .A1(n81), .A2(regs[1752]), .B1(n26), .B2(regs[728]), .ZN(
        n2005) );
  OAI211_X1 U2763 ( .C1(n65), .C2(n2007), .A(n2006), .B(n2005), .ZN(
        curr_proc_regs[728]) );
  AOI22_X1 U2764 ( .A1(n114), .A2(regs[217]), .B1(n73), .B2(regs[2265]), .ZN(
        n2009) );
  AOI22_X1 U2765 ( .A1(n82), .A2(regs[1753]), .B1(n45), .B2(regs[729]), .ZN(
        n2008) );
  OAI211_X1 U2766 ( .C1(n2207), .C2(n2010), .A(n2009), .B(n2008), .ZN(
        curr_proc_regs[729]) );
  AOI22_X1 U2767 ( .A1(n114), .A2(regs[2120]), .B1(n9), .B2(regs[1608]), .ZN(
        n2012) );
  AOI22_X1 U2768 ( .A1(n61), .A2(regs[584]), .B1(n46), .B2(regs[72]), .ZN(
        n2011) );
  OAI211_X1 U2769 ( .C1(n101), .C2(n2013), .A(n2012), .B(n2011), .ZN(
        curr_proc_regs[72]) );
  AOI22_X1 U2770 ( .A1(n114), .A2(regs[218]), .B1(n9), .B2(regs[2266]), .ZN(
        n2015) );
  AOI22_X1 U2771 ( .A1(n82), .A2(regs[1754]), .B1(n34), .B2(regs[730]), .ZN(
        n2014) );
  OAI211_X1 U2772 ( .C1(n65), .C2(n2016), .A(n2015), .B(n2014), .ZN(
        curr_proc_regs[730]) );
  AOI22_X1 U2773 ( .A1(n114), .A2(regs[219]), .B1(n9), .B2(regs[2267]), .ZN(
        n2018) );
  AOI22_X1 U2774 ( .A1(n2), .A2(regs[1243]), .B1(n19), .B2(regs[1755]), .ZN(
        n2017) );
  OAI211_X1 U2775 ( .C1(n25), .C2(n2019), .A(n2018), .B(n2017), .ZN(
        curr_proc_regs[731]) );
  AOI22_X1 U2776 ( .A1(n114), .A2(regs[220]), .B1(n9), .B2(regs[2268]), .ZN(
        n2021) );
  AOI22_X1 U2777 ( .A1(n59), .A2(regs[1244]), .B1(n19), .B2(regs[1756]), .ZN(
        n2020) );
  OAI211_X1 U2778 ( .C1(n25), .C2(n2022), .A(n2021), .B(n2020), .ZN(
        curr_proc_regs[732]) );
  AOI22_X1 U2779 ( .A1(n114), .A2(regs[221]), .B1(n9), .B2(regs[2269]), .ZN(
        n2024) );
  AOI22_X1 U2780 ( .A1(n82), .A2(regs[1757]), .B1(n45), .B2(regs[733]), .ZN(
        n2023) );
  OAI211_X1 U2781 ( .C1(n65), .C2(n2025), .A(n2024), .B(n2023), .ZN(
        curr_proc_regs[733]) );
  AOI22_X1 U2782 ( .A1(n114), .A2(regs[222]), .B1(n14), .B2(regs[2270]), .ZN(
        n2027) );
  AOI22_X1 U2783 ( .A1(n60), .A2(regs[1246]), .B1(n97), .B2(regs[1758]), .ZN(
        n2026) );
  OAI211_X1 U2784 ( .C1(n25), .C2(n2028), .A(n2027), .B(n2026), .ZN(
        curr_proc_regs[734]) );
  AOI22_X1 U2785 ( .A1(n114), .A2(regs[223]), .B1(n73), .B2(regs[2271]), .ZN(
        n2030) );
  AOI22_X1 U2786 ( .A1(n2), .A2(regs[1247]), .B1(n19), .B2(regs[1759]), .ZN(
        n2029) );
  OAI211_X1 U2787 ( .C1(n25), .C2(n2031), .A(n2030), .B(n2029), .ZN(
        curr_proc_regs[735]) );
  AOI22_X1 U2788 ( .A1(n113), .A2(regs[224]), .B1(n14), .B2(regs[2272]), .ZN(
        n2033) );
  AOI22_X1 U2789 ( .A1(n82), .A2(regs[1760]), .B1(n32), .B2(regs[736]), .ZN(
        n2032) );
  OAI211_X1 U2790 ( .C1(n65), .C2(n2034), .A(n2033), .B(n2032), .ZN(
        curr_proc_regs[736]) );
  AOI22_X1 U2791 ( .A1(n113), .A2(regs[225]), .B1(n14), .B2(regs[2273]), .ZN(
        n2036) );
  AOI22_X1 U2792 ( .A1(n82), .A2(regs[1761]), .B1(n32), .B2(regs[737]), .ZN(
        n2035) );
  OAI211_X1 U2793 ( .C1(n65), .C2(n2037), .A(n2036), .B(n2035), .ZN(
        curr_proc_regs[737]) );
  AOI22_X1 U2794 ( .A1(n113), .A2(regs[226]), .B1(n72), .B2(regs[2274]), .ZN(
        n2039) );
  AOI22_X1 U2795 ( .A1(n59), .A2(regs[1250]), .B1(n97), .B2(regs[1762]), .ZN(
        n2038) );
  OAI211_X1 U2796 ( .C1(n2134), .C2(n2040), .A(n2039), .B(n2038), .ZN(
        curr_proc_regs[738]) );
  AOI22_X1 U2797 ( .A1(n113), .A2(regs[227]), .B1(n72), .B2(regs[2275]), .ZN(
        n2042) );
  AOI22_X1 U2798 ( .A1(n82), .A2(regs[1763]), .B1(n32), .B2(regs[739]), .ZN(
        n2041) );
  OAI211_X1 U2799 ( .C1(n65), .C2(n2043), .A(n2042), .B(n2041), .ZN(
        curr_proc_regs[739]) );
  AOI22_X1 U2800 ( .A1(n113), .A2(regs[2121]), .B1(n14), .B2(regs[1609]), .ZN(
        n2045) );
  AOI22_X1 U2801 ( .A1(n2), .A2(regs[585]), .B1(n32), .B2(regs[73]), .ZN(n2044) );
  OAI211_X1 U2802 ( .C1(n100), .C2(n2046), .A(n2045), .B(n2044), .ZN(
        curr_proc_regs[73]) );
  AOI22_X1 U2803 ( .A1(n113), .A2(regs[228]), .B1(n77), .B2(regs[2276]), .ZN(
        n2048) );
  AOI22_X1 U2804 ( .A1(n82), .A2(regs[1764]), .B1(n32), .B2(regs[740]), .ZN(
        n2047) );
  OAI211_X1 U2805 ( .C1(n65), .C2(n2049), .A(n2048), .B(n2047), .ZN(
        curr_proc_regs[740]) );
  AOI22_X1 U2806 ( .A1(n113), .A2(regs[229]), .B1(n14), .B2(regs[2277]), .ZN(
        n2051) );
  AOI22_X1 U2807 ( .A1(n82), .A2(regs[1765]), .B1(n32), .B2(regs[741]), .ZN(
        n2050) );
  OAI211_X1 U2808 ( .C1(n65), .C2(n2052), .A(n2051), .B(n2050), .ZN(
        curr_proc_regs[741]) );
  AOI22_X1 U2809 ( .A1(n113), .A2(regs[230]), .B1(n14), .B2(regs[2278]), .ZN(
        n2054) );
  AOI22_X1 U2810 ( .A1(n82), .A2(regs[1766]), .B1(n32), .B2(regs[742]), .ZN(
        n2053) );
  OAI211_X1 U2811 ( .C1(n1), .C2(n2055), .A(n2054), .B(n2053), .ZN(
        curr_proc_regs[742]) );
  AOI22_X1 U2812 ( .A1(n113), .A2(regs[231]), .B1(n73), .B2(regs[2279]), .ZN(
        n2057) );
  AOI22_X1 U2813 ( .A1(n82), .A2(regs[1767]), .B1(n32), .B2(regs[743]), .ZN(
        n2056) );
  OAI211_X1 U2814 ( .C1(n65), .C2(n2058), .A(n2057), .B(n2056), .ZN(
        curr_proc_regs[743]) );
  AOI22_X1 U2815 ( .A1(n113), .A2(regs[232]), .B1(n14), .B2(regs[2280]), .ZN(
        n2060) );
  AOI22_X1 U2816 ( .A1(n82), .A2(regs[1768]), .B1(n32), .B2(regs[744]), .ZN(
        n2059) );
  OAI211_X1 U2817 ( .C1(n65), .C2(n2061), .A(n2060), .B(n2059), .ZN(
        curr_proc_regs[744]) );
  AOI22_X1 U2818 ( .A1(n113), .A2(regs[233]), .B1(n14), .B2(regs[2281]), .ZN(
        n2063) );
  AOI22_X1 U2819 ( .A1(n82), .A2(regs[1769]), .B1(n32), .B2(regs[745]), .ZN(
        n2062) );
  OAI211_X1 U2820 ( .C1(n1), .C2(n2064), .A(n2063), .B(n2062), .ZN(
        curr_proc_regs[745]) );
  AOI22_X1 U2821 ( .A1(n111), .A2(regs[234]), .B1(n15), .B2(regs[2282]), .ZN(
        n2066) );
  AOI22_X1 U2822 ( .A1(n78), .A2(regs[1770]), .B1(n32), .B2(regs[746]), .ZN(
        n2065) );
  OAI211_X1 U2823 ( .C1(n1), .C2(n2067), .A(n2066), .B(n2065), .ZN(
        curr_proc_regs[746]) );
  AOI22_X1 U2824 ( .A1(n110), .A2(regs[235]), .B1(n72), .B2(regs[2283]), .ZN(
        n2069) );
  AOI22_X1 U2825 ( .A1(n61), .A2(regs[1259]), .B1(n19), .B2(regs[1771]), .ZN(
        n2068) );
  OAI211_X1 U2826 ( .C1(n24), .C2(n2070), .A(n2069), .B(n2068), .ZN(
        curr_proc_regs[747]) );
  AOI22_X1 U2827 ( .A1(n112), .A2(regs[236]), .B1(n14), .B2(regs[2284]), .ZN(
        n2072) );
  AOI22_X1 U2828 ( .A1(n2), .A2(regs[1260]), .B1(n19), .B2(regs[1772]), .ZN(
        n2071) );
  OAI211_X1 U2829 ( .C1(n25), .C2(n2073), .A(n2072), .B(n2071), .ZN(
        curr_proc_regs[748]) );
  AOI22_X1 U2830 ( .A1(n112), .A2(regs[237]), .B1(n72), .B2(regs[2285]), .ZN(
        n2075) );
  AOI22_X1 U2831 ( .A1(n79), .A2(regs[1773]), .B1(n33), .B2(regs[749]), .ZN(
        n2074) );
  OAI211_X1 U2832 ( .C1(n65), .C2(n2076), .A(n2075), .B(n2074), .ZN(
        curr_proc_regs[749]) );
  AOI22_X1 U2833 ( .A1(n110), .A2(regs[2122]), .B1(n73), .B2(regs[1610]), .ZN(
        n2078) );
  AOI22_X1 U2834 ( .A1(n59), .A2(regs[586]), .B1(n33), .B2(regs[74]), .ZN(
        n2077) );
  OAI211_X1 U2835 ( .C1(n102), .C2(n2079), .A(n2078), .B(n2077), .ZN(
        curr_proc_regs[74]) );
  AOI22_X1 U2836 ( .A1(n111), .A2(regs[238]), .B1(n67), .B2(regs[2286]), .ZN(
        n2081) );
  AOI22_X1 U2837 ( .A1(n60), .A2(regs[1262]), .B1(n19), .B2(regs[1774]), .ZN(
        n2080) );
  OAI211_X1 U2838 ( .C1(n25), .C2(n2082), .A(n2081), .B(n2080), .ZN(
        curr_proc_regs[750]) );
  AOI22_X1 U2839 ( .A1(n110), .A2(regs[239]), .B1(n14), .B2(regs[2287]), .ZN(
        n2084) );
  AOI22_X1 U2840 ( .A1(n59), .A2(regs[1263]), .B1(n19), .B2(regs[1775]), .ZN(
        n2083) );
  OAI211_X1 U2841 ( .C1(n25), .C2(n2085), .A(n2084), .B(n2083), .ZN(
        curr_proc_regs[751]) );
  AOI22_X1 U2842 ( .A1(n112), .A2(regs[240]), .B1(n72), .B2(regs[2288]), .ZN(
        n2087) );
  AOI22_X1 U2843 ( .A1(n80), .A2(regs[1776]), .B1(n33), .B2(regs[752]), .ZN(
        n2086) );
  OAI211_X1 U2844 ( .C1(n1), .C2(n2088), .A(n2087), .B(n2086), .ZN(
        curr_proc_regs[752]) );
  AOI22_X1 U2845 ( .A1(n111), .A2(regs[241]), .B1(n72), .B2(regs[2289]), .ZN(
        n2090) );
  AOI22_X1 U2846 ( .A1(n2), .A2(regs[1265]), .B1(n19), .B2(regs[1777]), .ZN(
        n2089) );
  OAI211_X1 U2847 ( .C1(n24), .C2(n2091), .A(n2090), .B(n2089), .ZN(
        curr_proc_regs[753]) );
  AOI22_X1 U2848 ( .A1(n112), .A2(regs[242]), .B1(n69), .B2(regs[2290]), .ZN(
        n2093) );
  AOI22_X1 U2849 ( .A1(n83), .A2(regs[1778]), .B1(n33), .B2(regs[754]), .ZN(
        n2092) );
  OAI211_X1 U2850 ( .C1(n65), .C2(n2094), .A(n2093), .B(n2092), .ZN(
        curr_proc_regs[754]) );
  AOI22_X1 U2851 ( .A1(n111), .A2(regs[243]), .B1(n72), .B2(regs[2291]), .ZN(
        n2096) );
  AOI22_X1 U2852 ( .A1(n13), .A2(regs[1267]), .B1(n19), .B2(regs[1779]), .ZN(
        n2095) );
  OAI211_X1 U2853 ( .C1(n2134), .C2(n2097), .A(n2096), .B(n2095), .ZN(
        curr_proc_regs[755]) );
  AOI22_X1 U2854 ( .A1(n110), .A2(regs[244]), .B1(n72), .B2(regs[2292]), .ZN(
        n2099) );
  AOI22_X1 U2855 ( .A1(n13), .A2(regs[1268]), .B1(n97), .B2(regs[1780]), .ZN(
        n2098) );
  OAI211_X1 U2856 ( .C1(n25), .C2(n2100), .A(n2099), .B(n2098), .ZN(
        curr_proc_regs[756]) );
  AOI22_X1 U2857 ( .A1(n111), .A2(regs[245]), .B1(n73), .B2(regs[2293]), .ZN(
        n2102) );
  AOI22_X1 U2858 ( .A1(n84), .A2(regs[1781]), .B1(n33), .B2(regs[757]), .ZN(
        n2101) );
  OAI211_X1 U2859 ( .C1(n65), .C2(n2103), .A(n2102), .B(n2101), .ZN(
        curr_proc_regs[757]) );
  AOI22_X1 U2860 ( .A1(n110), .A2(regs[246]), .B1(n77), .B2(regs[2294]), .ZN(
        n2105) );
  AOI22_X1 U2861 ( .A1(n85), .A2(regs[1782]), .B1(n33), .B2(regs[758]), .ZN(
        n2104) );
  OAI211_X1 U2862 ( .C1(n65), .C2(n2106), .A(n2105), .B(n2104), .ZN(
        curr_proc_regs[758]) );
  AOI22_X1 U2863 ( .A1(n112), .A2(regs[247]), .B1(n72), .B2(regs[2295]), .ZN(
        n2108) );
  AOI22_X1 U2864 ( .A1(n2), .A2(regs[1271]), .B1(n97), .B2(regs[1783]), .ZN(
        n2107) );
  OAI211_X1 U2865 ( .C1(n25), .C2(n2109), .A(n2108), .B(n2107), .ZN(
        curr_proc_regs[759]) );
  INV_X1 U2866 ( .A(regs[1099]), .ZN(n2112) );
  AOI22_X1 U2867 ( .A1(n112), .A2(regs[2123]), .B1(n72), .B2(regs[1611]), .ZN(
        n2111) );
  AOI22_X1 U2868 ( .A1(n13), .A2(regs[587]), .B1(n33), .B2(regs[75]), .ZN(
        n2110) );
  OAI211_X1 U2869 ( .C1(n99), .C2(n2112), .A(n2111), .B(n2110), .ZN(
        curr_proc_regs[75]) );
  AOI22_X1 U2870 ( .A1(n111), .A2(regs[248]), .B1(n73), .B2(regs[2296]), .ZN(
        n2114) );
  AOI22_X1 U2871 ( .A1(n53), .A2(regs[1272]), .B1(n19), .B2(regs[1784]), .ZN(
        n2113) );
  OAI211_X1 U2872 ( .C1(n25), .C2(n2115), .A(n2114), .B(n2113), .ZN(
        curr_proc_regs[760]) );
  AOI22_X1 U2873 ( .A1(n110), .A2(regs[249]), .B1(n9), .B2(regs[2297]), .ZN(
        n2117) );
  AOI22_X1 U2874 ( .A1(n13), .A2(regs[1273]), .B1(n97), .B2(regs[1785]), .ZN(
        n2116) );
  OAI211_X1 U2875 ( .C1(n2134), .C2(n2118), .A(n2117), .B(n2116), .ZN(
        curr_proc_regs[761]) );
  AOI22_X1 U2876 ( .A1(n112), .A2(regs[250]), .B1(n72), .B2(regs[2298]), .ZN(
        n2120) );
  AOI22_X1 U2877 ( .A1(n60), .A2(regs[1274]), .B1(n19), .B2(regs[1786]), .ZN(
        n2119) );
  OAI211_X1 U2878 ( .C1(n25), .C2(n2121), .A(n2120), .B(n2119), .ZN(
        curr_proc_regs[762]) );
  AOI22_X1 U2879 ( .A1(n111), .A2(regs[251]), .B1(n72), .B2(regs[2299]), .ZN(
        n2123) );
  AOI22_X1 U2880 ( .A1(n86), .A2(regs[1787]), .B1(n33), .B2(regs[763]), .ZN(
        n2122) );
  OAI211_X1 U2881 ( .C1(n65), .C2(n2124), .A(n2123), .B(n2122), .ZN(
        curr_proc_regs[763]) );
  AOI22_X1 U2882 ( .A1(n111), .A2(regs[252]), .B1(n73), .B2(regs[2300]), .ZN(
        n2126) );
  AOI22_X1 U2883 ( .A1(n87), .A2(regs[1788]), .B1(n33), .B2(regs[764]), .ZN(
        n2125) );
  OAI211_X1 U2884 ( .C1(n65), .C2(n2127), .A(n2126), .B(n2125), .ZN(
        curr_proc_regs[764]) );
  AOI22_X1 U2885 ( .A1(n110), .A2(regs[253]), .B1(n14), .B2(regs[2301]), .ZN(
        n2129) );
  AOI22_X1 U2886 ( .A1(n61), .A2(regs[1277]), .B1(n97), .B2(regs[1789]), .ZN(
        n2128) );
  OAI211_X1 U2887 ( .C1(n25), .C2(n2130), .A(n2129), .B(n2128), .ZN(
        curr_proc_regs[765]) );
  AOI22_X1 U2888 ( .A1(n110), .A2(regs[254]), .B1(n66), .B2(regs[2302]), .ZN(
        n2132) );
  AOI22_X1 U2889 ( .A1(n61), .A2(regs[1278]), .B1(n97), .B2(regs[1790]), .ZN(
        n2131) );
  OAI211_X1 U2890 ( .C1(n25), .C2(n2133), .A(n2132), .B(n2131), .ZN(
        curr_proc_regs[766]) );
  AOI22_X1 U2891 ( .A1(n112), .A2(regs[255]), .B1(n72), .B2(regs[2303]), .ZN(
        n2136) );
  AOI22_X1 U2892 ( .A1(n83), .A2(regs[1791]), .B1(n33), .B2(regs[767]), .ZN(
        n2135) );
  OAI211_X1 U2893 ( .C1(n65), .C2(n2137), .A(n2136), .B(n2135), .ZN(
        curr_proc_regs[767]) );
  AOI22_X1 U2894 ( .A1(n111), .A2(regs[2124]), .B1(n14), .B2(regs[1612]), .ZN(
        n2139) );
  AOI22_X1 U2895 ( .A1(n2), .A2(regs[588]), .B1(n33), .B2(regs[76]), .ZN(n2138) );
  OAI211_X1 U2896 ( .C1(n5), .C2(n2140), .A(n2139), .B(n2138), .ZN(
        curr_proc_regs[76]) );
  INV_X1 U2897 ( .A(regs[589]), .ZN(n2143) );
  AOI22_X1 U2898 ( .A1(n110), .A2(regs[2125]), .B1(n14), .B2(regs[1613]), .ZN(
        n2142) );
  AOI22_X1 U2899 ( .A1(n95), .A2(regs[1101]), .B1(n34), .B2(regs[77]), .ZN(
        n2141) );
  OAI211_X1 U2900 ( .C1(n65), .C2(n2143), .A(n2142), .B(n2141), .ZN(
        curr_proc_regs[77]) );
  AOI22_X1 U2901 ( .A1(n112), .A2(regs[2126]), .B1(n72), .B2(regs[1614]), .ZN(
        n2145) );
  AOI22_X1 U2902 ( .A1(n59), .A2(regs[590]), .B1(n34), .B2(regs[78]), .ZN(
        n2144) );
  OAI211_X1 U2903 ( .C1(n16), .C2(n2146), .A(n2145), .B(n2144), .ZN(
        curr_proc_regs[78]) );
  AOI22_X1 U2904 ( .A1(n111), .A2(regs[2127]), .B1(n73), .B2(regs[1615]), .ZN(
        n2148) );
  AOI22_X1 U2905 ( .A1(n60), .A2(regs[591]), .B1(n34), .B2(regs[79]), .ZN(
        n2147) );
  OAI211_X1 U2906 ( .C1(n2221), .C2(n2149), .A(n2148), .B(n2147), .ZN(
        curr_proc_regs[79]) );
  AOI22_X1 U2907 ( .A1(n110), .A2(regs[2055]), .B1(n14), .B2(regs[1543]), .ZN(
        n2151) );
  AOI22_X1 U2908 ( .A1(n2), .A2(regs[519]), .B1(n34), .B2(regs[7]), .ZN(n2150)
         );
  OAI211_X1 U2909 ( .C1(n16), .C2(n2152), .A(n2151), .B(n2150), .ZN(
        curr_proc_regs[7]) );
  AOI22_X1 U2910 ( .A1(n112), .A2(regs[2128]), .B1(n14), .B2(regs[1616]), .ZN(
        n2154) );
  AOI22_X1 U2911 ( .A1(n13), .A2(regs[592]), .B1(n34), .B2(regs[80]), .ZN(
        n2153) );
  OAI211_X1 U2912 ( .C1(n102), .C2(n2155), .A(n2154), .B(n2153), .ZN(
        curr_proc_regs[80]) );
  AOI22_X1 U2913 ( .A1(n111), .A2(regs[2129]), .B1(n14), .B2(regs[1617]), .ZN(
        n2157) );
  AOI22_X1 U2914 ( .A1(n59), .A2(regs[593]), .B1(n34), .B2(regs[81]), .ZN(
        n2156) );
  OAI211_X1 U2915 ( .C1(n2221), .C2(n2158), .A(n2157), .B(n2156), .ZN(
        curr_proc_regs[81]) );
  INV_X1 U2916 ( .A(regs[1106]), .ZN(n2161) );
  AOI22_X1 U2917 ( .A1(n110), .A2(regs[2130]), .B1(n70), .B2(regs[1618]), .ZN(
        n2160) );
  AOI22_X1 U2918 ( .A1(n60), .A2(regs[594]), .B1(n34), .B2(regs[82]), .ZN(
        n2159) );
  OAI211_X1 U2919 ( .C1(n2221), .C2(n2161), .A(n2160), .B(n2159), .ZN(
        curr_proc_regs[82]) );
  INV_X1 U2920 ( .A(regs[1107]), .ZN(n2164) );
  AOI22_X1 U2921 ( .A1(n112), .A2(regs[2131]), .B1(n14), .B2(regs[1619]), .ZN(
        n2163) );
  AOI22_X1 U2922 ( .A1(n60), .A2(regs[595]), .B1(n34), .B2(regs[83]), .ZN(
        n2162) );
  OAI211_X1 U2923 ( .C1(n101), .C2(n2164), .A(n2163), .B(n2162), .ZN(
        curr_proc_regs[83]) );
  INV_X1 U2924 ( .A(regs[1108]), .ZN(n2167) );
  AOI22_X1 U2925 ( .A1(n112), .A2(regs[2132]), .B1(n14), .B2(regs[1620]), .ZN(
        n2166) );
  AOI22_X1 U2926 ( .A1(n60), .A2(regs[596]), .B1(n34), .B2(regs[84]), .ZN(
        n2165) );
  OAI211_X1 U2927 ( .C1(n2221), .C2(n2167), .A(n2166), .B(n2165), .ZN(
        curr_proc_regs[84]) );
  INV_X1 U2928 ( .A(regs[597]), .ZN(n2170) );
  AOI22_X1 U2929 ( .A1(n112), .A2(regs[2133]), .B1(n14), .B2(regs[1621]), .ZN(
        n2169) );
  AOI22_X1 U2930 ( .A1(n94), .A2(regs[1109]), .B1(n34), .B2(regs[85]), .ZN(
        n2168) );
  OAI211_X1 U2931 ( .C1(n1), .C2(n2170), .A(n2169), .B(n2168), .ZN(
        curr_proc_regs[85]) );
  AOI22_X1 U2932 ( .A1(n112), .A2(regs[2134]), .B1(n14), .B2(regs[1622]), .ZN(
        n2172) );
  AOI22_X1 U2933 ( .A1(n58), .A2(regs[598]), .B1(n34), .B2(regs[86]), .ZN(
        n2171) );
  OAI211_X1 U2934 ( .C1(n99), .C2(n2173), .A(n2172), .B(n2171), .ZN(
        curr_proc_regs[86]) );
  AOI22_X1 U2935 ( .A1(n112), .A2(regs[2135]), .B1(n66), .B2(regs[1623]), .ZN(
        n2175) );
  AOI22_X1 U2936 ( .A1(n60), .A2(regs[599]), .B1(n35), .B2(regs[87]), .ZN(
        n2174) );
  OAI211_X1 U2937 ( .C1(n16), .C2(n2176), .A(n2175), .B(n2174), .ZN(
        curr_proc_regs[87]) );
  AOI22_X1 U2938 ( .A1(n112), .A2(regs[2136]), .B1(n15), .B2(regs[1624]), .ZN(
        n2178) );
  AOI22_X1 U2939 ( .A1(n60), .A2(regs[600]), .B1(n35), .B2(regs[88]), .ZN(
        n2177) );
  OAI211_X1 U2940 ( .C1(n102), .C2(n2179), .A(n2178), .B(n2177), .ZN(
        curr_proc_regs[88]) );
  INV_X1 U2941 ( .A(regs[1113]), .ZN(n2182) );
  AOI22_X1 U2942 ( .A1(n112), .A2(regs[2137]), .B1(n14), .B2(regs[1625]), .ZN(
        n2181) );
  AOI22_X1 U2943 ( .A1(n60), .A2(regs[601]), .B1(n35), .B2(regs[89]), .ZN(
        n2180) );
  OAI211_X1 U2944 ( .C1(n100), .C2(n2182), .A(n2181), .B(n2180), .ZN(
        curr_proc_regs[89]) );
  AOI22_X1 U2945 ( .A1(n112), .A2(regs[2056]), .B1(n67), .B2(regs[1544]), .ZN(
        n2184) );
  AOI22_X1 U2946 ( .A1(n55), .A2(regs[520]), .B1(n35), .B2(regs[8]), .ZN(n2183) );
  OAI211_X1 U2947 ( .C1(n5), .C2(n2185), .A(n2184), .B(n2183), .ZN(
        curr_proc_regs[8]) );
  INV_X1 U2948 ( .A(regs[602]), .ZN(n2188) );
  AOI22_X1 U2949 ( .A1(n112), .A2(regs[2138]), .B1(n14), .B2(regs[1626]), .ZN(
        n2187) );
  AOI22_X1 U2950 ( .A1(n81), .A2(regs[1114]), .B1(n35), .B2(regs[90]), .ZN(
        n2186) );
  OAI211_X1 U2951 ( .C1(n65), .C2(n2188), .A(n2187), .B(n2186), .ZN(
        curr_proc_regs[90]) );
  INV_X1 U2952 ( .A(regs[603]), .ZN(n2191) );
  AOI22_X1 U2953 ( .A1(n112), .A2(regs[2139]), .B1(n14), .B2(regs[1627]), .ZN(
        n2190) );
  AOI22_X1 U2954 ( .A1(n84), .A2(regs[1115]), .B1(n35), .B2(regs[91]), .ZN(
        n2189) );
  OAI211_X1 U2955 ( .C1(n1), .C2(n2191), .A(n2190), .B(n2189), .ZN(
        curr_proc_regs[91]) );
  AOI22_X1 U2956 ( .A1(n112), .A2(regs[2140]), .B1(n14), .B2(regs[1628]), .ZN(
        n2193) );
  AOI22_X1 U2957 ( .A1(n60), .A2(regs[604]), .B1(n35), .B2(regs[92]), .ZN(
        n2192) );
  OAI211_X1 U2958 ( .C1(n102), .C2(n2194), .A(n2193), .B(n2192), .ZN(
        curr_proc_regs[92]) );
  INV_X1 U2959 ( .A(regs[1117]), .ZN(n2197) );
  AOI22_X1 U2960 ( .A1(n112), .A2(regs[2141]), .B1(n14), .B2(regs[1629]), .ZN(
        n2196) );
  AOI22_X1 U2961 ( .A1(n61), .A2(regs[605]), .B1(n35), .B2(regs[93]), .ZN(
        n2195) );
  OAI211_X1 U2962 ( .C1(n102), .C2(n2197), .A(n2196), .B(n2195), .ZN(
        curr_proc_regs[93]) );
  INV_X1 U2963 ( .A(regs[1118]), .ZN(n2200) );
  AOI22_X1 U2964 ( .A1(n111), .A2(regs[2142]), .B1(n4), .B2(regs[1630]), .ZN(
        n2199) );
  AOI22_X1 U2965 ( .A1(n56), .A2(regs[606]), .B1(n35), .B2(regs[94]), .ZN(
        n2198) );
  OAI211_X1 U2966 ( .C1(n99), .C2(n2200), .A(n2199), .B(n2198), .ZN(
        curr_proc_regs[94]) );
  AOI22_X1 U2967 ( .A1(n111), .A2(regs[2143]), .B1(n14), .B2(regs[1631]), .ZN(
        n2202) );
  AOI22_X1 U2968 ( .A1(n58), .A2(regs[607]), .B1(n35), .B2(regs[95]), .ZN(
        n2201) );
  OAI211_X1 U2969 ( .C1(n2221), .C2(n2203), .A(n2202), .B(n2201), .ZN(
        curr_proc_regs[95]) );
  INV_X1 U2970 ( .A(regs[608]), .ZN(n2206) );
  AOI22_X1 U2971 ( .A1(n111), .A2(regs[2144]), .B1(n2217), .B2(regs[1632]), 
        .ZN(n2205) );
  AOI22_X1 U2972 ( .A1(n83), .A2(regs[1120]), .B1(n35), .B2(regs[96]), .ZN(
        n2204) );
  OAI211_X1 U2973 ( .C1(n65), .C2(n2206), .A(n2205), .B(n2204), .ZN(
        curr_proc_regs[96]) );
  INV_X1 U2974 ( .A(regs[1121]), .ZN(n2210) );
  AOI22_X1 U2975 ( .A1(n111), .A2(regs[2145]), .B1(n17), .B2(regs[1633]), .ZN(
        n2209) );
  AOI22_X1 U2976 ( .A1(n62), .A2(regs[609]), .B1(n36), .B2(regs[97]), .ZN(
        n2208) );
  OAI211_X1 U2977 ( .C1(n102), .C2(n2210), .A(n2209), .B(n2208), .ZN(
        curr_proc_regs[97]) );
  INV_X1 U2978 ( .A(regs[1122]), .ZN(n2213) );
  AOI22_X1 U2979 ( .A1(n6), .A2(regs[2146]), .B1(n72), .B2(regs[1634]), .ZN(
        n2212) );
  AOI22_X1 U2980 ( .A1(n60), .A2(regs[610]), .B1(n36), .B2(regs[98]), .ZN(
        n2211) );
  OAI211_X1 U2981 ( .C1(n2221), .C2(n2213), .A(n2212), .B(n2211), .ZN(
        curr_proc_regs[98]) );
  AOI22_X1 U2982 ( .A1(n103), .A2(regs[2147]), .B1(n72), .B2(regs[1635]), .ZN(
        n2215) );
  AOI22_X1 U2983 ( .A1(n56), .A2(regs[611]), .B1(n36), .B2(regs[99]), .ZN(
        n2214) );
  OAI211_X1 U2984 ( .C1(n100), .C2(n2216), .A(n2215), .B(n2214), .ZN(
        curr_proc_regs[99]) );
  INV_X1 U2985 ( .A(regs[1033]), .ZN(n2220) );
  AOI22_X1 U2986 ( .A1(n119), .A2(regs[2057]), .B1(n72), .B2(regs[1545]), .ZN(
        n2219) );
  AOI22_X1 U2987 ( .A1(n54), .A2(regs[521]), .B1(n36), .B2(regs[9]), .ZN(n2218) );
  OAI211_X1 U2988 ( .C1(n2221), .C2(n2220), .A(n2219), .B(n2218), .ZN(
        curr_proc_regs[9]) );
endmodule


module mux_N32_M5_0 ( S, Q, Y );
  input [4:0] S;
  input [1023:0] Q;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687;

  AOI22_X1 U2 ( .A1(n673), .A2(Q[509]), .B1(n672), .B2(Q[573]), .ZN(n1) );
  AOI22_X1 U3 ( .A1(n675), .A2(Q[669]), .B1(n674), .B2(Q[477]), .ZN(n2) );
  AOI22_X1 U4 ( .A1(n677), .A2(Q[381]), .B1(n676), .B2(Q[317]), .ZN(n3) );
  AOI22_X1 U5 ( .A1(n679), .A2(Q[413]), .B1(n678), .B2(Q[285]), .ZN(n4) );
  NAND4_X1 U6 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(n5) );
  AOI22_X1 U7 ( .A1(n681), .A2(Q[349]), .B1(n680), .B2(Q[445]), .ZN(n6) );
  AOI22_X1 U8 ( .A1(n683), .A2(Q[253]), .B1(n682), .B2(Q[157]), .ZN(n7) );
  AOI22_X1 U9 ( .A1(n685), .A2(Q[93]), .B1(n684), .B2(Q[189]), .ZN(n8) );
  AOI22_X1 U10 ( .A1(n687), .A2(Q[221]), .B1(n686), .B2(Q[61]), .ZN(n9) );
  NAND4_X1 U11 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n10) );
  AOI22_X1 U12 ( .A1(n656), .A2(Q[1021]), .B1(n655), .B2(Q[957]), .ZN(n11) );
  AOI22_X1 U13 ( .A1(n658), .A2(Q[989]), .B1(n657), .B2(Q[925]), .ZN(n12) );
  AOI222_X1 U14 ( .A1(n660), .A2(Q[829]), .B1(n661), .B2(Q[125]), .C1(n659), 
        .C2(Q[765]), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n14) );
  AOI22_X1 U16 ( .A1(n663), .A2(Q[861]), .B1(n662), .B2(Q[733]), .ZN(n15) );
  AOI22_X1 U17 ( .A1(n665), .A2(Q[797]), .B1(n664), .B2(Q[893]), .ZN(n16) );
  NAND4_X1 U18 ( .A1(n635), .A2(n636), .A3(n15), .A4(n16), .ZN(n17) );
  OR4_X1 U19 ( .A1(n5), .A2(n10), .A3(n14), .A4(n17), .ZN(Y[29]) );
  AOI22_X1 U20 ( .A1(n673), .A2(Q[499]), .B1(n672), .B2(Q[563]), .ZN(n18) );
  AOI22_X1 U21 ( .A1(n675), .A2(Q[659]), .B1(n674), .B2(Q[467]), .ZN(n19) );
  AOI22_X1 U22 ( .A1(n677), .A2(Q[371]), .B1(n676), .B2(Q[307]), .ZN(n20) );
  AOI22_X1 U23 ( .A1(n679), .A2(Q[403]), .B1(n678), .B2(Q[275]), .ZN(n21) );
  NAND4_X1 U24 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .ZN(n22) );
  AOI22_X1 U25 ( .A1(n681), .A2(Q[339]), .B1(n680), .B2(Q[435]), .ZN(n23) );
  AOI22_X1 U26 ( .A1(n683), .A2(Q[243]), .B1(n682), .B2(Q[147]), .ZN(n24) );
  AOI22_X1 U27 ( .A1(n685), .A2(Q[83]), .B1(n684), .B2(Q[179]), .ZN(n25) );
  AOI22_X1 U28 ( .A1(n687), .A2(Q[211]), .B1(n686), .B2(Q[51]), .ZN(n26) );
  NAND4_X1 U29 ( .A1(n23), .A2(n24), .A3(n25), .A4(n26), .ZN(n27) );
  AOI22_X1 U30 ( .A1(n656), .A2(Q[1011]), .B1(n655), .B2(Q[947]), .ZN(n28) );
  AOI22_X1 U31 ( .A1(n658), .A2(Q[979]), .B1(n657), .B2(Q[915]), .ZN(n29) );
  AOI222_X1 U32 ( .A1(n660), .A2(Q[819]), .B1(n661), .B2(Q[115]), .C1(n659), 
        .C2(Q[755]), .ZN(n30) );
  NAND3_X1 U33 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n31) );
  AOI22_X1 U34 ( .A1(n663), .A2(Q[851]), .B1(n662), .B2(Q[723]), .ZN(n32) );
  AOI22_X1 U35 ( .A1(n665), .A2(Q[787]), .B1(n664), .B2(Q[883]), .ZN(n33) );
  NAND4_X1 U36 ( .A1(n613), .A2(n614), .A3(n32), .A4(n33), .ZN(n34) );
  OR4_X1 U37 ( .A1(n22), .A2(n27), .A3(n31), .A4(n34), .ZN(Y[19]) );
  AOI22_X1 U38 ( .A1(n673), .A2(Q[498]), .B1(n672), .B2(Q[562]), .ZN(n35) );
  AOI22_X1 U39 ( .A1(n675), .A2(Q[658]), .B1(n674), .B2(Q[466]), .ZN(n36) );
  AOI22_X1 U40 ( .A1(n677), .A2(Q[370]), .B1(n676), .B2(Q[306]), .ZN(n37) );
  AOI22_X1 U41 ( .A1(n679), .A2(Q[402]), .B1(n678), .B2(Q[274]), .ZN(n38) );
  NAND4_X1 U42 ( .A1(n35), .A2(n36), .A3(n37), .A4(n38), .ZN(n39) );
  AOI22_X1 U43 ( .A1(n681), .A2(Q[338]), .B1(n680), .B2(Q[434]), .ZN(n40) );
  AOI22_X1 U44 ( .A1(n683), .A2(Q[242]), .B1(n682), .B2(Q[146]), .ZN(n41) );
  AOI22_X1 U45 ( .A1(n685), .A2(Q[82]), .B1(n684), .B2(Q[178]), .ZN(n42) );
  AOI22_X1 U46 ( .A1(n687), .A2(Q[210]), .B1(n686), .B2(Q[50]), .ZN(n43) );
  NAND4_X1 U47 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n44) );
  AOI22_X1 U48 ( .A1(n656), .A2(Q[1010]), .B1(n655), .B2(Q[946]), .ZN(n45) );
  AOI22_X1 U49 ( .A1(n658), .A2(Q[978]), .B1(n657), .B2(Q[914]), .ZN(n46) );
  AOI222_X1 U50 ( .A1(n660), .A2(Q[818]), .B1(n661), .B2(Q[114]), .C1(n659), 
        .C2(Q[754]), .ZN(n47) );
  NAND3_X1 U51 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n48) );
  AOI22_X1 U52 ( .A1(n663), .A2(Q[850]), .B1(n662), .B2(Q[722]), .ZN(n49) );
  AOI22_X1 U53 ( .A1(n665), .A2(Q[786]), .B1(n664), .B2(Q[882]), .ZN(n50) );
  NAND4_X1 U54 ( .A1(n611), .A2(n612), .A3(n49), .A4(n50), .ZN(n51) );
  OR4_X1 U55 ( .A1(n39), .A2(n44), .A3(n48), .A4(n51), .ZN(Y[18]) );
  AOI22_X1 U56 ( .A1(n673), .A2(Q[497]), .B1(n672), .B2(Q[561]), .ZN(n52) );
  AOI22_X1 U57 ( .A1(n675), .A2(Q[657]), .B1(n674), .B2(Q[465]), .ZN(n53) );
  AOI22_X1 U58 ( .A1(n677), .A2(Q[369]), .B1(n676), .B2(Q[305]), .ZN(n54) );
  AOI22_X1 U59 ( .A1(n679), .A2(Q[401]), .B1(n678), .B2(Q[273]), .ZN(n55) );
  NAND4_X1 U60 ( .A1(n52), .A2(n53), .A3(n54), .A4(n55), .ZN(n56) );
  AOI22_X1 U61 ( .A1(n681), .A2(Q[337]), .B1(n680), .B2(Q[433]), .ZN(n57) );
  AOI22_X1 U62 ( .A1(n683), .A2(Q[241]), .B1(n682), .B2(Q[145]), .ZN(n58) );
  AOI22_X1 U63 ( .A1(n685), .A2(Q[81]), .B1(n684), .B2(Q[177]), .ZN(n59) );
  AOI22_X1 U64 ( .A1(n687), .A2(Q[209]), .B1(n686), .B2(Q[49]), .ZN(n60) );
  NAND4_X1 U65 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(n61) );
  AOI22_X1 U66 ( .A1(n656), .A2(Q[1009]), .B1(n655), .B2(Q[945]), .ZN(n62) );
  AOI22_X1 U67 ( .A1(n658), .A2(Q[977]), .B1(n657), .B2(Q[913]), .ZN(n63) );
  AOI222_X1 U68 ( .A1(n660), .A2(Q[817]), .B1(n661), .B2(Q[113]), .C1(n659), 
        .C2(Q[753]), .ZN(n64) );
  NAND3_X1 U69 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n65) );
  AOI22_X1 U70 ( .A1(n663), .A2(Q[849]), .B1(n662), .B2(Q[721]), .ZN(n66) );
  AOI22_X1 U71 ( .A1(n665), .A2(Q[785]), .B1(n664), .B2(Q[881]), .ZN(n67) );
  NAND4_X1 U72 ( .A1(n609), .A2(n610), .A3(n66), .A4(n67), .ZN(n68) );
  OR4_X1 U73 ( .A1(n56), .A2(n61), .A3(n65), .A4(n68), .ZN(Y[17]) );
  AOI22_X1 U74 ( .A1(n673), .A2(Q[496]), .B1(n672), .B2(Q[560]), .ZN(n69) );
  AOI22_X1 U75 ( .A1(n675), .A2(Q[656]), .B1(n674), .B2(Q[464]), .ZN(n70) );
  AOI22_X1 U76 ( .A1(n677), .A2(Q[368]), .B1(n676), .B2(Q[304]), .ZN(n71) );
  AOI22_X1 U77 ( .A1(n679), .A2(Q[400]), .B1(n678), .B2(Q[272]), .ZN(n72) );
  NAND4_X1 U78 ( .A1(n69), .A2(n70), .A3(n71), .A4(n72), .ZN(n73) );
  AOI22_X1 U79 ( .A1(n681), .A2(Q[336]), .B1(n680), .B2(Q[432]), .ZN(n74) );
  AOI22_X1 U80 ( .A1(n683), .A2(Q[240]), .B1(n682), .B2(Q[144]), .ZN(n75) );
  AOI22_X1 U81 ( .A1(n685), .A2(Q[80]), .B1(n684), .B2(Q[176]), .ZN(n76) );
  AOI22_X1 U82 ( .A1(n687), .A2(Q[208]), .B1(n686), .B2(Q[48]), .ZN(n77) );
  NAND4_X1 U83 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(n78) );
  AOI22_X1 U84 ( .A1(n656), .A2(Q[1008]), .B1(n655), .B2(Q[944]), .ZN(n79) );
  AOI22_X1 U85 ( .A1(n658), .A2(Q[976]), .B1(n657), .B2(Q[912]), .ZN(n80) );
  AOI222_X1 U86 ( .A1(n660), .A2(Q[816]), .B1(n661), .B2(Q[112]), .C1(n659), 
        .C2(Q[752]), .ZN(n81) );
  NAND3_X1 U87 ( .A1(n79), .A2(n80), .A3(n81), .ZN(n82) );
  AOI22_X1 U88 ( .A1(n663), .A2(Q[848]), .B1(n662), .B2(Q[720]), .ZN(n83) );
  AOI22_X1 U89 ( .A1(n665), .A2(Q[784]), .B1(n664), .B2(Q[880]), .ZN(n84) );
  NAND4_X1 U90 ( .A1(n607), .A2(n608), .A3(n83), .A4(n84), .ZN(n85) );
  OR4_X1 U91 ( .A1(n73), .A2(n78), .A3(n82), .A4(n85), .ZN(Y[16]) );
  AOI22_X1 U92 ( .A1(n673), .A2(Q[495]), .B1(n672), .B2(Q[559]), .ZN(n86) );
  AOI22_X1 U93 ( .A1(n675), .A2(Q[655]), .B1(n674), .B2(Q[463]), .ZN(n87) );
  AOI22_X1 U94 ( .A1(n677), .A2(Q[367]), .B1(n676), .B2(Q[303]), .ZN(n88) );
  AOI22_X1 U95 ( .A1(n679), .A2(Q[399]), .B1(n678), .B2(Q[271]), .ZN(n89) );
  NAND4_X1 U96 ( .A1(n86), .A2(n87), .A3(n88), .A4(n89), .ZN(n90) );
  AOI22_X1 U97 ( .A1(n681), .A2(Q[335]), .B1(n680), .B2(Q[431]), .ZN(n91) );
  AOI22_X1 U98 ( .A1(n683), .A2(Q[239]), .B1(n682), .B2(Q[143]), .ZN(n92) );
  AOI22_X1 U99 ( .A1(n685), .A2(Q[79]), .B1(n684), .B2(Q[175]), .ZN(n93) );
  AOI22_X1 U100 ( .A1(n687), .A2(Q[207]), .B1(n686), .B2(Q[47]), .ZN(n94) );
  NAND4_X1 U101 ( .A1(n91), .A2(n92), .A3(n93), .A4(n94), .ZN(n95) );
  AOI22_X1 U102 ( .A1(n656), .A2(Q[1007]), .B1(n655), .B2(Q[943]), .ZN(n96) );
  AOI22_X1 U103 ( .A1(n658), .A2(Q[975]), .B1(n657), .B2(Q[911]), .ZN(n97) );
  AOI222_X1 U104 ( .A1(n660), .A2(Q[815]), .B1(n661), .B2(Q[111]), .C1(n659), 
        .C2(Q[751]), .ZN(n98) );
  NAND3_X1 U105 ( .A1(n96), .A2(n97), .A3(n98), .ZN(n99) );
  AOI22_X1 U106 ( .A1(n663), .A2(Q[847]), .B1(n662), .B2(Q[719]), .ZN(n100) );
  AOI22_X1 U107 ( .A1(n665), .A2(Q[783]), .B1(n664), .B2(Q[879]), .ZN(n101) );
  NAND4_X1 U108 ( .A1(n605), .A2(n606), .A3(n100), .A4(n101), .ZN(n102) );
  OR4_X1 U109 ( .A1(n90), .A2(n95), .A3(n99), .A4(n102), .ZN(Y[15]) );
  AOI22_X1 U110 ( .A1(n673), .A2(Q[494]), .B1(n672), .B2(Q[558]), .ZN(n103) );
  AOI22_X1 U111 ( .A1(n675), .A2(Q[654]), .B1(n674), .B2(Q[462]), .ZN(n104) );
  AOI22_X1 U112 ( .A1(n677), .A2(Q[366]), .B1(n676), .B2(Q[302]), .ZN(n105) );
  AOI22_X1 U113 ( .A1(n679), .A2(Q[398]), .B1(n678), .B2(Q[270]), .ZN(n106) );
  NAND4_X1 U114 ( .A1(n103), .A2(n104), .A3(n105), .A4(n106), .ZN(n107) );
  AOI22_X1 U115 ( .A1(n681), .A2(Q[334]), .B1(n680), .B2(Q[430]), .ZN(n108) );
  AOI22_X1 U116 ( .A1(n683), .A2(Q[238]), .B1(n682), .B2(Q[142]), .ZN(n109) );
  AOI22_X1 U117 ( .A1(n685), .A2(Q[78]), .B1(n684), .B2(Q[174]), .ZN(n110) );
  AOI22_X1 U118 ( .A1(n687), .A2(Q[206]), .B1(n686), .B2(Q[46]), .ZN(n111) );
  NAND4_X1 U119 ( .A1(n108), .A2(n109), .A3(n110), .A4(n111), .ZN(n112) );
  AOI22_X1 U120 ( .A1(n656), .A2(Q[1006]), .B1(n655), .B2(Q[942]), .ZN(n113)
         );
  AOI22_X1 U121 ( .A1(n658), .A2(Q[974]), .B1(n657), .B2(Q[910]), .ZN(n114) );
  AOI222_X1 U122 ( .A1(n660), .A2(Q[814]), .B1(n661), .B2(Q[110]), .C1(n659), 
        .C2(Q[750]), .ZN(n115) );
  NAND3_X1 U123 ( .A1(n113), .A2(n114), .A3(n115), .ZN(n116) );
  AOI22_X1 U124 ( .A1(n663), .A2(Q[846]), .B1(n662), .B2(Q[718]), .ZN(n117) );
  AOI22_X1 U125 ( .A1(n665), .A2(Q[782]), .B1(n664), .B2(Q[878]), .ZN(n118) );
  NAND4_X1 U126 ( .A1(n603), .A2(n604), .A3(n117), .A4(n118), .ZN(n119) );
  OR4_X1 U127 ( .A1(n107), .A2(n112), .A3(n116), .A4(n119), .ZN(Y[14]) );
  AOI22_X1 U128 ( .A1(n673), .A2(Q[493]), .B1(n672), .B2(Q[557]), .ZN(n120) );
  AOI22_X1 U129 ( .A1(n675), .A2(Q[653]), .B1(n674), .B2(Q[461]), .ZN(n121) );
  AOI22_X1 U130 ( .A1(n677), .A2(Q[365]), .B1(n676), .B2(Q[301]), .ZN(n122) );
  AOI22_X1 U131 ( .A1(n679), .A2(Q[397]), .B1(n678), .B2(Q[269]), .ZN(n123) );
  NAND4_X1 U132 ( .A1(n120), .A2(n121), .A3(n122), .A4(n123), .ZN(n124) );
  AOI22_X1 U133 ( .A1(n681), .A2(Q[333]), .B1(n680), .B2(Q[429]), .ZN(n125) );
  AOI22_X1 U134 ( .A1(n683), .A2(Q[237]), .B1(n682), .B2(Q[141]), .ZN(n126) );
  AOI22_X1 U135 ( .A1(n685), .A2(Q[77]), .B1(n684), .B2(Q[173]), .ZN(n127) );
  AOI22_X1 U136 ( .A1(n687), .A2(Q[205]), .B1(n686), .B2(Q[45]), .ZN(n128) );
  NAND4_X1 U137 ( .A1(n125), .A2(n126), .A3(n127), .A4(n128), .ZN(n129) );
  AOI22_X1 U138 ( .A1(n656), .A2(Q[1005]), .B1(n655), .B2(Q[941]), .ZN(n130)
         );
  AOI22_X1 U139 ( .A1(n658), .A2(Q[973]), .B1(n657), .B2(Q[909]), .ZN(n131) );
  AOI222_X1 U140 ( .A1(n660), .A2(Q[813]), .B1(n661), .B2(Q[109]), .C1(n659), 
        .C2(Q[749]), .ZN(n132) );
  NAND3_X1 U141 ( .A1(n130), .A2(n131), .A3(n132), .ZN(n133) );
  AOI22_X1 U142 ( .A1(n663), .A2(Q[845]), .B1(n662), .B2(Q[717]), .ZN(n134) );
  AOI22_X1 U143 ( .A1(n665), .A2(Q[781]), .B1(n664), .B2(Q[877]), .ZN(n135) );
  NAND4_X1 U144 ( .A1(n601), .A2(n602), .A3(n134), .A4(n135), .ZN(n136) );
  OR4_X1 U145 ( .A1(n124), .A2(n129), .A3(n133), .A4(n136), .ZN(Y[13]) );
  AOI22_X1 U146 ( .A1(n673), .A2(Q[492]), .B1(n672), .B2(Q[556]), .ZN(n137) );
  AOI22_X1 U147 ( .A1(n675), .A2(Q[652]), .B1(n674), .B2(Q[460]), .ZN(n138) );
  AOI22_X1 U148 ( .A1(n677), .A2(Q[364]), .B1(n676), .B2(Q[300]), .ZN(n139) );
  AOI22_X1 U149 ( .A1(n679), .A2(Q[396]), .B1(n678), .B2(Q[268]), .ZN(n140) );
  NAND4_X1 U150 ( .A1(n137), .A2(n138), .A3(n139), .A4(n140), .ZN(n141) );
  AOI22_X1 U151 ( .A1(n681), .A2(Q[332]), .B1(n680), .B2(Q[428]), .ZN(n142) );
  AOI22_X1 U152 ( .A1(n683), .A2(Q[236]), .B1(n682), .B2(Q[140]), .ZN(n143) );
  AOI22_X1 U153 ( .A1(n685), .A2(Q[76]), .B1(n684), .B2(Q[172]), .ZN(n144) );
  AOI22_X1 U154 ( .A1(n687), .A2(Q[204]), .B1(n686), .B2(Q[44]), .ZN(n145) );
  NAND4_X1 U155 ( .A1(n142), .A2(n143), .A3(n144), .A4(n145), .ZN(n146) );
  AOI22_X1 U156 ( .A1(n656), .A2(Q[1004]), .B1(n655), .B2(Q[940]), .ZN(n147)
         );
  AOI22_X1 U157 ( .A1(n658), .A2(Q[972]), .B1(n657), .B2(Q[908]), .ZN(n148) );
  AOI222_X1 U158 ( .A1(n660), .A2(Q[812]), .B1(n661), .B2(Q[108]), .C1(n659), 
        .C2(Q[748]), .ZN(n149) );
  NAND3_X1 U159 ( .A1(n147), .A2(n148), .A3(n149), .ZN(n150) );
  AOI22_X1 U160 ( .A1(n663), .A2(Q[844]), .B1(n662), .B2(Q[716]), .ZN(n151) );
  AOI22_X1 U161 ( .A1(n665), .A2(Q[780]), .B1(n664), .B2(Q[876]), .ZN(n152) );
  NAND4_X1 U162 ( .A1(n599), .A2(n600), .A3(n151), .A4(n152), .ZN(n153) );
  OR4_X1 U163 ( .A1(n141), .A2(n146), .A3(n150), .A4(n153), .ZN(Y[12]) );
  AOI22_X1 U164 ( .A1(n561), .A2(Q[511]), .B1(n560), .B2(Q[575]), .ZN(n154) );
  AOI22_X1 U165 ( .A1(n563), .A2(Q[671]), .B1(n562), .B2(Q[479]), .ZN(n155) );
  AOI22_X1 U166 ( .A1(n565), .A2(Q[383]), .B1(n564), .B2(Q[319]), .ZN(n156) );
  AOI22_X1 U167 ( .A1(n567), .A2(Q[415]), .B1(n566), .B2(Q[287]), .ZN(n157) );
  NAND4_X1 U168 ( .A1(n154), .A2(n155), .A3(n156), .A4(n157), .ZN(n158) );
  AOI22_X1 U169 ( .A1(n569), .A2(Q[351]), .B1(n568), .B2(Q[447]), .ZN(n159) );
  AOI22_X1 U170 ( .A1(n571), .A2(Q[255]), .B1(n570), .B2(Q[159]), .ZN(n160) );
  AOI22_X1 U171 ( .A1(n573), .A2(Q[95]), .B1(n572), .B2(Q[191]), .ZN(n161) );
  AOI22_X1 U172 ( .A1(n575), .A2(Q[223]), .B1(n574), .B2(Q[63]), .ZN(n162) );
  NAND4_X1 U173 ( .A1(n159), .A2(n160), .A3(n161), .A4(n162), .ZN(n163) );
  AOI22_X1 U174 ( .A1(n546), .A2(Q[1023]), .B1(n545), .B2(Q[959]), .ZN(n164)
         );
  AOI22_X1 U175 ( .A1(n548), .A2(Q[991]), .B1(n547), .B2(Q[927]), .ZN(n165) );
  AOI222_X1 U176 ( .A1(n550), .A2(Q[831]), .B1(n551), .B2(Q[127]), .C1(n549), 
        .C2(Q[767]), .ZN(n166) );
  NAND3_X1 U177 ( .A1(n164), .A2(n165), .A3(n166), .ZN(n167) );
  AOI22_X1 U178 ( .A1(n553), .A2(Q[863]), .B1(n552), .B2(Q[735]), .ZN(n168) );
  AOI22_X1 U179 ( .A1(n555), .A2(Q[799]), .B1(n554), .B2(Q[895]), .ZN(n169) );
  NAND4_X1 U180 ( .A1(n641), .A2(n642), .A3(n168), .A4(n169), .ZN(n170) );
  OR4_X1 U181 ( .A1(n158), .A2(n163), .A3(n167), .A4(n170), .ZN(Y[31]) );
  AOI22_X1 U182 ( .A1(n561), .A2(Q[510]), .B1(n560), .B2(Q[574]), .ZN(n171) );
  AOI22_X1 U183 ( .A1(n563), .A2(Q[670]), .B1(n562), .B2(Q[478]), .ZN(n172) );
  AOI22_X1 U184 ( .A1(n565), .A2(Q[382]), .B1(n564), .B2(Q[318]), .ZN(n173) );
  AOI22_X1 U185 ( .A1(n567), .A2(Q[414]), .B1(n566), .B2(Q[286]), .ZN(n174) );
  NAND4_X1 U186 ( .A1(n171), .A2(n172), .A3(n173), .A4(n174), .ZN(n175) );
  AOI22_X1 U187 ( .A1(n569), .A2(Q[350]), .B1(n568), .B2(Q[446]), .ZN(n176) );
  AOI22_X1 U188 ( .A1(n571), .A2(Q[254]), .B1(n570), .B2(Q[158]), .ZN(n177) );
  AOI22_X1 U189 ( .A1(n573), .A2(Q[94]), .B1(n572), .B2(Q[190]), .ZN(n178) );
  AOI22_X1 U190 ( .A1(n575), .A2(Q[222]), .B1(n574), .B2(Q[62]), .ZN(n179) );
  NAND4_X1 U191 ( .A1(n176), .A2(n177), .A3(n178), .A4(n179), .ZN(n180) );
  AOI22_X1 U192 ( .A1(n546), .A2(Q[1022]), .B1(n545), .B2(Q[958]), .ZN(n181)
         );
  AOI22_X1 U193 ( .A1(n548), .A2(Q[990]), .B1(n547), .B2(Q[926]), .ZN(n182) );
  AOI222_X1 U194 ( .A1(n550), .A2(Q[830]), .B1(n551), .B2(Q[126]), .C1(n549), 
        .C2(Q[766]), .ZN(n183) );
  NAND3_X1 U195 ( .A1(n181), .A2(n182), .A3(n183), .ZN(n184) );
  AOI22_X1 U196 ( .A1(n553), .A2(Q[862]), .B1(n552), .B2(Q[734]), .ZN(n185) );
  AOI22_X1 U197 ( .A1(n555), .A2(Q[798]), .B1(n554), .B2(Q[894]), .ZN(n186) );
  NAND4_X1 U198 ( .A1(n639), .A2(n640), .A3(n185), .A4(n186), .ZN(n187) );
  OR4_X1 U199 ( .A1(n175), .A2(n180), .A3(n184), .A4(n187), .ZN(Y[30]) );
  AOI22_X1 U200 ( .A1(n561), .A2(Q[508]), .B1(n560), .B2(Q[572]), .ZN(n188) );
  AOI22_X1 U201 ( .A1(n563), .A2(Q[668]), .B1(n562), .B2(Q[476]), .ZN(n189) );
  AOI22_X1 U202 ( .A1(n565), .A2(Q[380]), .B1(n564), .B2(Q[316]), .ZN(n190) );
  AOI22_X1 U203 ( .A1(n567), .A2(Q[412]), .B1(n566), .B2(Q[284]), .ZN(n191) );
  NAND4_X1 U204 ( .A1(n188), .A2(n189), .A3(n190), .A4(n191), .ZN(n192) );
  AOI22_X1 U205 ( .A1(n569), .A2(Q[348]), .B1(n568), .B2(Q[444]), .ZN(n193) );
  AOI22_X1 U206 ( .A1(n571), .A2(Q[252]), .B1(n570), .B2(Q[156]), .ZN(n194) );
  AOI22_X1 U207 ( .A1(n573), .A2(Q[92]), .B1(n572), .B2(Q[188]), .ZN(n195) );
  AOI22_X1 U208 ( .A1(n575), .A2(Q[220]), .B1(n574), .B2(Q[60]), .ZN(n196) );
  NAND4_X1 U209 ( .A1(n193), .A2(n194), .A3(n195), .A4(n196), .ZN(n197) );
  AOI22_X1 U210 ( .A1(n546), .A2(Q[1020]), .B1(n545), .B2(Q[956]), .ZN(n198)
         );
  AOI22_X1 U211 ( .A1(n548), .A2(Q[988]), .B1(n547), .B2(Q[924]), .ZN(n199) );
  AOI222_X1 U212 ( .A1(n550), .A2(Q[828]), .B1(n551), .B2(Q[124]), .C1(n549), 
        .C2(Q[764]), .ZN(n200) );
  NAND3_X1 U213 ( .A1(n198), .A2(n199), .A3(n200), .ZN(n201) );
  AOI22_X1 U214 ( .A1(n553), .A2(Q[860]), .B1(n552), .B2(Q[732]), .ZN(n202) );
  AOI22_X1 U215 ( .A1(n555), .A2(Q[796]), .B1(n554), .B2(Q[892]), .ZN(n203) );
  NAND4_X1 U216 ( .A1(n633), .A2(n634), .A3(n202), .A4(n203), .ZN(n204) );
  OR4_X1 U217 ( .A1(n192), .A2(n197), .A3(n201), .A4(n204), .ZN(Y[28]) );
  AOI22_X1 U218 ( .A1(n561), .A2(Q[507]), .B1(n560), .B2(Q[571]), .ZN(n205) );
  AOI22_X1 U219 ( .A1(n563), .A2(Q[667]), .B1(n562), .B2(Q[475]), .ZN(n206) );
  AOI22_X1 U220 ( .A1(n565), .A2(Q[379]), .B1(n564), .B2(Q[315]), .ZN(n207) );
  AOI22_X1 U221 ( .A1(n567), .A2(Q[411]), .B1(n566), .B2(Q[283]), .ZN(n208) );
  NAND4_X1 U222 ( .A1(n205), .A2(n206), .A3(n207), .A4(n208), .ZN(n209) );
  AOI22_X1 U223 ( .A1(n569), .A2(Q[347]), .B1(n568), .B2(Q[443]), .ZN(n210) );
  AOI22_X1 U224 ( .A1(n571), .A2(Q[251]), .B1(n570), .B2(Q[155]), .ZN(n211) );
  AOI22_X1 U225 ( .A1(n573), .A2(Q[91]), .B1(n572), .B2(Q[187]), .ZN(n212) );
  AOI22_X1 U226 ( .A1(n575), .A2(Q[219]), .B1(n574), .B2(Q[59]), .ZN(n213) );
  NAND4_X1 U227 ( .A1(n210), .A2(n211), .A3(n212), .A4(n213), .ZN(n214) );
  AOI22_X1 U228 ( .A1(n546), .A2(Q[1019]), .B1(n545), .B2(Q[955]), .ZN(n215)
         );
  AOI22_X1 U229 ( .A1(n548), .A2(Q[987]), .B1(n547), .B2(Q[923]), .ZN(n216) );
  AOI222_X1 U230 ( .A1(n550), .A2(Q[827]), .B1(n551), .B2(Q[123]), .C1(n549), 
        .C2(Q[763]), .ZN(n217) );
  NAND3_X1 U231 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n218) );
  AOI22_X1 U232 ( .A1(n553), .A2(Q[859]), .B1(n552), .B2(Q[731]), .ZN(n219) );
  AOI22_X1 U233 ( .A1(n555), .A2(Q[795]), .B1(n554), .B2(Q[891]), .ZN(n220) );
  NAND4_X1 U234 ( .A1(n631), .A2(n632), .A3(n219), .A4(n220), .ZN(n221) );
  OR4_X1 U235 ( .A1(n209), .A2(n214), .A3(n218), .A4(n221), .ZN(Y[27]) );
  AOI22_X1 U236 ( .A1(n561), .A2(Q[506]), .B1(n560), .B2(Q[570]), .ZN(n222) );
  AOI22_X1 U237 ( .A1(n563), .A2(Q[666]), .B1(n562), .B2(Q[474]), .ZN(n223) );
  AOI22_X1 U238 ( .A1(n565), .A2(Q[378]), .B1(n564), .B2(Q[314]), .ZN(n224) );
  AOI22_X1 U239 ( .A1(n567), .A2(Q[410]), .B1(n566), .B2(Q[282]), .ZN(n225) );
  NAND4_X1 U240 ( .A1(n222), .A2(n223), .A3(n224), .A4(n225), .ZN(n226) );
  AOI22_X1 U241 ( .A1(n569), .A2(Q[346]), .B1(n568), .B2(Q[442]), .ZN(n227) );
  AOI22_X1 U242 ( .A1(n571), .A2(Q[250]), .B1(n570), .B2(Q[154]), .ZN(n228) );
  AOI22_X1 U243 ( .A1(n573), .A2(Q[90]), .B1(n572), .B2(Q[186]), .ZN(n229) );
  AOI22_X1 U244 ( .A1(n575), .A2(Q[218]), .B1(n574), .B2(Q[58]), .ZN(n230) );
  NAND4_X1 U245 ( .A1(n227), .A2(n228), .A3(n229), .A4(n230), .ZN(n231) );
  AOI22_X1 U246 ( .A1(n546), .A2(Q[1018]), .B1(n545), .B2(Q[954]), .ZN(n232)
         );
  AOI22_X1 U247 ( .A1(n548), .A2(Q[986]), .B1(n547), .B2(Q[922]), .ZN(n233) );
  AOI222_X1 U248 ( .A1(n550), .A2(Q[826]), .B1(n551), .B2(Q[122]), .C1(n549), 
        .C2(Q[762]), .ZN(n234) );
  NAND3_X1 U249 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n235) );
  AOI22_X1 U250 ( .A1(n553), .A2(Q[858]), .B1(n552), .B2(Q[730]), .ZN(n236) );
  AOI22_X1 U251 ( .A1(n555), .A2(Q[794]), .B1(n554), .B2(Q[890]), .ZN(n237) );
  NAND4_X1 U252 ( .A1(n629), .A2(n630), .A3(n236), .A4(n237), .ZN(n238) );
  OR4_X1 U253 ( .A1(n226), .A2(n231), .A3(n235), .A4(n238), .ZN(Y[26]) );
  AOI22_X1 U254 ( .A1(n561), .A2(Q[505]), .B1(n560), .B2(Q[569]), .ZN(n239) );
  AOI22_X1 U255 ( .A1(n563), .A2(Q[665]), .B1(n562), .B2(Q[473]), .ZN(n240) );
  AOI22_X1 U256 ( .A1(n565), .A2(Q[377]), .B1(n564), .B2(Q[313]), .ZN(n241) );
  AOI22_X1 U257 ( .A1(n567), .A2(Q[409]), .B1(n566), .B2(Q[281]), .ZN(n242) );
  NAND4_X1 U258 ( .A1(n239), .A2(n240), .A3(n241), .A4(n242), .ZN(n243) );
  AOI22_X1 U259 ( .A1(n569), .A2(Q[345]), .B1(n568), .B2(Q[441]), .ZN(n244) );
  AOI22_X1 U260 ( .A1(n571), .A2(Q[249]), .B1(n570), .B2(Q[153]), .ZN(n245) );
  AOI22_X1 U261 ( .A1(n573), .A2(Q[89]), .B1(n572), .B2(Q[185]), .ZN(n246) );
  AOI22_X1 U262 ( .A1(n575), .A2(Q[217]), .B1(n574), .B2(Q[57]), .ZN(n247) );
  NAND4_X1 U263 ( .A1(n244), .A2(n245), .A3(n246), .A4(n247), .ZN(n248) );
  AOI22_X1 U264 ( .A1(n546), .A2(Q[1017]), .B1(n545), .B2(Q[953]), .ZN(n249)
         );
  AOI22_X1 U265 ( .A1(n548), .A2(Q[985]), .B1(n547), .B2(Q[921]), .ZN(n250) );
  AOI222_X1 U266 ( .A1(n550), .A2(Q[825]), .B1(n551), .B2(Q[121]), .C1(n549), 
        .C2(Q[761]), .ZN(n251) );
  NAND3_X1 U267 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n252) );
  AOI22_X1 U268 ( .A1(n553), .A2(Q[857]), .B1(n552), .B2(Q[729]), .ZN(n253) );
  AOI22_X1 U269 ( .A1(n555), .A2(Q[793]), .B1(n554), .B2(Q[889]), .ZN(n254) );
  NAND4_X1 U270 ( .A1(n627), .A2(n628), .A3(n253), .A4(n254), .ZN(n255) );
  OR4_X1 U271 ( .A1(n243), .A2(n248), .A3(n252), .A4(n255), .ZN(Y[25]) );
  AOI22_X1 U272 ( .A1(n561), .A2(Q[504]), .B1(n560), .B2(Q[568]), .ZN(n256) );
  AOI22_X1 U273 ( .A1(n563), .A2(Q[664]), .B1(n562), .B2(Q[472]), .ZN(n257) );
  AOI22_X1 U274 ( .A1(n565), .A2(Q[376]), .B1(n564), .B2(Q[312]), .ZN(n258) );
  AOI22_X1 U275 ( .A1(n567), .A2(Q[408]), .B1(n566), .B2(Q[280]), .ZN(n259) );
  NAND4_X1 U276 ( .A1(n256), .A2(n257), .A3(n258), .A4(n259), .ZN(n260) );
  AOI22_X1 U277 ( .A1(n569), .A2(Q[344]), .B1(n568), .B2(Q[440]), .ZN(n261) );
  AOI22_X1 U278 ( .A1(n571), .A2(Q[248]), .B1(n570), .B2(Q[152]), .ZN(n262) );
  AOI22_X1 U279 ( .A1(n573), .A2(Q[88]), .B1(n572), .B2(Q[184]), .ZN(n263) );
  AOI22_X1 U280 ( .A1(n575), .A2(Q[216]), .B1(n574), .B2(Q[56]), .ZN(n264) );
  NAND4_X1 U281 ( .A1(n261), .A2(n262), .A3(n263), .A4(n264), .ZN(n265) );
  AOI22_X1 U282 ( .A1(n546), .A2(Q[1016]), .B1(n545), .B2(Q[952]), .ZN(n266)
         );
  AOI22_X1 U283 ( .A1(n548), .A2(Q[984]), .B1(n547), .B2(Q[920]), .ZN(n267) );
  AOI222_X1 U284 ( .A1(n550), .A2(Q[824]), .B1(n551), .B2(Q[120]), .C1(n549), 
        .C2(Q[760]), .ZN(n268) );
  NAND3_X1 U285 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n269) );
  AOI22_X1 U286 ( .A1(n553), .A2(Q[856]), .B1(n552), .B2(Q[728]), .ZN(n270) );
  AOI22_X1 U287 ( .A1(n555), .A2(Q[792]), .B1(n554), .B2(Q[888]), .ZN(n271) );
  NAND4_X1 U288 ( .A1(n625), .A2(n626), .A3(n270), .A4(n271), .ZN(n272) );
  OR4_X1 U289 ( .A1(n260), .A2(n265), .A3(n269), .A4(n272), .ZN(Y[24]) );
  AOI22_X1 U290 ( .A1(n561), .A2(Q[503]), .B1(n560), .B2(Q[567]), .ZN(n273) );
  AOI22_X1 U291 ( .A1(n563), .A2(Q[663]), .B1(n562), .B2(Q[471]), .ZN(n274) );
  AOI22_X1 U292 ( .A1(n565), .A2(Q[375]), .B1(n564), .B2(Q[311]), .ZN(n275) );
  AOI22_X1 U293 ( .A1(n567), .A2(Q[407]), .B1(n566), .B2(Q[279]), .ZN(n276) );
  NAND4_X1 U294 ( .A1(n273), .A2(n274), .A3(n275), .A4(n276), .ZN(n277) );
  AOI22_X1 U295 ( .A1(n569), .A2(Q[343]), .B1(n568), .B2(Q[439]), .ZN(n278) );
  AOI22_X1 U296 ( .A1(n571), .A2(Q[247]), .B1(n570), .B2(Q[151]), .ZN(n279) );
  AOI22_X1 U297 ( .A1(n573), .A2(Q[87]), .B1(n572), .B2(Q[183]), .ZN(n280) );
  AOI22_X1 U298 ( .A1(n575), .A2(Q[215]), .B1(n574), .B2(Q[55]), .ZN(n281) );
  NAND4_X1 U299 ( .A1(n278), .A2(n279), .A3(n280), .A4(n281), .ZN(n282) );
  AOI22_X1 U300 ( .A1(n546), .A2(Q[1015]), .B1(n545), .B2(Q[951]), .ZN(n283)
         );
  AOI22_X1 U301 ( .A1(n548), .A2(Q[983]), .B1(n547), .B2(Q[919]), .ZN(n284) );
  AOI222_X1 U302 ( .A1(n550), .A2(Q[823]), .B1(n551), .B2(Q[119]), .C1(n549), 
        .C2(Q[759]), .ZN(n285) );
  NAND3_X1 U303 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n286) );
  AOI22_X1 U304 ( .A1(n553), .A2(Q[855]), .B1(n552), .B2(Q[727]), .ZN(n287) );
  AOI22_X1 U305 ( .A1(n555), .A2(Q[791]), .B1(n554), .B2(Q[887]), .ZN(n288) );
  NAND4_X1 U306 ( .A1(n623), .A2(n624), .A3(n287), .A4(n288), .ZN(n289) );
  OR4_X1 U307 ( .A1(n277), .A2(n282), .A3(n286), .A4(n289), .ZN(Y[23]) );
  AOI22_X1 U308 ( .A1(n561), .A2(Q[502]), .B1(n560), .B2(Q[566]), .ZN(n290) );
  AOI22_X1 U309 ( .A1(n563), .A2(Q[662]), .B1(n562), .B2(Q[470]), .ZN(n291) );
  AOI22_X1 U310 ( .A1(n565), .A2(Q[374]), .B1(n564), .B2(Q[310]), .ZN(n292) );
  AOI22_X1 U311 ( .A1(n567), .A2(Q[406]), .B1(n566), .B2(Q[278]), .ZN(n293) );
  NAND4_X1 U312 ( .A1(n290), .A2(n291), .A3(n292), .A4(n293), .ZN(n294) );
  AOI22_X1 U313 ( .A1(n569), .A2(Q[342]), .B1(n568), .B2(Q[438]), .ZN(n295) );
  AOI22_X1 U314 ( .A1(n571), .A2(Q[246]), .B1(n570), .B2(Q[150]), .ZN(n296) );
  AOI22_X1 U315 ( .A1(n573), .A2(Q[86]), .B1(n572), .B2(Q[182]), .ZN(n297) );
  AOI22_X1 U316 ( .A1(n575), .A2(Q[214]), .B1(n574), .B2(Q[54]), .ZN(n298) );
  NAND4_X1 U317 ( .A1(n295), .A2(n296), .A3(n297), .A4(n298), .ZN(n299) );
  AOI22_X1 U318 ( .A1(n546), .A2(Q[1014]), .B1(n545), .B2(Q[950]), .ZN(n300)
         );
  AOI22_X1 U319 ( .A1(n548), .A2(Q[982]), .B1(n547), .B2(Q[918]), .ZN(n301) );
  AOI222_X1 U320 ( .A1(n550), .A2(Q[822]), .B1(n551), .B2(Q[118]), .C1(n549), 
        .C2(Q[758]), .ZN(n302) );
  NAND3_X1 U321 ( .A1(n300), .A2(n301), .A3(n302), .ZN(n303) );
  AOI22_X1 U322 ( .A1(n553), .A2(Q[854]), .B1(n552), .B2(Q[726]), .ZN(n304) );
  AOI22_X1 U323 ( .A1(n555), .A2(Q[790]), .B1(n554), .B2(Q[886]), .ZN(n305) );
  NAND4_X1 U324 ( .A1(n621), .A2(n622), .A3(n304), .A4(n305), .ZN(n306) );
  OR4_X1 U325 ( .A1(n294), .A2(n299), .A3(n303), .A4(n306), .ZN(Y[22]) );
  AOI22_X1 U326 ( .A1(n561), .A2(Q[501]), .B1(n560), .B2(Q[565]), .ZN(n307) );
  AOI22_X1 U327 ( .A1(n563), .A2(Q[661]), .B1(n562), .B2(Q[469]), .ZN(n308) );
  AOI22_X1 U328 ( .A1(n565), .A2(Q[373]), .B1(n564), .B2(Q[309]), .ZN(n309) );
  AOI22_X1 U329 ( .A1(n567), .A2(Q[405]), .B1(n566), .B2(Q[277]), .ZN(n310) );
  NAND4_X1 U330 ( .A1(n307), .A2(n308), .A3(n309), .A4(n310), .ZN(n311) );
  AOI22_X1 U331 ( .A1(n569), .A2(Q[341]), .B1(n568), .B2(Q[437]), .ZN(n312) );
  AOI22_X1 U332 ( .A1(n571), .A2(Q[245]), .B1(n570), .B2(Q[149]), .ZN(n313) );
  AOI22_X1 U333 ( .A1(n573), .A2(Q[85]), .B1(n572), .B2(Q[181]), .ZN(n314) );
  AOI22_X1 U334 ( .A1(n575), .A2(Q[213]), .B1(n574), .B2(Q[53]), .ZN(n315) );
  NAND4_X1 U335 ( .A1(n312), .A2(n313), .A3(n314), .A4(n315), .ZN(n316) );
  AOI22_X1 U336 ( .A1(n546), .A2(Q[1013]), .B1(n545), .B2(Q[949]), .ZN(n317)
         );
  AOI22_X1 U337 ( .A1(n548), .A2(Q[981]), .B1(n547), .B2(Q[917]), .ZN(n318) );
  AOI222_X1 U338 ( .A1(n550), .A2(Q[821]), .B1(n551), .B2(Q[117]), .C1(n549), 
        .C2(Q[757]), .ZN(n319) );
  NAND3_X1 U339 ( .A1(n317), .A2(n318), .A3(n319), .ZN(n320) );
  AOI22_X1 U340 ( .A1(n553), .A2(Q[853]), .B1(n552), .B2(Q[725]), .ZN(n321) );
  AOI22_X1 U341 ( .A1(n555), .A2(Q[789]), .B1(n554), .B2(Q[885]), .ZN(n322) );
  NAND4_X1 U342 ( .A1(n619), .A2(n620), .A3(n321), .A4(n322), .ZN(n323) );
  OR4_X1 U343 ( .A1(n311), .A2(n316), .A3(n320), .A4(n323), .ZN(Y[21]) );
  AOI22_X1 U344 ( .A1(n561), .A2(Q[500]), .B1(n560), .B2(Q[564]), .ZN(n324) );
  AOI22_X1 U345 ( .A1(n563), .A2(Q[660]), .B1(n562), .B2(Q[468]), .ZN(n325) );
  AOI22_X1 U346 ( .A1(n565), .A2(Q[372]), .B1(n564), .B2(Q[308]), .ZN(n326) );
  AOI22_X1 U347 ( .A1(n567), .A2(Q[404]), .B1(n566), .B2(Q[276]), .ZN(n327) );
  NAND4_X1 U348 ( .A1(n324), .A2(n325), .A3(n326), .A4(n327), .ZN(n328) );
  AOI22_X1 U349 ( .A1(n569), .A2(Q[340]), .B1(n568), .B2(Q[436]), .ZN(n329) );
  AOI22_X1 U350 ( .A1(n571), .A2(Q[244]), .B1(n570), .B2(Q[148]), .ZN(n330) );
  AOI22_X1 U351 ( .A1(n573), .A2(Q[84]), .B1(n572), .B2(Q[180]), .ZN(n331) );
  AOI22_X1 U352 ( .A1(n575), .A2(Q[212]), .B1(n574), .B2(Q[52]), .ZN(n332) );
  NAND4_X1 U353 ( .A1(n329), .A2(n330), .A3(n331), .A4(n332), .ZN(n333) );
  AOI22_X1 U354 ( .A1(n546), .A2(Q[1012]), .B1(n545), .B2(Q[948]), .ZN(n334)
         );
  AOI22_X1 U355 ( .A1(n548), .A2(Q[980]), .B1(n547), .B2(Q[916]), .ZN(n335) );
  AOI222_X1 U356 ( .A1(n550), .A2(Q[820]), .B1(n551), .B2(Q[116]), .C1(n549), 
        .C2(Q[756]), .ZN(n336) );
  NAND3_X1 U357 ( .A1(n334), .A2(n335), .A3(n336), .ZN(n337) );
  AOI22_X1 U358 ( .A1(n553), .A2(Q[852]), .B1(n552), .B2(Q[724]), .ZN(n338) );
  AOI22_X1 U359 ( .A1(n555), .A2(Q[788]), .B1(n554), .B2(Q[884]), .ZN(n339) );
  NAND4_X1 U360 ( .A1(n617), .A2(n618), .A3(n338), .A4(n339), .ZN(n340) );
  OR4_X1 U361 ( .A1(n328), .A2(n333), .A3(n337), .A4(n340), .ZN(Y[20]) );
  AOI22_X1 U362 ( .A1(n673), .A2(Q[491]), .B1(n672), .B2(Q[555]), .ZN(n341) );
  AOI22_X1 U363 ( .A1(n675), .A2(Q[651]), .B1(n674), .B2(Q[459]), .ZN(n342) );
  AOI22_X1 U364 ( .A1(n677), .A2(Q[363]), .B1(n676), .B2(Q[299]), .ZN(n343) );
  AOI22_X1 U365 ( .A1(n679), .A2(Q[395]), .B1(n678), .B2(Q[267]), .ZN(n344) );
  NAND4_X1 U366 ( .A1(n341), .A2(n342), .A3(n343), .A4(n344), .ZN(n345) );
  AOI22_X1 U367 ( .A1(n681), .A2(Q[331]), .B1(n680), .B2(Q[427]), .ZN(n346) );
  AOI22_X1 U368 ( .A1(n683), .A2(Q[235]), .B1(n682), .B2(Q[139]), .ZN(n347) );
  AOI22_X1 U369 ( .A1(n685), .A2(Q[75]), .B1(n684), .B2(Q[171]), .ZN(n348) );
  AOI22_X1 U370 ( .A1(n687), .A2(Q[203]), .B1(n686), .B2(Q[43]), .ZN(n349) );
  NAND4_X1 U371 ( .A1(n346), .A2(n347), .A3(n348), .A4(n349), .ZN(n350) );
  AOI22_X1 U372 ( .A1(n656), .A2(Q[1003]), .B1(n655), .B2(Q[939]), .ZN(n351)
         );
  AOI22_X1 U373 ( .A1(n658), .A2(Q[971]), .B1(n657), .B2(Q[907]), .ZN(n352) );
  AOI222_X1 U374 ( .A1(n660), .A2(Q[811]), .B1(n661), .B2(Q[107]), .C1(n659), 
        .C2(Q[747]), .ZN(n353) );
  NAND3_X1 U375 ( .A1(n351), .A2(n352), .A3(n353), .ZN(n354) );
  AOI22_X1 U376 ( .A1(n663), .A2(Q[843]), .B1(n662), .B2(Q[715]), .ZN(n355) );
  AOI22_X1 U377 ( .A1(n665), .A2(Q[779]), .B1(n664), .B2(Q[875]), .ZN(n356) );
  NAND4_X1 U378 ( .A1(n597), .A2(n598), .A3(n355), .A4(n356), .ZN(n357) );
  OR4_X1 U379 ( .A1(n345), .A2(n350), .A3(n354), .A4(n357), .ZN(Y[11]) );
  AOI22_X1 U380 ( .A1(n561), .A2(Q[490]), .B1(n560), .B2(Q[554]), .ZN(n358) );
  AOI22_X1 U381 ( .A1(n563), .A2(Q[650]), .B1(n562), .B2(Q[458]), .ZN(n359) );
  AOI22_X1 U382 ( .A1(n565), .A2(Q[362]), .B1(n564), .B2(Q[298]), .ZN(n360) );
  AOI22_X1 U383 ( .A1(n567), .A2(Q[394]), .B1(n566), .B2(Q[266]), .ZN(n361) );
  NAND4_X1 U384 ( .A1(n358), .A2(n359), .A3(n360), .A4(n361), .ZN(n362) );
  AOI22_X1 U385 ( .A1(n569), .A2(Q[330]), .B1(n568), .B2(Q[426]), .ZN(n363) );
  AOI22_X1 U386 ( .A1(n571), .A2(Q[234]), .B1(n570), .B2(Q[138]), .ZN(n364) );
  AOI22_X1 U387 ( .A1(n573), .A2(Q[74]), .B1(n572), .B2(Q[170]), .ZN(n365) );
  AOI22_X1 U388 ( .A1(n575), .A2(Q[202]), .B1(n574), .B2(Q[42]), .ZN(n366) );
  NAND4_X1 U389 ( .A1(n363), .A2(n364), .A3(n365), .A4(n366), .ZN(n367) );
  AOI22_X1 U390 ( .A1(n546), .A2(Q[1002]), .B1(n545), .B2(Q[938]), .ZN(n368)
         );
  AOI22_X1 U391 ( .A1(n548), .A2(Q[970]), .B1(n547), .B2(Q[906]), .ZN(n369) );
  AOI222_X1 U392 ( .A1(n550), .A2(Q[810]), .B1(n551), .B2(Q[106]), .C1(n549), 
        .C2(Q[746]), .ZN(n370) );
  NAND3_X1 U393 ( .A1(n368), .A2(n369), .A3(n370), .ZN(n371) );
  AOI22_X1 U394 ( .A1(n553), .A2(Q[842]), .B1(n552), .B2(Q[714]), .ZN(n372) );
  AOI22_X1 U395 ( .A1(n555), .A2(Q[778]), .B1(n554), .B2(Q[874]), .ZN(n373) );
  NAND4_X1 U396 ( .A1(n595), .A2(n596), .A3(n372), .A4(n373), .ZN(n374) );
  OR4_X1 U397 ( .A1(n362), .A2(n367), .A3(n371), .A4(n374), .ZN(Y[10]) );
  AOI22_X1 U398 ( .A1(n561), .A2(Q[489]), .B1(n560), .B2(Q[553]), .ZN(n375) );
  AOI22_X1 U399 ( .A1(n563), .A2(Q[649]), .B1(n562), .B2(Q[457]), .ZN(n376) );
  AOI22_X1 U400 ( .A1(n565), .A2(Q[361]), .B1(n564), .B2(Q[297]), .ZN(n377) );
  AOI22_X1 U401 ( .A1(n567), .A2(Q[393]), .B1(n566), .B2(Q[265]), .ZN(n378) );
  NAND4_X1 U402 ( .A1(n375), .A2(n376), .A3(n377), .A4(n378), .ZN(n379) );
  AOI22_X1 U403 ( .A1(n569), .A2(Q[329]), .B1(n568), .B2(Q[425]), .ZN(n380) );
  AOI22_X1 U404 ( .A1(n571), .A2(Q[233]), .B1(n570), .B2(Q[137]), .ZN(n381) );
  AOI22_X1 U405 ( .A1(n573), .A2(Q[73]), .B1(n572), .B2(Q[169]), .ZN(n382) );
  AOI22_X1 U406 ( .A1(n575), .A2(Q[201]), .B1(n574), .B2(Q[41]), .ZN(n383) );
  NAND4_X1 U407 ( .A1(n380), .A2(n381), .A3(n382), .A4(n383), .ZN(n384) );
  AOI22_X1 U408 ( .A1(n546), .A2(Q[1001]), .B1(n545), .B2(Q[937]), .ZN(n385)
         );
  AOI22_X1 U409 ( .A1(n548), .A2(Q[969]), .B1(n547), .B2(Q[905]), .ZN(n386) );
  AOI222_X1 U410 ( .A1(n550), .A2(Q[809]), .B1(n551), .B2(Q[105]), .C1(n549), 
        .C2(Q[745]), .ZN(n387) );
  NAND3_X1 U411 ( .A1(n385), .A2(n386), .A3(n387), .ZN(n388) );
  AOI22_X1 U412 ( .A1(n553), .A2(Q[841]), .B1(n552), .B2(Q[713]), .ZN(n389) );
  AOI22_X1 U413 ( .A1(n555), .A2(Q[777]), .B1(n554), .B2(Q[873]), .ZN(n390) );
  NAND4_X1 U414 ( .A1(n670), .A2(n671), .A3(n389), .A4(n390), .ZN(n391) );
  OR4_X1 U415 ( .A1(n379), .A2(n384), .A3(n388), .A4(n391), .ZN(Y[9]) );
  AOI22_X1 U416 ( .A1(n561), .A2(Q[488]), .B1(n560), .B2(Q[552]), .ZN(n392) );
  AOI22_X1 U417 ( .A1(n563), .A2(Q[648]), .B1(n562), .B2(Q[456]), .ZN(n393) );
  AOI22_X1 U418 ( .A1(n565), .A2(Q[360]), .B1(n564), .B2(Q[296]), .ZN(n394) );
  AOI22_X1 U419 ( .A1(n567), .A2(Q[392]), .B1(n566), .B2(Q[264]), .ZN(n395) );
  NAND4_X1 U420 ( .A1(n392), .A2(n393), .A3(n394), .A4(n395), .ZN(n396) );
  AOI22_X1 U421 ( .A1(n569), .A2(Q[328]), .B1(n568), .B2(Q[424]), .ZN(n397) );
  AOI22_X1 U422 ( .A1(n571), .A2(Q[232]), .B1(n570), .B2(Q[136]), .ZN(n398) );
  AOI22_X1 U423 ( .A1(n573), .A2(Q[72]), .B1(n572), .B2(Q[168]), .ZN(n399) );
  AOI22_X1 U424 ( .A1(n575), .A2(Q[200]), .B1(n574), .B2(Q[40]), .ZN(n400) );
  NAND4_X1 U425 ( .A1(n397), .A2(n398), .A3(n399), .A4(n400), .ZN(n401) );
  AOI22_X1 U426 ( .A1(n546), .A2(Q[1000]), .B1(n545), .B2(Q[936]), .ZN(n402)
         );
  AOI22_X1 U427 ( .A1(n548), .A2(Q[968]), .B1(n547), .B2(Q[904]), .ZN(n403) );
  AOI222_X1 U428 ( .A1(n550), .A2(Q[808]), .B1(n551), .B2(Q[104]), .C1(n549), 
        .C2(Q[744]), .ZN(n404) );
  NAND3_X1 U429 ( .A1(n402), .A2(n403), .A3(n404), .ZN(n405) );
  AOI22_X1 U430 ( .A1(n553), .A2(Q[840]), .B1(n552), .B2(Q[712]), .ZN(n406) );
  AOI22_X1 U431 ( .A1(n555), .A2(Q[776]), .B1(n554), .B2(Q[872]), .ZN(n407) );
  NAND4_X1 U432 ( .A1(n653), .A2(n654), .A3(n406), .A4(n407), .ZN(n408) );
  OR4_X1 U433 ( .A1(n396), .A2(n401), .A3(n405), .A4(n408), .ZN(Y[8]) );
  AOI22_X1 U434 ( .A1(n561), .A2(Q[487]), .B1(n560), .B2(Q[551]), .ZN(n409) );
  AOI22_X1 U435 ( .A1(n563), .A2(Q[647]), .B1(n562), .B2(Q[455]), .ZN(n410) );
  AOI22_X1 U436 ( .A1(n565), .A2(Q[359]), .B1(n564), .B2(Q[295]), .ZN(n411) );
  AOI22_X1 U437 ( .A1(n567), .A2(Q[391]), .B1(n566), .B2(Q[263]), .ZN(n412) );
  NAND4_X1 U438 ( .A1(n409), .A2(n410), .A3(n411), .A4(n412), .ZN(n413) );
  AOI22_X1 U439 ( .A1(n569), .A2(Q[327]), .B1(n568), .B2(Q[423]), .ZN(n414) );
  AOI22_X1 U440 ( .A1(n571), .A2(Q[231]), .B1(n570), .B2(Q[135]), .ZN(n415) );
  AOI22_X1 U441 ( .A1(n573), .A2(Q[71]), .B1(n572), .B2(Q[167]), .ZN(n416) );
  AOI22_X1 U442 ( .A1(n575), .A2(Q[199]), .B1(n574), .B2(Q[39]), .ZN(n417) );
  NAND4_X1 U443 ( .A1(n414), .A2(n415), .A3(n416), .A4(n417), .ZN(n418) );
  AOI22_X1 U444 ( .A1(n546), .A2(Q[999]), .B1(n545), .B2(Q[935]), .ZN(n419) );
  AOI22_X1 U445 ( .A1(n548), .A2(Q[967]), .B1(n547), .B2(Q[903]), .ZN(n420) );
  AOI222_X1 U446 ( .A1(n550), .A2(Q[807]), .B1(n551), .B2(Q[103]), .C1(n549), 
        .C2(Q[743]), .ZN(n421) );
  NAND3_X1 U447 ( .A1(n419), .A2(n420), .A3(n421), .ZN(n422) );
  AOI22_X1 U448 ( .A1(n553), .A2(Q[839]), .B1(n552), .B2(Q[711]), .ZN(n423) );
  AOI22_X1 U449 ( .A1(n555), .A2(Q[775]), .B1(n554), .B2(Q[871]), .ZN(n424) );
  NAND4_X1 U450 ( .A1(n651), .A2(n652), .A3(n423), .A4(n424), .ZN(n425) );
  OR4_X1 U451 ( .A1(n413), .A2(n418), .A3(n422), .A4(n425), .ZN(Y[7]) );
  AOI22_X1 U452 ( .A1(n561), .A2(Q[486]), .B1(n560), .B2(Q[550]), .ZN(n426) );
  AOI22_X1 U453 ( .A1(n563), .A2(Q[646]), .B1(n562), .B2(Q[454]), .ZN(n427) );
  AOI22_X1 U454 ( .A1(n565), .A2(Q[358]), .B1(n564), .B2(Q[294]), .ZN(n428) );
  AOI22_X1 U455 ( .A1(n567), .A2(Q[390]), .B1(n566), .B2(Q[262]), .ZN(n429) );
  NAND4_X1 U456 ( .A1(n426), .A2(n427), .A3(n428), .A4(n429), .ZN(n430) );
  AOI22_X1 U457 ( .A1(n569), .A2(Q[326]), .B1(n568), .B2(Q[422]), .ZN(n431) );
  AOI22_X1 U458 ( .A1(n571), .A2(Q[230]), .B1(n570), .B2(Q[134]), .ZN(n432) );
  AOI22_X1 U459 ( .A1(n573), .A2(Q[70]), .B1(n572), .B2(Q[166]), .ZN(n433) );
  AOI22_X1 U460 ( .A1(n575), .A2(Q[198]), .B1(n574), .B2(Q[38]), .ZN(n434) );
  NAND4_X1 U461 ( .A1(n431), .A2(n432), .A3(n433), .A4(n434), .ZN(n435) );
  AOI22_X1 U462 ( .A1(n546), .A2(Q[998]), .B1(n545), .B2(Q[934]), .ZN(n436) );
  AOI22_X1 U463 ( .A1(n548), .A2(Q[966]), .B1(n547), .B2(Q[902]), .ZN(n437) );
  AOI222_X1 U464 ( .A1(n550), .A2(Q[806]), .B1(n551), .B2(Q[102]), .C1(n549), 
        .C2(Q[742]), .ZN(n438) );
  NAND3_X1 U465 ( .A1(n436), .A2(n437), .A3(n438), .ZN(n439) );
  AOI22_X1 U466 ( .A1(n553), .A2(Q[838]), .B1(n552), .B2(Q[710]), .ZN(n440) );
  AOI22_X1 U467 ( .A1(n555), .A2(Q[774]), .B1(n554), .B2(Q[870]), .ZN(n441) );
  NAND4_X1 U468 ( .A1(n649), .A2(n650), .A3(n440), .A4(n441), .ZN(n442) );
  OR4_X1 U469 ( .A1(n430), .A2(n435), .A3(n439), .A4(n442), .ZN(Y[6]) );
  AOI22_X1 U470 ( .A1(n561), .A2(Q[485]), .B1(n560), .B2(Q[549]), .ZN(n443) );
  AOI22_X1 U471 ( .A1(n563), .A2(Q[645]), .B1(n562), .B2(Q[453]), .ZN(n444) );
  AOI22_X1 U472 ( .A1(n565), .A2(Q[357]), .B1(n564), .B2(Q[293]), .ZN(n445) );
  AOI22_X1 U473 ( .A1(n567), .A2(Q[389]), .B1(n566), .B2(Q[261]), .ZN(n446) );
  NAND4_X1 U474 ( .A1(n443), .A2(n444), .A3(n445), .A4(n446), .ZN(n447) );
  AOI22_X1 U475 ( .A1(n569), .A2(Q[325]), .B1(n568), .B2(Q[421]), .ZN(n448) );
  AOI22_X1 U476 ( .A1(n571), .A2(Q[229]), .B1(n570), .B2(Q[133]), .ZN(n449) );
  AOI22_X1 U477 ( .A1(n573), .A2(Q[69]), .B1(n572), .B2(Q[165]), .ZN(n450) );
  AOI22_X1 U478 ( .A1(n575), .A2(Q[197]), .B1(n574), .B2(Q[37]), .ZN(n451) );
  NAND4_X1 U479 ( .A1(n448), .A2(n449), .A3(n450), .A4(n451), .ZN(n452) );
  AOI22_X1 U480 ( .A1(n546), .A2(Q[997]), .B1(n545), .B2(Q[933]), .ZN(n453) );
  AOI22_X1 U481 ( .A1(n548), .A2(Q[965]), .B1(n547), .B2(Q[901]), .ZN(n454) );
  AOI222_X1 U482 ( .A1(n550), .A2(Q[805]), .B1(n551), .B2(Q[101]), .C1(n549), 
        .C2(Q[741]), .ZN(n455) );
  NAND3_X1 U483 ( .A1(n453), .A2(n454), .A3(n455), .ZN(n456) );
  AOI22_X1 U484 ( .A1(n553), .A2(Q[837]), .B1(n552), .B2(Q[709]), .ZN(n457) );
  AOI22_X1 U485 ( .A1(n555), .A2(Q[773]), .B1(n554), .B2(Q[869]), .ZN(n458) );
  NAND4_X1 U486 ( .A1(n647), .A2(n648), .A3(n457), .A4(n458), .ZN(n459) );
  OR4_X1 U487 ( .A1(n447), .A2(n452), .A3(n456), .A4(n459), .ZN(Y[5]) );
  AOI22_X1 U488 ( .A1(n561), .A2(Q[484]), .B1(n560), .B2(Q[548]), .ZN(n460) );
  AOI22_X1 U489 ( .A1(n563), .A2(Q[644]), .B1(n562), .B2(Q[452]), .ZN(n461) );
  AOI22_X1 U490 ( .A1(n565), .A2(Q[356]), .B1(n564), .B2(Q[292]), .ZN(n462) );
  AOI22_X1 U491 ( .A1(n567), .A2(Q[388]), .B1(n566), .B2(Q[260]), .ZN(n463) );
  NAND4_X1 U492 ( .A1(n460), .A2(n461), .A3(n462), .A4(n463), .ZN(n464) );
  AOI22_X1 U493 ( .A1(n569), .A2(Q[324]), .B1(n568), .B2(Q[420]), .ZN(n465) );
  AOI22_X1 U494 ( .A1(n571), .A2(Q[228]), .B1(n570), .B2(Q[132]), .ZN(n466) );
  AOI22_X1 U495 ( .A1(n573), .A2(Q[68]), .B1(n572), .B2(Q[164]), .ZN(n467) );
  AOI22_X1 U496 ( .A1(n575), .A2(Q[196]), .B1(n574), .B2(Q[36]), .ZN(n468) );
  NAND4_X1 U497 ( .A1(n465), .A2(n466), .A3(n467), .A4(n468), .ZN(n469) );
  AOI22_X1 U498 ( .A1(n546), .A2(Q[996]), .B1(n545), .B2(Q[932]), .ZN(n470) );
  AOI22_X1 U499 ( .A1(n548), .A2(Q[964]), .B1(n547), .B2(Q[900]), .ZN(n471) );
  AOI222_X1 U500 ( .A1(n550), .A2(Q[804]), .B1(n551), .B2(Q[100]), .C1(n549), 
        .C2(Q[740]), .ZN(n472) );
  NAND3_X1 U501 ( .A1(n470), .A2(n471), .A3(n472), .ZN(n473) );
  AOI22_X1 U502 ( .A1(n553), .A2(Q[836]), .B1(n552), .B2(Q[708]), .ZN(n474) );
  AOI22_X1 U503 ( .A1(n555), .A2(Q[772]), .B1(n554), .B2(Q[868]), .ZN(n475) );
  NAND4_X1 U504 ( .A1(n645), .A2(n646), .A3(n474), .A4(n475), .ZN(n476) );
  OR4_X1 U505 ( .A1(n464), .A2(n469), .A3(n473), .A4(n476), .ZN(Y[4]) );
  AOI22_X1 U506 ( .A1(n561), .A2(Q[483]), .B1(n560), .B2(Q[547]), .ZN(n477) );
  AOI22_X1 U507 ( .A1(n563), .A2(Q[643]), .B1(n562), .B2(Q[451]), .ZN(n478) );
  AOI22_X1 U508 ( .A1(n565), .A2(Q[355]), .B1(n564), .B2(Q[291]), .ZN(n479) );
  AOI22_X1 U509 ( .A1(n567), .A2(Q[387]), .B1(n566), .B2(Q[259]), .ZN(n480) );
  NAND4_X1 U510 ( .A1(n477), .A2(n478), .A3(n479), .A4(n480), .ZN(n481) );
  AOI22_X1 U511 ( .A1(n569), .A2(Q[323]), .B1(n568), .B2(Q[419]), .ZN(n482) );
  AOI22_X1 U512 ( .A1(n571), .A2(Q[227]), .B1(n570), .B2(Q[131]), .ZN(n483) );
  AOI22_X1 U513 ( .A1(n573), .A2(Q[67]), .B1(n572), .B2(Q[163]), .ZN(n484) );
  AOI22_X1 U514 ( .A1(n575), .A2(Q[195]), .B1(n574), .B2(Q[35]), .ZN(n485) );
  NAND4_X1 U515 ( .A1(n482), .A2(n483), .A3(n484), .A4(n485), .ZN(n486) );
  AOI22_X1 U516 ( .A1(n546), .A2(Q[995]), .B1(n545), .B2(Q[931]), .ZN(n487) );
  AOI22_X1 U517 ( .A1(n548), .A2(Q[963]), .B1(n547), .B2(Q[899]), .ZN(n488) );
  AOI222_X1 U518 ( .A1(n550), .A2(Q[803]), .B1(n551), .B2(Q[99]), .C1(n549), 
        .C2(Q[739]), .ZN(n489) );
  NAND3_X1 U519 ( .A1(n487), .A2(n488), .A3(n489), .ZN(n490) );
  AOI22_X1 U520 ( .A1(n553), .A2(Q[835]), .B1(n552), .B2(Q[707]), .ZN(n491) );
  AOI22_X1 U521 ( .A1(n555), .A2(Q[771]), .B1(n554), .B2(Q[867]), .ZN(n492) );
  NAND4_X1 U522 ( .A1(n643), .A2(n644), .A3(n491), .A4(n492), .ZN(n493) );
  OR4_X1 U523 ( .A1(n481), .A2(n486), .A3(n490), .A4(n493), .ZN(Y[3]) );
  AOI22_X1 U524 ( .A1(n561), .A2(Q[482]), .B1(n560), .B2(Q[546]), .ZN(n494) );
  AOI22_X1 U525 ( .A1(n563), .A2(Q[642]), .B1(n562), .B2(Q[450]), .ZN(n495) );
  AOI22_X1 U526 ( .A1(n565), .A2(Q[354]), .B1(n564), .B2(Q[290]), .ZN(n496) );
  AOI22_X1 U527 ( .A1(n567), .A2(Q[386]), .B1(n566), .B2(Q[258]), .ZN(n497) );
  NAND4_X1 U528 ( .A1(n494), .A2(n495), .A3(n496), .A4(n497), .ZN(n498) );
  AOI22_X1 U529 ( .A1(n569), .A2(Q[322]), .B1(n568), .B2(Q[418]), .ZN(n499) );
  AOI22_X1 U530 ( .A1(n571), .A2(Q[226]), .B1(n570), .B2(Q[130]), .ZN(n500) );
  AOI22_X1 U531 ( .A1(n573), .A2(Q[66]), .B1(n572), .B2(Q[162]), .ZN(n501) );
  AOI22_X1 U532 ( .A1(n575), .A2(Q[194]), .B1(n574), .B2(Q[34]), .ZN(n502) );
  NAND4_X1 U533 ( .A1(n499), .A2(n500), .A3(n501), .A4(n502), .ZN(n503) );
  AOI22_X1 U534 ( .A1(n546), .A2(Q[994]), .B1(n545), .B2(Q[930]), .ZN(n504) );
  AOI22_X1 U535 ( .A1(n548), .A2(Q[962]), .B1(n547), .B2(Q[898]), .ZN(n505) );
  AOI222_X1 U536 ( .A1(n550), .A2(Q[802]), .B1(n551), .B2(Q[98]), .C1(n549), 
        .C2(Q[738]), .ZN(n506) );
  NAND3_X1 U537 ( .A1(n504), .A2(n505), .A3(n506), .ZN(n507) );
  AOI22_X1 U538 ( .A1(n553), .A2(Q[834]), .B1(n552), .B2(Q[706]), .ZN(n508) );
  AOI22_X1 U539 ( .A1(n555), .A2(Q[770]), .B1(n554), .B2(Q[866]), .ZN(n509) );
  NAND4_X1 U540 ( .A1(n637), .A2(n638), .A3(n508), .A4(n509), .ZN(n510) );
  OR4_X1 U541 ( .A1(n498), .A2(n503), .A3(n507), .A4(n510), .ZN(Y[2]) );
  AOI22_X1 U542 ( .A1(n561), .A2(Q[481]), .B1(n560), .B2(Q[545]), .ZN(n511) );
  AOI22_X1 U543 ( .A1(n563), .A2(Q[641]), .B1(n562), .B2(Q[449]), .ZN(n512) );
  AOI22_X1 U544 ( .A1(n565), .A2(Q[353]), .B1(n564), .B2(Q[289]), .ZN(n513) );
  AOI22_X1 U545 ( .A1(n567), .A2(Q[385]), .B1(n566), .B2(Q[257]), .ZN(n514) );
  NAND4_X1 U546 ( .A1(n511), .A2(n512), .A3(n513), .A4(n514), .ZN(n515) );
  AOI22_X1 U547 ( .A1(n569), .A2(Q[321]), .B1(n568), .B2(Q[417]), .ZN(n516) );
  AOI22_X1 U548 ( .A1(n571), .A2(Q[225]), .B1(n570), .B2(Q[129]), .ZN(n517) );
  AOI22_X1 U549 ( .A1(n573), .A2(Q[65]), .B1(n572), .B2(Q[161]), .ZN(n518) );
  AOI22_X1 U550 ( .A1(n575), .A2(Q[193]), .B1(n574), .B2(Q[33]), .ZN(n519) );
  NAND4_X1 U551 ( .A1(n516), .A2(n517), .A3(n518), .A4(n519), .ZN(n520) );
  AOI22_X1 U552 ( .A1(n546), .A2(Q[993]), .B1(n545), .B2(Q[929]), .ZN(n521) );
  AOI22_X1 U553 ( .A1(n548), .A2(Q[961]), .B1(n547), .B2(Q[897]), .ZN(n522) );
  AOI222_X1 U554 ( .A1(n550), .A2(Q[801]), .B1(n551), .B2(Q[97]), .C1(n549), 
        .C2(Q[737]), .ZN(n523) );
  NAND3_X1 U555 ( .A1(n521), .A2(n522), .A3(n523), .ZN(n524) );
  AOI22_X1 U556 ( .A1(n553), .A2(Q[833]), .B1(n552), .B2(Q[705]), .ZN(n525) );
  AOI22_X1 U557 ( .A1(n555), .A2(Q[769]), .B1(n554), .B2(Q[865]), .ZN(n526) );
  NAND4_X1 U558 ( .A1(n615), .A2(n616), .A3(n525), .A4(n526), .ZN(n527) );
  OR4_X1 U559 ( .A1(n515), .A2(n520), .A3(n524), .A4(n527), .ZN(Y[1]) );
  AOI22_X1 U560 ( .A1(n561), .A2(Q[480]), .B1(n560), .B2(Q[544]), .ZN(n528) );
  AOI22_X1 U561 ( .A1(n563), .A2(Q[640]), .B1(n562), .B2(Q[448]), .ZN(n529) );
  AOI22_X1 U562 ( .A1(n565), .A2(Q[352]), .B1(n564), .B2(Q[288]), .ZN(n530) );
  AOI22_X1 U563 ( .A1(n567), .A2(Q[384]), .B1(n566), .B2(Q[256]), .ZN(n531) );
  NAND4_X1 U564 ( .A1(n528), .A2(n529), .A3(n530), .A4(n531), .ZN(n532) );
  AOI22_X1 U565 ( .A1(n569), .A2(Q[320]), .B1(n568), .B2(Q[416]), .ZN(n533) );
  AOI22_X1 U566 ( .A1(n571), .A2(Q[224]), .B1(n570), .B2(Q[128]), .ZN(n534) );
  AOI22_X1 U567 ( .A1(n573), .A2(Q[64]), .B1(n572), .B2(Q[160]), .ZN(n535) );
  AOI22_X1 U568 ( .A1(n575), .A2(Q[192]), .B1(n574), .B2(Q[32]), .ZN(n536) );
  NAND4_X1 U569 ( .A1(n533), .A2(n534), .A3(n535), .A4(n536), .ZN(n537) );
  AOI22_X1 U570 ( .A1(n546), .A2(Q[992]), .B1(n545), .B2(Q[928]), .ZN(n538) );
  AOI22_X1 U571 ( .A1(n548), .A2(Q[960]), .B1(n547), .B2(Q[896]), .ZN(n539) );
  AOI222_X1 U572 ( .A1(n550), .A2(Q[800]), .B1(n551), .B2(Q[96]), .C1(n549), 
        .C2(Q[736]), .ZN(n540) );
  NAND3_X1 U573 ( .A1(n538), .A2(n539), .A3(n540), .ZN(n541) );
  AOI22_X1 U574 ( .A1(n553), .A2(Q[832]), .B1(n552), .B2(Q[704]), .ZN(n542) );
  AOI22_X1 U575 ( .A1(n555), .A2(Q[768]), .B1(n554), .B2(Q[864]), .ZN(n543) );
  NAND4_X1 U576 ( .A1(n580), .A2(n581), .A3(n542), .A4(n543), .ZN(n544) );
  OR4_X1 U577 ( .A1(n532), .A2(n537), .A3(n541), .A4(n544), .ZN(Y[0]) );
  BUF_X1 U578 ( .A(n686), .Z(n574) );
  BUF_X1 U579 ( .A(n687), .Z(n575) );
  BUF_X1 U580 ( .A(n684), .Z(n572) );
  BUF_X1 U581 ( .A(n685), .Z(n573) );
  BUF_X1 U582 ( .A(n682), .Z(n570) );
  BUF_X1 U583 ( .A(n683), .Z(n571) );
  BUF_X1 U584 ( .A(n680), .Z(n568) );
  BUF_X1 U585 ( .A(n681), .Z(n569) );
  BUF_X1 U586 ( .A(n678), .Z(n566) );
  BUF_X1 U587 ( .A(n679), .Z(n567) );
  BUF_X1 U588 ( .A(n676), .Z(n564) );
  BUF_X1 U589 ( .A(n677), .Z(n565) );
  BUF_X1 U590 ( .A(n674), .Z(n562) );
  BUF_X1 U591 ( .A(n675), .Z(n563) );
  BUF_X1 U592 ( .A(n672), .Z(n560) );
  BUF_X1 U593 ( .A(n673), .Z(n561) );
  BUF_X1 U594 ( .A(n668), .Z(n558) );
  BUF_X1 U595 ( .A(n669), .Z(n559) );
  BUF_X1 U596 ( .A(n666), .Z(n556) );
  BUF_X1 U597 ( .A(n667), .Z(n557) );
  BUF_X1 U598 ( .A(n664), .Z(n554) );
  BUF_X1 U599 ( .A(n665), .Z(n555) );
  BUF_X1 U600 ( .A(n662), .Z(n552) );
  BUF_X1 U601 ( .A(n663), .Z(n553) );
  BUF_X1 U602 ( .A(n661), .Z(n551) );
  BUF_X1 U603 ( .A(n659), .Z(n549) );
  BUF_X1 U604 ( .A(n660), .Z(n550) );
  BUF_X1 U605 ( .A(n657), .Z(n547) );
  BUF_X1 U606 ( .A(n658), .Z(n548) );
  BUF_X1 U607 ( .A(n655), .Z(n545) );
  BUF_X1 U608 ( .A(n656), .Z(n546) );
  OR2_X1 U609 ( .A1(S[1]), .A2(S[2]), .ZN(n593) );
  OR2_X1 U610 ( .A1(n576), .A2(S[1]), .ZN(n590) );
  NAND2_X1 U611 ( .A1(S[1]), .A2(S[2]), .ZN(n592) );
  NAND3_X1 U612 ( .A1(S[3]), .A2(S[4]), .A3(S[0]), .ZN(n579) );
  NOR2_X1 U613 ( .A1(n592), .A2(n579), .ZN(n656) );
  INV_X1 U614 ( .A(S[2]), .ZN(n576) );
  NOR2_X1 U615 ( .A1(n579), .A2(n590), .ZN(n655) );
  INV_X1 U616 ( .A(S[0]), .ZN(n577) );
  NAND3_X1 U617 ( .A1(S[4]), .A2(S[3]), .A3(n577), .ZN(n578) );
  NOR2_X1 U618 ( .A1(n592), .A2(n578), .ZN(n658) );
  NOR2_X1 U619 ( .A1(n590), .A2(n578), .ZN(n657) );
  NOR2_X1 U620 ( .A1(n579), .A2(n593), .ZN(n660) );
  INV_X1 U621 ( .A(S[3]), .ZN(n587) );
  NAND3_X1 U622 ( .A1(S[4]), .A2(S[0]), .A3(n587), .ZN(n583) );
  NOR2_X1 U623 ( .A1(n592), .A2(n583), .ZN(n659) );
  NAND2_X1 U624 ( .A1(S[1]), .A2(n576), .ZN(n589) );
  INV_X1 U625 ( .A(S[4]), .ZN(n582) );
  NAND3_X1 U626 ( .A1(S[0]), .A2(n587), .A3(n582), .ZN(n594) );
  NOR2_X1 U627 ( .A1(n589), .A2(n594), .ZN(n661) );
  NOR2_X1 U628 ( .A1(n589), .A2(n578), .ZN(n663) );
  NAND3_X1 U629 ( .A1(S[4]), .A2(n587), .A3(n577), .ZN(n584) );
  NOR2_X1 U630 ( .A1(n592), .A2(n584), .ZN(n662) );
  NOR2_X1 U631 ( .A1(n578), .A2(n593), .ZN(n665) );
  NOR2_X1 U632 ( .A1(n589), .A2(n579), .ZN(n664) );
  NOR2_X1 U633 ( .A1(n590), .A2(n583), .ZN(n667) );
  NOR2_X1 U634 ( .A1(n589), .A2(n584), .ZN(n666) );
  AOI22_X1 U635 ( .A1(n557), .A2(Q[672]), .B1(n556), .B2(Q[576]), .ZN(n581) );
  NOR2_X1 U636 ( .A1(n593), .A2(n584), .ZN(n669) );
  NOR2_X1 U637 ( .A1(n589), .A2(n583), .ZN(n668) );
  AOI22_X1 U638 ( .A1(n559), .A2(Q[512]), .B1(n558), .B2(Q[608]), .ZN(n580) );
  NAND3_X1 U639 ( .A1(S[3]), .A2(S[0]), .A3(n582), .ZN(n586) );
  NOR2_X1 U640 ( .A1(n592), .A2(n586), .ZN(n673) );
  NOR2_X1 U641 ( .A1(n593), .A2(n583), .ZN(n672) );
  NOR2_X1 U642 ( .A1(n590), .A2(n584), .ZN(n675) );
  NOR2_X1 U643 ( .A1(S[4]), .A2(S[0]), .ZN(n588) );
  NAND2_X1 U644 ( .A1(S[3]), .A2(n588), .ZN(n585) );
  NOR2_X1 U645 ( .A1(n592), .A2(n585), .ZN(n674) );
  NOR2_X1 U646 ( .A1(n589), .A2(n586), .ZN(n677) );
  NOR2_X1 U647 ( .A1(n593), .A2(n586), .ZN(n676) );
  NOR2_X1 U648 ( .A1(n590), .A2(n585), .ZN(n679) );
  NOR2_X1 U649 ( .A1(n593), .A2(n585), .ZN(n678) );
  NOR2_X1 U650 ( .A1(n589), .A2(n585), .ZN(n681) );
  NOR2_X1 U651 ( .A1(n590), .A2(n586), .ZN(n680) );
  NOR2_X1 U652 ( .A1(n594), .A2(n592), .ZN(n683) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n590), .A2(n591), .ZN(n682) );
  NOR2_X1 U655 ( .A1(n589), .A2(n591), .ZN(n685) );
  NOR2_X1 U656 ( .A1(n594), .A2(n590), .ZN(n684) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n687) );
  NOR2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n686) );
  AOI22_X1 U659 ( .A1(n557), .A2(Q[682]), .B1(n556), .B2(Q[586]), .ZN(n596) );
  AOI22_X1 U660 ( .A1(n559), .A2(Q[522]), .B1(n558), .B2(Q[618]), .ZN(n595) );
  AOI22_X1 U661 ( .A1(n667), .A2(Q[683]), .B1(n666), .B2(Q[587]), .ZN(n598) );
  AOI22_X1 U662 ( .A1(n669), .A2(Q[523]), .B1(n668), .B2(Q[619]), .ZN(n597) );
  AOI22_X1 U663 ( .A1(n667), .A2(Q[684]), .B1(n666), .B2(Q[588]), .ZN(n600) );
  AOI22_X1 U664 ( .A1(n669), .A2(Q[524]), .B1(n668), .B2(Q[620]), .ZN(n599) );
  AOI22_X1 U665 ( .A1(n667), .A2(Q[685]), .B1(n666), .B2(Q[589]), .ZN(n602) );
  AOI22_X1 U666 ( .A1(n669), .A2(Q[525]), .B1(n668), .B2(Q[621]), .ZN(n601) );
  AOI22_X1 U667 ( .A1(n667), .A2(Q[686]), .B1(n666), .B2(Q[590]), .ZN(n604) );
  AOI22_X1 U668 ( .A1(n669), .A2(Q[526]), .B1(n668), .B2(Q[622]), .ZN(n603) );
  AOI22_X1 U669 ( .A1(n667), .A2(Q[687]), .B1(n666), .B2(Q[591]), .ZN(n606) );
  AOI22_X1 U670 ( .A1(n669), .A2(Q[527]), .B1(n668), .B2(Q[623]), .ZN(n605) );
  AOI22_X1 U671 ( .A1(n667), .A2(Q[688]), .B1(n666), .B2(Q[592]), .ZN(n608) );
  AOI22_X1 U672 ( .A1(n669), .A2(Q[528]), .B1(n668), .B2(Q[624]), .ZN(n607) );
  AOI22_X1 U673 ( .A1(n667), .A2(Q[689]), .B1(n666), .B2(Q[593]), .ZN(n610) );
  AOI22_X1 U674 ( .A1(n669), .A2(Q[529]), .B1(n668), .B2(Q[625]), .ZN(n609) );
  AOI22_X1 U675 ( .A1(n667), .A2(Q[690]), .B1(n666), .B2(Q[594]), .ZN(n612) );
  AOI22_X1 U676 ( .A1(n669), .A2(Q[530]), .B1(n668), .B2(Q[626]), .ZN(n611) );
  AOI22_X1 U677 ( .A1(n667), .A2(Q[691]), .B1(n666), .B2(Q[595]), .ZN(n614) );
  AOI22_X1 U678 ( .A1(n669), .A2(Q[531]), .B1(n668), .B2(Q[627]), .ZN(n613) );
  AOI22_X1 U679 ( .A1(n557), .A2(Q[673]), .B1(n556), .B2(Q[577]), .ZN(n616) );
  AOI22_X1 U680 ( .A1(n559), .A2(Q[513]), .B1(n558), .B2(Q[609]), .ZN(n615) );
  AOI22_X1 U681 ( .A1(n557), .A2(Q[692]), .B1(n556), .B2(Q[596]), .ZN(n618) );
  AOI22_X1 U682 ( .A1(n559), .A2(Q[532]), .B1(n558), .B2(Q[628]), .ZN(n617) );
  AOI22_X1 U683 ( .A1(n557), .A2(Q[693]), .B1(n556), .B2(Q[597]), .ZN(n620) );
  AOI22_X1 U684 ( .A1(n559), .A2(Q[533]), .B1(n558), .B2(Q[629]), .ZN(n619) );
  AOI22_X1 U685 ( .A1(n557), .A2(Q[694]), .B1(n556), .B2(Q[598]), .ZN(n622) );
  AOI22_X1 U686 ( .A1(n559), .A2(Q[534]), .B1(n558), .B2(Q[630]), .ZN(n621) );
  AOI22_X1 U687 ( .A1(n557), .A2(Q[695]), .B1(n556), .B2(Q[599]), .ZN(n624) );
  AOI22_X1 U688 ( .A1(n559), .A2(Q[535]), .B1(n558), .B2(Q[631]), .ZN(n623) );
  AOI22_X1 U689 ( .A1(n557), .A2(Q[696]), .B1(n556), .B2(Q[600]), .ZN(n626) );
  AOI22_X1 U690 ( .A1(n559), .A2(Q[536]), .B1(n558), .B2(Q[632]), .ZN(n625) );
  AOI22_X1 U691 ( .A1(n557), .A2(Q[697]), .B1(n556), .B2(Q[601]), .ZN(n628) );
  AOI22_X1 U692 ( .A1(n559), .A2(Q[537]), .B1(n558), .B2(Q[633]), .ZN(n627) );
  AOI22_X1 U693 ( .A1(n557), .A2(Q[698]), .B1(n556), .B2(Q[602]), .ZN(n630) );
  AOI22_X1 U694 ( .A1(n559), .A2(Q[538]), .B1(n558), .B2(Q[634]), .ZN(n629) );
  AOI22_X1 U695 ( .A1(n557), .A2(Q[699]), .B1(n556), .B2(Q[603]), .ZN(n632) );
  AOI22_X1 U696 ( .A1(n559), .A2(Q[539]), .B1(n558), .B2(Q[635]), .ZN(n631) );
  AOI22_X1 U697 ( .A1(n557), .A2(Q[700]), .B1(n556), .B2(Q[604]), .ZN(n634) );
  AOI22_X1 U698 ( .A1(n559), .A2(Q[540]), .B1(n558), .B2(Q[636]), .ZN(n633) );
  AOI22_X1 U699 ( .A1(n667), .A2(Q[701]), .B1(n666), .B2(Q[605]), .ZN(n636) );
  AOI22_X1 U700 ( .A1(n669), .A2(Q[541]), .B1(n668), .B2(Q[637]), .ZN(n635) );
  AOI22_X1 U701 ( .A1(n557), .A2(Q[674]), .B1(n556), .B2(Q[578]), .ZN(n638) );
  AOI22_X1 U702 ( .A1(n559), .A2(Q[514]), .B1(n558), .B2(Q[610]), .ZN(n637) );
  AOI22_X1 U703 ( .A1(n557), .A2(Q[702]), .B1(n556), .B2(Q[606]), .ZN(n640) );
  AOI22_X1 U704 ( .A1(n559), .A2(Q[542]), .B1(n558), .B2(Q[638]), .ZN(n639) );
  AOI22_X1 U705 ( .A1(n557), .A2(Q[703]), .B1(n556), .B2(Q[607]), .ZN(n642) );
  AOI22_X1 U706 ( .A1(n559), .A2(Q[543]), .B1(n558), .B2(Q[639]), .ZN(n641) );
  AOI22_X1 U707 ( .A1(n557), .A2(Q[675]), .B1(n556), .B2(Q[579]), .ZN(n644) );
  AOI22_X1 U708 ( .A1(n559), .A2(Q[515]), .B1(n558), .B2(Q[611]), .ZN(n643) );
  AOI22_X1 U709 ( .A1(n557), .A2(Q[676]), .B1(n556), .B2(Q[580]), .ZN(n646) );
  AOI22_X1 U710 ( .A1(n559), .A2(Q[516]), .B1(n558), .B2(Q[612]), .ZN(n645) );
  AOI22_X1 U711 ( .A1(n557), .A2(Q[677]), .B1(n556), .B2(Q[581]), .ZN(n648) );
  AOI22_X1 U712 ( .A1(n559), .A2(Q[517]), .B1(n558), .B2(Q[613]), .ZN(n647) );
  AOI22_X1 U713 ( .A1(n557), .A2(Q[678]), .B1(n556), .B2(Q[582]), .ZN(n650) );
  AOI22_X1 U714 ( .A1(n559), .A2(Q[518]), .B1(n558), .B2(Q[614]), .ZN(n649) );
  AOI22_X1 U715 ( .A1(n557), .A2(Q[679]), .B1(n556), .B2(Q[583]), .ZN(n652) );
  AOI22_X1 U716 ( .A1(n559), .A2(Q[519]), .B1(n558), .B2(Q[615]), .ZN(n651) );
  AOI22_X1 U717 ( .A1(n557), .A2(Q[680]), .B1(n556), .B2(Q[584]), .ZN(n654) );
  AOI22_X1 U718 ( .A1(n559), .A2(Q[520]), .B1(n558), .B2(Q[616]), .ZN(n653) );
  AOI22_X1 U719 ( .A1(n557), .A2(Q[681]), .B1(n556), .B2(Q[585]), .ZN(n671) );
  AOI22_X1 U720 ( .A1(n559), .A2(Q[521]), .B1(n558), .B2(Q[617]), .ZN(n670) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 ( CLK, RST, IRAM_ADDRESS, 
        IRAM_ISSUE, IRAM_READY, IRAM_DATA, DRAM_ADDRESS, DRAM_ISSUE, 
        DRAM_READNOTWRITE, DRAM_READY, DRAM_DATA_IN, DRAM_DATA_OUT, DATA_SIZE, 
        DRAMRF_ADDRESS, DRAMRF_ISSUE, DRAMRF_READNOTWRITE, DRAMRF_READY, 
        DRAMRF_DATA_IN, DRAMRF_DATA_OUT, DATA_SIZE_RF );
  output [31:0] IRAM_ADDRESS;
  input [31:0] IRAM_DATA;
  output [31:0] DRAM_ADDRESS;
  input [31:0] DRAM_DATA_IN;
  output [31:0] DRAM_DATA_OUT;
  output [1:0] DATA_SIZE;
  output [31:0] DRAMRF_ADDRESS;
  input [31:0] DRAMRF_DATA_IN;
  output [31:0] DRAMRF_DATA_OUT;
  output [1:0] DATA_SIZE_RF;
  input CLK, RST, IRAM_READY, DRAM_READY, DRAMRF_READY;
  output IRAM_ISSUE, DRAM_ISSUE, DRAM_READNOTWRITE, DRAMRF_ISSUE,
         DRAMRF_READNOTWRITE;
  wire   i_HAZARD_SIG_CU, i_BUSY_WINDOW, i_SEL_CMPB, i_NPC_SEL, i_S2,
         i_SEL_ALU_SETCMP, \i_SEL_LGET[1] , i_DATAMEM_RM, i_S3, i_WF, i_RF1,
         i_RF2, \CU_I/N315 , \CU_I/N314 , \CU_I/N302 , \CU_I/N301 ,
         \CU_I/i_FILL_delay , \CU_I/CW_MEM[WB_EN] , \CU_I/CW_MEM[WB_MUX_SEL] ,
         \CU_I/CW_MEM[MEM_EN] , \CU_I/CW_EX[WB_EN] , \CU_I/CW_EX[WB_MUX_SEL] ,
         \CU_I/CW_EX[EX_EN] , \CU_I/CW_ID[WB_EN] , \CU_I/CW_ID[WB_MUX_SEL] ,
         \CU_I/CW_ID[MEM_EN] , \CU_I/CW_ID[DATA_SIZE][0] ,
         \CU_I/CW_ID[DATA_SIZE][1] , \CU_I/CW_ID[DRAM_RE] ,
         \CU_I/CW_ID[DRAM_WE] , \CU_I/CW_ID[MUXB_SEL] , \CU_I/CW_ID[MUXA_SEL] ,
         \CU_I/CW_ID[EX_EN] , \CU_I/CW_ID[ID_EN] , \CU_I/CW_ID[UNSIGNED_ID] ,
         \CU_I/CW_IF[WB_EN] , \CU_I/CW[WB_MUX_SEL] , \CU_I/CW[DATA_SIZE][0] ,
         \CU_I/CW[DATA_SIZE][1] , \CU_I/CW[DRAM_WE] , \CU_I/CW[MUXB_SEL] ,
         \CU_I/CW[NPC_SEL] , \CU_I/CW[UNSIGNED_ID] , \CU_I/CW[SEL_CMPB] ,
         \CU_I/CW[RF_RD2_EN] , \CU_I/CW[RF_RD1_EN] ,
         \DECODEhw/i_tickcounter[31] , \DECODEhw/i_tickcounter[29] ,
         \DECODEhw/i_tickcounter[26] , \DECODEhw/i_tickcounter[24] ,
         \DECODEhw/i_tickcounter[22] , \DECODEhw/i_tickcounter[20] ,
         \DECODEhw/i_tickcounter[18] , \DECODEhw/i_tickcounter[16] ,
         \DECODEhw/i_tickcounter[14] , \DECODEhw/i_tickcounter[12] ,
         \DECODEhw/i_tickcounter[10] , \DECODEhw/i_tickcounter[8] ,
         \DECODEhw/i_tickcounter[6] , \DECODEhw/i_tickcounter[4] ,
         \DECODEhw/i_tickcounter[2] , \DECODEhw/i_WR1 ,
         \DataPath/i_PIPLIN_WRB2[4] , \DataPath/i_PIPLIN_WRB2[3] ,
         \DataPath/i_PIPLIN_WRB2[2] , \DataPath/i_PIPLIN_WRB2[1] ,
         \DataPath/i_PIPLIN_WRB2[0] , \DataPath/i_PIPLIN_WRB1[4] ,
         \DataPath/i_PIPLIN_WRB1[3] , \DataPath/i_PIPLIN_WRB1[2] ,
         \DataPath/i_PIPLIN_WRB1[1] , \DataPath/i_PIPLIN_WRB1[0] ,
         \DataPath/i_REG_MEM_ALUOUT[31] , \DataPath/i_REG_MEM_ALUOUT[30] ,
         \DataPath/i_REG_MEM_ALUOUT[29] , \DataPath/i_REG_MEM_ALUOUT[28] ,
         \DataPath/i_REG_MEM_ALUOUT[27] , \DataPath/i_REG_MEM_ALUOUT[26] ,
         \DataPath/i_REG_MEM_ALUOUT[25] , \DataPath/i_REG_MEM_ALUOUT[24] ,
         \DataPath/i_REG_MEM_ALUOUT[23] , \DataPath/i_REG_MEM_ALUOUT[22] ,
         \DataPath/i_REG_MEM_ALUOUT[21] , \DataPath/i_REG_MEM_ALUOUT[20] ,
         \DataPath/i_REG_MEM_ALUOUT[19] , \DataPath/i_REG_MEM_ALUOUT[18] ,
         \DataPath/i_REG_MEM_ALUOUT[17] , \DataPath/i_REG_MEM_ALUOUT[16] ,
         \DataPath/i_REG_MEM_ALUOUT[15] , \DataPath/i_REG_MEM_ALUOUT[14] ,
         \DataPath/i_REG_MEM_ALUOUT[13] , \DataPath/i_REG_MEM_ALUOUT[12] ,
         \DataPath/i_REG_MEM_ALUOUT[11] , \DataPath/i_REG_MEM_ALUOUT[10] ,
         \DataPath/i_REG_MEM_ALUOUT[9] , \DataPath/i_REG_MEM_ALUOUT[8] ,
         \DataPath/i_REG_MEM_ALUOUT[7] , \DataPath/i_REG_MEM_ALUOUT[6] ,
         \DataPath/i_REG_MEM_ALUOUT[5] , \DataPath/i_REG_MEM_ALUOUT[4] ,
         \DataPath/i_REG_MEM_ALUOUT[3] , \DataPath/i_REG_MEM_ALUOUT[2] ,
         \DataPath/i_REG_MEM_ALUOUT[1] , \DataPath/i_REG_MEM_ALUOUT[0] ,
         \DataPath/i_REG_LDSTR_OUT[31] , \DataPath/i_REG_LDSTR_OUT[30] ,
         \DataPath/i_REG_LDSTR_OUT[29] , \DataPath/i_REG_LDSTR_OUT[28] ,
         \DataPath/i_REG_LDSTR_OUT[27] , \DataPath/i_REG_LDSTR_OUT[26] ,
         \DataPath/i_REG_LDSTR_OUT[25] , \DataPath/i_REG_LDSTR_OUT[24] ,
         \DataPath/i_REG_LDSTR_OUT[23] , \DataPath/i_REG_LDSTR_OUT[22] ,
         \DataPath/i_REG_LDSTR_OUT[21] , \DataPath/i_REG_LDSTR_OUT[20] ,
         \DataPath/i_REG_LDSTR_OUT[19] , \DataPath/i_REG_LDSTR_OUT[18] ,
         \DataPath/i_REG_LDSTR_OUT[17] , \DataPath/i_REG_LDSTR_OUT[16] ,
         \DataPath/i_REG_LDSTR_OUT[15] , \DataPath/i_REG_LDSTR_OUT[14] ,
         \DataPath/i_REG_LDSTR_OUT[13] , \DataPath/i_REG_LDSTR_OUT[12] ,
         \DataPath/i_REG_LDSTR_OUT[11] , \DataPath/i_REG_LDSTR_OUT[10] ,
         \DataPath/i_REG_LDSTR_OUT[9] , \DataPath/i_REG_LDSTR_OUT[8] ,
         \DataPath/i_REG_LDSTR_OUT[7] , \DataPath/i_REG_LDSTR_OUT[6] ,
         \DataPath/i_REG_LDSTR_OUT[5] , \DataPath/i_REG_LDSTR_OUT[4] ,
         \DataPath/i_REG_LDSTR_OUT[3] , \DataPath/i_REG_LDSTR_OUT[2] ,
         \DataPath/i_REG_LDSTR_OUT[1] , \DataPath/i_REG_LDSTR_OUT[0] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[31] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[30] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[29] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[28] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[27] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[26] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[25] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[24] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[23] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[22] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[21] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[20] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[19] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[18] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[17] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[16] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[15] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[14] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[13] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[12] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[11] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[10] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[9] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[8] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[7] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[6] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[5] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[4] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[3] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[2] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[1] ,
         \DataPath/i_REG_ME_DATA_DATAMEM[0] , \DataPath/i_LGET[0] ,
         \DataPath/i_PIPLIN_IN2[31] , \DataPath/i_PIPLIN_IN2[30] ,
         \DataPath/i_PIPLIN_IN2[29] , \DataPath/i_PIPLIN_IN2[28] ,
         \DataPath/i_PIPLIN_IN2[27] , \DataPath/i_PIPLIN_IN2[26] ,
         \DataPath/i_PIPLIN_IN2[25] , \DataPath/i_PIPLIN_IN2[24] ,
         \DataPath/i_PIPLIN_IN2[23] , \DataPath/i_PIPLIN_IN2[22] ,
         \DataPath/i_PIPLIN_IN2[21] , \DataPath/i_PIPLIN_IN2[20] ,
         \DataPath/i_PIPLIN_IN2[19] , \DataPath/i_PIPLIN_IN2[18] ,
         \DataPath/i_PIPLIN_IN2[17] , \DataPath/i_PIPLIN_IN2[16] ,
         \DataPath/i_PIPLIN_IN2[15] , \DataPath/i_PIPLIN_IN2[14] ,
         \DataPath/i_PIPLIN_IN2[13] , \DataPath/i_PIPLIN_IN2[12] ,
         \DataPath/i_PIPLIN_IN2[11] , \DataPath/i_PIPLIN_IN2[10] ,
         \DataPath/i_PIPLIN_IN2[9] , \DataPath/i_PIPLIN_IN2[8] ,
         \DataPath/i_PIPLIN_IN2[7] , \DataPath/i_PIPLIN_IN2[5] ,
         \DataPath/i_PIPLIN_IN2[4] , \DataPath/i_PIPLIN_IN2[3] ,
         \DataPath/i_PIPLIN_IN2[2] , \DataPath/i_PIPLIN_IN2[1] ,
         \DataPath/i_PIPLIN_IN2[0] , \DataPath/i_PIPLIN_IN1[15] ,
         \DataPath/i_PIPLIN_IN1[14] , \DataPath/i_PIPLIN_IN1[13] ,
         \DataPath/i_PIPLIN_IN1[12] , \DataPath/i_PIPLIN_IN1[11] ,
         \DataPath/i_PIPLIN_IN1[10] , \DataPath/i_PIPLIN_IN1[9] ,
         \DataPath/i_PIPLIN_IN1[8] , \DataPath/i_PIPLIN_IN1[7] ,
         \DataPath/i_PIPLIN_IN1[6] , \DataPath/i_PIPLIN_IN1[5] ,
         \DataPath/i_PIPLIN_IN1[4] , \DataPath/i_PIPLIN_IN1[3] ,
         \DataPath/i_PIPLIN_IN1[2] , \DataPath/i_PIPLIN_IN1[1] ,
         \DataPath/i_PIPLIN_IN1[0] , \DataPath/i_PIPLIN_B[0] ,
         \DataPath/i_PIPLIN_B[1] , \DataPath/i_PIPLIN_B[2] ,
         \DataPath/i_PIPLIN_B[3] , \DataPath/i_PIPLIN_B[4] ,
         \DataPath/i_PIPLIN_B[5] , \DataPath/i_PIPLIN_B[7] ,
         \DataPath/i_PIPLIN_B[8] , \DataPath/i_PIPLIN_B[9] ,
         \DataPath/i_PIPLIN_B[10] , \DataPath/i_PIPLIN_B[11] ,
         \DataPath/i_PIPLIN_B[12] , \DataPath/i_PIPLIN_B[13] ,
         \DataPath/i_PIPLIN_B[14] , \DataPath/i_PIPLIN_B[15] ,
         \DataPath/i_PIPLIN_B[16] , \DataPath/i_PIPLIN_B[17] ,
         \DataPath/i_PIPLIN_B[18] , \DataPath/i_PIPLIN_B[19] ,
         \DataPath/i_PIPLIN_B[20] , \DataPath/i_PIPLIN_B[21] ,
         \DataPath/i_PIPLIN_B[22] , \DataPath/i_PIPLIN_B[23] ,
         \DataPath/i_PIPLIN_B[24] , \DataPath/i_PIPLIN_B[25] ,
         \DataPath/i_PIPLIN_B[26] , \DataPath/i_PIPLIN_B[27] ,
         \DataPath/i_PIPLIN_B[28] , \DataPath/i_PIPLIN_B[29] ,
         \DataPath/i_PIPLIN_B[30] , \DataPath/i_PIPLIN_B[31] ,
         \DataPath/i_PIPLIN_A[31] , \DataPath/i_PIPLIN_A[30] ,
         \DataPath/i_PIPLIN_A[29] , \DataPath/i_PIPLIN_A[28] ,
         \DataPath/i_PIPLIN_A[27] , \DataPath/i_PIPLIN_A[26] ,
         \DataPath/i_PIPLIN_A[25] , \DataPath/i_PIPLIN_A[24] ,
         \DataPath/i_PIPLIN_A[23] , \DataPath/i_PIPLIN_A[22] ,
         \DataPath/i_PIPLIN_A[21] , \DataPath/i_PIPLIN_A[20] ,
         \DataPath/i_PIPLIN_A[19] , \DataPath/i_PIPLIN_A[18] ,
         \DataPath/i_PIPLIN_A[17] , \DataPath/i_PIPLIN_A[16] ,
         \DataPath/i_PIPLIN_A[15] , \DataPath/i_PIPLIN_A[14] ,
         \DataPath/i_PIPLIN_A[13] , \DataPath/i_PIPLIN_A[12] ,
         \DataPath/i_PIPLIN_A[11] , \DataPath/i_PIPLIN_A[10] ,
         \DataPath/i_PIPLIN_A[9] , \DataPath/i_PIPLIN_A[8] ,
         \DataPath/i_PIPLIN_A[7] , \DataPath/i_PIPLIN_A[6] ,
         \DataPath/i_PIPLIN_A[5] , \DataPath/i_PIPLIN_A[4] ,
         \DataPath/i_PIPLIN_A[3] , \DataPath/i_PIPLIN_A[2] ,
         \DataPath/i_PIPLIN_A[1] , \DataPath/i_PIPLIN_A[0] ,
         \DataPath/RF/bus_sel_savedwin_data[511] ,
         \DataPath/RF/bus_sel_savedwin_data[510] ,
         \DataPath/RF/bus_sel_savedwin_data[509] ,
         \DataPath/RF/bus_sel_savedwin_data[508] ,
         \DataPath/RF/bus_sel_savedwin_data[507] ,
         \DataPath/RF/bus_sel_savedwin_data[506] ,
         \DataPath/RF/bus_sel_savedwin_data[505] ,
         \DataPath/RF/bus_sel_savedwin_data[504] ,
         \DataPath/RF/bus_sel_savedwin_data[503] ,
         \DataPath/RF/bus_sel_savedwin_data[502] ,
         \DataPath/RF/bus_sel_savedwin_data[501] ,
         \DataPath/RF/bus_sel_savedwin_data[500] ,
         \DataPath/RF/bus_sel_savedwin_data[499] ,
         \DataPath/RF/bus_sel_savedwin_data[498] ,
         \DataPath/RF/bus_sel_savedwin_data[497] ,
         \DataPath/RF/bus_sel_savedwin_data[496] ,
         \DataPath/RF/bus_sel_savedwin_data[495] ,
         \DataPath/RF/bus_sel_savedwin_data[494] ,
         \DataPath/RF/bus_sel_savedwin_data[493] ,
         \DataPath/RF/bus_sel_savedwin_data[492] ,
         \DataPath/RF/bus_sel_savedwin_data[491] ,
         \DataPath/RF/bus_sel_savedwin_data[490] ,
         \DataPath/RF/bus_sel_savedwin_data[489] ,
         \DataPath/RF/bus_sel_savedwin_data[488] ,
         \DataPath/RF/bus_sel_savedwin_data[487] ,
         \DataPath/RF/bus_sel_savedwin_data[486] ,
         \DataPath/RF/bus_sel_savedwin_data[485] ,
         \DataPath/RF/bus_sel_savedwin_data[484] ,
         \DataPath/RF/bus_sel_savedwin_data[483] ,
         \DataPath/RF/bus_sel_savedwin_data[482] ,
         \DataPath/RF/bus_sel_savedwin_data[481] ,
         \DataPath/RF/bus_sel_savedwin_data[480] ,
         \DataPath/RF/bus_sel_savedwin_data[479] ,
         \DataPath/RF/bus_sel_savedwin_data[478] ,
         \DataPath/RF/bus_sel_savedwin_data[477] ,
         \DataPath/RF/bus_sel_savedwin_data[476] ,
         \DataPath/RF/bus_sel_savedwin_data[475] ,
         \DataPath/RF/bus_sel_savedwin_data[474] ,
         \DataPath/RF/bus_sel_savedwin_data[473] ,
         \DataPath/RF/bus_sel_savedwin_data[472] ,
         \DataPath/RF/bus_sel_savedwin_data[471] ,
         \DataPath/RF/bus_sel_savedwin_data[470] ,
         \DataPath/RF/bus_sel_savedwin_data[469] ,
         \DataPath/RF/bus_sel_savedwin_data[468] ,
         \DataPath/RF/bus_sel_savedwin_data[467] ,
         \DataPath/RF/bus_sel_savedwin_data[466] ,
         \DataPath/RF/bus_sel_savedwin_data[465] ,
         \DataPath/RF/bus_sel_savedwin_data[464] ,
         \DataPath/RF/bus_sel_savedwin_data[463] ,
         \DataPath/RF/bus_sel_savedwin_data[462] ,
         \DataPath/RF/bus_sel_savedwin_data[461] ,
         \DataPath/RF/bus_sel_savedwin_data[460] ,
         \DataPath/RF/bus_sel_savedwin_data[459] ,
         \DataPath/RF/bus_sel_savedwin_data[458] ,
         \DataPath/RF/bus_sel_savedwin_data[457] ,
         \DataPath/RF/bus_sel_savedwin_data[456] ,
         \DataPath/RF/bus_sel_savedwin_data[455] ,
         \DataPath/RF/bus_sel_savedwin_data[454] ,
         \DataPath/RF/bus_sel_savedwin_data[453] ,
         \DataPath/RF/bus_sel_savedwin_data[452] ,
         \DataPath/RF/bus_sel_savedwin_data[451] ,
         \DataPath/RF/bus_sel_savedwin_data[450] ,
         \DataPath/RF/bus_sel_savedwin_data[449] ,
         \DataPath/RF/bus_sel_savedwin_data[448] ,
         \DataPath/RF/bus_sel_savedwin_data[447] ,
         \DataPath/RF/bus_sel_savedwin_data[446] ,
         \DataPath/RF/bus_sel_savedwin_data[445] ,
         \DataPath/RF/bus_sel_savedwin_data[444] ,
         \DataPath/RF/bus_sel_savedwin_data[443] ,
         \DataPath/RF/bus_sel_savedwin_data[442] ,
         \DataPath/RF/bus_sel_savedwin_data[441] ,
         \DataPath/RF/bus_sel_savedwin_data[440] ,
         \DataPath/RF/bus_sel_savedwin_data[439] ,
         \DataPath/RF/bus_sel_savedwin_data[438] ,
         \DataPath/RF/bus_sel_savedwin_data[437] ,
         \DataPath/RF/bus_sel_savedwin_data[436] ,
         \DataPath/RF/bus_sel_savedwin_data[435] ,
         \DataPath/RF/bus_sel_savedwin_data[434] ,
         \DataPath/RF/bus_sel_savedwin_data[433] ,
         \DataPath/RF/bus_sel_savedwin_data[432] ,
         \DataPath/RF/bus_sel_savedwin_data[431] ,
         \DataPath/RF/bus_sel_savedwin_data[430] ,
         \DataPath/RF/bus_sel_savedwin_data[429] ,
         \DataPath/RF/bus_sel_savedwin_data[428] ,
         \DataPath/RF/bus_sel_savedwin_data[427] ,
         \DataPath/RF/bus_sel_savedwin_data[426] ,
         \DataPath/RF/bus_sel_savedwin_data[425] ,
         \DataPath/RF/bus_sel_savedwin_data[424] ,
         \DataPath/RF/bus_sel_savedwin_data[423] ,
         \DataPath/RF/bus_sel_savedwin_data[422] ,
         \DataPath/RF/bus_sel_savedwin_data[421] ,
         \DataPath/RF/bus_sel_savedwin_data[420] ,
         \DataPath/RF/bus_sel_savedwin_data[419] ,
         \DataPath/RF/bus_sel_savedwin_data[418] ,
         \DataPath/RF/bus_sel_savedwin_data[417] ,
         \DataPath/RF/bus_sel_savedwin_data[416] ,
         \DataPath/RF/bus_sel_savedwin_data[415] ,
         \DataPath/RF/bus_sel_savedwin_data[414] ,
         \DataPath/RF/bus_sel_savedwin_data[413] ,
         \DataPath/RF/bus_sel_savedwin_data[412] ,
         \DataPath/RF/bus_sel_savedwin_data[411] ,
         \DataPath/RF/bus_sel_savedwin_data[410] ,
         \DataPath/RF/bus_sel_savedwin_data[409] ,
         \DataPath/RF/bus_sel_savedwin_data[408] ,
         \DataPath/RF/bus_sel_savedwin_data[407] ,
         \DataPath/RF/bus_sel_savedwin_data[406] ,
         \DataPath/RF/bus_sel_savedwin_data[405] ,
         \DataPath/RF/bus_sel_savedwin_data[404] ,
         \DataPath/RF/bus_sel_savedwin_data[403] ,
         \DataPath/RF/bus_sel_savedwin_data[402] ,
         \DataPath/RF/bus_sel_savedwin_data[401] ,
         \DataPath/RF/bus_sel_savedwin_data[400] ,
         \DataPath/RF/bus_sel_savedwin_data[399] ,
         \DataPath/RF/bus_sel_savedwin_data[398] ,
         \DataPath/RF/bus_sel_savedwin_data[397] ,
         \DataPath/RF/bus_sel_savedwin_data[396] ,
         \DataPath/RF/bus_sel_savedwin_data[395] ,
         \DataPath/RF/bus_sel_savedwin_data[394] ,
         \DataPath/RF/bus_sel_savedwin_data[393] ,
         \DataPath/RF/bus_sel_savedwin_data[392] ,
         \DataPath/RF/bus_sel_savedwin_data[391] ,
         \DataPath/RF/bus_sel_savedwin_data[390] ,
         \DataPath/RF/bus_sel_savedwin_data[389] ,
         \DataPath/RF/bus_sel_savedwin_data[388] ,
         \DataPath/RF/bus_sel_savedwin_data[387] ,
         \DataPath/RF/bus_sel_savedwin_data[386] ,
         \DataPath/RF/bus_sel_savedwin_data[385] ,
         \DataPath/RF/bus_sel_savedwin_data[384] ,
         \DataPath/RF/bus_sel_savedwin_data[383] ,
         \DataPath/RF/bus_sel_savedwin_data[382] ,
         \DataPath/RF/bus_sel_savedwin_data[381] ,
         \DataPath/RF/bus_sel_savedwin_data[380] ,
         \DataPath/RF/bus_sel_savedwin_data[379] ,
         \DataPath/RF/bus_sel_savedwin_data[378] ,
         \DataPath/RF/bus_sel_savedwin_data[377] ,
         \DataPath/RF/bus_sel_savedwin_data[376] ,
         \DataPath/RF/bus_sel_savedwin_data[375] ,
         \DataPath/RF/bus_sel_savedwin_data[374] ,
         \DataPath/RF/bus_sel_savedwin_data[373] ,
         \DataPath/RF/bus_sel_savedwin_data[372] ,
         \DataPath/RF/bus_sel_savedwin_data[371] ,
         \DataPath/RF/bus_sel_savedwin_data[370] ,
         \DataPath/RF/bus_sel_savedwin_data[369] ,
         \DataPath/RF/bus_sel_savedwin_data[368] ,
         \DataPath/RF/bus_sel_savedwin_data[367] ,
         \DataPath/RF/bus_sel_savedwin_data[366] ,
         \DataPath/RF/bus_sel_savedwin_data[365] ,
         \DataPath/RF/bus_sel_savedwin_data[364] ,
         \DataPath/RF/bus_sel_savedwin_data[363] ,
         \DataPath/RF/bus_sel_savedwin_data[362] ,
         \DataPath/RF/bus_sel_savedwin_data[361] ,
         \DataPath/RF/bus_sel_savedwin_data[360] ,
         \DataPath/RF/bus_sel_savedwin_data[359] ,
         \DataPath/RF/bus_sel_savedwin_data[358] ,
         \DataPath/RF/bus_sel_savedwin_data[357] ,
         \DataPath/RF/bus_sel_savedwin_data[356] ,
         \DataPath/RF/bus_sel_savedwin_data[355] ,
         \DataPath/RF/bus_sel_savedwin_data[354] ,
         \DataPath/RF/bus_sel_savedwin_data[353] ,
         \DataPath/RF/bus_sel_savedwin_data[352] ,
         \DataPath/RF/bus_sel_savedwin_data[351] ,
         \DataPath/RF/bus_sel_savedwin_data[350] ,
         \DataPath/RF/bus_sel_savedwin_data[349] ,
         \DataPath/RF/bus_sel_savedwin_data[348] ,
         \DataPath/RF/bus_sel_savedwin_data[347] ,
         \DataPath/RF/bus_sel_savedwin_data[346] ,
         \DataPath/RF/bus_sel_savedwin_data[345] ,
         \DataPath/RF/bus_sel_savedwin_data[344] ,
         \DataPath/RF/bus_sel_savedwin_data[343] ,
         \DataPath/RF/bus_sel_savedwin_data[342] ,
         \DataPath/RF/bus_sel_savedwin_data[341] ,
         \DataPath/RF/bus_sel_savedwin_data[340] ,
         \DataPath/RF/bus_sel_savedwin_data[339] ,
         \DataPath/RF/bus_sel_savedwin_data[338] ,
         \DataPath/RF/bus_sel_savedwin_data[337] ,
         \DataPath/RF/bus_sel_savedwin_data[336] ,
         \DataPath/RF/bus_sel_savedwin_data[335] ,
         \DataPath/RF/bus_sel_savedwin_data[334] ,
         \DataPath/RF/bus_sel_savedwin_data[333] ,
         \DataPath/RF/bus_sel_savedwin_data[332] ,
         \DataPath/RF/bus_sel_savedwin_data[331] ,
         \DataPath/RF/bus_sel_savedwin_data[330] ,
         \DataPath/RF/bus_sel_savedwin_data[329] ,
         \DataPath/RF/bus_sel_savedwin_data[328] ,
         \DataPath/RF/bus_sel_savedwin_data[327] ,
         \DataPath/RF/bus_sel_savedwin_data[326] ,
         \DataPath/RF/bus_sel_savedwin_data[325] ,
         \DataPath/RF/bus_sel_savedwin_data[324] ,
         \DataPath/RF/bus_sel_savedwin_data[323] ,
         \DataPath/RF/bus_sel_savedwin_data[322] ,
         \DataPath/RF/bus_sel_savedwin_data[321] ,
         \DataPath/RF/bus_sel_savedwin_data[320] ,
         \DataPath/RF/bus_sel_savedwin_data[319] ,
         \DataPath/RF/bus_sel_savedwin_data[318] ,
         \DataPath/RF/bus_sel_savedwin_data[317] ,
         \DataPath/RF/bus_sel_savedwin_data[316] ,
         \DataPath/RF/bus_sel_savedwin_data[315] ,
         \DataPath/RF/bus_sel_savedwin_data[314] ,
         \DataPath/RF/bus_sel_savedwin_data[313] ,
         \DataPath/RF/bus_sel_savedwin_data[312] ,
         \DataPath/RF/bus_sel_savedwin_data[311] ,
         \DataPath/RF/bus_sel_savedwin_data[310] ,
         \DataPath/RF/bus_sel_savedwin_data[309] ,
         \DataPath/RF/bus_sel_savedwin_data[308] ,
         \DataPath/RF/bus_sel_savedwin_data[307] ,
         \DataPath/RF/bus_sel_savedwin_data[306] ,
         \DataPath/RF/bus_sel_savedwin_data[305] ,
         \DataPath/RF/bus_sel_savedwin_data[304] ,
         \DataPath/RF/bus_sel_savedwin_data[303] ,
         \DataPath/RF/bus_sel_savedwin_data[302] ,
         \DataPath/RF/bus_sel_savedwin_data[301] ,
         \DataPath/RF/bus_sel_savedwin_data[300] ,
         \DataPath/RF/bus_sel_savedwin_data[299] ,
         \DataPath/RF/bus_sel_savedwin_data[298] ,
         \DataPath/RF/bus_sel_savedwin_data[297] ,
         \DataPath/RF/bus_sel_savedwin_data[296] ,
         \DataPath/RF/bus_sel_savedwin_data[295] ,
         \DataPath/RF/bus_sel_savedwin_data[294] ,
         \DataPath/RF/bus_sel_savedwin_data[293] ,
         \DataPath/RF/bus_sel_savedwin_data[292] ,
         \DataPath/RF/bus_sel_savedwin_data[291] ,
         \DataPath/RF/bus_sel_savedwin_data[290] ,
         \DataPath/RF/bus_sel_savedwin_data[289] ,
         \DataPath/RF/bus_sel_savedwin_data[288] ,
         \DataPath/RF/bus_sel_savedwin_data[287] ,
         \DataPath/RF/bus_sel_savedwin_data[286] ,
         \DataPath/RF/bus_sel_savedwin_data[285] ,
         \DataPath/RF/bus_sel_savedwin_data[284] ,
         \DataPath/RF/bus_sel_savedwin_data[283] ,
         \DataPath/RF/bus_sel_savedwin_data[282] ,
         \DataPath/RF/bus_sel_savedwin_data[281] ,
         \DataPath/RF/bus_sel_savedwin_data[280] ,
         \DataPath/RF/bus_sel_savedwin_data[279] ,
         \DataPath/RF/bus_sel_savedwin_data[278] ,
         \DataPath/RF/bus_sel_savedwin_data[277] ,
         \DataPath/RF/bus_sel_savedwin_data[276] ,
         \DataPath/RF/bus_sel_savedwin_data[275] ,
         \DataPath/RF/bus_sel_savedwin_data[274] ,
         \DataPath/RF/bus_sel_savedwin_data[273] ,
         \DataPath/RF/bus_sel_savedwin_data[272] ,
         \DataPath/RF/bus_sel_savedwin_data[271] ,
         \DataPath/RF/bus_sel_savedwin_data[270] ,
         \DataPath/RF/bus_sel_savedwin_data[269] ,
         \DataPath/RF/bus_sel_savedwin_data[268] ,
         \DataPath/RF/bus_sel_savedwin_data[267] ,
         \DataPath/RF/bus_sel_savedwin_data[266] ,
         \DataPath/RF/bus_sel_savedwin_data[265] ,
         \DataPath/RF/bus_sel_savedwin_data[264] ,
         \DataPath/RF/bus_sel_savedwin_data[263] ,
         \DataPath/RF/bus_sel_savedwin_data[262] ,
         \DataPath/RF/bus_sel_savedwin_data[261] ,
         \DataPath/RF/bus_sel_savedwin_data[260] ,
         \DataPath/RF/bus_sel_savedwin_data[259] ,
         \DataPath/RF/bus_sel_savedwin_data[258] ,
         \DataPath/RF/bus_sel_savedwin_data[257] ,
         \DataPath/RF/bus_sel_savedwin_data[256] ,
         \DataPath/RF/bus_sel_savedwin_data[255] ,
         \DataPath/RF/bus_sel_savedwin_data[254] ,
         \DataPath/RF/bus_sel_savedwin_data[253] ,
         \DataPath/RF/bus_sel_savedwin_data[252] ,
         \DataPath/RF/bus_sel_savedwin_data[251] ,
         \DataPath/RF/bus_sel_savedwin_data[250] ,
         \DataPath/RF/bus_sel_savedwin_data[249] ,
         \DataPath/RF/bus_sel_savedwin_data[248] ,
         \DataPath/RF/bus_sel_savedwin_data[247] ,
         \DataPath/RF/bus_sel_savedwin_data[246] ,
         \DataPath/RF/bus_sel_savedwin_data[245] ,
         \DataPath/RF/bus_sel_savedwin_data[244] ,
         \DataPath/RF/bus_sel_savedwin_data[243] ,
         \DataPath/RF/bus_sel_savedwin_data[242] ,
         \DataPath/RF/bus_sel_savedwin_data[241] ,
         \DataPath/RF/bus_sel_savedwin_data[240] ,
         \DataPath/RF/bus_sel_savedwin_data[239] ,
         \DataPath/RF/bus_sel_savedwin_data[238] ,
         \DataPath/RF/bus_sel_savedwin_data[237] ,
         \DataPath/RF/bus_sel_savedwin_data[236] ,
         \DataPath/RF/bus_sel_savedwin_data[235] ,
         \DataPath/RF/bus_sel_savedwin_data[234] ,
         \DataPath/RF/bus_sel_savedwin_data[233] ,
         \DataPath/RF/bus_sel_savedwin_data[232] ,
         \DataPath/RF/bus_sel_savedwin_data[231] ,
         \DataPath/RF/bus_sel_savedwin_data[230] ,
         \DataPath/RF/bus_sel_savedwin_data[229] ,
         \DataPath/RF/bus_sel_savedwin_data[228] ,
         \DataPath/RF/bus_sel_savedwin_data[227] ,
         \DataPath/RF/bus_sel_savedwin_data[226] ,
         \DataPath/RF/bus_sel_savedwin_data[225] ,
         \DataPath/RF/bus_sel_savedwin_data[224] ,
         \DataPath/RF/bus_sel_savedwin_data[223] ,
         \DataPath/RF/bus_sel_savedwin_data[222] ,
         \DataPath/RF/bus_sel_savedwin_data[221] ,
         \DataPath/RF/bus_sel_savedwin_data[220] ,
         \DataPath/RF/bus_sel_savedwin_data[219] ,
         \DataPath/RF/bus_sel_savedwin_data[218] ,
         \DataPath/RF/bus_sel_savedwin_data[217] ,
         \DataPath/RF/bus_sel_savedwin_data[216] ,
         \DataPath/RF/bus_sel_savedwin_data[215] ,
         \DataPath/RF/bus_sel_savedwin_data[214] ,
         \DataPath/RF/bus_sel_savedwin_data[213] ,
         \DataPath/RF/bus_sel_savedwin_data[212] ,
         \DataPath/RF/bus_sel_savedwin_data[211] ,
         \DataPath/RF/bus_sel_savedwin_data[210] ,
         \DataPath/RF/bus_sel_savedwin_data[209] ,
         \DataPath/RF/bus_sel_savedwin_data[208] ,
         \DataPath/RF/bus_sel_savedwin_data[207] ,
         \DataPath/RF/bus_sel_savedwin_data[206] ,
         \DataPath/RF/bus_sel_savedwin_data[205] ,
         \DataPath/RF/bus_sel_savedwin_data[204] ,
         \DataPath/RF/bus_sel_savedwin_data[203] ,
         \DataPath/RF/bus_sel_savedwin_data[202] ,
         \DataPath/RF/bus_sel_savedwin_data[201] ,
         \DataPath/RF/bus_sel_savedwin_data[200] ,
         \DataPath/RF/bus_sel_savedwin_data[199] ,
         \DataPath/RF/bus_sel_savedwin_data[198] ,
         \DataPath/RF/bus_sel_savedwin_data[197] ,
         \DataPath/RF/bus_sel_savedwin_data[196] ,
         \DataPath/RF/bus_sel_savedwin_data[195] ,
         \DataPath/RF/bus_sel_savedwin_data[194] ,
         \DataPath/RF/bus_sel_savedwin_data[193] ,
         \DataPath/RF/bus_sel_savedwin_data[192] ,
         \DataPath/RF/bus_sel_savedwin_data[191] ,
         \DataPath/RF/bus_sel_savedwin_data[190] ,
         \DataPath/RF/bus_sel_savedwin_data[189] ,
         \DataPath/RF/bus_sel_savedwin_data[188] ,
         \DataPath/RF/bus_sel_savedwin_data[187] ,
         \DataPath/RF/bus_sel_savedwin_data[186] ,
         \DataPath/RF/bus_sel_savedwin_data[185] ,
         \DataPath/RF/bus_sel_savedwin_data[184] ,
         \DataPath/RF/bus_sel_savedwin_data[183] ,
         \DataPath/RF/bus_sel_savedwin_data[182] ,
         \DataPath/RF/bus_sel_savedwin_data[181] ,
         \DataPath/RF/bus_sel_savedwin_data[180] ,
         \DataPath/RF/bus_sel_savedwin_data[179] ,
         \DataPath/RF/bus_sel_savedwin_data[178] ,
         \DataPath/RF/bus_sel_savedwin_data[177] ,
         \DataPath/RF/bus_sel_savedwin_data[176] ,
         \DataPath/RF/bus_sel_savedwin_data[175] ,
         \DataPath/RF/bus_sel_savedwin_data[174] ,
         \DataPath/RF/bus_sel_savedwin_data[173] ,
         \DataPath/RF/bus_sel_savedwin_data[172] ,
         \DataPath/RF/bus_sel_savedwin_data[171] ,
         \DataPath/RF/bus_sel_savedwin_data[170] ,
         \DataPath/RF/bus_sel_savedwin_data[169] ,
         \DataPath/RF/bus_sel_savedwin_data[168] ,
         \DataPath/RF/bus_sel_savedwin_data[167] ,
         \DataPath/RF/bus_sel_savedwin_data[166] ,
         \DataPath/RF/bus_sel_savedwin_data[165] ,
         \DataPath/RF/bus_sel_savedwin_data[164] ,
         \DataPath/RF/bus_sel_savedwin_data[163] ,
         \DataPath/RF/bus_sel_savedwin_data[162] ,
         \DataPath/RF/bus_sel_savedwin_data[161] ,
         \DataPath/RF/bus_sel_savedwin_data[160] ,
         \DataPath/RF/bus_sel_savedwin_data[159] ,
         \DataPath/RF/bus_sel_savedwin_data[158] ,
         \DataPath/RF/bus_sel_savedwin_data[157] ,
         \DataPath/RF/bus_sel_savedwin_data[156] ,
         \DataPath/RF/bus_sel_savedwin_data[155] ,
         \DataPath/RF/bus_sel_savedwin_data[154] ,
         \DataPath/RF/bus_sel_savedwin_data[153] ,
         \DataPath/RF/bus_sel_savedwin_data[152] ,
         \DataPath/RF/bus_sel_savedwin_data[151] ,
         \DataPath/RF/bus_sel_savedwin_data[150] ,
         \DataPath/RF/bus_sel_savedwin_data[149] ,
         \DataPath/RF/bus_sel_savedwin_data[148] ,
         \DataPath/RF/bus_sel_savedwin_data[147] ,
         \DataPath/RF/bus_sel_savedwin_data[146] ,
         \DataPath/RF/bus_sel_savedwin_data[145] ,
         \DataPath/RF/bus_sel_savedwin_data[144] ,
         \DataPath/RF/bus_sel_savedwin_data[143] ,
         \DataPath/RF/bus_sel_savedwin_data[142] ,
         \DataPath/RF/bus_sel_savedwin_data[141] ,
         \DataPath/RF/bus_sel_savedwin_data[140] ,
         \DataPath/RF/bus_sel_savedwin_data[139] ,
         \DataPath/RF/bus_sel_savedwin_data[138] ,
         \DataPath/RF/bus_sel_savedwin_data[137] ,
         \DataPath/RF/bus_sel_savedwin_data[136] ,
         \DataPath/RF/bus_sel_savedwin_data[135] ,
         \DataPath/RF/bus_sel_savedwin_data[134] ,
         \DataPath/RF/bus_sel_savedwin_data[133] ,
         \DataPath/RF/bus_sel_savedwin_data[132] ,
         \DataPath/RF/bus_sel_savedwin_data[131] ,
         \DataPath/RF/bus_sel_savedwin_data[130] ,
         \DataPath/RF/bus_sel_savedwin_data[129] ,
         \DataPath/RF/bus_sel_savedwin_data[128] ,
         \DataPath/RF/bus_sel_savedwin_data[127] ,
         \DataPath/RF/bus_sel_savedwin_data[126] ,
         \DataPath/RF/bus_sel_savedwin_data[125] ,
         \DataPath/RF/bus_sel_savedwin_data[124] ,
         \DataPath/RF/bus_sel_savedwin_data[123] ,
         \DataPath/RF/bus_sel_savedwin_data[122] ,
         \DataPath/RF/bus_sel_savedwin_data[121] ,
         \DataPath/RF/bus_sel_savedwin_data[120] ,
         \DataPath/RF/bus_sel_savedwin_data[119] ,
         \DataPath/RF/bus_sel_savedwin_data[118] ,
         \DataPath/RF/bus_sel_savedwin_data[117] ,
         \DataPath/RF/bus_sel_savedwin_data[116] ,
         \DataPath/RF/bus_sel_savedwin_data[115] ,
         \DataPath/RF/bus_sel_savedwin_data[114] ,
         \DataPath/RF/bus_sel_savedwin_data[113] ,
         \DataPath/RF/bus_sel_savedwin_data[112] ,
         \DataPath/RF/bus_sel_savedwin_data[111] ,
         \DataPath/RF/bus_sel_savedwin_data[110] ,
         \DataPath/RF/bus_sel_savedwin_data[109] ,
         \DataPath/RF/bus_sel_savedwin_data[108] ,
         \DataPath/RF/bus_sel_savedwin_data[107] ,
         \DataPath/RF/bus_sel_savedwin_data[106] ,
         \DataPath/RF/bus_sel_savedwin_data[105] ,
         \DataPath/RF/bus_sel_savedwin_data[104] ,
         \DataPath/RF/bus_sel_savedwin_data[103] ,
         \DataPath/RF/bus_sel_savedwin_data[102] ,
         \DataPath/RF/bus_sel_savedwin_data[101] ,
         \DataPath/RF/bus_sel_savedwin_data[100] ,
         \DataPath/RF/bus_sel_savedwin_data[99] ,
         \DataPath/RF/bus_sel_savedwin_data[98] ,
         \DataPath/RF/bus_sel_savedwin_data[97] ,
         \DataPath/RF/bus_sel_savedwin_data[96] ,
         \DataPath/RF/bus_sel_savedwin_data[95] ,
         \DataPath/RF/bus_sel_savedwin_data[94] ,
         \DataPath/RF/bus_sel_savedwin_data[93] ,
         \DataPath/RF/bus_sel_savedwin_data[92] ,
         \DataPath/RF/bus_sel_savedwin_data[91] ,
         \DataPath/RF/bus_sel_savedwin_data[90] ,
         \DataPath/RF/bus_sel_savedwin_data[89] ,
         \DataPath/RF/bus_sel_savedwin_data[88] ,
         \DataPath/RF/bus_sel_savedwin_data[87] ,
         \DataPath/RF/bus_sel_savedwin_data[86] ,
         \DataPath/RF/bus_sel_savedwin_data[85] ,
         \DataPath/RF/bus_sel_savedwin_data[84] ,
         \DataPath/RF/bus_sel_savedwin_data[83] ,
         \DataPath/RF/bus_sel_savedwin_data[82] ,
         \DataPath/RF/bus_sel_savedwin_data[81] ,
         \DataPath/RF/bus_sel_savedwin_data[80] ,
         \DataPath/RF/bus_sel_savedwin_data[79] ,
         \DataPath/RF/bus_sel_savedwin_data[78] ,
         \DataPath/RF/bus_sel_savedwin_data[77] ,
         \DataPath/RF/bus_sel_savedwin_data[76] ,
         \DataPath/RF/bus_sel_savedwin_data[75] ,
         \DataPath/RF/bus_sel_savedwin_data[74] ,
         \DataPath/RF/bus_sel_savedwin_data[73] ,
         \DataPath/RF/bus_sel_savedwin_data[72] ,
         \DataPath/RF/bus_sel_savedwin_data[71] ,
         \DataPath/RF/bus_sel_savedwin_data[70] ,
         \DataPath/RF/bus_sel_savedwin_data[69] ,
         \DataPath/RF/bus_sel_savedwin_data[68] ,
         \DataPath/RF/bus_sel_savedwin_data[67] ,
         \DataPath/RF/bus_sel_savedwin_data[66] ,
         \DataPath/RF/bus_sel_savedwin_data[65] ,
         \DataPath/RF/bus_sel_savedwin_data[64] ,
         \DataPath/RF/bus_sel_savedwin_data[63] ,
         \DataPath/RF/bus_sel_savedwin_data[62] ,
         \DataPath/RF/bus_sel_savedwin_data[61] ,
         \DataPath/RF/bus_sel_savedwin_data[60] ,
         \DataPath/RF/bus_sel_savedwin_data[59] ,
         \DataPath/RF/bus_sel_savedwin_data[58] ,
         \DataPath/RF/bus_sel_savedwin_data[57] ,
         \DataPath/RF/bus_sel_savedwin_data[56] ,
         \DataPath/RF/bus_sel_savedwin_data[55] ,
         \DataPath/RF/bus_sel_savedwin_data[54] ,
         \DataPath/RF/bus_sel_savedwin_data[53] ,
         \DataPath/RF/bus_sel_savedwin_data[52] ,
         \DataPath/RF/bus_sel_savedwin_data[51] ,
         \DataPath/RF/bus_sel_savedwin_data[50] ,
         \DataPath/RF/bus_sel_savedwin_data[49] ,
         \DataPath/RF/bus_sel_savedwin_data[48] ,
         \DataPath/RF/bus_sel_savedwin_data[47] ,
         \DataPath/RF/bus_sel_savedwin_data[46] ,
         \DataPath/RF/bus_sel_savedwin_data[45] ,
         \DataPath/RF/bus_sel_savedwin_data[44] ,
         \DataPath/RF/bus_sel_savedwin_data[43] ,
         \DataPath/RF/bus_sel_savedwin_data[42] ,
         \DataPath/RF/bus_sel_savedwin_data[41] ,
         \DataPath/RF/bus_sel_savedwin_data[40] ,
         \DataPath/RF/bus_sel_savedwin_data[39] ,
         \DataPath/RF/bus_sel_savedwin_data[38] ,
         \DataPath/RF/bus_sel_savedwin_data[37] ,
         \DataPath/RF/bus_sel_savedwin_data[36] ,
         \DataPath/RF/bus_sel_savedwin_data[35] ,
         \DataPath/RF/bus_sel_savedwin_data[34] ,
         \DataPath/RF/bus_sel_savedwin_data[33] ,
         \DataPath/RF/bus_sel_savedwin_data[32] ,
         \DataPath/RF/bus_sel_savedwin_data[31] ,
         \DataPath/RF/bus_sel_savedwin_data[30] ,
         \DataPath/RF/bus_sel_savedwin_data[29] ,
         \DataPath/RF/bus_sel_savedwin_data[28] ,
         \DataPath/RF/bus_sel_savedwin_data[27] ,
         \DataPath/RF/bus_sel_savedwin_data[26] ,
         \DataPath/RF/bus_sel_savedwin_data[25] ,
         \DataPath/RF/bus_sel_savedwin_data[24] ,
         \DataPath/RF/bus_sel_savedwin_data[23] ,
         \DataPath/RF/bus_sel_savedwin_data[22] ,
         \DataPath/RF/bus_sel_savedwin_data[21] ,
         \DataPath/RF/bus_sel_savedwin_data[20] ,
         \DataPath/RF/bus_sel_savedwin_data[19] ,
         \DataPath/RF/bus_sel_savedwin_data[18] ,
         \DataPath/RF/bus_sel_savedwin_data[17] ,
         \DataPath/RF/bus_sel_savedwin_data[16] ,
         \DataPath/RF/bus_sel_savedwin_data[15] ,
         \DataPath/RF/bus_sel_savedwin_data[14] ,
         \DataPath/RF/bus_sel_savedwin_data[13] ,
         \DataPath/RF/bus_sel_savedwin_data[12] ,
         \DataPath/RF/bus_sel_savedwin_data[11] ,
         \DataPath/RF/bus_sel_savedwin_data[10] ,
         \DataPath/RF/bus_sel_savedwin_data[9] ,
         \DataPath/RF/bus_sel_savedwin_data[8] ,
         \DataPath/RF/bus_sel_savedwin_data[7] ,
         \DataPath/RF/bus_sel_savedwin_data[6] ,
         \DataPath/RF/bus_sel_savedwin_data[5] ,
         \DataPath/RF/bus_sel_savedwin_data[4] ,
         \DataPath/RF/bus_sel_savedwin_data[3] ,
         \DataPath/RF/bus_sel_savedwin_data[2] ,
         \DataPath/RF/bus_sel_savedwin_data[1] ,
         \DataPath/RF/bus_sel_savedwin_data[0] , \DataPath/RF/c_swin[0] ,
         \DataPath/RF/c_swin[1] , \DataPath/RF/c_swin[2] ,
         \DataPath/RF/c_swin[3] , \DataPath/RF/internal_out2[31] ,
         \DataPath/RF/internal_out2[30] , \DataPath/RF/internal_out2[29] ,
         \DataPath/RF/internal_out2[28] , \DataPath/RF/internal_out2[27] ,
         \DataPath/RF/internal_out2[26] , \DataPath/RF/internal_out2[25] ,
         \DataPath/RF/internal_out2[24] , \DataPath/RF/internal_out2[23] ,
         \DataPath/RF/internal_out2[22] , \DataPath/RF/internal_out2[21] ,
         \DataPath/RF/internal_out2[20] , \DataPath/RF/internal_out2[19] ,
         \DataPath/RF/internal_out2[18] , \DataPath/RF/internal_out2[17] ,
         \DataPath/RF/internal_out2[16] , \DataPath/RF/internal_out2[15] ,
         \DataPath/RF/internal_out2[14] , \DataPath/RF/internal_out2[13] ,
         \DataPath/RF/internal_out2[12] , \DataPath/RF/internal_out2[11] ,
         \DataPath/RF/internal_out2[10] , \DataPath/RF/internal_out2[9] ,
         \DataPath/RF/internal_out2[8] , \DataPath/RF/internal_out2[7] ,
         \DataPath/RF/internal_out2[6] , \DataPath/RF/internal_out2[5] ,
         \DataPath/RF/internal_out2[4] , \DataPath/RF/internal_out2[3] ,
         \DataPath/RF/internal_out2[2] , \DataPath/RF/internal_out2[1] ,
         \DataPath/RF/internal_out2[0] , \DataPath/RF/internal_out1[31] ,
         \DataPath/RF/internal_out1[30] , \DataPath/RF/internal_out1[29] ,
         \DataPath/RF/internal_out1[28] , \DataPath/RF/internal_out1[27] ,
         \DataPath/RF/internal_out1[26] , \DataPath/RF/internal_out1[25] ,
         \DataPath/RF/internal_out1[24] , \DataPath/RF/internal_out1[23] ,
         \DataPath/RF/internal_out1[22] , \DataPath/RF/internal_out1[21] ,
         \DataPath/RF/internal_out1[20] , \DataPath/RF/internal_out1[19] ,
         \DataPath/RF/internal_out1[18] , \DataPath/RF/internal_out1[17] ,
         \DataPath/RF/internal_out1[16] , \DataPath/RF/internal_out1[15] ,
         \DataPath/RF/internal_out1[14] , \DataPath/RF/internal_out1[13] ,
         \DataPath/RF/internal_out1[12] , \DataPath/RF/internal_out1[11] ,
         \DataPath/RF/internal_out1[10] , \DataPath/RF/internal_out1[9] ,
         \DataPath/RF/internal_out1[8] , \DataPath/RF/internal_out1[7] ,
         \DataPath/RF/internal_out1[6] , \DataPath/RF/internal_out1[5] ,
         \DataPath/RF/internal_out1[4] , \DataPath/RF/internal_out1[3] ,
         \DataPath/RF/internal_out1[2] , \DataPath/RF/internal_out1[1] ,
         \DataPath/RF/internal_out1[0] ,
         \DataPath/RF/bus_complete_win_data[32] ,
         \DataPath/RF/bus_complete_win_data[33] ,
         \DataPath/RF/bus_complete_win_data[34] ,
         \DataPath/RF/bus_complete_win_data[35] ,
         \DataPath/RF/bus_complete_win_data[36] ,
         \DataPath/RF/bus_complete_win_data[37] ,
         \DataPath/RF/bus_complete_win_data[38] ,
         \DataPath/RF/bus_complete_win_data[39] ,
         \DataPath/RF/bus_complete_win_data[40] ,
         \DataPath/RF/bus_complete_win_data[41] ,
         \DataPath/RF/bus_complete_win_data[42] ,
         \DataPath/RF/bus_complete_win_data[43] ,
         \DataPath/RF/bus_complete_win_data[44] ,
         \DataPath/RF/bus_complete_win_data[45] ,
         \DataPath/RF/bus_complete_win_data[46] ,
         \DataPath/RF/bus_complete_win_data[47] ,
         \DataPath/RF/bus_complete_win_data[48] ,
         \DataPath/RF/bus_complete_win_data[49] ,
         \DataPath/RF/bus_complete_win_data[50] ,
         \DataPath/RF/bus_complete_win_data[51] ,
         \DataPath/RF/bus_complete_win_data[52] ,
         \DataPath/RF/bus_complete_win_data[53] ,
         \DataPath/RF/bus_complete_win_data[54] ,
         \DataPath/RF/bus_complete_win_data[55] ,
         \DataPath/RF/bus_complete_win_data[56] ,
         \DataPath/RF/bus_complete_win_data[57] ,
         \DataPath/RF/bus_complete_win_data[58] ,
         \DataPath/RF/bus_complete_win_data[59] ,
         \DataPath/RF/bus_complete_win_data[60] ,
         \DataPath/RF/bus_complete_win_data[61] ,
         \DataPath/RF/bus_complete_win_data[62] ,
         \DataPath/RF/bus_complete_win_data[63] ,
         \DataPath/RF/bus_complete_win_data[64] ,
         \DataPath/RF/bus_complete_win_data[65] ,
         \DataPath/RF/bus_complete_win_data[66] ,
         \DataPath/RF/bus_complete_win_data[67] ,
         \DataPath/RF/bus_complete_win_data[68] ,
         \DataPath/RF/bus_complete_win_data[69] ,
         \DataPath/RF/bus_complete_win_data[70] ,
         \DataPath/RF/bus_complete_win_data[71] ,
         \DataPath/RF/bus_complete_win_data[72] ,
         \DataPath/RF/bus_complete_win_data[73] ,
         \DataPath/RF/bus_complete_win_data[74] ,
         \DataPath/RF/bus_complete_win_data[75] ,
         \DataPath/RF/bus_complete_win_data[76] ,
         \DataPath/RF/bus_complete_win_data[77] ,
         \DataPath/RF/bus_complete_win_data[78] ,
         \DataPath/RF/bus_complete_win_data[79] ,
         \DataPath/RF/bus_complete_win_data[80] ,
         \DataPath/RF/bus_complete_win_data[81] ,
         \DataPath/RF/bus_complete_win_data[82] ,
         \DataPath/RF/bus_complete_win_data[83] ,
         \DataPath/RF/bus_complete_win_data[84] ,
         \DataPath/RF/bus_complete_win_data[85] ,
         \DataPath/RF/bus_complete_win_data[86] ,
         \DataPath/RF/bus_complete_win_data[87] ,
         \DataPath/RF/bus_complete_win_data[88] ,
         \DataPath/RF/bus_complete_win_data[89] ,
         \DataPath/RF/bus_complete_win_data[90] ,
         \DataPath/RF/bus_complete_win_data[91] ,
         \DataPath/RF/bus_complete_win_data[92] ,
         \DataPath/RF/bus_complete_win_data[93] ,
         \DataPath/RF/bus_complete_win_data[94] ,
         \DataPath/RF/bus_complete_win_data[95] ,
         \DataPath/RF/bus_complete_win_data[96] ,
         \DataPath/RF/bus_complete_win_data[97] ,
         \DataPath/RF/bus_complete_win_data[98] ,
         \DataPath/RF/bus_complete_win_data[99] ,
         \DataPath/RF/bus_complete_win_data[100] ,
         \DataPath/RF/bus_complete_win_data[101] ,
         \DataPath/RF/bus_complete_win_data[102] ,
         \DataPath/RF/bus_complete_win_data[103] ,
         \DataPath/RF/bus_complete_win_data[104] ,
         \DataPath/RF/bus_complete_win_data[105] ,
         \DataPath/RF/bus_complete_win_data[106] ,
         \DataPath/RF/bus_complete_win_data[107] ,
         \DataPath/RF/bus_complete_win_data[108] ,
         \DataPath/RF/bus_complete_win_data[109] ,
         \DataPath/RF/bus_complete_win_data[110] ,
         \DataPath/RF/bus_complete_win_data[111] ,
         \DataPath/RF/bus_complete_win_data[112] ,
         \DataPath/RF/bus_complete_win_data[113] ,
         \DataPath/RF/bus_complete_win_data[114] ,
         \DataPath/RF/bus_complete_win_data[115] ,
         \DataPath/RF/bus_complete_win_data[116] ,
         \DataPath/RF/bus_complete_win_data[117] ,
         \DataPath/RF/bus_complete_win_data[118] ,
         \DataPath/RF/bus_complete_win_data[119] ,
         \DataPath/RF/bus_complete_win_data[120] ,
         \DataPath/RF/bus_complete_win_data[121] ,
         \DataPath/RF/bus_complete_win_data[122] ,
         \DataPath/RF/bus_complete_win_data[123] ,
         \DataPath/RF/bus_complete_win_data[124] ,
         \DataPath/RF/bus_complete_win_data[125] ,
         \DataPath/RF/bus_complete_win_data[126] ,
         \DataPath/RF/bus_complete_win_data[127] ,
         \DataPath/RF/bus_complete_win_data[128] ,
         \DataPath/RF/bus_complete_win_data[129] ,
         \DataPath/RF/bus_complete_win_data[130] ,
         \DataPath/RF/bus_complete_win_data[131] ,
         \DataPath/RF/bus_complete_win_data[132] ,
         \DataPath/RF/bus_complete_win_data[133] ,
         \DataPath/RF/bus_complete_win_data[134] ,
         \DataPath/RF/bus_complete_win_data[135] ,
         \DataPath/RF/bus_complete_win_data[136] ,
         \DataPath/RF/bus_complete_win_data[137] ,
         \DataPath/RF/bus_complete_win_data[138] ,
         \DataPath/RF/bus_complete_win_data[139] ,
         \DataPath/RF/bus_complete_win_data[140] ,
         \DataPath/RF/bus_complete_win_data[141] ,
         \DataPath/RF/bus_complete_win_data[142] ,
         \DataPath/RF/bus_complete_win_data[143] ,
         \DataPath/RF/bus_complete_win_data[144] ,
         \DataPath/RF/bus_complete_win_data[145] ,
         \DataPath/RF/bus_complete_win_data[146] ,
         \DataPath/RF/bus_complete_win_data[147] ,
         \DataPath/RF/bus_complete_win_data[148] ,
         \DataPath/RF/bus_complete_win_data[149] ,
         \DataPath/RF/bus_complete_win_data[150] ,
         \DataPath/RF/bus_complete_win_data[151] ,
         \DataPath/RF/bus_complete_win_data[152] ,
         \DataPath/RF/bus_complete_win_data[153] ,
         \DataPath/RF/bus_complete_win_data[154] ,
         \DataPath/RF/bus_complete_win_data[155] ,
         \DataPath/RF/bus_complete_win_data[156] ,
         \DataPath/RF/bus_complete_win_data[157] ,
         \DataPath/RF/bus_complete_win_data[158] ,
         \DataPath/RF/bus_complete_win_data[159] ,
         \DataPath/RF/bus_complete_win_data[160] ,
         \DataPath/RF/bus_complete_win_data[161] ,
         \DataPath/RF/bus_complete_win_data[162] ,
         \DataPath/RF/bus_complete_win_data[163] ,
         \DataPath/RF/bus_complete_win_data[164] ,
         \DataPath/RF/bus_complete_win_data[165] ,
         \DataPath/RF/bus_complete_win_data[166] ,
         \DataPath/RF/bus_complete_win_data[167] ,
         \DataPath/RF/bus_complete_win_data[168] ,
         \DataPath/RF/bus_complete_win_data[169] ,
         \DataPath/RF/bus_complete_win_data[170] ,
         \DataPath/RF/bus_complete_win_data[171] ,
         \DataPath/RF/bus_complete_win_data[172] ,
         \DataPath/RF/bus_complete_win_data[173] ,
         \DataPath/RF/bus_complete_win_data[174] ,
         \DataPath/RF/bus_complete_win_data[175] ,
         \DataPath/RF/bus_complete_win_data[176] ,
         \DataPath/RF/bus_complete_win_data[177] ,
         \DataPath/RF/bus_complete_win_data[178] ,
         \DataPath/RF/bus_complete_win_data[179] ,
         \DataPath/RF/bus_complete_win_data[180] ,
         \DataPath/RF/bus_complete_win_data[181] ,
         \DataPath/RF/bus_complete_win_data[182] ,
         \DataPath/RF/bus_complete_win_data[183] ,
         \DataPath/RF/bus_complete_win_data[184] ,
         \DataPath/RF/bus_complete_win_data[185] ,
         \DataPath/RF/bus_complete_win_data[186] ,
         \DataPath/RF/bus_complete_win_data[187] ,
         \DataPath/RF/bus_complete_win_data[188] ,
         \DataPath/RF/bus_complete_win_data[189] ,
         \DataPath/RF/bus_complete_win_data[190] ,
         \DataPath/RF/bus_complete_win_data[191] ,
         \DataPath/RF/bus_complete_win_data[192] ,
         \DataPath/RF/bus_complete_win_data[193] ,
         \DataPath/RF/bus_complete_win_data[194] ,
         \DataPath/RF/bus_complete_win_data[195] ,
         \DataPath/RF/bus_complete_win_data[196] ,
         \DataPath/RF/bus_complete_win_data[197] ,
         \DataPath/RF/bus_complete_win_data[198] ,
         \DataPath/RF/bus_complete_win_data[199] ,
         \DataPath/RF/bus_complete_win_data[200] ,
         \DataPath/RF/bus_complete_win_data[201] ,
         \DataPath/RF/bus_complete_win_data[202] ,
         \DataPath/RF/bus_complete_win_data[203] ,
         \DataPath/RF/bus_complete_win_data[204] ,
         \DataPath/RF/bus_complete_win_data[205] ,
         \DataPath/RF/bus_complete_win_data[206] ,
         \DataPath/RF/bus_complete_win_data[207] ,
         \DataPath/RF/bus_complete_win_data[208] ,
         \DataPath/RF/bus_complete_win_data[209] ,
         \DataPath/RF/bus_complete_win_data[210] ,
         \DataPath/RF/bus_complete_win_data[211] ,
         \DataPath/RF/bus_complete_win_data[212] ,
         \DataPath/RF/bus_complete_win_data[213] ,
         \DataPath/RF/bus_complete_win_data[214] ,
         \DataPath/RF/bus_complete_win_data[215] ,
         \DataPath/RF/bus_complete_win_data[216] ,
         \DataPath/RF/bus_complete_win_data[217] ,
         \DataPath/RF/bus_complete_win_data[218] ,
         \DataPath/RF/bus_complete_win_data[219] ,
         \DataPath/RF/bus_complete_win_data[220] ,
         \DataPath/RF/bus_complete_win_data[221] ,
         \DataPath/RF/bus_complete_win_data[222] ,
         \DataPath/RF/bus_complete_win_data[223] ,
         \DataPath/RF/bus_complete_win_data[224] ,
         \DataPath/RF/bus_complete_win_data[225] ,
         \DataPath/RF/bus_complete_win_data[226] ,
         \DataPath/RF/bus_complete_win_data[227] ,
         \DataPath/RF/bus_complete_win_data[228] ,
         \DataPath/RF/bus_complete_win_data[229] ,
         \DataPath/RF/bus_complete_win_data[230] ,
         \DataPath/RF/bus_complete_win_data[231] ,
         \DataPath/RF/bus_complete_win_data[232] ,
         \DataPath/RF/bus_complete_win_data[233] ,
         \DataPath/RF/bus_complete_win_data[234] ,
         \DataPath/RF/bus_complete_win_data[235] ,
         \DataPath/RF/bus_complete_win_data[236] ,
         \DataPath/RF/bus_complete_win_data[237] ,
         \DataPath/RF/bus_complete_win_data[238] ,
         \DataPath/RF/bus_complete_win_data[239] ,
         \DataPath/RF/bus_complete_win_data[240] ,
         \DataPath/RF/bus_complete_win_data[241] ,
         \DataPath/RF/bus_complete_win_data[242] ,
         \DataPath/RF/bus_complete_win_data[243] ,
         \DataPath/RF/bus_complete_win_data[244] ,
         \DataPath/RF/bus_complete_win_data[245] ,
         \DataPath/RF/bus_complete_win_data[246] ,
         \DataPath/RF/bus_complete_win_data[247] ,
         \DataPath/RF/bus_complete_win_data[248] ,
         \DataPath/RF/bus_complete_win_data[249] ,
         \DataPath/RF/bus_complete_win_data[250] ,
         \DataPath/RF/bus_complete_win_data[251] ,
         \DataPath/RF/bus_complete_win_data[252] ,
         \DataPath/RF/bus_complete_win_data[253] ,
         \DataPath/RF/bus_complete_win_data[254] ,
         \DataPath/RF/bus_complete_win_data[255] ,
         \DataPath/RF/bus_selected_win_data[0] ,
         \DataPath/RF/bus_selected_win_data[1] ,
         \DataPath/RF/bus_selected_win_data[2] ,
         \DataPath/RF/bus_selected_win_data[3] ,
         \DataPath/RF/bus_selected_win_data[4] ,
         \DataPath/RF/bus_selected_win_data[5] ,
         \DataPath/RF/bus_selected_win_data[6] ,
         \DataPath/RF/bus_selected_win_data[7] ,
         \DataPath/RF/bus_selected_win_data[8] ,
         \DataPath/RF/bus_selected_win_data[9] ,
         \DataPath/RF/bus_selected_win_data[10] ,
         \DataPath/RF/bus_selected_win_data[11] ,
         \DataPath/RF/bus_selected_win_data[12] ,
         \DataPath/RF/bus_selected_win_data[13] ,
         \DataPath/RF/bus_selected_win_data[14] ,
         \DataPath/RF/bus_selected_win_data[15] ,
         \DataPath/RF/bus_selected_win_data[16] ,
         \DataPath/RF/bus_selected_win_data[17] ,
         \DataPath/RF/bus_selected_win_data[18] ,
         \DataPath/RF/bus_selected_win_data[19] ,
         \DataPath/RF/bus_selected_win_data[20] ,
         \DataPath/RF/bus_selected_win_data[21] ,
         \DataPath/RF/bus_selected_win_data[22] ,
         \DataPath/RF/bus_selected_win_data[23] ,
         \DataPath/RF/bus_selected_win_data[24] ,
         \DataPath/RF/bus_selected_win_data[25] ,
         \DataPath/RF/bus_selected_win_data[26] ,
         \DataPath/RF/bus_selected_win_data[27] ,
         \DataPath/RF/bus_selected_win_data[28] ,
         \DataPath/RF/bus_selected_win_data[29] ,
         \DataPath/RF/bus_selected_win_data[30] ,
         \DataPath/RF/bus_selected_win_data[31] ,
         \DataPath/RF/bus_selected_win_data[32] ,
         \DataPath/RF/bus_selected_win_data[33] ,
         \DataPath/RF/bus_selected_win_data[34] ,
         \DataPath/RF/bus_selected_win_data[35] ,
         \DataPath/RF/bus_selected_win_data[36] ,
         \DataPath/RF/bus_selected_win_data[37] ,
         \DataPath/RF/bus_selected_win_data[38] ,
         \DataPath/RF/bus_selected_win_data[39] ,
         \DataPath/RF/bus_selected_win_data[40] ,
         \DataPath/RF/bus_selected_win_data[41] ,
         \DataPath/RF/bus_selected_win_data[42] ,
         \DataPath/RF/bus_selected_win_data[43] ,
         \DataPath/RF/bus_selected_win_data[44] ,
         \DataPath/RF/bus_selected_win_data[45] ,
         \DataPath/RF/bus_selected_win_data[46] ,
         \DataPath/RF/bus_selected_win_data[47] ,
         \DataPath/RF/bus_selected_win_data[48] ,
         \DataPath/RF/bus_selected_win_data[49] ,
         \DataPath/RF/bus_selected_win_data[50] ,
         \DataPath/RF/bus_selected_win_data[51] ,
         \DataPath/RF/bus_selected_win_data[52] ,
         \DataPath/RF/bus_selected_win_data[53] ,
         \DataPath/RF/bus_selected_win_data[54] ,
         \DataPath/RF/bus_selected_win_data[55] ,
         \DataPath/RF/bus_selected_win_data[56] ,
         \DataPath/RF/bus_selected_win_data[57] ,
         \DataPath/RF/bus_selected_win_data[58] ,
         \DataPath/RF/bus_selected_win_data[59] ,
         \DataPath/RF/bus_selected_win_data[60] ,
         \DataPath/RF/bus_selected_win_data[61] ,
         \DataPath/RF/bus_selected_win_data[62] ,
         \DataPath/RF/bus_selected_win_data[63] ,
         \DataPath/RF/bus_selected_win_data[64] ,
         \DataPath/RF/bus_selected_win_data[65] ,
         \DataPath/RF/bus_selected_win_data[66] ,
         \DataPath/RF/bus_selected_win_data[67] ,
         \DataPath/RF/bus_selected_win_data[68] ,
         \DataPath/RF/bus_selected_win_data[69] ,
         \DataPath/RF/bus_selected_win_data[70] ,
         \DataPath/RF/bus_selected_win_data[71] ,
         \DataPath/RF/bus_selected_win_data[72] ,
         \DataPath/RF/bus_selected_win_data[73] ,
         \DataPath/RF/bus_selected_win_data[74] ,
         \DataPath/RF/bus_selected_win_data[75] ,
         \DataPath/RF/bus_selected_win_data[76] ,
         \DataPath/RF/bus_selected_win_data[77] ,
         \DataPath/RF/bus_selected_win_data[78] ,
         \DataPath/RF/bus_selected_win_data[79] ,
         \DataPath/RF/bus_selected_win_data[80] ,
         \DataPath/RF/bus_selected_win_data[81] ,
         \DataPath/RF/bus_selected_win_data[82] ,
         \DataPath/RF/bus_selected_win_data[83] ,
         \DataPath/RF/bus_selected_win_data[84] ,
         \DataPath/RF/bus_selected_win_data[85] ,
         \DataPath/RF/bus_selected_win_data[86] ,
         \DataPath/RF/bus_selected_win_data[87] ,
         \DataPath/RF/bus_selected_win_data[88] ,
         \DataPath/RF/bus_selected_win_data[89] ,
         \DataPath/RF/bus_selected_win_data[90] ,
         \DataPath/RF/bus_selected_win_data[91] ,
         \DataPath/RF/bus_selected_win_data[92] ,
         \DataPath/RF/bus_selected_win_data[93] ,
         \DataPath/RF/bus_selected_win_data[94] ,
         \DataPath/RF/bus_selected_win_data[95] ,
         \DataPath/RF/bus_selected_win_data[96] ,
         \DataPath/RF/bus_selected_win_data[97] ,
         \DataPath/RF/bus_selected_win_data[98] ,
         \DataPath/RF/bus_selected_win_data[99] ,
         \DataPath/RF/bus_selected_win_data[100] ,
         \DataPath/RF/bus_selected_win_data[101] ,
         \DataPath/RF/bus_selected_win_data[102] ,
         \DataPath/RF/bus_selected_win_data[103] ,
         \DataPath/RF/bus_selected_win_data[104] ,
         \DataPath/RF/bus_selected_win_data[105] ,
         \DataPath/RF/bus_selected_win_data[106] ,
         \DataPath/RF/bus_selected_win_data[107] ,
         \DataPath/RF/bus_selected_win_data[108] ,
         \DataPath/RF/bus_selected_win_data[109] ,
         \DataPath/RF/bus_selected_win_data[110] ,
         \DataPath/RF/bus_selected_win_data[111] ,
         \DataPath/RF/bus_selected_win_data[112] ,
         \DataPath/RF/bus_selected_win_data[113] ,
         \DataPath/RF/bus_selected_win_data[114] ,
         \DataPath/RF/bus_selected_win_data[115] ,
         \DataPath/RF/bus_selected_win_data[116] ,
         \DataPath/RF/bus_selected_win_data[117] ,
         \DataPath/RF/bus_selected_win_data[118] ,
         \DataPath/RF/bus_selected_win_data[119] ,
         \DataPath/RF/bus_selected_win_data[120] ,
         \DataPath/RF/bus_selected_win_data[121] ,
         \DataPath/RF/bus_selected_win_data[122] ,
         \DataPath/RF/bus_selected_win_data[123] ,
         \DataPath/RF/bus_selected_win_data[124] ,
         \DataPath/RF/bus_selected_win_data[125] ,
         \DataPath/RF/bus_selected_win_data[126] ,
         \DataPath/RF/bus_selected_win_data[127] ,
         \DataPath/RF/bus_selected_win_data[128] ,
         \DataPath/RF/bus_selected_win_data[129] ,
         \DataPath/RF/bus_selected_win_data[130] ,
         \DataPath/RF/bus_selected_win_data[131] ,
         \DataPath/RF/bus_selected_win_data[132] ,
         \DataPath/RF/bus_selected_win_data[133] ,
         \DataPath/RF/bus_selected_win_data[134] ,
         \DataPath/RF/bus_selected_win_data[135] ,
         \DataPath/RF/bus_selected_win_data[136] ,
         \DataPath/RF/bus_selected_win_data[137] ,
         \DataPath/RF/bus_selected_win_data[138] ,
         \DataPath/RF/bus_selected_win_data[139] ,
         \DataPath/RF/bus_selected_win_data[140] ,
         \DataPath/RF/bus_selected_win_data[141] ,
         \DataPath/RF/bus_selected_win_data[142] ,
         \DataPath/RF/bus_selected_win_data[143] ,
         \DataPath/RF/bus_selected_win_data[144] ,
         \DataPath/RF/bus_selected_win_data[145] ,
         \DataPath/RF/bus_selected_win_data[146] ,
         \DataPath/RF/bus_selected_win_data[147] ,
         \DataPath/RF/bus_selected_win_data[148] ,
         \DataPath/RF/bus_selected_win_data[149] ,
         \DataPath/RF/bus_selected_win_data[150] ,
         \DataPath/RF/bus_selected_win_data[151] ,
         \DataPath/RF/bus_selected_win_data[152] ,
         \DataPath/RF/bus_selected_win_data[153] ,
         \DataPath/RF/bus_selected_win_data[154] ,
         \DataPath/RF/bus_selected_win_data[155] ,
         \DataPath/RF/bus_selected_win_data[156] ,
         \DataPath/RF/bus_selected_win_data[157] ,
         \DataPath/RF/bus_selected_win_data[158] ,
         \DataPath/RF/bus_selected_win_data[159] ,
         \DataPath/RF/bus_selected_win_data[160] ,
         \DataPath/RF/bus_selected_win_data[161] ,
         \DataPath/RF/bus_selected_win_data[162] ,
         \DataPath/RF/bus_selected_win_data[163] ,
         \DataPath/RF/bus_selected_win_data[164] ,
         \DataPath/RF/bus_selected_win_data[165] ,
         \DataPath/RF/bus_selected_win_data[166] ,
         \DataPath/RF/bus_selected_win_data[167] ,
         \DataPath/RF/bus_selected_win_data[168] ,
         \DataPath/RF/bus_selected_win_data[169] ,
         \DataPath/RF/bus_selected_win_data[170] ,
         \DataPath/RF/bus_selected_win_data[171] ,
         \DataPath/RF/bus_selected_win_data[172] ,
         \DataPath/RF/bus_selected_win_data[173] ,
         \DataPath/RF/bus_selected_win_data[174] ,
         \DataPath/RF/bus_selected_win_data[175] ,
         \DataPath/RF/bus_selected_win_data[176] ,
         \DataPath/RF/bus_selected_win_data[177] ,
         \DataPath/RF/bus_selected_win_data[178] ,
         \DataPath/RF/bus_selected_win_data[179] ,
         \DataPath/RF/bus_selected_win_data[180] ,
         \DataPath/RF/bus_selected_win_data[181] ,
         \DataPath/RF/bus_selected_win_data[182] ,
         \DataPath/RF/bus_selected_win_data[183] ,
         \DataPath/RF/bus_selected_win_data[184] ,
         \DataPath/RF/bus_selected_win_data[185] ,
         \DataPath/RF/bus_selected_win_data[186] ,
         \DataPath/RF/bus_selected_win_data[187] ,
         \DataPath/RF/bus_selected_win_data[188] ,
         \DataPath/RF/bus_selected_win_data[189] ,
         \DataPath/RF/bus_selected_win_data[190] ,
         \DataPath/RF/bus_selected_win_data[191] ,
         \DataPath/RF/bus_selected_win_data[192] ,
         \DataPath/RF/bus_selected_win_data[193] ,
         \DataPath/RF/bus_selected_win_data[194] ,
         \DataPath/RF/bus_selected_win_data[195] ,
         \DataPath/RF/bus_selected_win_data[196] ,
         \DataPath/RF/bus_selected_win_data[197] ,
         \DataPath/RF/bus_selected_win_data[198] ,
         \DataPath/RF/bus_selected_win_data[199] ,
         \DataPath/RF/bus_selected_win_data[200] ,
         \DataPath/RF/bus_selected_win_data[201] ,
         \DataPath/RF/bus_selected_win_data[202] ,
         \DataPath/RF/bus_selected_win_data[203] ,
         \DataPath/RF/bus_selected_win_data[204] ,
         \DataPath/RF/bus_selected_win_data[205] ,
         \DataPath/RF/bus_selected_win_data[206] ,
         \DataPath/RF/bus_selected_win_data[207] ,
         \DataPath/RF/bus_selected_win_data[208] ,
         \DataPath/RF/bus_selected_win_data[209] ,
         \DataPath/RF/bus_selected_win_data[210] ,
         \DataPath/RF/bus_selected_win_data[211] ,
         \DataPath/RF/bus_selected_win_data[212] ,
         \DataPath/RF/bus_selected_win_data[213] ,
         \DataPath/RF/bus_selected_win_data[214] ,
         \DataPath/RF/bus_selected_win_data[215] ,
         \DataPath/RF/bus_selected_win_data[216] ,
         \DataPath/RF/bus_selected_win_data[217] ,
         \DataPath/RF/bus_selected_win_data[218] ,
         \DataPath/RF/bus_selected_win_data[219] ,
         \DataPath/RF/bus_selected_win_data[220] ,
         \DataPath/RF/bus_selected_win_data[221] ,
         \DataPath/RF/bus_selected_win_data[222] ,
         \DataPath/RF/bus_selected_win_data[223] ,
         \DataPath/RF/bus_selected_win_data[224] ,
         \DataPath/RF/bus_selected_win_data[225] ,
         \DataPath/RF/bus_selected_win_data[226] ,
         \DataPath/RF/bus_selected_win_data[227] ,
         \DataPath/RF/bus_selected_win_data[228] ,
         \DataPath/RF/bus_selected_win_data[229] ,
         \DataPath/RF/bus_selected_win_data[230] ,
         \DataPath/RF/bus_selected_win_data[231] ,
         \DataPath/RF/bus_selected_win_data[232] ,
         \DataPath/RF/bus_selected_win_data[233] ,
         \DataPath/RF/bus_selected_win_data[234] ,
         \DataPath/RF/bus_selected_win_data[235] ,
         \DataPath/RF/bus_selected_win_data[236] ,
         \DataPath/RF/bus_selected_win_data[237] ,
         \DataPath/RF/bus_selected_win_data[238] ,
         \DataPath/RF/bus_selected_win_data[239] ,
         \DataPath/RF/bus_selected_win_data[240] ,
         \DataPath/RF/bus_selected_win_data[241] ,
         \DataPath/RF/bus_selected_win_data[242] ,
         \DataPath/RF/bus_selected_win_data[243] ,
         \DataPath/RF/bus_selected_win_data[244] ,
         \DataPath/RF/bus_selected_win_data[245] ,
         \DataPath/RF/bus_selected_win_data[246] ,
         \DataPath/RF/bus_selected_win_data[247] ,
         \DataPath/RF/bus_selected_win_data[248] ,
         \DataPath/RF/bus_selected_win_data[249] ,
         \DataPath/RF/bus_selected_win_data[250] ,
         \DataPath/RF/bus_selected_win_data[251] ,
         \DataPath/RF/bus_selected_win_data[252] ,
         \DataPath/RF/bus_selected_win_data[253] ,
         \DataPath/RF/bus_selected_win_data[254] ,
         \DataPath/RF/bus_selected_win_data[255] ,
         \DataPath/RF/bus_selected_win_data[256] ,
         \DataPath/RF/bus_selected_win_data[257] ,
         \DataPath/RF/bus_selected_win_data[258] ,
         \DataPath/RF/bus_selected_win_data[259] ,
         \DataPath/RF/bus_selected_win_data[260] ,
         \DataPath/RF/bus_selected_win_data[261] ,
         \DataPath/RF/bus_selected_win_data[262] ,
         \DataPath/RF/bus_selected_win_data[263] ,
         \DataPath/RF/bus_selected_win_data[264] ,
         \DataPath/RF/bus_selected_win_data[265] ,
         \DataPath/RF/bus_selected_win_data[266] ,
         \DataPath/RF/bus_selected_win_data[267] ,
         \DataPath/RF/bus_selected_win_data[268] ,
         \DataPath/RF/bus_selected_win_data[269] ,
         \DataPath/RF/bus_selected_win_data[270] ,
         \DataPath/RF/bus_selected_win_data[271] ,
         \DataPath/RF/bus_selected_win_data[272] ,
         \DataPath/RF/bus_selected_win_data[273] ,
         \DataPath/RF/bus_selected_win_data[274] ,
         \DataPath/RF/bus_selected_win_data[275] ,
         \DataPath/RF/bus_selected_win_data[276] ,
         \DataPath/RF/bus_selected_win_data[277] ,
         \DataPath/RF/bus_selected_win_data[278] ,
         \DataPath/RF/bus_selected_win_data[279] ,
         \DataPath/RF/bus_selected_win_data[280] ,
         \DataPath/RF/bus_selected_win_data[281] ,
         \DataPath/RF/bus_selected_win_data[282] ,
         \DataPath/RF/bus_selected_win_data[283] ,
         \DataPath/RF/bus_selected_win_data[284] ,
         \DataPath/RF/bus_selected_win_data[285] ,
         \DataPath/RF/bus_selected_win_data[286] ,
         \DataPath/RF/bus_selected_win_data[287] ,
         \DataPath/RF/bus_selected_win_data[288] ,
         \DataPath/RF/bus_selected_win_data[289] ,
         \DataPath/RF/bus_selected_win_data[290] ,
         \DataPath/RF/bus_selected_win_data[291] ,
         \DataPath/RF/bus_selected_win_data[292] ,
         \DataPath/RF/bus_selected_win_data[293] ,
         \DataPath/RF/bus_selected_win_data[294] ,
         \DataPath/RF/bus_selected_win_data[295] ,
         \DataPath/RF/bus_selected_win_data[296] ,
         \DataPath/RF/bus_selected_win_data[297] ,
         \DataPath/RF/bus_selected_win_data[298] ,
         \DataPath/RF/bus_selected_win_data[299] ,
         \DataPath/RF/bus_selected_win_data[300] ,
         \DataPath/RF/bus_selected_win_data[301] ,
         \DataPath/RF/bus_selected_win_data[302] ,
         \DataPath/RF/bus_selected_win_data[303] ,
         \DataPath/RF/bus_selected_win_data[304] ,
         \DataPath/RF/bus_selected_win_data[305] ,
         \DataPath/RF/bus_selected_win_data[306] ,
         \DataPath/RF/bus_selected_win_data[307] ,
         \DataPath/RF/bus_selected_win_data[308] ,
         \DataPath/RF/bus_selected_win_data[309] ,
         \DataPath/RF/bus_selected_win_data[310] ,
         \DataPath/RF/bus_selected_win_data[311] ,
         \DataPath/RF/bus_selected_win_data[312] ,
         \DataPath/RF/bus_selected_win_data[313] ,
         \DataPath/RF/bus_selected_win_data[314] ,
         \DataPath/RF/bus_selected_win_data[315] ,
         \DataPath/RF/bus_selected_win_data[316] ,
         \DataPath/RF/bus_selected_win_data[317] ,
         \DataPath/RF/bus_selected_win_data[318] ,
         \DataPath/RF/bus_selected_win_data[319] ,
         \DataPath/RF/bus_selected_win_data[320] ,
         \DataPath/RF/bus_selected_win_data[321] ,
         \DataPath/RF/bus_selected_win_data[322] ,
         \DataPath/RF/bus_selected_win_data[323] ,
         \DataPath/RF/bus_selected_win_data[324] ,
         \DataPath/RF/bus_selected_win_data[325] ,
         \DataPath/RF/bus_selected_win_data[326] ,
         \DataPath/RF/bus_selected_win_data[327] ,
         \DataPath/RF/bus_selected_win_data[328] ,
         \DataPath/RF/bus_selected_win_data[329] ,
         \DataPath/RF/bus_selected_win_data[330] ,
         \DataPath/RF/bus_selected_win_data[331] ,
         \DataPath/RF/bus_selected_win_data[332] ,
         \DataPath/RF/bus_selected_win_data[333] ,
         \DataPath/RF/bus_selected_win_data[334] ,
         \DataPath/RF/bus_selected_win_data[335] ,
         \DataPath/RF/bus_selected_win_data[336] ,
         \DataPath/RF/bus_selected_win_data[337] ,
         \DataPath/RF/bus_selected_win_data[338] ,
         \DataPath/RF/bus_selected_win_data[339] ,
         \DataPath/RF/bus_selected_win_data[340] ,
         \DataPath/RF/bus_selected_win_data[341] ,
         \DataPath/RF/bus_selected_win_data[342] ,
         \DataPath/RF/bus_selected_win_data[343] ,
         \DataPath/RF/bus_selected_win_data[344] ,
         \DataPath/RF/bus_selected_win_data[345] ,
         \DataPath/RF/bus_selected_win_data[346] ,
         \DataPath/RF/bus_selected_win_data[347] ,
         \DataPath/RF/bus_selected_win_data[348] ,
         \DataPath/RF/bus_selected_win_data[349] ,
         \DataPath/RF/bus_selected_win_data[350] ,
         \DataPath/RF/bus_selected_win_data[351] ,
         \DataPath/RF/bus_selected_win_data[352] ,
         \DataPath/RF/bus_selected_win_data[353] ,
         \DataPath/RF/bus_selected_win_data[354] ,
         \DataPath/RF/bus_selected_win_data[355] ,
         \DataPath/RF/bus_selected_win_data[356] ,
         \DataPath/RF/bus_selected_win_data[357] ,
         \DataPath/RF/bus_selected_win_data[358] ,
         \DataPath/RF/bus_selected_win_data[359] ,
         \DataPath/RF/bus_selected_win_data[360] ,
         \DataPath/RF/bus_selected_win_data[361] ,
         \DataPath/RF/bus_selected_win_data[362] ,
         \DataPath/RF/bus_selected_win_data[363] ,
         \DataPath/RF/bus_selected_win_data[364] ,
         \DataPath/RF/bus_selected_win_data[365] ,
         \DataPath/RF/bus_selected_win_data[366] ,
         \DataPath/RF/bus_selected_win_data[367] ,
         \DataPath/RF/bus_selected_win_data[368] ,
         \DataPath/RF/bus_selected_win_data[369] ,
         \DataPath/RF/bus_selected_win_data[370] ,
         \DataPath/RF/bus_selected_win_data[371] ,
         \DataPath/RF/bus_selected_win_data[372] ,
         \DataPath/RF/bus_selected_win_data[373] ,
         \DataPath/RF/bus_selected_win_data[374] ,
         \DataPath/RF/bus_selected_win_data[375] ,
         \DataPath/RF/bus_selected_win_data[376] ,
         \DataPath/RF/bus_selected_win_data[377] ,
         \DataPath/RF/bus_selected_win_data[378] ,
         \DataPath/RF/bus_selected_win_data[379] ,
         \DataPath/RF/bus_selected_win_data[380] ,
         \DataPath/RF/bus_selected_win_data[381] ,
         \DataPath/RF/bus_selected_win_data[382] ,
         \DataPath/RF/bus_selected_win_data[383] ,
         \DataPath/RF/bus_selected_win_data[384] ,
         \DataPath/RF/bus_selected_win_data[385] ,
         \DataPath/RF/bus_selected_win_data[386] ,
         \DataPath/RF/bus_selected_win_data[387] ,
         \DataPath/RF/bus_selected_win_data[388] ,
         \DataPath/RF/bus_selected_win_data[389] ,
         \DataPath/RF/bus_selected_win_data[390] ,
         \DataPath/RF/bus_selected_win_data[391] ,
         \DataPath/RF/bus_selected_win_data[392] ,
         \DataPath/RF/bus_selected_win_data[393] ,
         \DataPath/RF/bus_selected_win_data[394] ,
         \DataPath/RF/bus_selected_win_data[395] ,
         \DataPath/RF/bus_selected_win_data[396] ,
         \DataPath/RF/bus_selected_win_data[397] ,
         \DataPath/RF/bus_selected_win_data[398] ,
         \DataPath/RF/bus_selected_win_data[399] ,
         \DataPath/RF/bus_selected_win_data[400] ,
         \DataPath/RF/bus_selected_win_data[401] ,
         \DataPath/RF/bus_selected_win_data[402] ,
         \DataPath/RF/bus_selected_win_data[403] ,
         \DataPath/RF/bus_selected_win_data[404] ,
         \DataPath/RF/bus_selected_win_data[405] ,
         \DataPath/RF/bus_selected_win_data[406] ,
         \DataPath/RF/bus_selected_win_data[407] ,
         \DataPath/RF/bus_selected_win_data[408] ,
         \DataPath/RF/bus_selected_win_data[409] ,
         \DataPath/RF/bus_selected_win_data[410] ,
         \DataPath/RF/bus_selected_win_data[411] ,
         \DataPath/RF/bus_selected_win_data[412] ,
         \DataPath/RF/bus_selected_win_data[413] ,
         \DataPath/RF/bus_selected_win_data[414] ,
         \DataPath/RF/bus_selected_win_data[415] ,
         \DataPath/RF/bus_selected_win_data[416] ,
         \DataPath/RF/bus_selected_win_data[417] ,
         \DataPath/RF/bus_selected_win_data[418] ,
         \DataPath/RF/bus_selected_win_data[419] ,
         \DataPath/RF/bus_selected_win_data[420] ,
         \DataPath/RF/bus_selected_win_data[421] ,
         \DataPath/RF/bus_selected_win_data[422] ,
         \DataPath/RF/bus_selected_win_data[423] ,
         \DataPath/RF/bus_selected_win_data[424] ,
         \DataPath/RF/bus_selected_win_data[425] ,
         \DataPath/RF/bus_selected_win_data[426] ,
         \DataPath/RF/bus_selected_win_data[427] ,
         \DataPath/RF/bus_selected_win_data[428] ,
         \DataPath/RF/bus_selected_win_data[429] ,
         \DataPath/RF/bus_selected_win_data[430] ,
         \DataPath/RF/bus_selected_win_data[431] ,
         \DataPath/RF/bus_selected_win_data[432] ,
         \DataPath/RF/bus_selected_win_data[433] ,
         \DataPath/RF/bus_selected_win_data[434] ,
         \DataPath/RF/bus_selected_win_data[435] ,
         \DataPath/RF/bus_selected_win_data[436] ,
         \DataPath/RF/bus_selected_win_data[437] ,
         \DataPath/RF/bus_selected_win_data[438] ,
         \DataPath/RF/bus_selected_win_data[439] ,
         \DataPath/RF/bus_selected_win_data[440] ,
         \DataPath/RF/bus_selected_win_data[441] ,
         \DataPath/RF/bus_selected_win_data[442] ,
         \DataPath/RF/bus_selected_win_data[443] ,
         \DataPath/RF/bus_selected_win_data[444] ,
         \DataPath/RF/bus_selected_win_data[445] ,
         \DataPath/RF/bus_selected_win_data[446] ,
         \DataPath/RF/bus_selected_win_data[447] ,
         \DataPath/RF/bus_selected_win_data[448] ,
         \DataPath/RF/bus_selected_win_data[449] ,
         \DataPath/RF/bus_selected_win_data[450] ,
         \DataPath/RF/bus_selected_win_data[451] ,
         \DataPath/RF/bus_selected_win_data[452] ,
         \DataPath/RF/bus_selected_win_data[453] ,
         \DataPath/RF/bus_selected_win_data[454] ,
         \DataPath/RF/bus_selected_win_data[455] ,
         \DataPath/RF/bus_selected_win_data[456] ,
         \DataPath/RF/bus_selected_win_data[457] ,
         \DataPath/RF/bus_selected_win_data[458] ,
         \DataPath/RF/bus_selected_win_data[459] ,
         \DataPath/RF/bus_selected_win_data[460] ,
         \DataPath/RF/bus_selected_win_data[461] ,
         \DataPath/RF/bus_selected_win_data[462] ,
         \DataPath/RF/bus_selected_win_data[463] ,
         \DataPath/RF/bus_selected_win_data[464] ,
         \DataPath/RF/bus_selected_win_data[465] ,
         \DataPath/RF/bus_selected_win_data[466] ,
         \DataPath/RF/bus_selected_win_data[467] ,
         \DataPath/RF/bus_selected_win_data[468] ,
         \DataPath/RF/bus_selected_win_data[469] ,
         \DataPath/RF/bus_selected_win_data[470] ,
         \DataPath/RF/bus_selected_win_data[471] ,
         \DataPath/RF/bus_selected_win_data[472] ,
         \DataPath/RF/bus_selected_win_data[473] ,
         \DataPath/RF/bus_selected_win_data[474] ,
         \DataPath/RF/bus_selected_win_data[475] ,
         \DataPath/RF/bus_selected_win_data[476] ,
         \DataPath/RF/bus_selected_win_data[477] ,
         \DataPath/RF/bus_selected_win_data[478] ,
         \DataPath/RF/bus_selected_win_data[479] ,
         \DataPath/RF/bus_selected_win_data[480] ,
         \DataPath/RF/bus_selected_win_data[481] ,
         \DataPath/RF/bus_selected_win_data[482] ,
         \DataPath/RF/bus_selected_win_data[483] ,
         \DataPath/RF/bus_selected_win_data[484] ,
         \DataPath/RF/bus_selected_win_data[485] ,
         \DataPath/RF/bus_selected_win_data[486] ,
         \DataPath/RF/bus_selected_win_data[487] ,
         \DataPath/RF/bus_selected_win_data[488] ,
         \DataPath/RF/bus_selected_win_data[489] ,
         \DataPath/RF/bus_selected_win_data[490] ,
         \DataPath/RF/bus_selected_win_data[491] ,
         \DataPath/RF/bus_selected_win_data[492] ,
         \DataPath/RF/bus_selected_win_data[493] ,
         \DataPath/RF/bus_selected_win_data[494] ,
         \DataPath/RF/bus_selected_win_data[495] ,
         \DataPath/RF/bus_selected_win_data[496] ,
         \DataPath/RF/bus_selected_win_data[497] ,
         \DataPath/RF/bus_selected_win_data[498] ,
         \DataPath/RF/bus_selected_win_data[499] ,
         \DataPath/RF/bus_selected_win_data[500] ,
         \DataPath/RF/bus_selected_win_data[501] ,
         \DataPath/RF/bus_selected_win_data[502] ,
         \DataPath/RF/bus_selected_win_data[503] ,
         \DataPath/RF/bus_selected_win_data[504] ,
         \DataPath/RF/bus_selected_win_data[505] ,
         \DataPath/RF/bus_selected_win_data[506] ,
         \DataPath/RF/bus_selected_win_data[507] ,
         \DataPath/RF/bus_selected_win_data[508] ,
         \DataPath/RF/bus_selected_win_data[509] ,
         \DataPath/RF/bus_selected_win_data[510] ,
         \DataPath/RF/bus_selected_win_data[511] ,
         \DataPath/RF/bus_selected_win_data[512] ,
         \DataPath/RF/bus_selected_win_data[513] ,
         \DataPath/RF/bus_selected_win_data[514] ,
         \DataPath/RF/bus_selected_win_data[515] ,
         \DataPath/RF/bus_selected_win_data[516] ,
         \DataPath/RF/bus_selected_win_data[517] ,
         \DataPath/RF/bus_selected_win_data[518] ,
         \DataPath/RF/bus_selected_win_data[519] ,
         \DataPath/RF/bus_selected_win_data[520] ,
         \DataPath/RF/bus_selected_win_data[521] ,
         \DataPath/RF/bus_selected_win_data[522] ,
         \DataPath/RF/bus_selected_win_data[523] ,
         \DataPath/RF/bus_selected_win_data[524] ,
         \DataPath/RF/bus_selected_win_data[525] ,
         \DataPath/RF/bus_selected_win_data[526] ,
         \DataPath/RF/bus_selected_win_data[527] ,
         \DataPath/RF/bus_selected_win_data[528] ,
         \DataPath/RF/bus_selected_win_data[529] ,
         \DataPath/RF/bus_selected_win_data[530] ,
         \DataPath/RF/bus_selected_win_data[531] ,
         \DataPath/RF/bus_selected_win_data[532] ,
         \DataPath/RF/bus_selected_win_data[533] ,
         \DataPath/RF/bus_selected_win_data[534] ,
         \DataPath/RF/bus_selected_win_data[535] ,
         \DataPath/RF/bus_selected_win_data[536] ,
         \DataPath/RF/bus_selected_win_data[537] ,
         \DataPath/RF/bus_selected_win_data[538] ,
         \DataPath/RF/bus_selected_win_data[539] ,
         \DataPath/RF/bus_selected_win_data[540] ,
         \DataPath/RF/bus_selected_win_data[541] ,
         \DataPath/RF/bus_selected_win_data[542] ,
         \DataPath/RF/bus_selected_win_data[543] ,
         \DataPath/RF/bus_selected_win_data[544] ,
         \DataPath/RF/bus_selected_win_data[545] ,
         \DataPath/RF/bus_selected_win_data[546] ,
         \DataPath/RF/bus_selected_win_data[547] ,
         \DataPath/RF/bus_selected_win_data[548] ,
         \DataPath/RF/bus_selected_win_data[549] ,
         \DataPath/RF/bus_selected_win_data[550] ,
         \DataPath/RF/bus_selected_win_data[551] ,
         \DataPath/RF/bus_selected_win_data[552] ,
         \DataPath/RF/bus_selected_win_data[553] ,
         \DataPath/RF/bus_selected_win_data[554] ,
         \DataPath/RF/bus_selected_win_data[555] ,
         \DataPath/RF/bus_selected_win_data[556] ,
         \DataPath/RF/bus_selected_win_data[557] ,
         \DataPath/RF/bus_selected_win_data[558] ,
         \DataPath/RF/bus_selected_win_data[559] ,
         \DataPath/RF/bus_selected_win_data[560] ,
         \DataPath/RF/bus_selected_win_data[561] ,
         \DataPath/RF/bus_selected_win_data[562] ,
         \DataPath/RF/bus_selected_win_data[563] ,
         \DataPath/RF/bus_selected_win_data[564] ,
         \DataPath/RF/bus_selected_win_data[565] ,
         \DataPath/RF/bus_selected_win_data[566] ,
         \DataPath/RF/bus_selected_win_data[567] ,
         \DataPath/RF/bus_selected_win_data[568] ,
         \DataPath/RF/bus_selected_win_data[569] ,
         \DataPath/RF/bus_selected_win_data[570] ,
         \DataPath/RF/bus_selected_win_data[571] ,
         \DataPath/RF/bus_selected_win_data[572] ,
         \DataPath/RF/bus_selected_win_data[573] ,
         \DataPath/RF/bus_selected_win_data[574] ,
         \DataPath/RF/bus_selected_win_data[575] ,
         \DataPath/RF/bus_selected_win_data[576] ,
         \DataPath/RF/bus_selected_win_data[577] ,
         \DataPath/RF/bus_selected_win_data[578] ,
         \DataPath/RF/bus_selected_win_data[579] ,
         \DataPath/RF/bus_selected_win_data[580] ,
         \DataPath/RF/bus_selected_win_data[581] ,
         \DataPath/RF/bus_selected_win_data[582] ,
         \DataPath/RF/bus_selected_win_data[583] ,
         \DataPath/RF/bus_selected_win_data[584] ,
         \DataPath/RF/bus_selected_win_data[585] ,
         \DataPath/RF/bus_selected_win_data[586] ,
         \DataPath/RF/bus_selected_win_data[587] ,
         \DataPath/RF/bus_selected_win_data[588] ,
         \DataPath/RF/bus_selected_win_data[589] ,
         \DataPath/RF/bus_selected_win_data[590] ,
         \DataPath/RF/bus_selected_win_data[591] ,
         \DataPath/RF/bus_selected_win_data[592] ,
         \DataPath/RF/bus_selected_win_data[593] ,
         \DataPath/RF/bus_selected_win_data[594] ,
         \DataPath/RF/bus_selected_win_data[595] ,
         \DataPath/RF/bus_selected_win_data[596] ,
         \DataPath/RF/bus_selected_win_data[597] ,
         \DataPath/RF/bus_selected_win_data[598] ,
         \DataPath/RF/bus_selected_win_data[599] ,
         \DataPath/RF/bus_selected_win_data[600] ,
         \DataPath/RF/bus_selected_win_data[601] ,
         \DataPath/RF/bus_selected_win_data[602] ,
         \DataPath/RF/bus_selected_win_data[603] ,
         \DataPath/RF/bus_selected_win_data[604] ,
         \DataPath/RF/bus_selected_win_data[605] ,
         \DataPath/RF/bus_selected_win_data[606] ,
         \DataPath/RF/bus_selected_win_data[607] ,
         \DataPath/RF/bus_selected_win_data[608] ,
         \DataPath/RF/bus_selected_win_data[609] ,
         \DataPath/RF/bus_selected_win_data[610] ,
         \DataPath/RF/bus_selected_win_data[611] ,
         \DataPath/RF/bus_selected_win_data[612] ,
         \DataPath/RF/bus_selected_win_data[613] ,
         \DataPath/RF/bus_selected_win_data[614] ,
         \DataPath/RF/bus_selected_win_data[615] ,
         \DataPath/RF/bus_selected_win_data[616] ,
         \DataPath/RF/bus_selected_win_data[617] ,
         \DataPath/RF/bus_selected_win_data[618] ,
         \DataPath/RF/bus_selected_win_data[619] ,
         \DataPath/RF/bus_selected_win_data[620] ,
         \DataPath/RF/bus_selected_win_data[621] ,
         \DataPath/RF/bus_selected_win_data[622] ,
         \DataPath/RF/bus_selected_win_data[623] ,
         \DataPath/RF/bus_selected_win_data[624] ,
         \DataPath/RF/bus_selected_win_data[625] ,
         \DataPath/RF/bus_selected_win_data[626] ,
         \DataPath/RF/bus_selected_win_data[627] ,
         \DataPath/RF/bus_selected_win_data[628] ,
         \DataPath/RF/bus_selected_win_data[629] ,
         \DataPath/RF/bus_selected_win_data[630] ,
         \DataPath/RF/bus_selected_win_data[631] ,
         \DataPath/RF/bus_selected_win_data[632] ,
         \DataPath/RF/bus_selected_win_data[633] ,
         \DataPath/RF/bus_selected_win_data[634] ,
         \DataPath/RF/bus_selected_win_data[635] ,
         \DataPath/RF/bus_selected_win_data[636] ,
         \DataPath/RF/bus_selected_win_data[637] ,
         \DataPath/RF/bus_selected_win_data[638] ,
         \DataPath/RF/bus_selected_win_data[639] ,
         \DataPath/RF/bus_selected_win_data[640] ,
         \DataPath/RF/bus_selected_win_data[641] ,
         \DataPath/RF/bus_selected_win_data[642] ,
         \DataPath/RF/bus_selected_win_data[643] ,
         \DataPath/RF/bus_selected_win_data[644] ,
         \DataPath/RF/bus_selected_win_data[645] ,
         \DataPath/RF/bus_selected_win_data[646] ,
         \DataPath/RF/bus_selected_win_data[647] ,
         \DataPath/RF/bus_selected_win_data[648] ,
         \DataPath/RF/bus_selected_win_data[649] ,
         \DataPath/RF/bus_selected_win_data[650] ,
         \DataPath/RF/bus_selected_win_data[651] ,
         \DataPath/RF/bus_selected_win_data[652] ,
         \DataPath/RF/bus_selected_win_data[653] ,
         \DataPath/RF/bus_selected_win_data[654] ,
         \DataPath/RF/bus_selected_win_data[655] ,
         \DataPath/RF/bus_selected_win_data[656] ,
         \DataPath/RF/bus_selected_win_data[657] ,
         \DataPath/RF/bus_selected_win_data[658] ,
         \DataPath/RF/bus_selected_win_data[659] ,
         \DataPath/RF/bus_selected_win_data[660] ,
         \DataPath/RF/bus_selected_win_data[661] ,
         \DataPath/RF/bus_selected_win_data[662] ,
         \DataPath/RF/bus_selected_win_data[663] ,
         \DataPath/RF/bus_selected_win_data[664] ,
         \DataPath/RF/bus_selected_win_data[665] ,
         \DataPath/RF/bus_selected_win_data[666] ,
         \DataPath/RF/bus_selected_win_data[667] ,
         \DataPath/RF/bus_selected_win_data[668] ,
         \DataPath/RF/bus_selected_win_data[669] ,
         \DataPath/RF/bus_selected_win_data[670] ,
         \DataPath/RF/bus_selected_win_data[671] ,
         \DataPath/RF/bus_selected_win_data[672] ,
         \DataPath/RF/bus_selected_win_data[673] ,
         \DataPath/RF/bus_selected_win_data[674] ,
         \DataPath/RF/bus_selected_win_data[675] ,
         \DataPath/RF/bus_selected_win_data[676] ,
         \DataPath/RF/bus_selected_win_data[677] ,
         \DataPath/RF/bus_selected_win_data[678] ,
         \DataPath/RF/bus_selected_win_data[679] ,
         \DataPath/RF/bus_selected_win_data[680] ,
         \DataPath/RF/bus_selected_win_data[681] ,
         \DataPath/RF/bus_selected_win_data[682] ,
         \DataPath/RF/bus_selected_win_data[683] ,
         \DataPath/RF/bus_selected_win_data[684] ,
         \DataPath/RF/bus_selected_win_data[685] ,
         \DataPath/RF/bus_selected_win_data[686] ,
         \DataPath/RF/bus_selected_win_data[687] ,
         \DataPath/RF/bus_selected_win_data[688] ,
         \DataPath/RF/bus_selected_win_data[689] ,
         \DataPath/RF/bus_selected_win_data[690] ,
         \DataPath/RF/bus_selected_win_data[691] ,
         \DataPath/RF/bus_selected_win_data[692] ,
         \DataPath/RF/bus_selected_win_data[693] ,
         \DataPath/RF/bus_selected_win_data[694] ,
         \DataPath/RF/bus_selected_win_data[695] ,
         \DataPath/RF/bus_selected_win_data[696] ,
         \DataPath/RF/bus_selected_win_data[697] ,
         \DataPath/RF/bus_selected_win_data[698] ,
         \DataPath/RF/bus_selected_win_data[699] ,
         \DataPath/RF/bus_selected_win_data[700] ,
         \DataPath/RF/bus_selected_win_data[701] ,
         \DataPath/RF/bus_selected_win_data[702] ,
         \DataPath/RF/bus_selected_win_data[703] ,
         \DataPath/RF/bus_selected_win_data[704] ,
         \DataPath/RF/bus_selected_win_data[705] ,
         \DataPath/RF/bus_selected_win_data[706] ,
         \DataPath/RF/bus_selected_win_data[707] ,
         \DataPath/RF/bus_selected_win_data[708] ,
         \DataPath/RF/bus_selected_win_data[709] ,
         \DataPath/RF/bus_selected_win_data[710] ,
         \DataPath/RF/bus_selected_win_data[711] ,
         \DataPath/RF/bus_selected_win_data[712] ,
         \DataPath/RF/bus_selected_win_data[713] ,
         \DataPath/RF/bus_selected_win_data[714] ,
         \DataPath/RF/bus_selected_win_data[715] ,
         \DataPath/RF/bus_selected_win_data[716] ,
         \DataPath/RF/bus_selected_win_data[717] ,
         \DataPath/RF/bus_selected_win_data[718] ,
         \DataPath/RF/bus_selected_win_data[719] ,
         \DataPath/RF/bus_selected_win_data[720] ,
         \DataPath/RF/bus_selected_win_data[721] ,
         \DataPath/RF/bus_selected_win_data[722] ,
         \DataPath/RF/bus_selected_win_data[723] ,
         \DataPath/RF/bus_selected_win_data[724] ,
         \DataPath/RF/bus_selected_win_data[725] ,
         \DataPath/RF/bus_selected_win_data[726] ,
         \DataPath/RF/bus_selected_win_data[727] ,
         \DataPath/RF/bus_selected_win_data[728] ,
         \DataPath/RF/bus_selected_win_data[729] ,
         \DataPath/RF/bus_selected_win_data[730] ,
         \DataPath/RF/bus_selected_win_data[731] ,
         \DataPath/RF/bus_selected_win_data[732] ,
         \DataPath/RF/bus_selected_win_data[733] ,
         \DataPath/RF/bus_selected_win_data[734] ,
         \DataPath/RF/bus_selected_win_data[735] ,
         \DataPath/RF/bus_selected_win_data[736] ,
         \DataPath/RF/bus_selected_win_data[737] ,
         \DataPath/RF/bus_selected_win_data[738] ,
         \DataPath/RF/bus_selected_win_data[739] ,
         \DataPath/RF/bus_selected_win_data[740] ,
         \DataPath/RF/bus_selected_win_data[741] ,
         \DataPath/RF/bus_selected_win_data[742] ,
         \DataPath/RF/bus_selected_win_data[743] ,
         \DataPath/RF/bus_selected_win_data[744] ,
         \DataPath/RF/bus_selected_win_data[745] ,
         \DataPath/RF/bus_selected_win_data[746] ,
         \DataPath/RF/bus_selected_win_data[747] ,
         \DataPath/RF/bus_selected_win_data[748] ,
         \DataPath/RF/bus_selected_win_data[749] ,
         \DataPath/RF/bus_selected_win_data[750] ,
         \DataPath/RF/bus_selected_win_data[751] ,
         \DataPath/RF/bus_selected_win_data[752] ,
         \DataPath/RF/bus_selected_win_data[753] ,
         \DataPath/RF/bus_selected_win_data[754] ,
         \DataPath/RF/bus_selected_win_data[755] ,
         \DataPath/RF/bus_selected_win_data[756] ,
         \DataPath/RF/bus_selected_win_data[757] ,
         \DataPath/RF/bus_selected_win_data[758] ,
         \DataPath/RF/bus_selected_win_data[759] ,
         \DataPath/RF/bus_selected_win_data[760] ,
         \DataPath/RF/bus_selected_win_data[761] ,
         \DataPath/RF/bus_selected_win_data[762] ,
         \DataPath/RF/bus_selected_win_data[763] ,
         \DataPath/RF/bus_selected_win_data[764] ,
         \DataPath/RF/bus_selected_win_data[765] ,
         \DataPath/RF/bus_selected_win_data[766] ,
         \DataPath/RF/bus_selected_win_data[767] ,
         \DataPath/RF/bus_reg_dataout[0] , \DataPath/RF/bus_reg_dataout[1] ,
         \DataPath/RF/bus_reg_dataout[2] , \DataPath/RF/bus_reg_dataout[3] ,
         \DataPath/RF/bus_reg_dataout[4] , \DataPath/RF/bus_reg_dataout[5] ,
         \DataPath/RF/bus_reg_dataout[6] , \DataPath/RF/bus_reg_dataout[7] ,
         \DataPath/RF/bus_reg_dataout[8] , \DataPath/RF/bus_reg_dataout[9] ,
         \DataPath/RF/bus_reg_dataout[10] , \DataPath/RF/bus_reg_dataout[11] ,
         \DataPath/RF/bus_reg_dataout[12] , \DataPath/RF/bus_reg_dataout[13] ,
         \DataPath/RF/bus_reg_dataout[14] , \DataPath/RF/bus_reg_dataout[15] ,
         \DataPath/RF/bus_reg_dataout[16] , \DataPath/RF/bus_reg_dataout[17] ,
         \DataPath/RF/bus_reg_dataout[18] , \DataPath/RF/bus_reg_dataout[19] ,
         \DataPath/RF/bus_reg_dataout[20] , \DataPath/RF/bus_reg_dataout[21] ,
         \DataPath/RF/bus_reg_dataout[22] , \DataPath/RF/bus_reg_dataout[23] ,
         \DataPath/RF/bus_reg_dataout[24] , \DataPath/RF/bus_reg_dataout[25] ,
         \DataPath/RF/bus_reg_dataout[26] , \DataPath/RF/bus_reg_dataout[27] ,
         \DataPath/RF/bus_reg_dataout[28] , \DataPath/RF/bus_reg_dataout[29] ,
         \DataPath/RF/bus_reg_dataout[30] , \DataPath/RF/bus_reg_dataout[31] ,
         \DataPath/RF/bus_reg_dataout[32] , \DataPath/RF/bus_reg_dataout[33] ,
         \DataPath/RF/bus_reg_dataout[34] , \DataPath/RF/bus_reg_dataout[35] ,
         \DataPath/RF/bus_reg_dataout[36] , \DataPath/RF/bus_reg_dataout[37] ,
         \DataPath/RF/bus_reg_dataout[38] , \DataPath/RF/bus_reg_dataout[39] ,
         \DataPath/RF/bus_reg_dataout[40] , \DataPath/RF/bus_reg_dataout[41] ,
         \DataPath/RF/bus_reg_dataout[42] , \DataPath/RF/bus_reg_dataout[43] ,
         \DataPath/RF/bus_reg_dataout[44] , \DataPath/RF/bus_reg_dataout[45] ,
         \DataPath/RF/bus_reg_dataout[46] , \DataPath/RF/bus_reg_dataout[47] ,
         \DataPath/RF/bus_reg_dataout[48] , \DataPath/RF/bus_reg_dataout[49] ,
         \DataPath/RF/bus_reg_dataout[50] , \DataPath/RF/bus_reg_dataout[51] ,
         \DataPath/RF/bus_reg_dataout[52] , \DataPath/RF/bus_reg_dataout[53] ,
         \DataPath/RF/bus_reg_dataout[54] , \DataPath/RF/bus_reg_dataout[55] ,
         \DataPath/RF/bus_reg_dataout[56] , \DataPath/RF/bus_reg_dataout[57] ,
         \DataPath/RF/bus_reg_dataout[58] , \DataPath/RF/bus_reg_dataout[59] ,
         \DataPath/RF/bus_reg_dataout[60] , \DataPath/RF/bus_reg_dataout[61] ,
         \DataPath/RF/bus_reg_dataout[62] , \DataPath/RF/bus_reg_dataout[63] ,
         \DataPath/RF/bus_reg_dataout[64] , \DataPath/RF/bus_reg_dataout[65] ,
         \DataPath/RF/bus_reg_dataout[66] , \DataPath/RF/bus_reg_dataout[67] ,
         \DataPath/RF/bus_reg_dataout[68] , \DataPath/RF/bus_reg_dataout[69] ,
         \DataPath/RF/bus_reg_dataout[70] , \DataPath/RF/bus_reg_dataout[71] ,
         \DataPath/RF/bus_reg_dataout[72] , \DataPath/RF/bus_reg_dataout[73] ,
         \DataPath/RF/bus_reg_dataout[74] , \DataPath/RF/bus_reg_dataout[75] ,
         \DataPath/RF/bus_reg_dataout[76] , \DataPath/RF/bus_reg_dataout[77] ,
         \DataPath/RF/bus_reg_dataout[78] , \DataPath/RF/bus_reg_dataout[79] ,
         \DataPath/RF/bus_reg_dataout[80] , \DataPath/RF/bus_reg_dataout[81] ,
         \DataPath/RF/bus_reg_dataout[82] , \DataPath/RF/bus_reg_dataout[83] ,
         \DataPath/RF/bus_reg_dataout[84] , \DataPath/RF/bus_reg_dataout[85] ,
         \DataPath/RF/bus_reg_dataout[86] , \DataPath/RF/bus_reg_dataout[87] ,
         \DataPath/RF/bus_reg_dataout[88] , \DataPath/RF/bus_reg_dataout[89] ,
         \DataPath/RF/bus_reg_dataout[90] , \DataPath/RF/bus_reg_dataout[91] ,
         \DataPath/RF/bus_reg_dataout[92] , \DataPath/RF/bus_reg_dataout[93] ,
         \DataPath/RF/bus_reg_dataout[94] , \DataPath/RF/bus_reg_dataout[95] ,
         \DataPath/RF/bus_reg_dataout[96] , \DataPath/RF/bus_reg_dataout[97] ,
         \DataPath/RF/bus_reg_dataout[98] , \DataPath/RF/bus_reg_dataout[99] ,
         \DataPath/RF/bus_reg_dataout[100] ,
         \DataPath/RF/bus_reg_dataout[101] ,
         \DataPath/RF/bus_reg_dataout[102] ,
         \DataPath/RF/bus_reg_dataout[103] ,
         \DataPath/RF/bus_reg_dataout[104] ,
         \DataPath/RF/bus_reg_dataout[105] ,
         \DataPath/RF/bus_reg_dataout[106] ,
         \DataPath/RF/bus_reg_dataout[107] ,
         \DataPath/RF/bus_reg_dataout[108] ,
         \DataPath/RF/bus_reg_dataout[109] ,
         \DataPath/RF/bus_reg_dataout[110] ,
         \DataPath/RF/bus_reg_dataout[111] ,
         \DataPath/RF/bus_reg_dataout[112] ,
         \DataPath/RF/bus_reg_dataout[113] ,
         \DataPath/RF/bus_reg_dataout[114] ,
         \DataPath/RF/bus_reg_dataout[115] ,
         \DataPath/RF/bus_reg_dataout[116] ,
         \DataPath/RF/bus_reg_dataout[117] ,
         \DataPath/RF/bus_reg_dataout[118] ,
         \DataPath/RF/bus_reg_dataout[119] ,
         \DataPath/RF/bus_reg_dataout[120] ,
         \DataPath/RF/bus_reg_dataout[121] ,
         \DataPath/RF/bus_reg_dataout[122] ,
         \DataPath/RF/bus_reg_dataout[123] ,
         \DataPath/RF/bus_reg_dataout[124] ,
         \DataPath/RF/bus_reg_dataout[125] ,
         \DataPath/RF/bus_reg_dataout[126] ,
         \DataPath/RF/bus_reg_dataout[127] ,
         \DataPath/RF/bus_reg_dataout[128] ,
         \DataPath/RF/bus_reg_dataout[129] ,
         \DataPath/RF/bus_reg_dataout[130] ,
         \DataPath/RF/bus_reg_dataout[131] ,
         \DataPath/RF/bus_reg_dataout[132] ,
         \DataPath/RF/bus_reg_dataout[133] ,
         \DataPath/RF/bus_reg_dataout[134] ,
         \DataPath/RF/bus_reg_dataout[135] ,
         \DataPath/RF/bus_reg_dataout[136] ,
         \DataPath/RF/bus_reg_dataout[137] ,
         \DataPath/RF/bus_reg_dataout[138] ,
         \DataPath/RF/bus_reg_dataout[139] ,
         \DataPath/RF/bus_reg_dataout[140] ,
         \DataPath/RF/bus_reg_dataout[141] ,
         \DataPath/RF/bus_reg_dataout[142] ,
         \DataPath/RF/bus_reg_dataout[143] ,
         \DataPath/RF/bus_reg_dataout[144] ,
         \DataPath/RF/bus_reg_dataout[145] ,
         \DataPath/RF/bus_reg_dataout[146] ,
         \DataPath/RF/bus_reg_dataout[147] ,
         \DataPath/RF/bus_reg_dataout[148] ,
         \DataPath/RF/bus_reg_dataout[149] ,
         \DataPath/RF/bus_reg_dataout[150] ,
         \DataPath/RF/bus_reg_dataout[151] ,
         \DataPath/RF/bus_reg_dataout[152] ,
         \DataPath/RF/bus_reg_dataout[153] ,
         \DataPath/RF/bus_reg_dataout[154] ,
         \DataPath/RF/bus_reg_dataout[155] ,
         \DataPath/RF/bus_reg_dataout[156] ,
         \DataPath/RF/bus_reg_dataout[157] ,
         \DataPath/RF/bus_reg_dataout[158] ,
         \DataPath/RF/bus_reg_dataout[159] ,
         \DataPath/RF/bus_reg_dataout[160] ,
         \DataPath/RF/bus_reg_dataout[161] ,
         \DataPath/RF/bus_reg_dataout[162] ,
         \DataPath/RF/bus_reg_dataout[163] ,
         \DataPath/RF/bus_reg_dataout[164] ,
         \DataPath/RF/bus_reg_dataout[165] ,
         \DataPath/RF/bus_reg_dataout[166] ,
         \DataPath/RF/bus_reg_dataout[167] ,
         \DataPath/RF/bus_reg_dataout[168] ,
         \DataPath/RF/bus_reg_dataout[169] ,
         \DataPath/RF/bus_reg_dataout[170] ,
         \DataPath/RF/bus_reg_dataout[171] ,
         \DataPath/RF/bus_reg_dataout[172] ,
         \DataPath/RF/bus_reg_dataout[173] ,
         \DataPath/RF/bus_reg_dataout[174] ,
         \DataPath/RF/bus_reg_dataout[175] ,
         \DataPath/RF/bus_reg_dataout[176] ,
         \DataPath/RF/bus_reg_dataout[177] ,
         \DataPath/RF/bus_reg_dataout[178] ,
         \DataPath/RF/bus_reg_dataout[179] ,
         \DataPath/RF/bus_reg_dataout[180] ,
         \DataPath/RF/bus_reg_dataout[181] ,
         \DataPath/RF/bus_reg_dataout[182] ,
         \DataPath/RF/bus_reg_dataout[183] ,
         \DataPath/RF/bus_reg_dataout[184] ,
         \DataPath/RF/bus_reg_dataout[185] ,
         \DataPath/RF/bus_reg_dataout[186] ,
         \DataPath/RF/bus_reg_dataout[187] ,
         \DataPath/RF/bus_reg_dataout[188] ,
         \DataPath/RF/bus_reg_dataout[189] ,
         \DataPath/RF/bus_reg_dataout[190] ,
         \DataPath/RF/bus_reg_dataout[191] ,
         \DataPath/RF/bus_reg_dataout[192] ,
         \DataPath/RF/bus_reg_dataout[193] ,
         \DataPath/RF/bus_reg_dataout[194] ,
         \DataPath/RF/bus_reg_dataout[195] ,
         \DataPath/RF/bus_reg_dataout[196] ,
         \DataPath/RF/bus_reg_dataout[197] ,
         \DataPath/RF/bus_reg_dataout[198] ,
         \DataPath/RF/bus_reg_dataout[199] ,
         \DataPath/RF/bus_reg_dataout[200] ,
         \DataPath/RF/bus_reg_dataout[201] ,
         \DataPath/RF/bus_reg_dataout[202] ,
         \DataPath/RF/bus_reg_dataout[203] ,
         \DataPath/RF/bus_reg_dataout[204] ,
         \DataPath/RF/bus_reg_dataout[205] ,
         \DataPath/RF/bus_reg_dataout[206] ,
         \DataPath/RF/bus_reg_dataout[207] ,
         \DataPath/RF/bus_reg_dataout[208] ,
         \DataPath/RF/bus_reg_dataout[209] ,
         \DataPath/RF/bus_reg_dataout[210] ,
         \DataPath/RF/bus_reg_dataout[211] ,
         \DataPath/RF/bus_reg_dataout[212] ,
         \DataPath/RF/bus_reg_dataout[213] ,
         \DataPath/RF/bus_reg_dataout[214] ,
         \DataPath/RF/bus_reg_dataout[215] ,
         \DataPath/RF/bus_reg_dataout[216] ,
         \DataPath/RF/bus_reg_dataout[217] ,
         \DataPath/RF/bus_reg_dataout[218] ,
         \DataPath/RF/bus_reg_dataout[219] ,
         \DataPath/RF/bus_reg_dataout[220] ,
         \DataPath/RF/bus_reg_dataout[221] ,
         \DataPath/RF/bus_reg_dataout[222] ,
         \DataPath/RF/bus_reg_dataout[223] ,
         \DataPath/RF/bus_reg_dataout[224] ,
         \DataPath/RF/bus_reg_dataout[225] ,
         \DataPath/RF/bus_reg_dataout[226] ,
         \DataPath/RF/bus_reg_dataout[227] ,
         \DataPath/RF/bus_reg_dataout[228] ,
         \DataPath/RF/bus_reg_dataout[229] ,
         \DataPath/RF/bus_reg_dataout[230] ,
         \DataPath/RF/bus_reg_dataout[231] ,
         \DataPath/RF/bus_reg_dataout[232] ,
         \DataPath/RF/bus_reg_dataout[233] ,
         \DataPath/RF/bus_reg_dataout[234] ,
         \DataPath/RF/bus_reg_dataout[235] ,
         \DataPath/RF/bus_reg_dataout[236] ,
         \DataPath/RF/bus_reg_dataout[237] ,
         \DataPath/RF/bus_reg_dataout[238] ,
         \DataPath/RF/bus_reg_dataout[239] ,
         \DataPath/RF/bus_reg_dataout[240] ,
         \DataPath/RF/bus_reg_dataout[241] ,
         \DataPath/RF/bus_reg_dataout[242] ,
         \DataPath/RF/bus_reg_dataout[243] ,
         \DataPath/RF/bus_reg_dataout[244] ,
         \DataPath/RF/bus_reg_dataout[245] ,
         \DataPath/RF/bus_reg_dataout[246] ,
         \DataPath/RF/bus_reg_dataout[247] ,
         \DataPath/RF/bus_reg_dataout[248] ,
         \DataPath/RF/bus_reg_dataout[249] ,
         \DataPath/RF/bus_reg_dataout[250] ,
         \DataPath/RF/bus_reg_dataout[251] ,
         \DataPath/RF/bus_reg_dataout[252] ,
         \DataPath/RF/bus_reg_dataout[253] ,
         \DataPath/RF/bus_reg_dataout[254] ,
         \DataPath/RF/bus_reg_dataout[255] ,
         \DataPath/RF/bus_reg_dataout[256] ,
         \DataPath/RF/bus_reg_dataout[257] ,
         \DataPath/RF/bus_reg_dataout[258] ,
         \DataPath/RF/bus_reg_dataout[259] ,
         \DataPath/RF/bus_reg_dataout[260] ,
         \DataPath/RF/bus_reg_dataout[261] ,
         \DataPath/RF/bus_reg_dataout[262] ,
         \DataPath/RF/bus_reg_dataout[263] ,
         \DataPath/RF/bus_reg_dataout[264] ,
         \DataPath/RF/bus_reg_dataout[265] ,
         \DataPath/RF/bus_reg_dataout[266] ,
         \DataPath/RF/bus_reg_dataout[267] ,
         \DataPath/RF/bus_reg_dataout[268] ,
         \DataPath/RF/bus_reg_dataout[269] ,
         \DataPath/RF/bus_reg_dataout[270] ,
         \DataPath/RF/bus_reg_dataout[271] ,
         \DataPath/RF/bus_reg_dataout[272] ,
         \DataPath/RF/bus_reg_dataout[273] ,
         \DataPath/RF/bus_reg_dataout[274] ,
         \DataPath/RF/bus_reg_dataout[275] ,
         \DataPath/RF/bus_reg_dataout[276] ,
         \DataPath/RF/bus_reg_dataout[277] ,
         \DataPath/RF/bus_reg_dataout[278] ,
         \DataPath/RF/bus_reg_dataout[279] ,
         \DataPath/RF/bus_reg_dataout[280] ,
         \DataPath/RF/bus_reg_dataout[281] ,
         \DataPath/RF/bus_reg_dataout[282] ,
         \DataPath/RF/bus_reg_dataout[283] ,
         \DataPath/RF/bus_reg_dataout[284] ,
         \DataPath/RF/bus_reg_dataout[285] ,
         \DataPath/RF/bus_reg_dataout[286] ,
         \DataPath/RF/bus_reg_dataout[287] ,
         \DataPath/RF/bus_reg_dataout[288] ,
         \DataPath/RF/bus_reg_dataout[289] ,
         \DataPath/RF/bus_reg_dataout[290] ,
         \DataPath/RF/bus_reg_dataout[291] ,
         \DataPath/RF/bus_reg_dataout[292] ,
         \DataPath/RF/bus_reg_dataout[293] ,
         \DataPath/RF/bus_reg_dataout[294] ,
         \DataPath/RF/bus_reg_dataout[295] ,
         \DataPath/RF/bus_reg_dataout[296] ,
         \DataPath/RF/bus_reg_dataout[297] ,
         \DataPath/RF/bus_reg_dataout[298] ,
         \DataPath/RF/bus_reg_dataout[299] ,
         \DataPath/RF/bus_reg_dataout[300] ,
         \DataPath/RF/bus_reg_dataout[301] ,
         \DataPath/RF/bus_reg_dataout[302] ,
         \DataPath/RF/bus_reg_dataout[303] ,
         \DataPath/RF/bus_reg_dataout[304] ,
         \DataPath/RF/bus_reg_dataout[305] ,
         \DataPath/RF/bus_reg_dataout[306] ,
         \DataPath/RF/bus_reg_dataout[307] ,
         \DataPath/RF/bus_reg_dataout[308] ,
         \DataPath/RF/bus_reg_dataout[309] ,
         \DataPath/RF/bus_reg_dataout[310] ,
         \DataPath/RF/bus_reg_dataout[311] ,
         \DataPath/RF/bus_reg_dataout[312] ,
         \DataPath/RF/bus_reg_dataout[313] ,
         \DataPath/RF/bus_reg_dataout[314] ,
         \DataPath/RF/bus_reg_dataout[315] ,
         \DataPath/RF/bus_reg_dataout[316] ,
         \DataPath/RF/bus_reg_dataout[317] ,
         \DataPath/RF/bus_reg_dataout[318] ,
         \DataPath/RF/bus_reg_dataout[319] ,
         \DataPath/RF/bus_reg_dataout[320] ,
         \DataPath/RF/bus_reg_dataout[321] ,
         \DataPath/RF/bus_reg_dataout[322] ,
         \DataPath/RF/bus_reg_dataout[323] ,
         \DataPath/RF/bus_reg_dataout[324] ,
         \DataPath/RF/bus_reg_dataout[325] ,
         \DataPath/RF/bus_reg_dataout[326] ,
         \DataPath/RF/bus_reg_dataout[327] ,
         \DataPath/RF/bus_reg_dataout[328] ,
         \DataPath/RF/bus_reg_dataout[329] ,
         \DataPath/RF/bus_reg_dataout[330] ,
         \DataPath/RF/bus_reg_dataout[331] ,
         \DataPath/RF/bus_reg_dataout[332] ,
         \DataPath/RF/bus_reg_dataout[333] ,
         \DataPath/RF/bus_reg_dataout[334] ,
         \DataPath/RF/bus_reg_dataout[335] ,
         \DataPath/RF/bus_reg_dataout[336] ,
         \DataPath/RF/bus_reg_dataout[337] ,
         \DataPath/RF/bus_reg_dataout[338] ,
         \DataPath/RF/bus_reg_dataout[339] ,
         \DataPath/RF/bus_reg_dataout[340] ,
         \DataPath/RF/bus_reg_dataout[341] ,
         \DataPath/RF/bus_reg_dataout[342] ,
         \DataPath/RF/bus_reg_dataout[343] ,
         \DataPath/RF/bus_reg_dataout[344] ,
         \DataPath/RF/bus_reg_dataout[345] ,
         \DataPath/RF/bus_reg_dataout[346] ,
         \DataPath/RF/bus_reg_dataout[347] ,
         \DataPath/RF/bus_reg_dataout[348] ,
         \DataPath/RF/bus_reg_dataout[349] ,
         \DataPath/RF/bus_reg_dataout[350] ,
         \DataPath/RF/bus_reg_dataout[351] ,
         \DataPath/RF/bus_reg_dataout[352] ,
         \DataPath/RF/bus_reg_dataout[353] ,
         \DataPath/RF/bus_reg_dataout[354] ,
         \DataPath/RF/bus_reg_dataout[355] ,
         \DataPath/RF/bus_reg_dataout[356] ,
         \DataPath/RF/bus_reg_dataout[357] ,
         \DataPath/RF/bus_reg_dataout[358] ,
         \DataPath/RF/bus_reg_dataout[359] ,
         \DataPath/RF/bus_reg_dataout[360] ,
         \DataPath/RF/bus_reg_dataout[361] ,
         \DataPath/RF/bus_reg_dataout[362] ,
         \DataPath/RF/bus_reg_dataout[363] ,
         \DataPath/RF/bus_reg_dataout[364] ,
         \DataPath/RF/bus_reg_dataout[365] ,
         \DataPath/RF/bus_reg_dataout[366] ,
         \DataPath/RF/bus_reg_dataout[367] ,
         \DataPath/RF/bus_reg_dataout[368] ,
         \DataPath/RF/bus_reg_dataout[369] ,
         \DataPath/RF/bus_reg_dataout[370] ,
         \DataPath/RF/bus_reg_dataout[371] ,
         \DataPath/RF/bus_reg_dataout[372] ,
         \DataPath/RF/bus_reg_dataout[373] ,
         \DataPath/RF/bus_reg_dataout[374] ,
         \DataPath/RF/bus_reg_dataout[375] ,
         \DataPath/RF/bus_reg_dataout[376] ,
         \DataPath/RF/bus_reg_dataout[377] ,
         \DataPath/RF/bus_reg_dataout[378] ,
         \DataPath/RF/bus_reg_dataout[379] ,
         \DataPath/RF/bus_reg_dataout[380] ,
         \DataPath/RF/bus_reg_dataout[381] ,
         \DataPath/RF/bus_reg_dataout[382] ,
         \DataPath/RF/bus_reg_dataout[383] ,
         \DataPath/RF/bus_reg_dataout[384] ,
         \DataPath/RF/bus_reg_dataout[385] ,
         \DataPath/RF/bus_reg_dataout[386] ,
         \DataPath/RF/bus_reg_dataout[387] ,
         \DataPath/RF/bus_reg_dataout[388] ,
         \DataPath/RF/bus_reg_dataout[389] ,
         \DataPath/RF/bus_reg_dataout[390] ,
         \DataPath/RF/bus_reg_dataout[391] ,
         \DataPath/RF/bus_reg_dataout[392] ,
         \DataPath/RF/bus_reg_dataout[393] ,
         \DataPath/RF/bus_reg_dataout[394] ,
         \DataPath/RF/bus_reg_dataout[395] ,
         \DataPath/RF/bus_reg_dataout[396] ,
         \DataPath/RF/bus_reg_dataout[397] ,
         \DataPath/RF/bus_reg_dataout[398] ,
         \DataPath/RF/bus_reg_dataout[399] ,
         \DataPath/RF/bus_reg_dataout[400] ,
         \DataPath/RF/bus_reg_dataout[401] ,
         \DataPath/RF/bus_reg_dataout[402] ,
         \DataPath/RF/bus_reg_dataout[403] ,
         \DataPath/RF/bus_reg_dataout[404] ,
         \DataPath/RF/bus_reg_dataout[405] ,
         \DataPath/RF/bus_reg_dataout[406] ,
         \DataPath/RF/bus_reg_dataout[407] ,
         \DataPath/RF/bus_reg_dataout[408] ,
         \DataPath/RF/bus_reg_dataout[409] ,
         \DataPath/RF/bus_reg_dataout[410] ,
         \DataPath/RF/bus_reg_dataout[411] ,
         \DataPath/RF/bus_reg_dataout[412] ,
         \DataPath/RF/bus_reg_dataout[413] ,
         \DataPath/RF/bus_reg_dataout[414] ,
         \DataPath/RF/bus_reg_dataout[415] ,
         \DataPath/RF/bus_reg_dataout[416] ,
         \DataPath/RF/bus_reg_dataout[417] ,
         \DataPath/RF/bus_reg_dataout[418] ,
         \DataPath/RF/bus_reg_dataout[419] ,
         \DataPath/RF/bus_reg_dataout[420] ,
         \DataPath/RF/bus_reg_dataout[421] ,
         \DataPath/RF/bus_reg_dataout[422] ,
         \DataPath/RF/bus_reg_dataout[423] ,
         \DataPath/RF/bus_reg_dataout[424] ,
         \DataPath/RF/bus_reg_dataout[425] ,
         \DataPath/RF/bus_reg_dataout[426] ,
         \DataPath/RF/bus_reg_dataout[427] ,
         \DataPath/RF/bus_reg_dataout[428] ,
         \DataPath/RF/bus_reg_dataout[429] ,
         \DataPath/RF/bus_reg_dataout[430] ,
         \DataPath/RF/bus_reg_dataout[431] ,
         \DataPath/RF/bus_reg_dataout[432] ,
         \DataPath/RF/bus_reg_dataout[433] ,
         \DataPath/RF/bus_reg_dataout[434] ,
         \DataPath/RF/bus_reg_dataout[435] ,
         \DataPath/RF/bus_reg_dataout[436] ,
         \DataPath/RF/bus_reg_dataout[437] ,
         \DataPath/RF/bus_reg_dataout[438] ,
         \DataPath/RF/bus_reg_dataout[439] ,
         \DataPath/RF/bus_reg_dataout[440] ,
         \DataPath/RF/bus_reg_dataout[441] ,
         \DataPath/RF/bus_reg_dataout[442] ,
         \DataPath/RF/bus_reg_dataout[443] ,
         \DataPath/RF/bus_reg_dataout[444] ,
         \DataPath/RF/bus_reg_dataout[445] ,
         \DataPath/RF/bus_reg_dataout[446] ,
         \DataPath/RF/bus_reg_dataout[447] ,
         \DataPath/RF/bus_reg_dataout[448] ,
         \DataPath/RF/bus_reg_dataout[449] ,
         \DataPath/RF/bus_reg_dataout[450] ,
         \DataPath/RF/bus_reg_dataout[451] ,
         \DataPath/RF/bus_reg_dataout[452] ,
         \DataPath/RF/bus_reg_dataout[453] ,
         \DataPath/RF/bus_reg_dataout[454] ,
         \DataPath/RF/bus_reg_dataout[455] ,
         \DataPath/RF/bus_reg_dataout[456] ,
         \DataPath/RF/bus_reg_dataout[457] ,
         \DataPath/RF/bus_reg_dataout[458] ,
         \DataPath/RF/bus_reg_dataout[459] ,
         \DataPath/RF/bus_reg_dataout[460] ,
         \DataPath/RF/bus_reg_dataout[461] ,
         \DataPath/RF/bus_reg_dataout[462] ,
         \DataPath/RF/bus_reg_dataout[463] ,
         \DataPath/RF/bus_reg_dataout[464] ,
         \DataPath/RF/bus_reg_dataout[465] ,
         \DataPath/RF/bus_reg_dataout[466] ,
         \DataPath/RF/bus_reg_dataout[467] ,
         \DataPath/RF/bus_reg_dataout[468] ,
         \DataPath/RF/bus_reg_dataout[469] ,
         \DataPath/RF/bus_reg_dataout[470] ,
         \DataPath/RF/bus_reg_dataout[471] ,
         \DataPath/RF/bus_reg_dataout[472] ,
         \DataPath/RF/bus_reg_dataout[473] ,
         \DataPath/RF/bus_reg_dataout[474] ,
         \DataPath/RF/bus_reg_dataout[475] ,
         \DataPath/RF/bus_reg_dataout[476] ,
         \DataPath/RF/bus_reg_dataout[477] ,
         \DataPath/RF/bus_reg_dataout[478] ,
         \DataPath/RF/bus_reg_dataout[479] ,
         \DataPath/RF/bus_reg_dataout[480] ,
         \DataPath/RF/bus_reg_dataout[481] ,
         \DataPath/RF/bus_reg_dataout[482] ,
         \DataPath/RF/bus_reg_dataout[483] ,
         \DataPath/RF/bus_reg_dataout[484] ,
         \DataPath/RF/bus_reg_dataout[485] ,
         \DataPath/RF/bus_reg_dataout[486] ,
         \DataPath/RF/bus_reg_dataout[487] ,
         \DataPath/RF/bus_reg_dataout[488] ,
         \DataPath/RF/bus_reg_dataout[489] ,
         \DataPath/RF/bus_reg_dataout[490] ,
         \DataPath/RF/bus_reg_dataout[491] ,
         \DataPath/RF/bus_reg_dataout[492] ,
         \DataPath/RF/bus_reg_dataout[493] ,
         \DataPath/RF/bus_reg_dataout[494] ,
         \DataPath/RF/bus_reg_dataout[495] ,
         \DataPath/RF/bus_reg_dataout[496] ,
         \DataPath/RF/bus_reg_dataout[497] ,
         \DataPath/RF/bus_reg_dataout[498] ,
         \DataPath/RF/bus_reg_dataout[499] ,
         \DataPath/RF/bus_reg_dataout[500] ,
         \DataPath/RF/bus_reg_dataout[501] ,
         \DataPath/RF/bus_reg_dataout[502] ,
         \DataPath/RF/bus_reg_dataout[503] ,
         \DataPath/RF/bus_reg_dataout[504] ,
         \DataPath/RF/bus_reg_dataout[505] ,
         \DataPath/RF/bus_reg_dataout[506] ,
         \DataPath/RF/bus_reg_dataout[507] ,
         \DataPath/RF/bus_reg_dataout[508] ,
         \DataPath/RF/bus_reg_dataout[509] ,
         \DataPath/RF/bus_reg_dataout[510] ,
         \DataPath/RF/bus_reg_dataout[511] ,
         \DataPath/RF/bus_reg_dataout[512] ,
         \DataPath/RF/bus_reg_dataout[513] ,
         \DataPath/RF/bus_reg_dataout[514] ,
         \DataPath/RF/bus_reg_dataout[515] ,
         \DataPath/RF/bus_reg_dataout[516] ,
         \DataPath/RF/bus_reg_dataout[517] ,
         \DataPath/RF/bus_reg_dataout[518] ,
         \DataPath/RF/bus_reg_dataout[519] ,
         \DataPath/RF/bus_reg_dataout[520] ,
         \DataPath/RF/bus_reg_dataout[521] ,
         \DataPath/RF/bus_reg_dataout[522] ,
         \DataPath/RF/bus_reg_dataout[523] ,
         \DataPath/RF/bus_reg_dataout[524] ,
         \DataPath/RF/bus_reg_dataout[525] ,
         \DataPath/RF/bus_reg_dataout[526] ,
         \DataPath/RF/bus_reg_dataout[527] ,
         \DataPath/RF/bus_reg_dataout[528] ,
         \DataPath/RF/bus_reg_dataout[529] ,
         \DataPath/RF/bus_reg_dataout[530] ,
         \DataPath/RF/bus_reg_dataout[531] ,
         \DataPath/RF/bus_reg_dataout[532] ,
         \DataPath/RF/bus_reg_dataout[533] ,
         \DataPath/RF/bus_reg_dataout[534] ,
         \DataPath/RF/bus_reg_dataout[535] ,
         \DataPath/RF/bus_reg_dataout[536] ,
         \DataPath/RF/bus_reg_dataout[537] ,
         \DataPath/RF/bus_reg_dataout[538] ,
         \DataPath/RF/bus_reg_dataout[539] ,
         \DataPath/RF/bus_reg_dataout[540] ,
         \DataPath/RF/bus_reg_dataout[541] ,
         \DataPath/RF/bus_reg_dataout[542] ,
         \DataPath/RF/bus_reg_dataout[543] ,
         \DataPath/RF/bus_reg_dataout[544] ,
         \DataPath/RF/bus_reg_dataout[545] ,
         \DataPath/RF/bus_reg_dataout[546] ,
         \DataPath/RF/bus_reg_dataout[547] ,
         \DataPath/RF/bus_reg_dataout[548] ,
         \DataPath/RF/bus_reg_dataout[549] ,
         \DataPath/RF/bus_reg_dataout[550] ,
         \DataPath/RF/bus_reg_dataout[551] ,
         \DataPath/RF/bus_reg_dataout[552] ,
         \DataPath/RF/bus_reg_dataout[553] ,
         \DataPath/RF/bus_reg_dataout[554] ,
         \DataPath/RF/bus_reg_dataout[555] ,
         \DataPath/RF/bus_reg_dataout[556] ,
         \DataPath/RF/bus_reg_dataout[557] ,
         \DataPath/RF/bus_reg_dataout[558] ,
         \DataPath/RF/bus_reg_dataout[559] ,
         \DataPath/RF/bus_reg_dataout[560] ,
         \DataPath/RF/bus_reg_dataout[561] ,
         \DataPath/RF/bus_reg_dataout[562] ,
         \DataPath/RF/bus_reg_dataout[563] ,
         \DataPath/RF/bus_reg_dataout[564] ,
         \DataPath/RF/bus_reg_dataout[565] ,
         \DataPath/RF/bus_reg_dataout[566] ,
         \DataPath/RF/bus_reg_dataout[567] ,
         \DataPath/RF/bus_reg_dataout[568] ,
         \DataPath/RF/bus_reg_dataout[569] ,
         \DataPath/RF/bus_reg_dataout[570] ,
         \DataPath/RF/bus_reg_dataout[571] ,
         \DataPath/RF/bus_reg_dataout[572] ,
         \DataPath/RF/bus_reg_dataout[573] ,
         \DataPath/RF/bus_reg_dataout[574] ,
         \DataPath/RF/bus_reg_dataout[575] ,
         \DataPath/RF/bus_reg_dataout[576] ,
         \DataPath/RF/bus_reg_dataout[577] ,
         \DataPath/RF/bus_reg_dataout[578] ,
         \DataPath/RF/bus_reg_dataout[579] ,
         \DataPath/RF/bus_reg_dataout[580] ,
         \DataPath/RF/bus_reg_dataout[581] ,
         \DataPath/RF/bus_reg_dataout[582] ,
         \DataPath/RF/bus_reg_dataout[583] ,
         \DataPath/RF/bus_reg_dataout[584] ,
         \DataPath/RF/bus_reg_dataout[585] ,
         \DataPath/RF/bus_reg_dataout[586] ,
         \DataPath/RF/bus_reg_dataout[587] ,
         \DataPath/RF/bus_reg_dataout[588] ,
         \DataPath/RF/bus_reg_dataout[589] ,
         \DataPath/RF/bus_reg_dataout[590] ,
         \DataPath/RF/bus_reg_dataout[591] ,
         \DataPath/RF/bus_reg_dataout[592] ,
         \DataPath/RF/bus_reg_dataout[593] ,
         \DataPath/RF/bus_reg_dataout[594] ,
         \DataPath/RF/bus_reg_dataout[595] ,
         \DataPath/RF/bus_reg_dataout[596] ,
         \DataPath/RF/bus_reg_dataout[597] ,
         \DataPath/RF/bus_reg_dataout[598] ,
         \DataPath/RF/bus_reg_dataout[599] ,
         \DataPath/RF/bus_reg_dataout[600] ,
         \DataPath/RF/bus_reg_dataout[601] ,
         \DataPath/RF/bus_reg_dataout[602] ,
         \DataPath/RF/bus_reg_dataout[603] ,
         \DataPath/RF/bus_reg_dataout[604] ,
         \DataPath/RF/bus_reg_dataout[605] ,
         \DataPath/RF/bus_reg_dataout[606] ,
         \DataPath/RF/bus_reg_dataout[607] ,
         \DataPath/RF/bus_reg_dataout[608] ,
         \DataPath/RF/bus_reg_dataout[609] ,
         \DataPath/RF/bus_reg_dataout[610] ,
         \DataPath/RF/bus_reg_dataout[611] ,
         \DataPath/RF/bus_reg_dataout[612] ,
         \DataPath/RF/bus_reg_dataout[613] ,
         \DataPath/RF/bus_reg_dataout[614] ,
         \DataPath/RF/bus_reg_dataout[615] ,
         \DataPath/RF/bus_reg_dataout[616] ,
         \DataPath/RF/bus_reg_dataout[617] ,
         \DataPath/RF/bus_reg_dataout[618] ,
         \DataPath/RF/bus_reg_dataout[619] ,
         \DataPath/RF/bus_reg_dataout[620] ,
         \DataPath/RF/bus_reg_dataout[621] ,
         \DataPath/RF/bus_reg_dataout[622] ,
         \DataPath/RF/bus_reg_dataout[623] ,
         \DataPath/RF/bus_reg_dataout[624] ,
         \DataPath/RF/bus_reg_dataout[625] ,
         \DataPath/RF/bus_reg_dataout[626] ,
         \DataPath/RF/bus_reg_dataout[627] ,
         \DataPath/RF/bus_reg_dataout[628] ,
         \DataPath/RF/bus_reg_dataout[629] ,
         \DataPath/RF/bus_reg_dataout[630] ,
         \DataPath/RF/bus_reg_dataout[631] ,
         \DataPath/RF/bus_reg_dataout[632] ,
         \DataPath/RF/bus_reg_dataout[633] ,
         \DataPath/RF/bus_reg_dataout[634] ,
         \DataPath/RF/bus_reg_dataout[635] ,
         \DataPath/RF/bus_reg_dataout[636] ,
         \DataPath/RF/bus_reg_dataout[637] ,
         \DataPath/RF/bus_reg_dataout[638] ,
         \DataPath/RF/bus_reg_dataout[639] ,
         \DataPath/RF/bus_reg_dataout[640] ,
         \DataPath/RF/bus_reg_dataout[641] ,
         \DataPath/RF/bus_reg_dataout[642] ,
         \DataPath/RF/bus_reg_dataout[643] ,
         \DataPath/RF/bus_reg_dataout[644] ,
         \DataPath/RF/bus_reg_dataout[645] ,
         \DataPath/RF/bus_reg_dataout[646] ,
         \DataPath/RF/bus_reg_dataout[647] ,
         \DataPath/RF/bus_reg_dataout[648] ,
         \DataPath/RF/bus_reg_dataout[649] ,
         \DataPath/RF/bus_reg_dataout[650] ,
         \DataPath/RF/bus_reg_dataout[651] ,
         \DataPath/RF/bus_reg_dataout[652] ,
         \DataPath/RF/bus_reg_dataout[653] ,
         \DataPath/RF/bus_reg_dataout[654] ,
         \DataPath/RF/bus_reg_dataout[655] ,
         \DataPath/RF/bus_reg_dataout[656] ,
         \DataPath/RF/bus_reg_dataout[657] ,
         \DataPath/RF/bus_reg_dataout[658] ,
         \DataPath/RF/bus_reg_dataout[659] ,
         \DataPath/RF/bus_reg_dataout[660] ,
         \DataPath/RF/bus_reg_dataout[661] ,
         \DataPath/RF/bus_reg_dataout[662] ,
         \DataPath/RF/bus_reg_dataout[663] ,
         \DataPath/RF/bus_reg_dataout[664] ,
         \DataPath/RF/bus_reg_dataout[665] ,
         \DataPath/RF/bus_reg_dataout[666] ,
         \DataPath/RF/bus_reg_dataout[667] ,
         \DataPath/RF/bus_reg_dataout[668] ,
         \DataPath/RF/bus_reg_dataout[669] ,
         \DataPath/RF/bus_reg_dataout[670] ,
         \DataPath/RF/bus_reg_dataout[671] ,
         \DataPath/RF/bus_reg_dataout[672] ,
         \DataPath/RF/bus_reg_dataout[673] ,
         \DataPath/RF/bus_reg_dataout[674] ,
         \DataPath/RF/bus_reg_dataout[675] ,
         \DataPath/RF/bus_reg_dataout[676] ,
         \DataPath/RF/bus_reg_dataout[677] ,
         \DataPath/RF/bus_reg_dataout[678] ,
         \DataPath/RF/bus_reg_dataout[679] ,
         \DataPath/RF/bus_reg_dataout[680] ,
         \DataPath/RF/bus_reg_dataout[681] ,
         \DataPath/RF/bus_reg_dataout[682] ,
         \DataPath/RF/bus_reg_dataout[683] ,
         \DataPath/RF/bus_reg_dataout[684] ,
         \DataPath/RF/bus_reg_dataout[685] ,
         \DataPath/RF/bus_reg_dataout[686] ,
         \DataPath/RF/bus_reg_dataout[687] ,
         \DataPath/RF/bus_reg_dataout[688] ,
         \DataPath/RF/bus_reg_dataout[689] ,
         \DataPath/RF/bus_reg_dataout[690] ,
         \DataPath/RF/bus_reg_dataout[691] ,
         \DataPath/RF/bus_reg_dataout[692] ,
         \DataPath/RF/bus_reg_dataout[693] ,
         \DataPath/RF/bus_reg_dataout[694] ,
         \DataPath/RF/bus_reg_dataout[695] ,
         \DataPath/RF/bus_reg_dataout[696] ,
         \DataPath/RF/bus_reg_dataout[697] ,
         \DataPath/RF/bus_reg_dataout[698] ,
         \DataPath/RF/bus_reg_dataout[699] ,
         \DataPath/RF/bus_reg_dataout[700] ,
         \DataPath/RF/bus_reg_dataout[701] ,
         \DataPath/RF/bus_reg_dataout[702] ,
         \DataPath/RF/bus_reg_dataout[703] ,
         \DataPath/RF/bus_reg_dataout[704] ,
         \DataPath/RF/bus_reg_dataout[705] ,
         \DataPath/RF/bus_reg_dataout[706] ,
         \DataPath/RF/bus_reg_dataout[707] ,
         \DataPath/RF/bus_reg_dataout[708] ,
         \DataPath/RF/bus_reg_dataout[709] ,
         \DataPath/RF/bus_reg_dataout[710] ,
         \DataPath/RF/bus_reg_dataout[711] ,
         \DataPath/RF/bus_reg_dataout[712] ,
         \DataPath/RF/bus_reg_dataout[713] ,
         \DataPath/RF/bus_reg_dataout[714] ,
         \DataPath/RF/bus_reg_dataout[715] ,
         \DataPath/RF/bus_reg_dataout[716] ,
         \DataPath/RF/bus_reg_dataout[717] ,
         \DataPath/RF/bus_reg_dataout[718] ,
         \DataPath/RF/bus_reg_dataout[719] ,
         \DataPath/RF/bus_reg_dataout[720] ,
         \DataPath/RF/bus_reg_dataout[721] ,
         \DataPath/RF/bus_reg_dataout[722] ,
         \DataPath/RF/bus_reg_dataout[723] ,
         \DataPath/RF/bus_reg_dataout[724] ,
         \DataPath/RF/bus_reg_dataout[725] ,
         \DataPath/RF/bus_reg_dataout[726] ,
         \DataPath/RF/bus_reg_dataout[727] ,
         \DataPath/RF/bus_reg_dataout[728] ,
         \DataPath/RF/bus_reg_dataout[729] ,
         \DataPath/RF/bus_reg_dataout[730] ,
         \DataPath/RF/bus_reg_dataout[731] ,
         \DataPath/RF/bus_reg_dataout[732] ,
         \DataPath/RF/bus_reg_dataout[733] ,
         \DataPath/RF/bus_reg_dataout[734] ,
         \DataPath/RF/bus_reg_dataout[735] ,
         \DataPath/RF/bus_reg_dataout[736] ,
         \DataPath/RF/bus_reg_dataout[737] ,
         \DataPath/RF/bus_reg_dataout[738] ,
         \DataPath/RF/bus_reg_dataout[739] ,
         \DataPath/RF/bus_reg_dataout[740] ,
         \DataPath/RF/bus_reg_dataout[741] ,
         \DataPath/RF/bus_reg_dataout[742] ,
         \DataPath/RF/bus_reg_dataout[743] ,
         \DataPath/RF/bus_reg_dataout[744] ,
         \DataPath/RF/bus_reg_dataout[745] ,
         \DataPath/RF/bus_reg_dataout[746] ,
         \DataPath/RF/bus_reg_dataout[747] ,
         \DataPath/RF/bus_reg_dataout[748] ,
         \DataPath/RF/bus_reg_dataout[749] ,
         \DataPath/RF/bus_reg_dataout[750] ,
         \DataPath/RF/bus_reg_dataout[751] ,
         \DataPath/RF/bus_reg_dataout[752] ,
         \DataPath/RF/bus_reg_dataout[753] ,
         \DataPath/RF/bus_reg_dataout[754] ,
         \DataPath/RF/bus_reg_dataout[755] ,
         \DataPath/RF/bus_reg_dataout[756] ,
         \DataPath/RF/bus_reg_dataout[757] ,
         \DataPath/RF/bus_reg_dataout[758] ,
         \DataPath/RF/bus_reg_dataout[759] ,
         \DataPath/RF/bus_reg_dataout[760] ,
         \DataPath/RF/bus_reg_dataout[761] ,
         \DataPath/RF/bus_reg_dataout[762] ,
         \DataPath/RF/bus_reg_dataout[763] ,
         \DataPath/RF/bus_reg_dataout[764] ,
         \DataPath/RF/bus_reg_dataout[765] ,
         \DataPath/RF/bus_reg_dataout[766] ,
         \DataPath/RF/bus_reg_dataout[767] ,
         \DataPath/RF/bus_reg_dataout[768] ,
         \DataPath/RF/bus_reg_dataout[769] ,
         \DataPath/RF/bus_reg_dataout[770] ,
         \DataPath/RF/bus_reg_dataout[771] ,
         \DataPath/RF/bus_reg_dataout[772] ,
         \DataPath/RF/bus_reg_dataout[773] ,
         \DataPath/RF/bus_reg_dataout[774] ,
         \DataPath/RF/bus_reg_dataout[775] ,
         \DataPath/RF/bus_reg_dataout[776] ,
         \DataPath/RF/bus_reg_dataout[777] ,
         \DataPath/RF/bus_reg_dataout[778] ,
         \DataPath/RF/bus_reg_dataout[779] ,
         \DataPath/RF/bus_reg_dataout[780] ,
         \DataPath/RF/bus_reg_dataout[781] ,
         \DataPath/RF/bus_reg_dataout[782] ,
         \DataPath/RF/bus_reg_dataout[783] ,
         \DataPath/RF/bus_reg_dataout[784] ,
         \DataPath/RF/bus_reg_dataout[785] ,
         \DataPath/RF/bus_reg_dataout[786] ,
         \DataPath/RF/bus_reg_dataout[787] ,
         \DataPath/RF/bus_reg_dataout[788] ,
         \DataPath/RF/bus_reg_dataout[789] ,
         \DataPath/RF/bus_reg_dataout[790] ,
         \DataPath/RF/bus_reg_dataout[791] ,
         \DataPath/RF/bus_reg_dataout[792] ,
         \DataPath/RF/bus_reg_dataout[793] ,
         \DataPath/RF/bus_reg_dataout[794] ,
         \DataPath/RF/bus_reg_dataout[795] ,
         \DataPath/RF/bus_reg_dataout[796] ,
         \DataPath/RF/bus_reg_dataout[797] ,
         \DataPath/RF/bus_reg_dataout[798] ,
         \DataPath/RF/bus_reg_dataout[799] ,
         \DataPath/RF/bus_reg_dataout[800] ,
         \DataPath/RF/bus_reg_dataout[801] ,
         \DataPath/RF/bus_reg_dataout[802] ,
         \DataPath/RF/bus_reg_dataout[803] ,
         \DataPath/RF/bus_reg_dataout[804] ,
         \DataPath/RF/bus_reg_dataout[805] ,
         \DataPath/RF/bus_reg_dataout[806] ,
         \DataPath/RF/bus_reg_dataout[807] ,
         \DataPath/RF/bus_reg_dataout[808] ,
         \DataPath/RF/bus_reg_dataout[809] ,
         \DataPath/RF/bus_reg_dataout[810] ,
         \DataPath/RF/bus_reg_dataout[811] ,
         \DataPath/RF/bus_reg_dataout[812] ,
         \DataPath/RF/bus_reg_dataout[813] ,
         \DataPath/RF/bus_reg_dataout[814] ,
         \DataPath/RF/bus_reg_dataout[815] ,
         \DataPath/RF/bus_reg_dataout[816] ,
         \DataPath/RF/bus_reg_dataout[817] ,
         \DataPath/RF/bus_reg_dataout[818] ,
         \DataPath/RF/bus_reg_dataout[819] ,
         \DataPath/RF/bus_reg_dataout[820] ,
         \DataPath/RF/bus_reg_dataout[821] ,
         \DataPath/RF/bus_reg_dataout[822] ,
         \DataPath/RF/bus_reg_dataout[823] ,
         \DataPath/RF/bus_reg_dataout[824] ,
         \DataPath/RF/bus_reg_dataout[825] ,
         \DataPath/RF/bus_reg_dataout[826] ,
         \DataPath/RF/bus_reg_dataout[827] ,
         \DataPath/RF/bus_reg_dataout[828] ,
         \DataPath/RF/bus_reg_dataout[829] ,
         \DataPath/RF/bus_reg_dataout[830] ,
         \DataPath/RF/bus_reg_dataout[831] ,
         \DataPath/RF/bus_reg_dataout[832] ,
         \DataPath/RF/bus_reg_dataout[833] ,
         \DataPath/RF/bus_reg_dataout[834] ,
         \DataPath/RF/bus_reg_dataout[835] ,
         \DataPath/RF/bus_reg_dataout[836] ,
         \DataPath/RF/bus_reg_dataout[837] ,
         \DataPath/RF/bus_reg_dataout[838] ,
         \DataPath/RF/bus_reg_dataout[839] ,
         \DataPath/RF/bus_reg_dataout[840] ,
         \DataPath/RF/bus_reg_dataout[841] ,
         \DataPath/RF/bus_reg_dataout[842] ,
         \DataPath/RF/bus_reg_dataout[843] ,
         \DataPath/RF/bus_reg_dataout[844] ,
         \DataPath/RF/bus_reg_dataout[845] ,
         \DataPath/RF/bus_reg_dataout[846] ,
         \DataPath/RF/bus_reg_dataout[847] ,
         \DataPath/RF/bus_reg_dataout[848] ,
         \DataPath/RF/bus_reg_dataout[849] ,
         \DataPath/RF/bus_reg_dataout[850] ,
         \DataPath/RF/bus_reg_dataout[851] ,
         \DataPath/RF/bus_reg_dataout[852] ,
         \DataPath/RF/bus_reg_dataout[853] ,
         \DataPath/RF/bus_reg_dataout[854] ,
         \DataPath/RF/bus_reg_dataout[855] ,
         \DataPath/RF/bus_reg_dataout[856] ,
         \DataPath/RF/bus_reg_dataout[857] ,
         \DataPath/RF/bus_reg_dataout[858] ,
         \DataPath/RF/bus_reg_dataout[859] ,
         \DataPath/RF/bus_reg_dataout[860] ,
         \DataPath/RF/bus_reg_dataout[861] ,
         \DataPath/RF/bus_reg_dataout[862] ,
         \DataPath/RF/bus_reg_dataout[863] ,
         \DataPath/RF/bus_reg_dataout[864] ,
         \DataPath/RF/bus_reg_dataout[865] ,
         \DataPath/RF/bus_reg_dataout[866] ,
         \DataPath/RF/bus_reg_dataout[867] ,
         \DataPath/RF/bus_reg_dataout[868] ,
         \DataPath/RF/bus_reg_dataout[869] ,
         \DataPath/RF/bus_reg_dataout[870] ,
         \DataPath/RF/bus_reg_dataout[871] ,
         \DataPath/RF/bus_reg_dataout[872] ,
         \DataPath/RF/bus_reg_dataout[873] ,
         \DataPath/RF/bus_reg_dataout[874] ,
         \DataPath/RF/bus_reg_dataout[875] ,
         \DataPath/RF/bus_reg_dataout[876] ,
         \DataPath/RF/bus_reg_dataout[877] ,
         \DataPath/RF/bus_reg_dataout[878] ,
         \DataPath/RF/bus_reg_dataout[879] ,
         \DataPath/RF/bus_reg_dataout[880] ,
         \DataPath/RF/bus_reg_dataout[881] ,
         \DataPath/RF/bus_reg_dataout[882] ,
         \DataPath/RF/bus_reg_dataout[883] ,
         \DataPath/RF/bus_reg_dataout[884] ,
         \DataPath/RF/bus_reg_dataout[885] ,
         \DataPath/RF/bus_reg_dataout[886] ,
         \DataPath/RF/bus_reg_dataout[887] ,
         \DataPath/RF/bus_reg_dataout[888] ,
         \DataPath/RF/bus_reg_dataout[889] ,
         \DataPath/RF/bus_reg_dataout[890] ,
         \DataPath/RF/bus_reg_dataout[891] ,
         \DataPath/RF/bus_reg_dataout[892] ,
         \DataPath/RF/bus_reg_dataout[893] ,
         \DataPath/RF/bus_reg_dataout[894] ,
         \DataPath/RF/bus_reg_dataout[895] ,
         \DataPath/RF/bus_reg_dataout[896] ,
         \DataPath/RF/bus_reg_dataout[897] ,
         \DataPath/RF/bus_reg_dataout[898] ,
         \DataPath/RF/bus_reg_dataout[899] ,
         \DataPath/RF/bus_reg_dataout[900] ,
         \DataPath/RF/bus_reg_dataout[901] ,
         \DataPath/RF/bus_reg_dataout[902] ,
         \DataPath/RF/bus_reg_dataout[903] ,
         \DataPath/RF/bus_reg_dataout[904] ,
         \DataPath/RF/bus_reg_dataout[905] ,
         \DataPath/RF/bus_reg_dataout[906] ,
         \DataPath/RF/bus_reg_dataout[907] ,
         \DataPath/RF/bus_reg_dataout[908] ,
         \DataPath/RF/bus_reg_dataout[909] ,
         \DataPath/RF/bus_reg_dataout[910] ,
         \DataPath/RF/bus_reg_dataout[911] ,
         \DataPath/RF/bus_reg_dataout[912] ,
         \DataPath/RF/bus_reg_dataout[913] ,
         \DataPath/RF/bus_reg_dataout[914] ,
         \DataPath/RF/bus_reg_dataout[915] ,
         \DataPath/RF/bus_reg_dataout[916] ,
         \DataPath/RF/bus_reg_dataout[917] ,
         \DataPath/RF/bus_reg_dataout[918] ,
         \DataPath/RF/bus_reg_dataout[919] ,
         \DataPath/RF/bus_reg_dataout[920] ,
         \DataPath/RF/bus_reg_dataout[921] ,
         \DataPath/RF/bus_reg_dataout[922] ,
         \DataPath/RF/bus_reg_dataout[923] ,
         \DataPath/RF/bus_reg_dataout[924] ,
         \DataPath/RF/bus_reg_dataout[925] ,
         \DataPath/RF/bus_reg_dataout[926] ,
         \DataPath/RF/bus_reg_dataout[927] ,
         \DataPath/RF/bus_reg_dataout[928] ,
         \DataPath/RF/bus_reg_dataout[929] ,
         \DataPath/RF/bus_reg_dataout[930] ,
         \DataPath/RF/bus_reg_dataout[931] ,
         \DataPath/RF/bus_reg_dataout[932] ,
         \DataPath/RF/bus_reg_dataout[933] ,
         \DataPath/RF/bus_reg_dataout[934] ,
         \DataPath/RF/bus_reg_dataout[935] ,
         \DataPath/RF/bus_reg_dataout[936] ,
         \DataPath/RF/bus_reg_dataout[937] ,
         \DataPath/RF/bus_reg_dataout[938] ,
         \DataPath/RF/bus_reg_dataout[939] ,
         \DataPath/RF/bus_reg_dataout[940] ,
         \DataPath/RF/bus_reg_dataout[941] ,
         \DataPath/RF/bus_reg_dataout[942] ,
         \DataPath/RF/bus_reg_dataout[943] ,
         \DataPath/RF/bus_reg_dataout[944] ,
         \DataPath/RF/bus_reg_dataout[945] ,
         \DataPath/RF/bus_reg_dataout[946] ,
         \DataPath/RF/bus_reg_dataout[947] ,
         \DataPath/RF/bus_reg_dataout[948] ,
         \DataPath/RF/bus_reg_dataout[949] ,
         \DataPath/RF/bus_reg_dataout[950] ,
         \DataPath/RF/bus_reg_dataout[951] ,
         \DataPath/RF/bus_reg_dataout[952] ,
         \DataPath/RF/bus_reg_dataout[953] ,
         \DataPath/RF/bus_reg_dataout[954] ,
         \DataPath/RF/bus_reg_dataout[955] ,
         \DataPath/RF/bus_reg_dataout[956] ,
         \DataPath/RF/bus_reg_dataout[957] ,
         \DataPath/RF/bus_reg_dataout[958] ,
         \DataPath/RF/bus_reg_dataout[959] ,
         \DataPath/RF/bus_reg_dataout[960] ,
         \DataPath/RF/bus_reg_dataout[961] ,
         \DataPath/RF/bus_reg_dataout[962] ,
         \DataPath/RF/bus_reg_dataout[963] ,
         \DataPath/RF/bus_reg_dataout[964] ,
         \DataPath/RF/bus_reg_dataout[965] ,
         \DataPath/RF/bus_reg_dataout[966] ,
         \DataPath/RF/bus_reg_dataout[967] ,
         \DataPath/RF/bus_reg_dataout[968] ,
         \DataPath/RF/bus_reg_dataout[969] ,
         \DataPath/RF/bus_reg_dataout[970] ,
         \DataPath/RF/bus_reg_dataout[971] ,
         \DataPath/RF/bus_reg_dataout[972] ,
         \DataPath/RF/bus_reg_dataout[973] ,
         \DataPath/RF/bus_reg_dataout[974] ,
         \DataPath/RF/bus_reg_dataout[975] ,
         \DataPath/RF/bus_reg_dataout[976] ,
         \DataPath/RF/bus_reg_dataout[977] ,
         \DataPath/RF/bus_reg_dataout[978] ,
         \DataPath/RF/bus_reg_dataout[979] ,
         \DataPath/RF/bus_reg_dataout[980] ,
         \DataPath/RF/bus_reg_dataout[981] ,
         \DataPath/RF/bus_reg_dataout[982] ,
         \DataPath/RF/bus_reg_dataout[983] ,
         \DataPath/RF/bus_reg_dataout[984] ,
         \DataPath/RF/bus_reg_dataout[985] ,
         \DataPath/RF/bus_reg_dataout[986] ,
         \DataPath/RF/bus_reg_dataout[987] ,
         \DataPath/RF/bus_reg_dataout[988] ,
         \DataPath/RF/bus_reg_dataout[989] ,
         \DataPath/RF/bus_reg_dataout[990] ,
         \DataPath/RF/bus_reg_dataout[991] ,
         \DataPath/RF/bus_reg_dataout[992] ,
         \DataPath/RF/bus_reg_dataout[993] ,
         \DataPath/RF/bus_reg_dataout[994] ,
         \DataPath/RF/bus_reg_dataout[995] ,
         \DataPath/RF/bus_reg_dataout[996] ,
         \DataPath/RF/bus_reg_dataout[997] ,
         \DataPath/RF/bus_reg_dataout[998] ,
         \DataPath/RF/bus_reg_dataout[999] ,
         \DataPath/RF/bus_reg_dataout[1000] ,
         \DataPath/RF/bus_reg_dataout[1001] ,
         \DataPath/RF/bus_reg_dataout[1002] ,
         \DataPath/RF/bus_reg_dataout[1003] ,
         \DataPath/RF/bus_reg_dataout[1004] ,
         \DataPath/RF/bus_reg_dataout[1005] ,
         \DataPath/RF/bus_reg_dataout[1006] ,
         \DataPath/RF/bus_reg_dataout[1007] ,
         \DataPath/RF/bus_reg_dataout[1008] ,
         \DataPath/RF/bus_reg_dataout[1009] ,
         \DataPath/RF/bus_reg_dataout[1010] ,
         \DataPath/RF/bus_reg_dataout[1011] ,
         \DataPath/RF/bus_reg_dataout[1012] ,
         \DataPath/RF/bus_reg_dataout[1013] ,
         \DataPath/RF/bus_reg_dataout[1014] ,
         \DataPath/RF/bus_reg_dataout[1015] ,
         \DataPath/RF/bus_reg_dataout[1016] ,
         \DataPath/RF/bus_reg_dataout[1017] ,
         \DataPath/RF/bus_reg_dataout[1018] ,
         \DataPath/RF/bus_reg_dataout[1019] ,
         \DataPath/RF/bus_reg_dataout[1020] ,
         \DataPath/RF/bus_reg_dataout[1021] ,
         \DataPath/RF/bus_reg_dataout[1022] ,
         \DataPath/RF/bus_reg_dataout[1023] ,
         \DataPath/RF/bus_reg_dataout[1024] ,
         \DataPath/RF/bus_reg_dataout[1025] ,
         \DataPath/RF/bus_reg_dataout[1026] ,
         \DataPath/RF/bus_reg_dataout[1027] ,
         \DataPath/RF/bus_reg_dataout[1028] ,
         \DataPath/RF/bus_reg_dataout[1029] ,
         \DataPath/RF/bus_reg_dataout[1030] ,
         \DataPath/RF/bus_reg_dataout[1031] ,
         \DataPath/RF/bus_reg_dataout[1032] ,
         \DataPath/RF/bus_reg_dataout[1033] ,
         \DataPath/RF/bus_reg_dataout[1034] ,
         \DataPath/RF/bus_reg_dataout[1035] ,
         \DataPath/RF/bus_reg_dataout[1036] ,
         \DataPath/RF/bus_reg_dataout[1037] ,
         \DataPath/RF/bus_reg_dataout[1038] ,
         \DataPath/RF/bus_reg_dataout[1039] ,
         \DataPath/RF/bus_reg_dataout[1040] ,
         \DataPath/RF/bus_reg_dataout[1041] ,
         \DataPath/RF/bus_reg_dataout[1042] ,
         \DataPath/RF/bus_reg_dataout[1043] ,
         \DataPath/RF/bus_reg_dataout[1044] ,
         \DataPath/RF/bus_reg_dataout[1045] ,
         \DataPath/RF/bus_reg_dataout[1046] ,
         \DataPath/RF/bus_reg_dataout[1047] ,
         \DataPath/RF/bus_reg_dataout[1048] ,
         \DataPath/RF/bus_reg_dataout[1049] ,
         \DataPath/RF/bus_reg_dataout[1050] ,
         \DataPath/RF/bus_reg_dataout[1051] ,
         \DataPath/RF/bus_reg_dataout[1052] ,
         \DataPath/RF/bus_reg_dataout[1053] ,
         \DataPath/RF/bus_reg_dataout[1054] ,
         \DataPath/RF/bus_reg_dataout[1055] ,
         \DataPath/RF/bus_reg_dataout[1056] ,
         \DataPath/RF/bus_reg_dataout[1057] ,
         \DataPath/RF/bus_reg_dataout[1058] ,
         \DataPath/RF/bus_reg_dataout[1059] ,
         \DataPath/RF/bus_reg_dataout[1060] ,
         \DataPath/RF/bus_reg_dataout[1061] ,
         \DataPath/RF/bus_reg_dataout[1062] ,
         \DataPath/RF/bus_reg_dataout[1063] ,
         \DataPath/RF/bus_reg_dataout[1064] ,
         \DataPath/RF/bus_reg_dataout[1065] ,
         \DataPath/RF/bus_reg_dataout[1066] ,
         \DataPath/RF/bus_reg_dataout[1067] ,
         \DataPath/RF/bus_reg_dataout[1068] ,
         \DataPath/RF/bus_reg_dataout[1069] ,
         \DataPath/RF/bus_reg_dataout[1070] ,
         \DataPath/RF/bus_reg_dataout[1071] ,
         \DataPath/RF/bus_reg_dataout[1072] ,
         \DataPath/RF/bus_reg_dataout[1073] ,
         \DataPath/RF/bus_reg_dataout[1074] ,
         \DataPath/RF/bus_reg_dataout[1075] ,
         \DataPath/RF/bus_reg_dataout[1076] ,
         \DataPath/RF/bus_reg_dataout[1077] ,
         \DataPath/RF/bus_reg_dataout[1078] ,
         \DataPath/RF/bus_reg_dataout[1079] ,
         \DataPath/RF/bus_reg_dataout[1080] ,
         \DataPath/RF/bus_reg_dataout[1081] ,
         \DataPath/RF/bus_reg_dataout[1082] ,
         \DataPath/RF/bus_reg_dataout[1083] ,
         \DataPath/RF/bus_reg_dataout[1084] ,
         \DataPath/RF/bus_reg_dataout[1085] ,
         \DataPath/RF/bus_reg_dataout[1086] ,
         \DataPath/RF/bus_reg_dataout[1087] ,
         \DataPath/RF/bus_reg_dataout[1088] ,
         \DataPath/RF/bus_reg_dataout[1089] ,
         \DataPath/RF/bus_reg_dataout[1090] ,
         \DataPath/RF/bus_reg_dataout[1091] ,
         \DataPath/RF/bus_reg_dataout[1092] ,
         \DataPath/RF/bus_reg_dataout[1093] ,
         \DataPath/RF/bus_reg_dataout[1094] ,
         \DataPath/RF/bus_reg_dataout[1095] ,
         \DataPath/RF/bus_reg_dataout[1096] ,
         \DataPath/RF/bus_reg_dataout[1097] ,
         \DataPath/RF/bus_reg_dataout[1098] ,
         \DataPath/RF/bus_reg_dataout[1099] ,
         \DataPath/RF/bus_reg_dataout[1100] ,
         \DataPath/RF/bus_reg_dataout[1101] ,
         \DataPath/RF/bus_reg_dataout[1102] ,
         \DataPath/RF/bus_reg_dataout[1103] ,
         \DataPath/RF/bus_reg_dataout[1104] ,
         \DataPath/RF/bus_reg_dataout[1105] ,
         \DataPath/RF/bus_reg_dataout[1106] ,
         \DataPath/RF/bus_reg_dataout[1107] ,
         \DataPath/RF/bus_reg_dataout[1108] ,
         \DataPath/RF/bus_reg_dataout[1109] ,
         \DataPath/RF/bus_reg_dataout[1110] ,
         \DataPath/RF/bus_reg_dataout[1111] ,
         \DataPath/RF/bus_reg_dataout[1112] ,
         \DataPath/RF/bus_reg_dataout[1113] ,
         \DataPath/RF/bus_reg_dataout[1114] ,
         \DataPath/RF/bus_reg_dataout[1115] ,
         \DataPath/RF/bus_reg_dataout[1116] ,
         \DataPath/RF/bus_reg_dataout[1117] ,
         \DataPath/RF/bus_reg_dataout[1118] ,
         \DataPath/RF/bus_reg_dataout[1119] ,
         \DataPath/RF/bus_reg_dataout[1120] ,
         \DataPath/RF/bus_reg_dataout[1121] ,
         \DataPath/RF/bus_reg_dataout[1122] ,
         \DataPath/RF/bus_reg_dataout[1123] ,
         \DataPath/RF/bus_reg_dataout[1124] ,
         \DataPath/RF/bus_reg_dataout[1125] ,
         \DataPath/RF/bus_reg_dataout[1126] ,
         \DataPath/RF/bus_reg_dataout[1127] ,
         \DataPath/RF/bus_reg_dataout[1128] ,
         \DataPath/RF/bus_reg_dataout[1129] ,
         \DataPath/RF/bus_reg_dataout[1130] ,
         \DataPath/RF/bus_reg_dataout[1131] ,
         \DataPath/RF/bus_reg_dataout[1132] ,
         \DataPath/RF/bus_reg_dataout[1133] ,
         \DataPath/RF/bus_reg_dataout[1134] ,
         \DataPath/RF/bus_reg_dataout[1135] ,
         \DataPath/RF/bus_reg_dataout[1136] ,
         \DataPath/RF/bus_reg_dataout[1137] ,
         \DataPath/RF/bus_reg_dataout[1138] ,
         \DataPath/RF/bus_reg_dataout[1139] ,
         \DataPath/RF/bus_reg_dataout[1140] ,
         \DataPath/RF/bus_reg_dataout[1141] ,
         \DataPath/RF/bus_reg_dataout[1142] ,
         \DataPath/RF/bus_reg_dataout[1143] ,
         \DataPath/RF/bus_reg_dataout[1144] ,
         \DataPath/RF/bus_reg_dataout[1145] ,
         \DataPath/RF/bus_reg_dataout[1146] ,
         \DataPath/RF/bus_reg_dataout[1147] ,
         \DataPath/RF/bus_reg_dataout[1148] ,
         \DataPath/RF/bus_reg_dataout[1149] ,
         \DataPath/RF/bus_reg_dataout[1150] ,
         \DataPath/RF/bus_reg_dataout[1151] ,
         \DataPath/RF/bus_reg_dataout[1152] ,
         \DataPath/RF/bus_reg_dataout[1153] ,
         \DataPath/RF/bus_reg_dataout[1154] ,
         \DataPath/RF/bus_reg_dataout[1155] ,
         \DataPath/RF/bus_reg_dataout[1156] ,
         \DataPath/RF/bus_reg_dataout[1157] ,
         \DataPath/RF/bus_reg_dataout[1158] ,
         \DataPath/RF/bus_reg_dataout[1159] ,
         \DataPath/RF/bus_reg_dataout[1160] ,
         \DataPath/RF/bus_reg_dataout[1161] ,
         \DataPath/RF/bus_reg_dataout[1162] ,
         \DataPath/RF/bus_reg_dataout[1163] ,
         \DataPath/RF/bus_reg_dataout[1164] ,
         \DataPath/RF/bus_reg_dataout[1165] ,
         \DataPath/RF/bus_reg_dataout[1166] ,
         \DataPath/RF/bus_reg_dataout[1167] ,
         \DataPath/RF/bus_reg_dataout[1168] ,
         \DataPath/RF/bus_reg_dataout[1169] ,
         \DataPath/RF/bus_reg_dataout[1170] ,
         \DataPath/RF/bus_reg_dataout[1171] ,
         \DataPath/RF/bus_reg_dataout[1172] ,
         \DataPath/RF/bus_reg_dataout[1173] ,
         \DataPath/RF/bus_reg_dataout[1174] ,
         \DataPath/RF/bus_reg_dataout[1175] ,
         \DataPath/RF/bus_reg_dataout[1176] ,
         \DataPath/RF/bus_reg_dataout[1177] ,
         \DataPath/RF/bus_reg_dataout[1178] ,
         \DataPath/RF/bus_reg_dataout[1179] ,
         \DataPath/RF/bus_reg_dataout[1180] ,
         \DataPath/RF/bus_reg_dataout[1181] ,
         \DataPath/RF/bus_reg_dataout[1182] ,
         \DataPath/RF/bus_reg_dataout[1183] ,
         \DataPath/RF/bus_reg_dataout[1184] ,
         \DataPath/RF/bus_reg_dataout[1185] ,
         \DataPath/RF/bus_reg_dataout[1186] ,
         \DataPath/RF/bus_reg_dataout[1187] ,
         \DataPath/RF/bus_reg_dataout[1188] ,
         \DataPath/RF/bus_reg_dataout[1189] ,
         \DataPath/RF/bus_reg_dataout[1190] ,
         \DataPath/RF/bus_reg_dataout[1191] ,
         \DataPath/RF/bus_reg_dataout[1192] ,
         \DataPath/RF/bus_reg_dataout[1193] ,
         \DataPath/RF/bus_reg_dataout[1194] ,
         \DataPath/RF/bus_reg_dataout[1195] ,
         \DataPath/RF/bus_reg_dataout[1196] ,
         \DataPath/RF/bus_reg_dataout[1197] ,
         \DataPath/RF/bus_reg_dataout[1198] ,
         \DataPath/RF/bus_reg_dataout[1199] ,
         \DataPath/RF/bus_reg_dataout[1200] ,
         \DataPath/RF/bus_reg_dataout[1201] ,
         \DataPath/RF/bus_reg_dataout[1202] ,
         \DataPath/RF/bus_reg_dataout[1203] ,
         \DataPath/RF/bus_reg_dataout[1204] ,
         \DataPath/RF/bus_reg_dataout[1205] ,
         \DataPath/RF/bus_reg_dataout[1206] ,
         \DataPath/RF/bus_reg_dataout[1207] ,
         \DataPath/RF/bus_reg_dataout[1208] ,
         \DataPath/RF/bus_reg_dataout[1209] ,
         \DataPath/RF/bus_reg_dataout[1210] ,
         \DataPath/RF/bus_reg_dataout[1211] ,
         \DataPath/RF/bus_reg_dataout[1212] ,
         \DataPath/RF/bus_reg_dataout[1213] ,
         \DataPath/RF/bus_reg_dataout[1214] ,
         \DataPath/RF/bus_reg_dataout[1215] ,
         \DataPath/RF/bus_reg_dataout[1216] ,
         \DataPath/RF/bus_reg_dataout[1217] ,
         \DataPath/RF/bus_reg_dataout[1218] ,
         \DataPath/RF/bus_reg_dataout[1219] ,
         \DataPath/RF/bus_reg_dataout[1220] ,
         \DataPath/RF/bus_reg_dataout[1221] ,
         \DataPath/RF/bus_reg_dataout[1222] ,
         \DataPath/RF/bus_reg_dataout[1223] ,
         \DataPath/RF/bus_reg_dataout[1224] ,
         \DataPath/RF/bus_reg_dataout[1225] ,
         \DataPath/RF/bus_reg_dataout[1226] ,
         \DataPath/RF/bus_reg_dataout[1227] ,
         \DataPath/RF/bus_reg_dataout[1228] ,
         \DataPath/RF/bus_reg_dataout[1229] ,
         \DataPath/RF/bus_reg_dataout[1230] ,
         \DataPath/RF/bus_reg_dataout[1231] ,
         \DataPath/RF/bus_reg_dataout[1232] ,
         \DataPath/RF/bus_reg_dataout[1233] ,
         \DataPath/RF/bus_reg_dataout[1234] ,
         \DataPath/RF/bus_reg_dataout[1235] ,
         \DataPath/RF/bus_reg_dataout[1236] ,
         \DataPath/RF/bus_reg_dataout[1237] ,
         \DataPath/RF/bus_reg_dataout[1238] ,
         \DataPath/RF/bus_reg_dataout[1239] ,
         \DataPath/RF/bus_reg_dataout[1240] ,
         \DataPath/RF/bus_reg_dataout[1241] ,
         \DataPath/RF/bus_reg_dataout[1242] ,
         \DataPath/RF/bus_reg_dataout[1243] ,
         \DataPath/RF/bus_reg_dataout[1244] ,
         \DataPath/RF/bus_reg_dataout[1245] ,
         \DataPath/RF/bus_reg_dataout[1246] ,
         \DataPath/RF/bus_reg_dataout[1247] ,
         \DataPath/RF/bus_reg_dataout[1248] ,
         \DataPath/RF/bus_reg_dataout[1249] ,
         \DataPath/RF/bus_reg_dataout[1250] ,
         \DataPath/RF/bus_reg_dataout[1251] ,
         \DataPath/RF/bus_reg_dataout[1252] ,
         \DataPath/RF/bus_reg_dataout[1253] ,
         \DataPath/RF/bus_reg_dataout[1254] ,
         \DataPath/RF/bus_reg_dataout[1255] ,
         \DataPath/RF/bus_reg_dataout[1256] ,
         \DataPath/RF/bus_reg_dataout[1257] ,
         \DataPath/RF/bus_reg_dataout[1258] ,
         \DataPath/RF/bus_reg_dataout[1259] ,
         \DataPath/RF/bus_reg_dataout[1260] ,
         \DataPath/RF/bus_reg_dataout[1261] ,
         \DataPath/RF/bus_reg_dataout[1262] ,
         \DataPath/RF/bus_reg_dataout[1263] ,
         \DataPath/RF/bus_reg_dataout[1264] ,
         \DataPath/RF/bus_reg_dataout[1265] ,
         \DataPath/RF/bus_reg_dataout[1266] ,
         \DataPath/RF/bus_reg_dataout[1267] ,
         \DataPath/RF/bus_reg_dataout[1268] ,
         \DataPath/RF/bus_reg_dataout[1269] ,
         \DataPath/RF/bus_reg_dataout[1270] ,
         \DataPath/RF/bus_reg_dataout[1271] ,
         \DataPath/RF/bus_reg_dataout[1272] ,
         \DataPath/RF/bus_reg_dataout[1273] ,
         \DataPath/RF/bus_reg_dataout[1274] ,
         \DataPath/RF/bus_reg_dataout[1275] ,
         \DataPath/RF/bus_reg_dataout[1276] ,
         \DataPath/RF/bus_reg_dataout[1277] ,
         \DataPath/RF/bus_reg_dataout[1278] ,
         \DataPath/RF/bus_reg_dataout[1279] ,
         \DataPath/RF/bus_reg_dataout[1280] ,
         \DataPath/RF/bus_reg_dataout[1281] ,
         \DataPath/RF/bus_reg_dataout[1282] ,
         \DataPath/RF/bus_reg_dataout[1283] ,
         \DataPath/RF/bus_reg_dataout[1284] ,
         \DataPath/RF/bus_reg_dataout[1285] ,
         \DataPath/RF/bus_reg_dataout[1286] ,
         \DataPath/RF/bus_reg_dataout[1287] ,
         \DataPath/RF/bus_reg_dataout[1288] ,
         \DataPath/RF/bus_reg_dataout[1289] ,
         \DataPath/RF/bus_reg_dataout[1290] ,
         \DataPath/RF/bus_reg_dataout[1291] ,
         \DataPath/RF/bus_reg_dataout[1292] ,
         \DataPath/RF/bus_reg_dataout[1293] ,
         \DataPath/RF/bus_reg_dataout[1294] ,
         \DataPath/RF/bus_reg_dataout[1295] ,
         \DataPath/RF/bus_reg_dataout[1296] ,
         \DataPath/RF/bus_reg_dataout[1297] ,
         \DataPath/RF/bus_reg_dataout[1298] ,
         \DataPath/RF/bus_reg_dataout[1299] ,
         \DataPath/RF/bus_reg_dataout[1300] ,
         \DataPath/RF/bus_reg_dataout[1301] ,
         \DataPath/RF/bus_reg_dataout[1302] ,
         \DataPath/RF/bus_reg_dataout[1303] ,
         \DataPath/RF/bus_reg_dataout[1304] ,
         \DataPath/RF/bus_reg_dataout[1305] ,
         \DataPath/RF/bus_reg_dataout[1306] ,
         \DataPath/RF/bus_reg_dataout[1307] ,
         \DataPath/RF/bus_reg_dataout[1308] ,
         \DataPath/RF/bus_reg_dataout[1309] ,
         \DataPath/RF/bus_reg_dataout[1310] ,
         \DataPath/RF/bus_reg_dataout[1311] ,
         \DataPath/RF/bus_reg_dataout[1312] ,
         \DataPath/RF/bus_reg_dataout[1313] ,
         \DataPath/RF/bus_reg_dataout[1314] ,
         \DataPath/RF/bus_reg_dataout[1315] ,
         \DataPath/RF/bus_reg_dataout[1316] ,
         \DataPath/RF/bus_reg_dataout[1317] ,
         \DataPath/RF/bus_reg_dataout[1318] ,
         \DataPath/RF/bus_reg_dataout[1319] ,
         \DataPath/RF/bus_reg_dataout[1320] ,
         \DataPath/RF/bus_reg_dataout[1321] ,
         \DataPath/RF/bus_reg_dataout[1322] ,
         \DataPath/RF/bus_reg_dataout[1323] ,
         \DataPath/RF/bus_reg_dataout[1324] ,
         \DataPath/RF/bus_reg_dataout[1325] ,
         \DataPath/RF/bus_reg_dataout[1326] ,
         \DataPath/RF/bus_reg_dataout[1327] ,
         \DataPath/RF/bus_reg_dataout[1328] ,
         \DataPath/RF/bus_reg_dataout[1329] ,
         \DataPath/RF/bus_reg_dataout[1330] ,
         \DataPath/RF/bus_reg_dataout[1331] ,
         \DataPath/RF/bus_reg_dataout[1332] ,
         \DataPath/RF/bus_reg_dataout[1333] ,
         \DataPath/RF/bus_reg_dataout[1334] ,
         \DataPath/RF/bus_reg_dataout[1335] ,
         \DataPath/RF/bus_reg_dataout[1336] ,
         \DataPath/RF/bus_reg_dataout[1337] ,
         \DataPath/RF/bus_reg_dataout[1338] ,
         \DataPath/RF/bus_reg_dataout[1339] ,
         \DataPath/RF/bus_reg_dataout[1340] ,
         \DataPath/RF/bus_reg_dataout[1341] ,
         \DataPath/RF/bus_reg_dataout[1342] ,
         \DataPath/RF/bus_reg_dataout[1343] ,
         \DataPath/RF/bus_reg_dataout[1344] ,
         \DataPath/RF/bus_reg_dataout[1345] ,
         \DataPath/RF/bus_reg_dataout[1346] ,
         \DataPath/RF/bus_reg_dataout[1347] ,
         \DataPath/RF/bus_reg_dataout[1348] ,
         \DataPath/RF/bus_reg_dataout[1349] ,
         \DataPath/RF/bus_reg_dataout[1350] ,
         \DataPath/RF/bus_reg_dataout[1351] ,
         \DataPath/RF/bus_reg_dataout[1352] ,
         \DataPath/RF/bus_reg_dataout[1353] ,
         \DataPath/RF/bus_reg_dataout[1354] ,
         \DataPath/RF/bus_reg_dataout[1355] ,
         \DataPath/RF/bus_reg_dataout[1356] ,
         \DataPath/RF/bus_reg_dataout[1357] ,
         \DataPath/RF/bus_reg_dataout[1358] ,
         \DataPath/RF/bus_reg_dataout[1359] ,
         \DataPath/RF/bus_reg_dataout[1360] ,
         \DataPath/RF/bus_reg_dataout[1361] ,
         \DataPath/RF/bus_reg_dataout[1362] ,
         \DataPath/RF/bus_reg_dataout[1363] ,
         \DataPath/RF/bus_reg_dataout[1364] ,
         \DataPath/RF/bus_reg_dataout[1365] ,
         \DataPath/RF/bus_reg_dataout[1366] ,
         \DataPath/RF/bus_reg_dataout[1367] ,
         \DataPath/RF/bus_reg_dataout[1368] ,
         \DataPath/RF/bus_reg_dataout[1369] ,
         \DataPath/RF/bus_reg_dataout[1370] ,
         \DataPath/RF/bus_reg_dataout[1371] ,
         \DataPath/RF/bus_reg_dataout[1372] ,
         \DataPath/RF/bus_reg_dataout[1373] ,
         \DataPath/RF/bus_reg_dataout[1374] ,
         \DataPath/RF/bus_reg_dataout[1375] ,
         \DataPath/RF/bus_reg_dataout[1376] ,
         \DataPath/RF/bus_reg_dataout[1377] ,
         \DataPath/RF/bus_reg_dataout[1378] ,
         \DataPath/RF/bus_reg_dataout[1379] ,
         \DataPath/RF/bus_reg_dataout[1380] ,
         \DataPath/RF/bus_reg_dataout[1381] ,
         \DataPath/RF/bus_reg_dataout[1382] ,
         \DataPath/RF/bus_reg_dataout[1383] ,
         \DataPath/RF/bus_reg_dataout[1384] ,
         \DataPath/RF/bus_reg_dataout[1385] ,
         \DataPath/RF/bus_reg_dataout[1386] ,
         \DataPath/RF/bus_reg_dataout[1387] ,
         \DataPath/RF/bus_reg_dataout[1388] ,
         \DataPath/RF/bus_reg_dataout[1389] ,
         \DataPath/RF/bus_reg_dataout[1390] ,
         \DataPath/RF/bus_reg_dataout[1391] ,
         \DataPath/RF/bus_reg_dataout[1392] ,
         \DataPath/RF/bus_reg_dataout[1393] ,
         \DataPath/RF/bus_reg_dataout[1394] ,
         \DataPath/RF/bus_reg_dataout[1395] ,
         \DataPath/RF/bus_reg_dataout[1396] ,
         \DataPath/RF/bus_reg_dataout[1397] ,
         \DataPath/RF/bus_reg_dataout[1398] ,
         \DataPath/RF/bus_reg_dataout[1399] ,
         \DataPath/RF/bus_reg_dataout[1400] ,
         \DataPath/RF/bus_reg_dataout[1401] ,
         \DataPath/RF/bus_reg_dataout[1402] ,
         \DataPath/RF/bus_reg_dataout[1403] ,
         \DataPath/RF/bus_reg_dataout[1404] ,
         \DataPath/RF/bus_reg_dataout[1405] ,
         \DataPath/RF/bus_reg_dataout[1406] ,
         \DataPath/RF/bus_reg_dataout[1407] ,
         \DataPath/RF/bus_reg_dataout[1408] ,
         \DataPath/RF/bus_reg_dataout[1409] ,
         \DataPath/RF/bus_reg_dataout[1410] ,
         \DataPath/RF/bus_reg_dataout[1411] ,
         \DataPath/RF/bus_reg_dataout[1412] ,
         \DataPath/RF/bus_reg_dataout[1413] ,
         \DataPath/RF/bus_reg_dataout[1414] ,
         \DataPath/RF/bus_reg_dataout[1415] ,
         \DataPath/RF/bus_reg_dataout[1416] ,
         \DataPath/RF/bus_reg_dataout[1417] ,
         \DataPath/RF/bus_reg_dataout[1418] ,
         \DataPath/RF/bus_reg_dataout[1419] ,
         \DataPath/RF/bus_reg_dataout[1420] ,
         \DataPath/RF/bus_reg_dataout[1421] ,
         \DataPath/RF/bus_reg_dataout[1422] ,
         \DataPath/RF/bus_reg_dataout[1423] ,
         \DataPath/RF/bus_reg_dataout[1424] ,
         \DataPath/RF/bus_reg_dataout[1425] ,
         \DataPath/RF/bus_reg_dataout[1426] ,
         \DataPath/RF/bus_reg_dataout[1427] ,
         \DataPath/RF/bus_reg_dataout[1428] ,
         \DataPath/RF/bus_reg_dataout[1429] ,
         \DataPath/RF/bus_reg_dataout[1430] ,
         \DataPath/RF/bus_reg_dataout[1431] ,
         \DataPath/RF/bus_reg_dataout[1432] ,
         \DataPath/RF/bus_reg_dataout[1433] ,
         \DataPath/RF/bus_reg_dataout[1434] ,
         \DataPath/RF/bus_reg_dataout[1435] ,
         \DataPath/RF/bus_reg_dataout[1436] ,
         \DataPath/RF/bus_reg_dataout[1437] ,
         \DataPath/RF/bus_reg_dataout[1438] ,
         \DataPath/RF/bus_reg_dataout[1439] ,
         \DataPath/RF/bus_reg_dataout[1440] ,
         \DataPath/RF/bus_reg_dataout[1441] ,
         \DataPath/RF/bus_reg_dataout[1442] ,
         \DataPath/RF/bus_reg_dataout[1443] ,
         \DataPath/RF/bus_reg_dataout[1444] ,
         \DataPath/RF/bus_reg_dataout[1445] ,
         \DataPath/RF/bus_reg_dataout[1446] ,
         \DataPath/RF/bus_reg_dataout[1447] ,
         \DataPath/RF/bus_reg_dataout[1448] ,
         \DataPath/RF/bus_reg_dataout[1449] ,
         \DataPath/RF/bus_reg_dataout[1450] ,
         \DataPath/RF/bus_reg_dataout[1451] ,
         \DataPath/RF/bus_reg_dataout[1452] ,
         \DataPath/RF/bus_reg_dataout[1453] ,
         \DataPath/RF/bus_reg_dataout[1454] ,
         \DataPath/RF/bus_reg_dataout[1455] ,
         \DataPath/RF/bus_reg_dataout[1456] ,
         \DataPath/RF/bus_reg_dataout[1457] ,
         \DataPath/RF/bus_reg_dataout[1458] ,
         \DataPath/RF/bus_reg_dataout[1459] ,
         \DataPath/RF/bus_reg_dataout[1460] ,
         \DataPath/RF/bus_reg_dataout[1461] ,
         \DataPath/RF/bus_reg_dataout[1462] ,
         \DataPath/RF/bus_reg_dataout[1463] ,
         \DataPath/RF/bus_reg_dataout[1464] ,
         \DataPath/RF/bus_reg_dataout[1465] ,
         \DataPath/RF/bus_reg_dataout[1466] ,
         \DataPath/RF/bus_reg_dataout[1467] ,
         \DataPath/RF/bus_reg_dataout[1468] ,
         \DataPath/RF/bus_reg_dataout[1469] ,
         \DataPath/RF/bus_reg_dataout[1470] ,
         \DataPath/RF/bus_reg_dataout[1471] ,
         \DataPath/RF/bus_reg_dataout[1472] ,
         \DataPath/RF/bus_reg_dataout[1473] ,
         \DataPath/RF/bus_reg_dataout[1474] ,
         \DataPath/RF/bus_reg_dataout[1475] ,
         \DataPath/RF/bus_reg_dataout[1476] ,
         \DataPath/RF/bus_reg_dataout[1477] ,
         \DataPath/RF/bus_reg_dataout[1478] ,
         \DataPath/RF/bus_reg_dataout[1479] ,
         \DataPath/RF/bus_reg_dataout[1480] ,
         \DataPath/RF/bus_reg_dataout[1481] ,
         \DataPath/RF/bus_reg_dataout[1482] ,
         \DataPath/RF/bus_reg_dataout[1483] ,
         \DataPath/RF/bus_reg_dataout[1484] ,
         \DataPath/RF/bus_reg_dataout[1485] ,
         \DataPath/RF/bus_reg_dataout[1486] ,
         \DataPath/RF/bus_reg_dataout[1487] ,
         \DataPath/RF/bus_reg_dataout[1488] ,
         \DataPath/RF/bus_reg_dataout[1489] ,
         \DataPath/RF/bus_reg_dataout[1490] ,
         \DataPath/RF/bus_reg_dataout[1491] ,
         \DataPath/RF/bus_reg_dataout[1492] ,
         \DataPath/RF/bus_reg_dataout[1493] ,
         \DataPath/RF/bus_reg_dataout[1494] ,
         \DataPath/RF/bus_reg_dataout[1495] ,
         \DataPath/RF/bus_reg_dataout[1496] ,
         \DataPath/RF/bus_reg_dataout[1497] ,
         \DataPath/RF/bus_reg_dataout[1498] ,
         \DataPath/RF/bus_reg_dataout[1499] ,
         \DataPath/RF/bus_reg_dataout[1500] ,
         \DataPath/RF/bus_reg_dataout[1501] ,
         \DataPath/RF/bus_reg_dataout[1502] ,
         \DataPath/RF/bus_reg_dataout[1503] ,
         \DataPath/RF/bus_reg_dataout[1504] ,
         \DataPath/RF/bus_reg_dataout[1505] ,
         \DataPath/RF/bus_reg_dataout[1506] ,
         \DataPath/RF/bus_reg_dataout[1507] ,
         \DataPath/RF/bus_reg_dataout[1508] ,
         \DataPath/RF/bus_reg_dataout[1509] ,
         \DataPath/RF/bus_reg_dataout[1510] ,
         \DataPath/RF/bus_reg_dataout[1511] ,
         \DataPath/RF/bus_reg_dataout[1512] ,
         \DataPath/RF/bus_reg_dataout[1513] ,
         \DataPath/RF/bus_reg_dataout[1514] ,
         \DataPath/RF/bus_reg_dataout[1515] ,
         \DataPath/RF/bus_reg_dataout[1516] ,
         \DataPath/RF/bus_reg_dataout[1517] ,
         \DataPath/RF/bus_reg_dataout[1518] ,
         \DataPath/RF/bus_reg_dataout[1519] ,
         \DataPath/RF/bus_reg_dataout[1520] ,
         \DataPath/RF/bus_reg_dataout[1521] ,
         \DataPath/RF/bus_reg_dataout[1522] ,
         \DataPath/RF/bus_reg_dataout[1523] ,
         \DataPath/RF/bus_reg_dataout[1524] ,
         \DataPath/RF/bus_reg_dataout[1525] ,
         \DataPath/RF/bus_reg_dataout[1526] ,
         \DataPath/RF/bus_reg_dataout[1527] ,
         \DataPath/RF/bus_reg_dataout[1528] ,
         \DataPath/RF/bus_reg_dataout[1529] ,
         \DataPath/RF/bus_reg_dataout[1530] ,
         \DataPath/RF/bus_reg_dataout[1531] ,
         \DataPath/RF/bus_reg_dataout[1532] ,
         \DataPath/RF/bus_reg_dataout[1533] ,
         \DataPath/RF/bus_reg_dataout[1534] ,
         \DataPath/RF/bus_reg_dataout[1535] ,
         \DataPath/RF/bus_reg_dataout[1536] ,
         \DataPath/RF/bus_reg_dataout[1537] ,
         \DataPath/RF/bus_reg_dataout[1538] ,
         \DataPath/RF/bus_reg_dataout[1539] ,
         \DataPath/RF/bus_reg_dataout[1540] ,
         \DataPath/RF/bus_reg_dataout[1541] ,
         \DataPath/RF/bus_reg_dataout[1542] ,
         \DataPath/RF/bus_reg_dataout[1543] ,
         \DataPath/RF/bus_reg_dataout[1544] ,
         \DataPath/RF/bus_reg_dataout[1545] ,
         \DataPath/RF/bus_reg_dataout[1546] ,
         \DataPath/RF/bus_reg_dataout[1547] ,
         \DataPath/RF/bus_reg_dataout[1548] ,
         \DataPath/RF/bus_reg_dataout[1549] ,
         \DataPath/RF/bus_reg_dataout[1550] ,
         \DataPath/RF/bus_reg_dataout[1551] ,
         \DataPath/RF/bus_reg_dataout[1552] ,
         \DataPath/RF/bus_reg_dataout[1553] ,
         \DataPath/RF/bus_reg_dataout[1554] ,
         \DataPath/RF/bus_reg_dataout[1555] ,
         \DataPath/RF/bus_reg_dataout[1556] ,
         \DataPath/RF/bus_reg_dataout[1557] ,
         \DataPath/RF/bus_reg_dataout[1558] ,
         \DataPath/RF/bus_reg_dataout[1559] ,
         \DataPath/RF/bus_reg_dataout[1560] ,
         \DataPath/RF/bus_reg_dataout[1561] ,
         \DataPath/RF/bus_reg_dataout[1562] ,
         \DataPath/RF/bus_reg_dataout[1563] ,
         \DataPath/RF/bus_reg_dataout[1564] ,
         \DataPath/RF/bus_reg_dataout[1565] ,
         \DataPath/RF/bus_reg_dataout[1566] ,
         \DataPath/RF/bus_reg_dataout[1567] ,
         \DataPath/RF/bus_reg_dataout[1568] ,
         \DataPath/RF/bus_reg_dataout[1569] ,
         \DataPath/RF/bus_reg_dataout[1570] ,
         \DataPath/RF/bus_reg_dataout[1571] ,
         \DataPath/RF/bus_reg_dataout[1572] ,
         \DataPath/RF/bus_reg_dataout[1573] ,
         \DataPath/RF/bus_reg_dataout[1574] ,
         \DataPath/RF/bus_reg_dataout[1575] ,
         \DataPath/RF/bus_reg_dataout[1576] ,
         \DataPath/RF/bus_reg_dataout[1577] ,
         \DataPath/RF/bus_reg_dataout[1578] ,
         \DataPath/RF/bus_reg_dataout[1579] ,
         \DataPath/RF/bus_reg_dataout[1580] ,
         \DataPath/RF/bus_reg_dataout[1581] ,
         \DataPath/RF/bus_reg_dataout[1582] ,
         \DataPath/RF/bus_reg_dataout[1583] ,
         \DataPath/RF/bus_reg_dataout[1584] ,
         \DataPath/RF/bus_reg_dataout[1585] ,
         \DataPath/RF/bus_reg_dataout[1586] ,
         \DataPath/RF/bus_reg_dataout[1587] ,
         \DataPath/RF/bus_reg_dataout[1588] ,
         \DataPath/RF/bus_reg_dataout[1589] ,
         \DataPath/RF/bus_reg_dataout[1590] ,
         \DataPath/RF/bus_reg_dataout[1591] ,
         \DataPath/RF/bus_reg_dataout[1592] ,
         \DataPath/RF/bus_reg_dataout[1593] ,
         \DataPath/RF/bus_reg_dataout[1594] ,
         \DataPath/RF/bus_reg_dataout[1595] ,
         \DataPath/RF/bus_reg_dataout[1596] ,
         \DataPath/RF/bus_reg_dataout[1597] ,
         \DataPath/RF/bus_reg_dataout[1598] ,
         \DataPath/RF/bus_reg_dataout[1599] ,
         \DataPath/RF/bus_reg_dataout[1600] ,
         \DataPath/RF/bus_reg_dataout[1601] ,
         \DataPath/RF/bus_reg_dataout[1602] ,
         \DataPath/RF/bus_reg_dataout[1603] ,
         \DataPath/RF/bus_reg_dataout[1604] ,
         \DataPath/RF/bus_reg_dataout[1605] ,
         \DataPath/RF/bus_reg_dataout[1606] ,
         \DataPath/RF/bus_reg_dataout[1607] ,
         \DataPath/RF/bus_reg_dataout[1608] ,
         \DataPath/RF/bus_reg_dataout[1609] ,
         \DataPath/RF/bus_reg_dataout[1610] ,
         \DataPath/RF/bus_reg_dataout[1611] ,
         \DataPath/RF/bus_reg_dataout[1612] ,
         \DataPath/RF/bus_reg_dataout[1613] ,
         \DataPath/RF/bus_reg_dataout[1614] ,
         \DataPath/RF/bus_reg_dataout[1615] ,
         \DataPath/RF/bus_reg_dataout[1616] ,
         \DataPath/RF/bus_reg_dataout[1617] ,
         \DataPath/RF/bus_reg_dataout[1618] ,
         \DataPath/RF/bus_reg_dataout[1619] ,
         \DataPath/RF/bus_reg_dataout[1620] ,
         \DataPath/RF/bus_reg_dataout[1621] ,
         \DataPath/RF/bus_reg_dataout[1622] ,
         \DataPath/RF/bus_reg_dataout[1623] ,
         \DataPath/RF/bus_reg_dataout[1624] ,
         \DataPath/RF/bus_reg_dataout[1625] ,
         \DataPath/RF/bus_reg_dataout[1626] ,
         \DataPath/RF/bus_reg_dataout[1627] ,
         \DataPath/RF/bus_reg_dataout[1628] ,
         \DataPath/RF/bus_reg_dataout[1629] ,
         \DataPath/RF/bus_reg_dataout[1630] ,
         \DataPath/RF/bus_reg_dataout[1631] ,
         \DataPath/RF/bus_reg_dataout[1632] ,
         \DataPath/RF/bus_reg_dataout[1633] ,
         \DataPath/RF/bus_reg_dataout[1634] ,
         \DataPath/RF/bus_reg_dataout[1635] ,
         \DataPath/RF/bus_reg_dataout[1636] ,
         \DataPath/RF/bus_reg_dataout[1637] ,
         \DataPath/RF/bus_reg_dataout[1638] ,
         \DataPath/RF/bus_reg_dataout[1639] ,
         \DataPath/RF/bus_reg_dataout[1640] ,
         \DataPath/RF/bus_reg_dataout[1641] ,
         \DataPath/RF/bus_reg_dataout[1642] ,
         \DataPath/RF/bus_reg_dataout[1643] ,
         \DataPath/RF/bus_reg_dataout[1644] ,
         \DataPath/RF/bus_reg_dataout[1645] ,
         \DataPath/RF/bus_reg_dataout[1646] ,
         \DataPath/RF/bus_reg_dataout[1647] ,
         \DataPath/RF/bus_reg_dataout[1648] ,
         \DataPath/RF/bus_reg_dataout[1649] ,
         \DataPath/RF/bus_reg_dataout[1650] ,
         \DataPath/RF/bus_reg_dataout[1651] ,
         \DataPath/RF/bus_reg_dataout[1652] ,
         \DataPath/RF/bus_reg_dataout[1653] ,
         \DataPath/RF/bus_reg_dataout[1654] ,
         \DataPath/RF/bus_reg_dataout[1655] ,
         \DataPath/RF/bus_reg_dataout[1656] ,
         \DataPath/RF/bus_reg_dataout[1657] ,
         \DataPath/RF/bus_reg_dataout[1658] ,
         \DataPath/RF/bus_reg_dataout[1659] ,
         \DataPath/RF/bus_reg_dataout[1660] ,
         \DataPath/RF/bus_reg_dataout[1661] ,
         \DataPath/RF/bus_reg_dataout[1662] ,
         \DataPath/RF/bus_reg_dataout[1663] ,
         \DataPath/RF/bus_reg_dataout[1664] ,
         \DataPath/RF/bus_reg_dataout[1665] ,
         \DataPath/RF/bus_reg_dataout[1666] ,
         \DataPath/RF/bus_reg_dataout[1667] ,
         \DataPath/RF/bus_reg_dataout[1668] ,
         \DataPath/RF/bus_reg_dataout[1669] ,
         \DataPath/RF/bus_reg_dataout[1670] ,
         \DataPath/RF/bus_reg_dataout[1671] ,
         \DataPath/RF/bus_reg_dataout[1672] ,
         \DataPath/RF/bus_reg_dataout[1673] ,
         \DataPath/RF/bus_reg_dataout[1674] ,
         \DataPath/RF/bus_reg_dataout[1675] ,
         \DataPath/RF/bus_reg_dataout[1676] ,
         \DataPath/RF/bus_reg_dataout[1677] ,
         \DataPath/RF/bus_reg_dataout[1678] ,
         \DataPath/RF/bus_reg_dataout[1679] ,
         \DataPath/RF/bus_reg_dataout[1680] ,
         \DataPath/RF/bus_reg_dataout[1681] ,
         \DataPath/RF/bus_reg_dataout[1682] ,
         \DataPath/RF/bus_reg_dataout[1683] ,
         \DataPath/RF/bus_reg_dataout[1684] ,
         \DataPath/RF/bus_reg_dataout[1685] ,
         \DataPath/RF/bus_reg_dataout[1686] ,
         \DataPath/RF/bus_reg_dataout[1687] ,
         \DataPath/RF/bus_reg_dataout[1688] ,
         \DataPath/RF/bus_reg_dataout[1689] ,
         \DataPath/RF/bus_reg_dataout[1690] ,
         \DataPath/RF/bus_reg_dataout[1691] ,
         \DataPath/RF/bus_reg_dataout[1692] ,
         \DataPath/RF/bus_reg_dataout[1693] ,
         \DataPath/RF/bus_reg_dataout[1694] ,
         \DataPath/RF/bus_reg_dataout[1695] ,
         \DataPath/RF/bus_reg_dataout[1696] ,
         \DataPath/RF/bus_reg_dataout[1697] ,
         \DataPath/RF/bus_reg_dataout[1698] ,
         \DataPath/RF/bus_reg_dataout[1699] ,
         \DataPath/RF/bus_reg_dataout[1700] ,
         \DataPath/RF/bus_reg_dataout[1701] ,
         \DataPath/RF/bus_reg_dataout[1702] ,
         \DataPath/RF/bus_reg_dataout[1703] ,
         \DataPath/RF/bus_reg_dataout[1704] ,
         \DataPath/RF/bus_reg_dataout[1705] ,
         \DataPath/RF/bus_reg_dataout[1706] ,
         \DataPath/RF/bus_reg_dataout[1707] ,
         \DataPath/RF/bus_reg_dataout[1708] ,
         \DataPath/RF/bus_reg_dataout[1709] ,
         \DataPath/RF/bus_reg_dataout[1710] ,
         \DataPath/RF/bus_reg_dataout[1711] ,
         \DataPath/RF/bus_reg_dataout[1712] ,
         \DataPath/RF/bus_reg_dataout[1713] ,
         \DataPath/RF/bus_reg_dataout[1714] ,
         \DataPath/RF/bus_reg_dataout[1715] ,
         \DataPath/RF/bus_reg_dataout[1716] ,
         \DataPath/RF/bus_reg_dataout[1717] ,
         \DataPath/RF/bus_reg_dataout[1718] ,
         \DataPath/RF/bus_reg_dataout[1719] ,
         \DataPath/RF/bus_reg_dataout[1720] ,
         \DataPath/RF/bus_reg_dataout[1721] ,
         \DataPath/RF/bus_reg_dataout[1722] ,
         \DataPath/RF/bus_reg_dataout[1723] ,
         \DataPath/RF/bus_reg_dataout[1724] ,
         \DataPath/RF/bus_reg_dataout[1725] ,
         \DataPath/RF/bus_reg_dataout[1726] ,
         \DataPath/RF/bus_reg_dataout[1727] ,
         \DataPath/RF/bus_reg_dataout[1728] ,
         \DataPath/RF/bus_reg_dataout[1729] ,
         \DataPath/RF/bus_reg_dataout[1730] ,
         \DataPath/RF/bus_reg_dataout[1731] ,
         \DataPath/RF/bus_reg_dataout[1732] ,
         \DataPath/RF/bus_reg_dataout[1733] ,
         \DataPath/RF/bus_reg_dataout[1734] ,
         \DataPath/RF/bus_reg_dataout[1735] ,
         \DataPath/RF/bus_reg_dataout[1736] ,
         \DataPath/RF/bus_reg_dataout[1737] ,
         \DataPath/RF/bus_reg_dataout[1738] ,
         \DataPath/RF/bus_reg_dataout[1739] ,
         \DataPath/RF/bus_reg_dataout[1740] ,
         \DataPath/RF/bus_reg_dataout[1741] ,
         \DataPath/RF/bus_reg_dataout[1742] ,
         \DataPath/RF/bus_reg_dataout[1743] ,
         \DataPath/RF/bus_reg_dataout[1744] ,
         \DataPath/RF/bus_reg_dataout[1745] ,
         \DataPath/RF/bus_reg_dataout[1746] ,
         \DataPath/RF/bus_reg_dataout[1747] ,
         \DataPath/RF/bus_reg_dataout[1748] ,
         \DataPath/RF/bus_reg_dataout[1749] ,
         \DataPath/RF/bus_reg_dataout[1750] ,
         \DataPath/RF/bus_reg_dataout[1751] ,
         \DataPath/RF/bus_reg_dataout[1752] ,
         \DataPath/RF/bus_reg_dataout[1753] ,
         \DataPath/RF/bus_reg_dataout[1754] ,
         \DataPath/RF/bus_reg_dataout[1755] ,
         \DataPath/RF/bus_reg_dataout[1756] ,
         \DataPath/RF/bus_reg_dataout[1757] ,
         \DataPath/RF/bus_reg_dataout[1758] ,
         \DataPath/RF/bus_reg_dataout[1759] ,
         \DataPath/RF/bus_reg_dataout[1760] ,
         \DataPath/RF/bus_reg_dataout[1761] ,
         \DataPath/RF/bus_reg_dataout[1762] ,
         \DataPath/RF/bus_reg_dataout[1763] ,
         \DataPath/RF/bus_reg_dataout[1764] ,
         \DataPath/RF/bus_reg_dataout[1765] ,
         \DataPath/RF/bus_reg_dataout[1766] ,
         \DataPath/RF/bus_reg_dataout[1767] ,
         \DataPath/RF/bus_reg_dataout[1768] ,
         \DataPath/RF/bus_reg_dataout[1769] ,
         \DataPath/RF/bus_reg_dataout[1770] ,
         \DataPath/RF/bus_reg_dataout[1771] ,
         \DataPath/RF/bus_reg_dataout[1772] ,
         \DataPath/RF/bus_reg_dataout[1773] ,
         \DataPath/RF/bus_reg_dataout[1774] ,
         \DataPath/RF/bus_reg_dataout[1775] ,
         \DataPath/RF/bus_reg_dataout[1776] ,
         \DataPath/RF/bus_reg_dataout[1777] ,
         \DataPath/RF/bus_reg_dataout[1778] ,
         \DataPath/RF/bus_reg_dataout[1779] ,
         \DataPath/RF/bus_reg_dataout[1780] ,
         \DataPath/RF/bus_reg_dataout[1781] ,
         \DataPath/RF/bus_reg_dataout[1782] ,
         \DataPath/RF/bus_reg_dataout[1783] ,
         \DataPath/RF/bus_reg_dataout[1784] ,
         \DataPath/RF/bus_reg_dataout[1785] ,
         \DataPath/RF/bus_reg_dataout[1786] ,
         \DataPath/RF/bus_reg_dataout[1787] ,
         \DataPath/RF/bus_reg_dataout[1788] ,
         \DataPath/RF/bus_reg_dataout[1789] ,
         \DataPath/RF/bus_reg_dataout[1790] ,
         \DataPath/RF/bus_reg_dataout[1791] ,
         \DataPath/RF/bus_reg_dataout[1792] ,
         \DataPath/RF/bus_reg_dataout[1793] ,
         \DataPath/RF/bus_reg_dataout[1794] ,
         \DataPath/RF/bus_reg_dataout[1795] ,
         \DataPath/RF/bus_reg_dataout[1796] ,
         \DataPath/RF/bus_reg_dataout[1797] ,
         \DataPath/RF/bus_reg_dataout[1798] ,
         \DataPath/RF/bus_reg_dataout[1799] ,
         \DataPath/RF/bus_reg_dataout[1800] ,
         \DataPath/RF/bus_reg_dataout[1801] ,
         \DataPath/RF/bus_reg_dataout[1802] ,
         \DataPath/RF/bus_reg_dataout[1803] ,
         \DataPath/RF/bus_reg_dataout[1804] ,
         \DataPath/RF/bus_reg_dataout[1805] ,
         \DataPath/RF/bus_reg_dataout[1806] ,
         \DataPath/RF/bus_reg_dataout[1807] ,
         \DataPath/RF/bus_reg_dataout[1808] ,
         \DataPath/RF/bus_reg_dataout[1809] ,
         \DataPath/RF/bus_reg_dataout[1810] ,
         \DataPath/RF/bus_reg_dataout[1811] ,
         \DataPath/RF/bus_reg_dataout[1812] ,
         \DataPath/RF/bus_reg_dataout[1813] ,
         \DataPath/RF/bus_reg_dataout[1814] ,
         \DataPath/RF/bus_reg_dataout[1815] ,
         \DataPath/RF/bus_reg_dataout[1816] ,
         \DataPath/RF/bus_reg_dataout[1817] ,
         \DataPath/RF/bus_reg_dataout[1818] ,
         \DataPath/RF/bus_reg_dataout[1819] ,
         \DataPath/RF/bus_reg_dataout[1820] ,
         \DataPath/RF/bus_reg_dataout[1821] ,
         \DataPath/RF/bus_reg_dataout[1822] ,
         \DataPath/RF/bus_reg_dataout[1823] ,
         \DataPath/RF/bus_reg_dataout[1824] ,
         \DataPath/RF/bus_reg_dataout[1825] ,
         \DataPath/RF/bus_reg_dataout[1826] ,
         \DataPath/RF/bus_reg_dataout[1827] ,
         \DataPath/RF/bus_reg_dataout[1828] ,
         \DataPath/RF/bus_reg_dataout[1829] ,
         \DataPath/RF/bus_reg_dataout[1830] ,
         \DataPath/RF/bus_reg_dataout[1831] ,
         \DataPath/RF/bus_reg_dataout[1832] ,
         \DataPath/RF/bus_reg_dataout[1833] ,
         \DataPath/RF/bus_reg_dataout[1834] ,
         \DataPath/RF/bus_reg_dataout[1835] ,
         \DataPath/RF/bus_reg_dataout[1836] ,
         \DataPath/RF/bus_reg_dataout[1837] ,
         \DataPath/RF/bus_reg_dataout[1838] ,
         \DataPath/RF/bus_reg_dataout[1839] ,
         \DataPath/RF/bus_reg_dataout[1840] ,
         \DataPath/RF/bus_reg_dataout[1841] ,
         \DataPath/RF/bus_reg_dataout[1842] ,
         \DataPath/RF/bus_reg_dataout[1843] ,
         \DataPath/RF/bus_reg_dataout[1844] ,
         \DataPath/RF/bus_reg_dataout[1845] ,
         \DataPath/RF/bus_reg_dataout[1846] ,
         \DataPath/RF/bus_reg_dataout[1847] ,
         \DataPath/RF/bus_reg_dataout[1848] ,
         \DataPath/RF/bus_reg_dataout[1849] ,
         \DataPath/RF/bus_reg_dataout[1850] ,
         \DataPath/RF/bus_reg_dataout[1851] ,
         \DataPath/RF/bus_reg_dataout[1852] ,
         \DataPath/RF/bus_reg_dataout[1853] ,
         \DataPath/RF/bus_reg_dataout[1854] ,
         \DataPath/RF/bus_reg_dataout[1855] ,
         \DataPath/RF/bus_reg_dataout[1856] ,
         \DataPath/RF/bus_reg_dataout[1857] ,
         \DataPath/RF/bus_reg_dataout[1858] ,
         \DataPath/RF/bus_reg_dataout[1859] ,
         \DataPath/RF/bus_reg_dataout[1860] ,
         \DataPath/RF/bus_reg_dataout[1861] ,
         \DataPath/RF/bus_reg_dataout[1862] ,
         \DataPath/RF/bus_reg_dataout[1863] ,
         \DataPath/RF/bus_reg_dataout[1864] ,
         \DataPath/RF/bus_reg_dataout[1865] ,
         \DataPath/RF/bus_reg_dataout[1866] ,
         \DataPath/RF/bus_reg_dataout[1867] ,
         \DataPath/RF/bus_reg_dataout[1868] ,
         \DataPath/RF/bus_reg_dataout[1869] ,
         \DataPath/RF/bus_reg_dataout[1870] ,
         \DataPath/RF/bus_reg_dataout[1871] ,
         \DataPath/RF/bus_reg_dataout[1872] ,
         \DataPath/RF/bus_reg_dataout[1873] ,
         \DataPath/RF/bus_reg_dataout[1874] ,
         \DataPath/RF/bus_reg_dataout[1875] ,
         \DataPath/RF/bus_reg_dataout[1876] ,
         \DataPath/RF/bus_reg_dataout[1877] ,
         \DataPath/RF/bus_reg_dataout[1878] ,
         \DataPath/RF/bus_reg_dataout[1879] ,
         \DataPath/RF/bus_reg_dataout[1880] ,
         \DataPath/RF/bus_reg_dataout[1881] ,
         \DataPath/RF/bus_reg_dataout[1882] ,
         \DataPath/RF/bus_reg_dataout[1883] ,
         \DataPath/RF/bus_reg_dataout[1884] ,
         \DataPath/RF/bus_reg_dataout[1885] ,
         \DataPath/RF/bus_reg_dataout[1886] ,
         \DataPath/RF/bus_reg_dataout[1887] ,
         \DataPath/RF/bus_reg_dataout[1888] ,
         \DataPath/RF/bus_reg_dataout[1889] ,
         \DataPath/RF/bus_reg_dataout[1890] ,
         \DataPath/RF/bus_reg_dataout[1891] ,
         \DataPath/RF/bus_reg_dataout[1892] ,
         \DataPath/RF/bus_reg_dataout[1893] ,
         \DataPath/RF/bus_reg_dataout[1894] ,
         \DataPath/RF/bus_reg_dataout[1895] ,
         \DataPath/RF/bus_reg_dataout[1896] ,
         \DataPath/RF/bus_reg_dataout[1897] ,
         \DataPath/RF/bus_reg_dataout[1898] ,
         \DataPath/RF/bus_reg_dataout[1899] ,
         \DataPath/RF/bus_reg_dataout[1900] ,
         \DataPath/RF/bus_reg_dataout[1901] ,
         \DataPath/RF/bus_reg_dataout[1902] ,
         \DataPath/RF/bus_reg_dataout[1903] ,
         \DataPath/RF/bus_reg_dataout[1904] ,
         \DataPath/RF/bus_reg_dataout[1905] ,
         \DataPath/RF/bus_reg_dataout[1906] ,
         \DataPath/RF/bus_reg_dataout[1907] ,
         \DataPath/RF/bus_reg_dataout[1908] ,
         \DataPath/RF/bus_reg_dataout[1909] ,
         \DataPath/RF/bus_reg_dataout[1910] ,
         \DataPath/RF/bus_reg_dataout[1911] ,
         \DataPath/RF/bus_reg_dataout[1912] ,
         \DataPath/RF/bus_reg_dataout[1913] ,
         \DataPath/RF/bus_reg_dataout[1914] ,
         \DataPath/RF/bus_reg_dataout[1915] ,
         \DataPath/RF/bus_reg_dataout[1916] ,
         \DataPath/RF/bus_reg_dataout[1917] ,
         \DataPath/RF/bus_reg_dataout[1918] ,
         \DataPath/RF/bus_reg_dataout[1919] ,
         \DataPath/RF/bus_reg_dataout[1920] ,
         \DataPath/RF/bus_reg_dataout[1921] ,
         \DataPath/RF/bus_reg_dataout[1922] ,
         \DataPath/RF/bus_reg_dataout[1923] ,
         \DataPath/RF/bus_reg_dataout[1924] ,
         \DataPath/RF/bus_reg_dataout[1925] ,
         \DataPath/RF/bus_reg_dataout[1926] ,
         \DataPath/RF/bus_reg_dataout[1927] ,
         \DataPath/RF/bus_reg_dataout[1928] ,
         \DataPath/RF/bus_reg_dataout[1929] ,
         \DataPath/RF/bus_reg_dataout[1930] ,
         \DataPath/RF/bus_reg_dataout[1931] ,
         \DataPath/RF/bus_reg_dataout[1932] ,
         \DataPath/RF/bus_reg_dataout[1933] ,
         \DataPath/RF/bus_reg_dataout[1934] ,
         \DataPath/RF/bus_reg_dataout[1935] ,
         \DataPath/RF/bus_reg_dataout[1936] ,
         \DataPath/RF/bus_reg_dataout[1937] ,
         \DataPath/RF/bus_reg_dataout[1938] ,
         \DataPath/RF/bus_reg_dataout[1939] ,
         \DataPath/RF/bus_reg_dataout[1940] ,
         \DataPath/RF/bus_reg_dataout[1941] ,
         \DataPath/RF/bus_reg_dataout[1942] ,
         \DataPath/RF/bus_reg_dataout[1943] ,
         \DataPath/RF/bus_reg_dataout[1944] ,
         \DataPath/RF/bus_reg_dataout[1945] ,
         \DataPath/RF/bus_reg_dataout[1946] ,
         \DataPath/RF/bus_reg_dataout[1947] ,
         \DataPath/RF/bus_reg_dataout[1948] ,
         \DataPath/RF/bus_reg_dataout[1949] ,
         \DataPath/RF/bus_reg_dataout[1950] ,
         \DataPath/RF/bus_reg_dataout[1951] ,
         \DataPath/RF/bus_reg_dataout[1952] ,
         \DataPath/RF/bus_reg_dataout[1953] ,
         \DataPath/RF/bus_reg_dataout[1954] ,
         \DataPath/RF/bus_reg_dataout[1955] ,
         \DataPath/RF/bus_reg_dataout[1956] ,
         \DataPath/RF/bus_reg_dataout[1957] ,
         \DataPath/RF/bus_reg_dataout[1958] ,
         \DataPath/RF/bus_reg_dataout[1959] ,
         \DataPath/RF/bus_reg_dataout[1960] ,
         \DataPath/RF/bus_reg_dataout[1961] ,
         \DataPath/RF/bus_reg_dataout[1962] ,
         \DataPath/RF/bus_reg_dataout[1963] ,
         \DataPath/RF/bus_reg_dataout[1964] ,
         \DataPath/RF/bus_reg_dataout[1965] ,
         \DataPath/RF/bus_reg_dataout[1966] ,
         \DataPath/RF/bus_reg_dataout[1967] ,
         \DataPath/RF/bus_reg_dataout[1968] ,
         \DataPath/RF/bus_reg_dataout[1969] ,
         \DataPath/RF/bus_reg_dataout[1970] ,
         \DataPath/RF/bus_reg_dataout[1971] ,
         \DataPath/RF/bus_reg_dataout[1972] ,
         \DataPath/RF/bus_reg_dataout[1973] ,
         \DataPath/RF/bus_reg_dataout[1974] ,
         \DataPath/RF/bus_reg_dataout[1975] ,
         \DataPath/RF/bus_reg_dataout[1976] ,
         \DataPath/RF/bus_reg_dataout[1977] ,
         \DataPath/RF/bus_reg_dataout[1978] ,
         \DataPath/RF/bus_reg_dataout[1979] ,
         \DataPath/RF/bus_reg_dataout[1980] ,
         \DataPath/RF/bus_reg_dataout[1981] ,
         \DataPath/RF/bus_reg_dataout[1982] ,
         \DataPath/RF/bus_reg_dataout[1983] ,
         \DataPath/RF/bus_reg_dataout[1984] ,
         \DataPath/RF/bus_reg_dataout[1985] ,
         \DataPath/RF/bus_reg_dataout[1986] ,
         \DataPath/RF/bus_reg_dataout[1987] ,
         \DataPath/RF/bus_reg_dataout[1988] ,
         \DataPath/RF/bus_reg_dataout[1989] ,
         \DataPath/RF/bus_reg_dataout[1990] ,
         \DataPath/RF/bus_reg_dataout[1991] ,
         \DataPath/RF/bus_reg_dataout[1992] ,
         \DataPath/RF/bus_reg_dataout[1993] ,
         \DataPath/RF/bus_reg_dataout[1994] ,
         \DataPath/RF/bus_reg_dataout[1995] ,
         \DataPath/RF/bus_reg_dataout[1996] ,
         \DataPath/RF/bus_reg_dataout[1997] ,
         \DataPath/RF/bus_reg_dataout[1998] ,
         \DataPath/RF/bus_reg_dataout[1999] ,
         \DataPath/RF/bus_reg_dataout[2000] ,
         \DataPath/RF/bus_reg_dataout[2001] ,
         \DataPath/RF/bus_reg_dataout[2002] ,
         \DataPath/RF/bus_reg_dataout[2003] ,
         \DataPath/RF/bus_reg_dataout[2004] ,
         \DataPath/RF/bus_reg_dataout[2005] ,
         \DataPath/RF/bus_reg_dataout[2006] ,
         \DataPath/RF/bus_reg_dataout[2007] ,
         \DataPath/RF/bus_reg_dataout[2008] ,
         \DataPath/RF/bus_reg_dataout[2009] ,
         \DataPath/RF/bus_reg_dataout[2010] ,
         \DataPath/RF/bus_reg_dataout[2011] ,
         \DataPath/RF/bus_reg_dataout[2012] ,
         \DataPath/RF/bus_reg_dataout[2013] ,
         \DataPath/RF/bus_reg_dataout[2014] ,
         \DataPath/RF/bus_reg_dataout[2015] ,
         \DataPath/RF/bus_reg_dataout[2016] ,
         \DataPath/RF/bus_reg_dataout[2017] ,
         \DataPath/RF/bus_reg_dataout[2018] ,
         \DataPath/RF/bus_reg_dataout[2019] ,
         \DataPath/RF/bus_reg_dataout[2020] ,
         \DataPath/RF/bus_reg_dataout[2021] ,
         \DataPath/RF/bus_reg_dataout[2022] ,
         \DataPath/RF/bus_reg_dataout[2023] ,
         \DataPath/RF/bus_reg_dataout[2024] ,
         \DataPath/RF/bus_reg_dataout[2025] ,
         \DataPath/RF/bus_reg_dataout[2026] ,
         \DataPath/RF/bus_reg_dataout[2027] ,
         \DataPath/RF/bus_reg_dataout[2028] ,
         \DataPath/RF/bus_reg_dataout[2029] ,
         \DataPath/RF/bus_reg_dataout[2030] ,
         \DataPath/RF/bus_reg_dataout[2031] ,
         \DataPath/RF/bus_reg_dataout[2032] ,
         \DataPath/RF/bus_reg_dataout[2033] ,
         \DataPath/RF/bus_reg_dataout[2034] ,
         \DataPath/RF/bus_reg_dataout[2035] ,
         \DataPath/RF/bus_reg_dataout[2036] ,
         \DataPath/RF/bus_reg_dataout[2037] ,
         \DataPath/RF/bus_reg_dataout[2038] ,
         \DataPath/RF/bus_reg_dataout[2039] ,
         \DataPath/RF/bus_reg_dataout[2040] ,
         \DataPath/RF/bus_reg_dataout[2041] ,
         \DataPath/RF/bus_reg_dataout[2042] ,
         \DataPath/RF/bus_reg_dataout[2043] ,
         \DataPath/RF/bus_reg_dataout[2044] ,
         \DataPath/RF/bus_reg_dataout[2045] ,
         \DataPath/RF/bus_reg_dataout[2046] ,
         \DataPath/RF/bus_reg_dataout[2047] ,
         \DataPath/RF/bus_reg_dataout[2048] ,
         \DataPath/RF/bus_reg_dataout[2049] ,
         \DataPath/RF/bus_reg_dataout[2050] ,
         \DataPath/RF/bus_reg_dataout[2051] ,
         \DataPath/RF/bus_reg_dataout[2052] ,
         \DataPath/RF/bus_reg_dataout[2053] ,
         \DataPath/RF/bus_reg_dataout[2054] ,
         \DataPath/RF/bus_reg_dataout[2055] ,
         \DataPath/RF/bus_reg_dataout[2056] ,
         \DataPath/RF/bus_reg_dataout[2057] ,
         \DataPath/RF/bus_reg_dataout[2058] ,
         \DataPath/RF/bus_reg_dataout[2059] ,
         \DataPath/RF/bus_reg_dataout[2060] ,
         \DataPath/RF/bus_reg_dataout[2061] ,
         \DataPath/RF/bus_reg_dataout[2062] ,
         \DataPath/RF/bus_reg_dataout[2063] ,
         \DataPath/RF/bus_reg_dataout[2064] ,
         \DataPath/RF/bus_reg_dataout[2065] ,
         \DataPath/RF/bus_reg_dataout[2066] ,
         \DataPath/RF/bus_reg_dataout[2067] ,
         \DataPath/RF/bus_reg_dataout[2068] ,
         \DataPath/RF/bus_reg_dataout[2069] ,
         \DataPath/RF/bus_reg_dataout[2070] ,
         \DataPath/RF/bus_reg_dataout[2071] ,
         \DataPath/RF/bus_reg_dataout[2072] ,
         \DataPath/RF/bus_reg_dataout[2073] ,
         \DataPath/RF/bus_reg_dataout[2074] ,
         \DataPath/RF/bus_reg_dataout[2075] ,
         \DataPath/RF/bus_reg_dataout[2076] ,
         \DataPath/RF/bus_reg_dataout[2077] ,
         \DataPath/RF/bus_reg_dataout[2078] ,
         \DataPath/RF/bus_reg_dataout[2079] ,
         \DataPath/RF/bus_reg_dataout[2080] ,
         \DataPath/RF/bus_reg_dataout[2081] ,
         \DataPath/RF/bus_reg_dataout[2082] ,
         \DataPath/RF/bus_reg_dataout[2083] ,
         \DataPath/RF/bus_reg_dataout[2084] ,
         \DataPath/RF/bus_reg_dataout[2085] ,
         \DataPath/RF/bus_reg_dataout[2086] ,
         \DataPath/RF/bus_reg_dataout[2087] ,
         \DataPath/RF/bus_reg_dataout[2088] ,
         \DataPath/RF/bus_reg_dataout[2089] ,
         \DataPath/RF/bus_reg_dataout[2090] ,
         \DataPath/RF/bus_reg_dataout[2091] ,
         \DataPath/RF/bus_reg_dataout[2092] ,
         \DataPath/RF/bus_reg_dataout[2093] ,
         \DataPath/RF/bus_reg_dataout[2094] ,
         \DataPath/RF/bus_reg_dataout[2095] ,
         \DataPath/RF/bus_reg_dataout[2096] ,
         \DataPath/RF/bus_reg_dataout[2097] ,
         \DataPath/RF/bus_reg_dataout[2098] ,
         \DataPath/RF/bus_reg_dataout[2099] ,
         \DataPath/RF/bus_reg_dataout[2100] ,
         \DataPath/RF/bus_reg_dataout[2101] ,
         \DataPath/RF/bus_reg_dataout[2102] ,
         \DataPath/RF/bus_reg_dataout[2103] ,
         \DataPath/RF/bus_reg_dataout[2104] ,
         \DataPath/RF/bus_reg_dataout[2105] ,
         \DataPath/RF/bus_reg_dataout[2106] ,
         \DataPath/RF/bus_reg_dataout[2107] ,
         \DataPath/RF/bus_reg_dataout[2108] ,
         \DataPath/RF/bus_reg_dataout[2109] ,
         \DataPath/RF/bus_reg_dataout[2110] ,
         \DataPath/RF/bus_reg_dataout[2111] ,
         \DataPath/RF/bus_reg_dataout[2112] ,
         \DataPath/RF/bus_reg_dataout[2113] ,
         \DataPath/RF/bus_reg_dataout[2114] ,
         \DataPath/RF/bus_reg_dataout[2115] ,
         \DataPath/RF/bus_reg_dataout[2116] ,
         \DataPath/RF/bus_reg_dataout[2117] ,
         \DataPath/RF/bus_reg_dataout[2118] ,
         \DataPath/RF/bus_reg_dataout[2119] ,
         \DataPath/RF/bus_reg_dataout[2120] ,
         \DataPath/RF/bus_reg_dataout[2121] ,
         \DataPath/RF/bus_reg_dataout[2122] ,
         \DataPath/RF/bus_reg_dataout[2123] ,
         \DataPath/RF/bus_reg_dataout[2124] ,
         \DataPath/RF/bus_reg_dataout[2125] ,
         \DataPath/RF/bus_reg_dataout[2126] ,
         \DataPath/RF/bus_reg_dataout[2127] ,
         \DataPath/RF/bus_reg_dataout[2128] ,
         \DataPath/RF/bus_reg_dataout[2129] ,
         \DataPath/RF/bus_reg_dataout[2130] ,
         \DataPath/RF/bus_reg_dataout[2131] ,
         \DataPath/RF/bus_reg_dataout[2132] ,
         \DataPath/RF/bus_reg_dataout[2133] ,
         \DataPath/RF/bus_reg_dataout[2134] ,
         \DataPath/RF/bus_reg_dataout[2135] ,
         \DataPath/RF/bus_reg_dataout[2136] ,
         \DataPath/RF/bus_reg_dataout[2137] ,
         \DataPath/RF/bus_reg_dataout[2138] ,
         \DataPath/RF/bus_reg_dataout[2139] ,
         \DataPath/RF/bus_reg_dataout[2140] ,
         \DataPath/RF/bus_reg_dataout[2141] ,
         \DataPath/RF/bus_reg_dataout[2142] ,
         \DataPath/RF/bus_reg_dataout[2143] ,
         \DataPath/RF/bus_reg_dataout[2144] ,
         \DataPath/RF/bus_reg_dataout[2145] ,
         \DataPath/RF/bus_reg_dataout[2146] ,
         \DataPath/RF/bus_reg_dataout[2147] ,
         \DataPath/RF/bus_reg_dataout[2148] ,
         \DataPath/RF/bus_reg_dataout[2149] ,
         \DataPath/RF/bus_reg_dataout[2150] ,
         \DataPath/RF/bus_reg_dataout[2151] ,
         \DataPath/RF/bus_reg_dataout[2152] ,
         \DataPath/RF/bus_reg_dataout[2153] ,
         \DataPath/RF/bus_reg_dataout[2154] ,
         \DataPath/RF/bus_reg_dataout[2155] ,
         \DataPath/RF/bus_reg_dataout[2156] ,
         \DataPath/RF/bus_reg_dataout[2157] ,
         \DataPath/RF/bus_reg_dataout[2158] ,
         \DataPath/RF/bus_reg_dataout[2159] ,
         \DataPath/RF/bus_reg_dataout[2160] ,
         \DataPath/RF/bus_reg_dataout[2161] ,
         \DataPath/RF/bus_reg_dataout[2162] ,
         \DataPath/RF/bus_reg_dataout[2163] ,
         \DataPath/RF/bus_reg_dataout[2164] ,
         \DataPath/RF/bus_reg_dataout[2165] ,
         \DataPath/RF/bus_reg_dataout[2166] ,
         \DataPath/RF/bus_reg_dataout[2167] ,
         \DataPath/RF/bus_reg_dataout[2168] ,
         \DataPath/RF/bus_reg_dataout[2169] ,
         \DataPath/RF/bus_reg_dataout[2170] ,
         \DataPath/RF/bus_reg_dataout[2171] ,
         \DataPath/RF/bus_reg_dataout[2172] ,
         \DataPath/RF/bus_reg_dataout[2173] ,
         \DataPath/RF/bus_reg_dataout[2174] ,
         \DataPath/RF/bus_reg_dataout[2175] ,
         \DataPath/RF/bus_reg_dataout[2176] ,
         \DataPath/RF/bus_reg_dataout[2177] ,
         \DataPath/RF/bus_reg_dataout[2178] ,
         \DataPath/RF/bus_reg_dataout[2179] ,
         \DataPath/RF/bus_reg_dataout[2180] ,
         \DataPath/RF/bus_reg_dataout[2181] ,
         \DataPath/RF/bus_reg_dataout[2182] ,
         \DataPath/RF/bus_reg_dataout[2183] ,
         \DataPath/RF/bus_reg_dataout[2184] ,
         \DataPath/RF/bus_reg_dataout[2185] ,
         \DataPath/RF/bus_reg_dataout[2186] ,
         \DataPath/RF/bus_reg_dataout[2187] ,
         \DataPath/RF/bus_reg_dataout[2188] ,
         \DataPath/RF/bus_reg_dataout[2189] ,
         \DataPath/RF/bus_reg_dataout[2190] ,
         \DataPath/RF/bus_reg_dataout[2191] ,
         \DataPath/RF/bus_reg_dataout[2192] ,
         \DataPath/RF/bus_reg_dataout[2193] ,
         \DataPath/RF/bus_reg_dataout[2194] ,
         \DataPath/RF/bus_reg_dataout[2195] ,
         \DataPath/RF/bus_reg_dataout[2196] ,
         \DataPath/RF/bus_reg_dataout[2197] ,
         \DataPath/RF/bus_reg_dataout[2198] ,
         \DataPath/RF/bus_reg_dataout[2199] ,
         \DataPath/RF/bus_reg_dataout[2200] ,
         \DataPath/RF/bus_reg_dataout[2201] ,
         \DataPath/RF/bus_reg_dataout[2202] ,
         \DataPath/RF/bus_reg_dataout[2203] ,
         \DataPath/RF/bus_reg_dataout[2204] ,
         \DataPath/RF/bus_reg_dataout[2205] ,
         \DataPath/RF/bus_reg_dataout[2206] ,
         \DataPath/RF/bus_reg_dataout[2207] ,
         \DataPath/RF/bus_reg_dataout[2208] ,
         \DataPath/RF/bus_reg_dataout[2209] ,
         \DataPath/RF/bus_reg_dataout[2210] ,
         \DataPath/RF/bus_reg_dataout[2211] ,
         \DataPath/RF/bus_reg_dataout[2212] ,
         \DataPath/RF/bus_reg_dataout[2213] ,
         \DataPath/RF/bus_reg_dataout[2214] ,
         \DataPath/RF/bus_reg_dataout[2215] ,
         \DataPath/RF/bus_reg_dataout[2216] ,
         \DataPath/RF/bus_reg_dataout[2217] ,
         \DataPath/RF/bus_reg_dataout[2218] ,
         \DataPath/RF/bus_reg_dataout[2219] ,
         \DataPath/RF/bus_reg_dataout[2220] ,
         \DataPath/RF/bus_reg_dataout[2221] ,
         \DataPath/RF/bus_reg_dataout[2222] ,
         \DataPath/RF/bus_reg_dataout[2223] ,
         \DataPath/RF/bus_reg_dataout[2224] ,
         \DataPath/RF/bus_reg_dataout[2225] ,
         \DataPath/RF/bus_reg_dataout[2226] ,
         \DataPath/RF/bus_reg_dataout[2227] ,
         \DataPath/RF/bus_reg_dataout[2228] ,
         \DataPath/RF/bus_reg_dataout[2229] ,
         \DataPath/RF/bus_reg_dataout[2230] ,
         \DataPath/RF/bus_reg_dataout[2231] ,
         \DataPath/RF/bus_reg_dataout[2232] ,
         \DataPath/RF/bus_reg_dataout[2233] ,
         \DataPath/RF/bus_reg_dataout[2234] ,
         \DataPath/RF/bus_reg_dataout[2235] ,
         \DataPath/RF/bus_reg_dataout[2236] ,
         \DataPath/RF/bus_reg_dataout[2237] ,
         \DataPath/RF/bus_reg_dataout[2238] ,
         \DataPath/RF/bus_reg_dataout[2239] ,
         \DataPath/RF/bus_reg_dataout[2240] ,
         \DataPath/RF/bus_reg_dataout[2241] ,
         \DataPath/RF/bus_reg_dataout[2242] ,
         \DataPath/RF/bus_reg_dataout[2243] ,
         \DataPath/RF/bus_reg_dataout[2244] ,
         \DataPath/RF/bus_reg_dataout[2245] ,
         \DataPath/RF/bus_reg_dataout[2246] ,
         \DataPath/RF/bus_reg_dataout[2247] ,
         \DataPath/RF/bus_reg_dataout[2248] ,
         \DataPath/RF/bus_reg_dataout[2249] ,
         \DataPath/RF/bus_reg_dataout[2250] ,
         \DataPath/RF/bus_reg_dataout[2251] ,
         \DataPath/RF/bus_reg_dataout[2252] ,
         \DataPath/RF/bus_reg_dataout[2253] ,
         \DataPath/RF/bus_reg_dataout[2254] ,
         \DataPath/RF/bus_reg_dataout[2255] ,
         \DataPath/RF/bus_reg_dataout[2256] ,
         \DataPath/RF/bus_reg_dataout[2257] ,
         \DataPath/RF/bus_reg_dataout[2258] ,
         \DataPath/RF/bus_reg_dataout[2259] ,
         \DataPath/RF/bus_reg_dataout[2260] ,
         \DataPath/RF/bus_reg_dataout[2261] ,
         \DataPath/RF/bus_reg_dataout[2262] ,
         \DataPath/RF/bus_reg_dataout[2263] ,
         \DataPath/RF/bus_reg_dataout[2264] ,
         \DataPath/RF/bus_reg_dataout[2265] ,
         \DataPath/RF/bus_reg_dataout[2266] ,
         \DataPath/RF/bus_reg_dataout[2267] ,
         \DataPath/RF/bus_reg_dataout[2268] ,
         \DataPath/RF/bus_reg_dataout[2269] ,
         \DataPath/RF/bus_reg_dataout[2270] ,
         \DataPath/RF/bus_reg_dataout[2271] ,
         \DataPath/RF/bus_reg_dataout[2272] ,
         \DataPath/RF/bus_reg_dataout[2273] ,
         \DataPath/RF/bus_reg_dataout[2274] ,
         \DataPath/RF/bus_reg_dataout[2275] ,
         \DataPath/RF/bus_reg_dataout[2276] ,
         \DataPath/RF/bus_reg_dataout[2277] ,
         \DataPath/RF/bus_reg_dataout[2278] ,
         \DataPath/RF/bus_reg_dataout[2279] ,
         \DataPath/RF/bus_reg_dataout[2280] ,
         \DataPath/RF/bus_reg_dataout[2281] ,
         \DataPath/RF/bus_reg_dataout[2282] ,
         \DataPath/RF/bus_reg_dataout[2283] ,
         \DataPath/RF/bus_reg_dataout[2284] ,
         \DataPath/RF/bus_reg_dataout[2285] ,
         \DataPath/RF/bus_reg_dataout[2286] ,
         \DataPath/RF/bus_reg_dataout[2287] ,
         \DataPath/RF/bus_reg_dataout[2288] ,
         \DataPath/RF/bus_reg_dataout[2289] ,
         \DataPath/RF/bus_reg_dataout[2290] ,
         \DataPath/RF/bus_reg_dataout[2291] ,
         \DataPath/RF/bus_reg_dataout[2292] ,
         \DataPath/RF/bus_reg_dataout[2293] ,
         \DataPath/RF/bus_reg_dataout[2294] ,
         \DataPath/RF/bus_reg_dataout[2295] ,
         \DataPath/RF/bus_reg_dataout[2296] ,
         \DataPath/RF/bus_reg_dataout[2297] ,
         \DataPath/RF/bus_reg_dataout[2298] ,
         \DataPath/RF/bus_reg_dataout[2299] ,
         \DataPath/RF/bus_reg_dataout[2300] ,
         \DataPath/RF/bus_reg_dataout[2301] ,
         \DataPath/RF/bus_reg_dataout[2302] ,
         \DataPath/RF/bus_reg_dataout[2303] ,
         \DataPath/RF/bus_reg_dataout[2304] ,
         \DataPath/RF/bus_reg_dataout[2305] ,
         \DataPath/RF/bus_reg_dataout[2306] ,
         \DataPath/RF/bus_reg_dataout[2307] ,
         \DataPath/RF/bus_reg_dataout[2308] ,
         \DataPath/RF/bus_reg_dataout[2309] ,
         \DataPath/RF/bus_reg_dataout[2310] ,
         \DataPath/RF/bus_reg_dataout[2311] ,
         \DataPath/RF/bus_reg_dataout[2312] ,
         \DataPath/RF/bus_reg_dataout[2313] ,
         \DataPath/RF/bus_reg_dataout[2314] ,
         \DataPath/RF/bus_reg_dataout[2315] ,
         \DataPath/RF/bus_reg_dataout[2316] ,
         \DataPath/RF/bus_reg_dataout[2317] ,
         \DataPath/RF/bus_reg_dataout[2318] ,
         \DataPath/RF/bus_reg_dataout[2319] ,
         \DataPath/RF/bus_reg_dataout[2320] ,
         \DataPath/RF/bus_reg_dataout[2321] ,
         \DataPath/RF/bus_reg_dataout[2322] ,
         \DataPath/RF/bus_reg_dataout[2323] ,
         \DataPath/RF/bus_reg_dataout[2324] ,
         \DataPath/RF/bus_reg_dataout[2325] ,
         \DataPath/RF/bus_reg_dataout[2326] ,
         \DataPath/RF/bus_reg_dataout[2327] ,
         \DataPath/RF/bus_reg_dataout[2328] ,
         \DataPath/RF/bus_reg_dataout[2329] ,
         \DataPath/RF/bus_reg_dataout[2330] ,
         \DataPath/RF/bus_reg_dataout[2331] ,
         \DataPath/RF/bus_reg_dataout[2332] ,
         \DataPath/RF/bus_reg_dataout[2333] ,
         \DataPath/RF/bus_reg_dataout[2334] ,
         \DataPath/RF/bus_reg_dataout[2335] ,
         \DataPath/RF/bus_reg_dataout[2336] ,
         \DataPath/RF/bus_reg_dataout[2337] ,
         \DataPath/RF/bus_reg_dataout[2338] ,
         \DataPath/RF/bus_reg_dataout[2339] ,
         \DataPath/RF/bus_reg_dataout[2340] ,
         \DataPath/RF/bus_reg_dataout[2341] ,
         \DataPath/RF/bus_reg_dataout[2342] ,
         \DataPath/RF/bus_reg_dataout[2343] ,
         \DataPath/RF/bus_reg_dataout[2344] ,
         \DataPath/RF/bus_reg_dataout[2345] ,
         \DataPath/RF/bus_reg_dataout[2346] ,
         \DataPath/RF/bus_reg_dataout[2347] ,
         \DataPath/RF/bus_reg_dataout[2348] ,
         \DataPath/RF/bus_reg_dataout[2349] ,
         \DataPath/RF/bus_reg_dataout[2350] ,
         \DataPath/RF/bus_reg_dataout[2351] ,
         \DataPath/RF/bus_reg_dataout[2352] ,
         \DataPath/RF/bus_reg_dataout[2353] ,
         \DataPath/RF/bus_reg_dataout[2354] ,
         \DataPath/RF/bus_reg_dataout[2355] ,
         \DataPath/RF/bus_reg_dataout[2356] ,
         \DataPath/RF/bus_reg_dataout[2357] ,
         \DataPath/RF/bus_reg_dataout[2358] ,
         \DataPath/RF/bus_reg_dataout[2359] ,
         \DataPath/RF/bus_reg_dataout[2360] ,
         \DataPath/RF/bus_reg_dataout[2361] ,
         \DataPath/RF/bus_reg_dataout[2362] ,
         \DataPath/RF/bus_reg_dataout[2363] ,
         \DataPath/RF/bus_reg_dataout[2364] ,
         \DataPath/RF/bus_reg_dataout[2365] ,
         \DataPath/RF/bus_reg_dataout[2366] ,
         \DataPath/RF/bus_reg_dataout[2367] ,
         \DataPath/RF/bus_reg_dataout[2368] ,
         \DataPath/RF/bus_reg_dataout[2369] ,
         \DataPath/RF/bus_reg_dataout[2370] ,
         \DataPath/RF/bus_reg_dataout[2371] ,
         \DataPath/RF/bus_reg_dataout[2372] ,
         \DataPath/RF/bus_reg_dataout[2373] ,
         \DataPath/RF/bus_reg_dataout[2374] ,
         \DataPath/RF/bus_reg_dataout[2375] ,
         \DataPath/RF/bus_reg_dataout[2376] ,
         \DataPath/RF/bus_reg_dataout[2377] ,
         \DataPath/RF/bus_reg_dataout[2378] ,
         \DataPath/RF/bus_reg_dataout[2379] ,
         \DataPath/RF/bus_reg_dataout[2380] ,
         \DataPath/RF/bus_reg_dataout[2381] ,
         \DataPath/RF/bus_reg_dataout[2382] ,
         \DataPath/RF/bus_reg_dataout[2383] ,
         \DataPath/RF/bus_reg_dataout[2384] ,
         \DataPath/RF/bus_reg_dataout[2385] ,
         \DataPath/RF/bus_reg_dataout[2386] ,
         \DataPath/RF/bus_reg_dataout[2387] ,
         \DataPath/RF/bus_reg_dataout[2388] ,
         \DataPath/RF/bus_reg_dataout[2389] ,
         \DataPath/RF/bus_reg_dataout[2390] ,
         \DataPath/RF/bus_reg_dataout[2391] ,
         \DataPath/RF/bus_reg_dataout[2392] ,
         \DataPath/RF/bus_reg_dataout[2393] ,
         \DataPath/RF/bus_reg_dataout[2394] ,
         \DataPath/RF/bus_reg_dataout[2395] ,
         \DataPath/RF/bus_reg_dataout[2396] ,
         \DataPath/RF/bus_reg_dataout[2397] ,
         \DataPath/RF/bus_reg_dataout[2398] ,
         \DataPath/RF/bus_reg_dataout[2399] ,
         \DataPath/RF/bus_reg_dataout[2400] ,
         \DataPath/RF/bus_reg_dataout[2401] ,
         \DataPath/RF/bus_reg_dataout[2402] ,
         \DataPath/RF/bus_reg_dataout[2403] ,
         \DataPath/RF/bus_reg_dataout[2404] ,
         \DataPath/RF/bus_reg_dataout[2405] ,
         \DataPath/RF/bus_reg_dataout[2406] ,
         \DataPath/RF/bus_reg_dataout[2407] ,
         \DataPath/RF/bus_reg_dataout[2408] ,
         \DataPath/RF/bus_reg_dataout[2409] ,
         \DataPath/RF/bus_reg_dataout[2410] ,
         \DataPath/RF/bus_reg_dataout[2411] ,
         \DataPath/RF/bus_reg_dataout[2412] ,
         \DataPath/RF/bus_reg_dataout[2413] ,
         \DataPath/RF/bus_reg_dataout[2414] ,
         \DataPath/RF/bus_reg_dataout[2415] ,
         \DataPath/RF/bus_reg_dataout[2416] ,
         \DataPath/RF/bus_reg_dataout[2417] ,
         \DataPath/RF/bus_reg_dataout[2418] ,
         \DataPath/RF/bus_reg_dataout[2419] ,
         \DataPath/RF/bus_reg_dataout[2420] ,
         \DataPath/RF/bus_reg_dataout[2421] ,
         \DataPath/RF/bus_reg_dataout[2422] ,
         \DataPath/RF/bus_reg_dataout[2423] ,
         \DataPath/RF/bus_reg_dataout[2424] ,
         \DataPath/RF/bus_reg_dataout[2425] ,
         \DataPath/RF/bus_reg_dataout[2426] ,
         \DataPath/RF/bus_reg_dataout[2427] ,
         \DataPath/RF/bus_reg_dataout[2428] ,
         \DataPath/RF/bus_reg_dataout[2429] ,
         \DataPath/RF/bus_reg_dataout[2430] ,
         \DataPath/RF/bus_reg_dataout[2431] ,
         \DataPath/RF/bus_reg_dataout[2432] ,
         \DataPath/RF/bus_reg_dataout[2433] ,
         \DataPath/RF/bus_reg_dataout[2434] ,
         \DataPath/RF/bus_reg_dataout[2435] ,
         \DataPath/RF/bus_reg_dataout[2436] ,
         \DataPath/RF/bus_reg_dataout[2437] ,
         \DataPath/RF/bus_reg_dataout[2438] ,
         \DataPath/RF/bus_reg_dataout[2439] ,
         \DataPath/RF/bus_reg_dataout[2440] ,
         \DataPath/RF/bus_reg_dataout[2441] ,
         \DataPath/RF/bus_reg_dataout[2442] ,
         \DataPath/RF/bus_reg_dataout[2443] ,
         \DataPath/RF/bus_reg_dataout[2444] ,
         \DataPath/RF/bus_reg_dataout[2445] ,
         \DataPath/RF/bus_reg_dataout[2446] ,
         \DataPath/RF/bus_reg_dataout[2447] ,
         \DataPath/RF/bus_reg_dataout[2448] ,
         \DataPath/RF/bus_reg_dataout[2449] ,
         \DataPath/RF/bus_reg_dataout[2450] ,
         \DataPath/RF/bus_reg_dataout[2451] ,
         \DataPath/RF/bus_reg_dataout[2452] ,
         \DataPath/RF/bus_reg_dataout[2453] ,
         \DataPath/RF/bus_reg_dataout[2454] ,
         \DataPath/RF/bus_reg_dataout[2455] ,
         \DataPath/RF/bus_reg_dataout[2456] ,
         \DataPath/RF/bus_reg_dataout[2457] ,
         \DataPath/RF/bus_reg_dataout[2458] ,
         \DataPath/RF/bus_reg_dataout[2459] ,
         \DataPath/RF/bus_reg_dataout[2460] ,
         \DataPath/RF/bus_reg_dataout[2461] ,
         \DataPath/RF/bus_reg_dataout[2462] ,
         \DataPath/RF/bus_reg_dataout[2463] ,
         \DataPath/RF/bus_reg_dataout[2464] ,
         \DataPath/RF/bus_reg_dataout[2465] ,
         \DataPath/RF/bus_reg_dataout[2466] ,
         \DataPath/RF/bus_reg_dataout[2467] ,
         \DataPath/RF/bus_reg_dataout[2468] ,
         \DataPath/RF/bus_reg_dataout[2469] ,
         \DataPath/RF/bus_reg_dataout[2470] ,
         \DataPath/RF/bus_reg_dataout[2471] ,
         \DataPath/RF/bus_reg_dataout[2472] ,
         \DataPath/RF/bus_reg_dataout[2473] ,
         \DataPath/RF/bus_reg_dataout[2474] ,
         \DataPath/RF/bus_reg_dataout[2475] ,
         \DataPath/RF/bus_reg_dataout[2476] ,
         \DataPath/RF/bus_reg_dataout[2477] ,
         \DataPath/RF/bus_reg_dataout[2478] ,
         \DataPath/RF/bus_reg_dataout[2479] ,
         \DataPath/RF/bus_reg_dataout[2480] ,
         \DataPath/RF/bus_reg_dataout[2481] ,
         \DataPath/RF/bus_reg_dataout[2482] ,
         \DataPath/RF/bus_reg_dataout[2483] ,
         \DataPath/RF/bus_reg_dataout[2484] ,
         \DataPath/RF/bus_reg_dataout[2485] ,
         \DataPath/RF/bus_reg_dataout[2486] ,
         \DataPath/RF/bus_reg_dataout[2487] ,
         \DataPath/RF/bus_reg_dataout[2488] ,
         \DataPath/RF/bus_reg_dataout[2489] ,
         \DataPath/RF/bus_reg_dataout[2490] ,
         \DataPath/RF/bus_reg_dataout[2491] ,
         \DataPath/RF/bus_reg_dataout[2492] ,
         \DataPath/RF/bus_reg_dataout[2493] ,
         \DataPath/RF/bus_reg_dataout[2494] ,
         \DataPath/RF/bus_reg_dataout[2495] ,
         \DataPath/RF/bus_reg_dataout[2496] ,
         \DataPath/RF/bus_reg_dataout[2497] ,
         \DataPath/RF/bus_reg_dataout[2498] ,
         \DataPath/RF/bus_reg_dataout[2499] ,
         \DataPath/RF/bus_reg_dataout[2500] ,
         \DataPath/RF/bus_reg_dataout[2501] ,
         \DataPath/RF/bus_reg_dataout[2502] ,
         \DataPath/RF/bus_reg_dataout[2503] ,
         \DataPath/RF/bus_reg_dataout[2504] ,
         \DataPath/RF/bus_reg_dataout[2505] ,
         \DataPath/RF/bus_reg_dataout[2506] ,
         \DataPath/RF/bus_reg_dataout[2507] ,
         \DataPath/RF/bus_reg_dataout[2508] ,
         \DataPath/RF/bus_reg_dataout[2509] ,
         \DataPath/RF/bus_reg_dataout[2510] ,
         \DataPath/RF/bus_reg_dataout[2511] ,
         \DataPath/RF/bus_reg_dataout[2512] ,
         \DataPath/RF/bus_reg_dataout[2513] ,
         \DataPath/RF/bus_reg_dataout[2514] ,
         \DataPath/RF/bus_reg_dataout[2515] ,
         \DataPath/RF/bus_reg_dataout[2516] ,
         \DataPath/RF/bus_reg_dataout[2517] ,
         \DataPath/RF/bus_reg_dataout[2518] ,
         \DataPath/RF/bus_reg_dataout[2519] ,
         \DataPath/RF/bus_reg_dataout[2520] ,
         \DataPath/RF/bus_reg_dataout[2521] ,
         \DataPath/RF/bus_reg_dataout[2522] ,
         \DataPath/RF/bus_reg_dataout[2523] ,
         \DataPath/RF/bus_reg_dataout[2524] ,
         \DataPath/RF/bus_reg_dataout[2525] ,
         \DataPath/RF/bus_reg_dataout[2526] ,
         \DataPath/RF/bus_reg_dataout[2527] ,
         \DataPath/RF/bus_reg_dataout[2528] ,
         \DataPath/RF/bus_reg_dataout[2529] ,
         \DataPath/RF/bus_reg_dataout[2530] ,
         \DataPath/RF/bus_reg_dataout[2531] ,
         \DataPath/RF/bus_reg_dataout[2532] ,
         \DataPath/RF/bus_reg_dataout[2533] ,
         \DataPath/RF/bus_reg_dataout[2534] ,
         \DataPath/RF/bus_reg_dataout[2535] ,
         \DataPath/RF/bus_reg_dataout[2536] ,
         \DataPath/RF/bus_reg_dataout[2537] ,
         \DataPath/RF/bus_reg_dataout[2538] ,
         \DataPath/RF/bus_reg_dataout[2539] ,
         \DataPath/RF/bus_reg_dataout[2540] ,
         \DataPath/RF/bus_reg_dataout[2541] ,
         \DataPath/RF/bus_reg_dataout[2542] ,
         \DataPath/RF/bus_reg_dataout[2543] ,
         \DataPath/RF/bus_reg_dataout[2544] ,
         \DataPath/RF/bus_reg_dataout[2545] ,
         \DataPath/RF/bus_reg_dataout[2546] ,
         \DataPath/RF/bus_reg_dataout[2547] ,
         \DataPath/RF/bus_reg_dataout[2548] ,
         \DataPath/RF/bus_reg_dataout[2549] ,
         \DataPath/RF/bus_reg_dataout[2550] ,
         \DataPath/RF/bus_reg_dataout[2551] ,
         \DataPath/RF/bus_reg_dataout[2552] ,
         \DataPath/RF/bus_reg_dataout[2553] ,
         \DataPath/RF/bus_reg_dataout[2554] ,
         \DataPath/RF/bus_reg_dataout[2555] ,
         \DataPath/RF/bus_reg_dataout[2556] ,
         \DataPath/RF/bus_reg_dataout[2557] ,
         \DataPath/RF/bus_reg_dataout[2558] ,
         \DataPath/RF/bus_reg_dataout[2559] , \DataPath/RF/c_win[0] ,
         \DataPath/RF/c_win[1] , \DataPath/RF/c_win[2] ,
         \DataPath/RF/c_win[3] , \DataPath/WRF_CUhw/N145 ,
         \DataPath/WRF_CUhw/curr_addr[2] , \DataPath/WRF_CUhw/curr_addr[3] ,
         \DataPath/WRF_CUhw/curr_addr[4] , \DataPath/WRF_CUhw/curr_addr[5] ,
         \DataPath/WRF_CUhw/curr_addr[6] , \DataPath/WRF_CUhw/curr_addr[7] ,
         \DataPath/WRF_CUhw/curr_addr[8] , \DataPath/WRF_CUhw/curr_addr[9] ,
         \DataPath/WRF_CUhw/curr_addr[10] , \DataPath/WRF_CUhw/curr_addr[11] ,
         \DataPath/WRF_CUhw/curr_addr[12] , \DataPath/WRF_CUhw/curr_addr[13] ,
         \DataPath/WRF_CUhw/curr_addr[14] , \DataPath/WRF_CUhw/curr_addr[15] ,
         \DataPath/WRF_CUhw/curr_addr[16] , \DataPath/WRF_CUhw/curr_addr[17] ,
         \DataPath/WRF_CUhw/curr_addr[18] , \DataPath/WRF_CUhw/curr_addr[19] ,
         \DataPath/WRF_CUhw/curr_addr[20] , \DataPath/WRF_CUhw/curr_addr[21] ,
         \DataPath/WRF_CUhw/curr_addr[22] , \DataPath/WRF_CUhw/curr_addr[23] ,
         \DataPath/WRF_CUhw/curr_addr[24] , \DataPath/WRF_CUhw/curr_addr[25] ,
         \DataPath/WRF_CUhw/curr_addr[26] , \DataPath/WRF_CUhw/curr_addr[27] ,
         \DataPath/WRF_CUhw/curr_addr[28] , \DataPath/WRF_CUhw/curr_addr[29] ,
         \DataPath/WRF_CUhw/curr_addr[30] , \DataPath/WRF_CUhw/curr_addr[31] ,
         \DataPath/WRF_CUhw/curr_data[31] , \DataPath/WRF_CUhw/curr_data[30] ,
         \DataPath/WRF_CUhw/curr_data[29] , \DataPath/WRF_CUhw/curr_data[28] ,
         \DataPath/WRF_CUhw/curr_data[27] , \DataPath/WRF_CUhw/curr_data[26] ,
         \DataPath/WRF_CUhw/curr_data[25] , \DataPath/WRF_CUhw/curr_data[24] ,
         \DataPath/WRF_CUhw/curr_data[23] , \DataPath/WRF_CUhw/curr_data[22] ,
         \DataPath/WRF_CUhw/curr_data[21] , \DataPath/WRF_CUhw/curr_data[20] ,
         \DataPath/WRF_CUhw/curr_data[19] , \DataPath/WRF_CUhw/curr_data[18] ,
         \DataPath/WRF_CUhw/curr_data[17] , \DataPath/WRF_CUhw/curr_data[16] ,
         \DataPath/WRF_CUhw/curr_data[15] , \DataPath/WRF_CUhw/curr_data[14] ,
         \DataPath/WRF_CUhw/curr_data[13] , \DataPath/WRF_CUhw/curr_data[12] ,
         \DataPath/WRF_CUhw/curr_data[11] , \DataPath/WRF_CUhw/curr_data[10] ,
         \DataPath/WRF_CUhw/curr_data[9] , \DataPath/WRF_CUhw/curr_data[8] ,
         \DataPath/WRF_CUhw/curr_data[7] , \DataPath/WRF_CUhw/curr_data[6] ,
         \DataPath/WRF_CUhw/curr_data[5] , \DataPath/WRF_CUhw/curr_data[4] ,
         \DataPath/WRF_CUhw/curr_data[3] , \DataPath/WRF_CUhw/curr_data[2] ,
         \DataPath/WRF_CUhw/curr_data[1] , \DataPath/WRF_CUhw/curr_data[0] ,
         \DataPath/ALUhw/i_Q_EXTENDED[61] , \DataPath/ALUhw/i_Q_EXTENDED[60] ,
         \DataPath/ALUhw/i_Q_EXTENDED[59] , \DataPath/ALUhw/i_Q_EXTENDED[58] ,
         \DataPath/ALUhw/i_Q_EXTENDED[57] , \DataPath/ALUhw/i_Q_EXTENDED[56] ,
         \DataPath/ALUhw/i_Q_EXTENDED[55] , \DataPath/ALUhw/i_Q_EXTENDED[54] ,
         \DataPath/ALUhw/i_Q_EXTENDED[53] , \DataPath/ALUhw/i_Q_EXTENDED[52] ,
         \DataPath/ALUhw/i_Q_EXTENDED[51] , \DataPath/ALUhw/i_Q_EXTENDED[50] ,
         \DataPath/ALUhw/i_Q_EXTENDED[49] , \DataPath/ALUhw/i_Q_EXTENDED[48] ,
         \DataPath/ALUhw/i_Q_EXTENDED[45] , \DataPath/ALUhw/i_Q_EXTENDED[42] ,
         \DataPath/ALUhw/i_Q_EXTENDED[41] , \DataPath/ALUhw/i_Q_EXTENDED[40] ,
         \DataPath/ALUhw/i_Q_EXTENDED[38] , \DataPath/ALUhw/i_Q_EXTENDED[36] ,
         \DataPath/ALUhw/i_Q_EXTENDED[32] , \DataPath/RF/RDPORT0_OUTLATCH/N35 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N34 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N33 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N32 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N31 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N30 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N29 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N28 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N27 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N26 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N25 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N24 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N23 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N22 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N21 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N20 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N19 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N18 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N17 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N16 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N15 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N14 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N13 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N12 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N11 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N10 , \DataPath/RF/RDPORT0_OUTLATCH/N9 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N8 , \DataPath/RF/RDPORT0_OUTLATCH/N7 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N6 , \DataPath/RF/RDPORT0_OUTLATCH/N5 ,
         \DataPath/RF/RDPORT0_OUTLATCH/N4 , \DataPath/RF/RDPORT0_OUTLATCH/N3 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N35 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N34 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N33 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N32 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N31 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N30 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N29 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N28 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N27 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N26 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N25 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N24 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N23 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N22 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N21 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N20 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N19 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N18 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N17 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N16 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N15 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N14 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N13 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N12 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N11 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N10 , \DataPath/RF/RDPORT1_OUTLATCH/N9 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N8 , \DataPath/RF/RDPORT1_OUTLATCH/N7 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N6 , \DataPath/RF/RDPORT1_OUTLATCH/N5 ,
         \DataPath/RF/RDPORT1_OUTLATCH/N4 , \DataPath/RF/RDPORT1_OUTLATCH/N3 ,
         \DataPath/RF/PUSH_ADDRGEN/N61 , \DataPath/RF/PUSH_ADDRGEN/N60 ,
         \DataPath/RF/PUSH_ADDRGEN/N59 , \DataPath/RF/PUSH_ADDRGEN/N58 ,
         \DataPath/RF/PUSH_ADDRGEN/N57 , \DataPath/RF/PUSH_ADDRGEN/N56 ,
         \DataPath/RF/PUSH_ADDRGEN/N55 , \DataPath/RF/PUSH_ADDRGEN/N54 ,
         \DataPath/RF/PUSH_ADDRGEN/N53 , \DataPath/RF/PUSH_ADDRGEN/N52 ,
         \DataPath/RF/PUSH_ADDRGEN/N51 , \DataPath/RF/PUSH_ADDRGEN/N50 ,
         \DataPath/RF/PUSH_ADDRGEN/N49 , \DataPath/RF/PUSH_ADDRGEN/N48 ,
         \DataPath/RF/PUSH_ADDRGEN/N47 , \DataPath/RF/PUSH_ADDRGEN/N46 ,
         \DataPath/RF/PUSH_ADDRGEN/curr_state[0] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[0] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[1] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[2] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[3] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[4] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[5] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[6] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[7] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[8] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[9] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[10] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[11] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[12] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[13] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[14] ,
         \DataPath/RF/PUSH_ADDRGEN/curr_addr[15] ,
         \DataPath/RF/POP_ADDRGEN/N61 , \DataPath/RF/POP_ADDRGEN/N60 ,
         \DataPath/RF/POP_ADDRGEN/N59 , \DataPath/RF/POP_ADDRGEN/N58 ,
         \DataPath/RF/POP_ADDRGEN/N57 , \DataPath/RF/POP_ADDRGEN/N56 ,
         \DataPath/RF/POP_ADDRGEN/N55 , \DataPath/RF/POP_ADDRGEN/N54 ,
         \DataPath/RF/POP_ADDRGEN/N53 , \DataPath/RF/POP_ADDRGEN/N52 ,
         \DataPath/RF/POP_ADDRGEN/N51 , \DataPath/RF/POP_ADDRGEN/N50 ,
         \DataPath/RF/POP_ADDRGEN/N49 , \DataPath/RF/POP_ADDRGEN/N48 ,
         \DataPath/RF/POP_ADDRGEN/N47 , \DataPath/RF/POP_ADDRGEN/N46 ,
         \DataPath/RF/POP_ADDRGEN/curr_state[1] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[0] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[1] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[2] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[3] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[4] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[5] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[6] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[7] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[8] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[9] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[10] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[11] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[12] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[13] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[14] ,
         \DataPath/RF/POP_ADDRGEN/curr_addr[15] ,
         \DataPath/ALUhw/MULT/mux_out[15][30] ,
         \DataPath/ALUhw/MULT/mux_out[15][31] ,
         \DataPath/ALUhw/MULT/mux_out[14][28] ,
         \DataPath/ALUhw/MULT/mux_out[14][29] ,
         \DataPath/ALUhw/MULT/mux_out[14][30] ,
         \DataPath/ALUhw/MULT/mux_out[14][31] ,
         \DataPath/ALUhw/MULT/mux_out[13][26] ,
         \DataPath/ALUhw/MULT/mux_out[13][27] ,
         \DataPath/ALUhw/MULT/mux_out[13][28] ,
         \DataPath/ALUhw/MULT/mux_out[13][29] ,
         \DataPath/ALUhw/MULT/mux_out[13][30] ,
         \DataPath/ALUhw/MULT/mux_out[13][31] ,
         \DataPath/ALUhw/MULT/mux_out[12][24] ,
         \DataPath/ALUhw/MULT/mux_out[12][25] ,
         \DataPath/ALUhw/MULT/mux_out[12][26] ,
         \DataPath/ALUhw/MULT/mux_out[12][27] ,
         \DataPath/ALUhw/MULT/mux_out[12][28] ,
         \DataPath/ALUhw/MULT/mux_out[12][29] ,
         \DataPath/ALUhw/MULT/mux_out[12][30] ,
         \DataPath/ALUhw/MULT/mux_out[12][31] ,
         \DataPath/ALUhw/MULT/mux_out[11][22] ,
         \DataPath/ALUhw/MULT/mux_out[11][23] ,
         \DataPath/ALUhw/MULT/mux_out[11][24] ,
         \DataPath/ALUhw/MULT/mux_out[11][25] ,
         \DataPath/ALUhw/MULT/mux_out[11][26] ,
         \DataPath/ALUhw/MULT/mux_out[11][27] ,
         \DataPath/ALUhw/MULT/mux_out[11][28] ,
         \DataPath/ALUhw/MULT/mux_out[11][29] ,
         \DataPath/ALUhw/MULT/mux_out[11][30] ,
         \DataPath/ALUhw/MULT/mux_out[11][31] ,
         \DataPath/ALUhw/MULT/mux_out[10][20] ,
         \DataPath/ALUhw/MULT/mux_out[10][21] ,
         \DataPath/ALUhw/MULT/mux_out[10][22] ,
         \DataPath/ALUhw/MULT/mux_out[10][23] ,
         \DataPath/ALUhw/MULT/mux_out[10][24] ,
         \DataPath/ALUhw/MULT/mux_out[10][25] ,
         \DataPath/ALUhw/MULT/mux_out[10][26] ,
         \DataPath/ALUhw/MULT/mux_out[10][27] ,
         \DataPath/ALUhw/MULT/mux_out[10][28] ,
         \DataPath/ALUhw/MULT/mux_out[10][29] ,
         \DataPath/ALUhw/MULT/mux_out[10][30] ,
         \DataPath/ALUhw/MULT/mux_out[10][31] ,
         \DataPath/ALUhw/MULT/mux_out[9][18] ,
         \DataPath/ALUhw/MULT/mux_out[9][19] ,
         \DataPath/ALUhw/MULT/mux_out[9][20] ,
         \DataPath/ALUhw/MULT/mux_out[9][21] ,
         \DataPath/ALUhw/MULT/mux_out[9][22] ,
         \DataPath/ALUhw/MULT/mux_out[9][23] ,
         \DataPath/ALUhw/MULT/mux_out[9][24] ,
         \DataPath/ALUhw/MULT/mux_out[9][25] ,
         \DataPath/ALUhw/MULT/mux_out[9][26] ,
         \DataPath/ALUhw/MULT/mux_out[9][27] ,
         \DataPath/ALUhw/MULT/mux_out[9][28] ,
         \DataPath/ALUhw/MULT/mux_out[9][29] ,
         \DataPath/ALUhw/MULT/mux_out[9][30] ,
         \DataPath/ALUhw/MULT/mux_out[9][31] ,
         \DataPath/ALUhw/MULT/mux_out[8][16] ,
         \DataPath/ALUhw/MULT/mux_out[8][17] ,
         \DataPath/ALUhw/MULT/mux_out[8][18] ,
         \DataPath/ALUhw/MULT/mux_out[8][19] ,
         \DataPath/ALUhw/MULT/mux_out[8][20] ,
         \DataPath/ALUhw/MULT/mux_out[8][21] ,
         \DataPath/ALUhw/MULT/mux_out[8][22] ,
         \DataPath/ALUhw/MULT/mux_out[8][23] ,
         \DataPath/ALUhw/MULT/mux_out[8][24] ,
         \DataPath/ALUhw/MULT/mux_out[8][25] ,
         \DataPath/ALUhw/MULT/mux_out[8][26] ,
         \DataPath/ALUhw/MULT/mux_out[8][27] ,
         \DataPath/ALUhw/MULT/mux_out[8][28] ,
         \DataPath/ALUhw/MULT/mux_out[8][29] ,
         \DataPath/ALUhw/MULT/mux_out[8][30] ,
         \DataPath/ALUhw/MULT/mux_out[8][31] ,
         \DataPath/ALUhw/MULT/mux_out[7][14] ,
         \DataPath/ALUhw/MULT/mux_out[7][15] ,
         \DataPath/ALUhw/MULT/mux_out[7][16] ,
         \DataPath/ALUhw/MULT/mux_out[7][17] ,
         \DataPath/ALUhw/MULT/mux_out[7][18] ,
         \DataPath/ALUhw/MULT/mux_out[7][19] ,
         \DataPath/ALUhw/MULT/mux_out[7][20] ,
         \DataPath/ALUhw/MULT/mux_out[7][21] ,
         \DataPath/ALUhw/MULT/mux_out[7][22] ,
         \DataPath/ALUhw/MULT/mux_out[7][23] ,
         \DataPath/ALUhw/MULT/mux_out[7][24] ,
         \DataPath/ALUhw/MULT/mux_out[7][25] ,
         \DataPath/ALUhw/MULT/mux_out[7][26] ,
         \DataPath/ALUhw/MULT/mux_out[7][27] ,
         \DataPath/ALUhw/MULT/mux_out[7][28] ,
         \DataPath/ALUhw/MULT/mux_out[7][29] ,
         \DataPath/ALUhw/MULT/mux_out[7][30] ,
         \DataPath/ALUhw/MULT/mux_out[7][31] ,
         \DataPath/ALUhw/MULT/mux_out[6][12] ,
         \DataPath/ALUhw/MULT/mux_out[6][13] ,
         \DataPath/ALUhw/MULT/mux_out[6][14] ,
         \DataPath/ALUhw/MULT/mux_out[6][15] ,
         \DataPath/ALUhw/MULT/mux_out[6][16] ,
         \DataPath/ALUhw/MULT/mux_out[6][17] ,
         \DataPath/ALUhw/MULT/mux_out[6][18] ,
         \DataPath/ALUhw/MULT/mux_out[6][19] ,
         \DataPath/ALUhw/MULT/mux_out[6][20] ,
         \DataPath/ALUhw/MULT/mux_out[6][21] ,
         \DataPath/ALUhw/MULT/mux_out[6][22] ,
         \DataPath/ALUhw/MULT/mux_out[6][23] ,
         \DataPath/ALUhw/MULT/mux_out[6][24] ,
         \DataPath/ALUhw/MULT/mux_out[6][25] ,
         \DataPath/ALUhw/MULT/mux_out[6][26] ,
         \DataPath/ALUhw/MULT/mux_out[6][27] ,
         \DataPath/ALUhw/MULT/mux_out[6][28] ,
         \DataPath/ALUhw/MULT/mux_out[6][29] ,
         \DataPath/ALUhw/MULT/mux_out[6][30] ,
         \DataPath/ALUhw/MULT/mux_out[6][31] ,
         \DataPath/ALUhw/MULT/mux_out[5][10] ,
         \DataPath/ALUhw/MULT/mux_out[5][11] ,
         \DataPath/ALUhw/MULT/mux_out[5][12] ,
         \DataPath/ALUhw/MULT/mux_out[5][13] ,
         \DataPath/ALUhw/MULT/mux_out[5][14] ,
         \DataPath/ALUhw/MULT/mux_out[5][15] ,
         \DataPath/ALUhw/MULT/mux_out[5][16] ,
         \DataPath/ALUhw/MULT/mux_out[5][17] ,
         \DataPath/ALUhw/MULT/mux_out[5][18] ,
         \DataPath/ALUhw/MULT/mux_out[5][19] ,
         \DataPath/ALUhw/MULT/mux_out[5][20] ,
         \DataPath/ALUhw/MULT/mux_out[5][21] ,
         \DataPath/ALUhw/MULT/mux_out[5][22] ,
         \DataPath/ALUhw/MULT/mux_out[5][23] ,
         \DataPath/ALUhw/MULT/mux_out[5][24] ,
         \DataPath/ALUhw/MULT/mux_out[5][25] ,
         \DataPath/ALUhw/MULT/mux_out[5][26] ,
         \DataPath/ALUhw/MULT/mux_out[5][27] ,
         \DataPath/ALUhw/MULT/mux_out[5][28] ,
         \DataPath/ALUhw/MULT/mux_out[5][29] ,
         \DataPath/ALUhw/MULT/mux_out[5][30] ,
         \DataPath/ALUhw/MULT/mux_out[5][31] ,
         \DataPath/ALUhw/MULT/mux_out[4][9] ,
         \DataPath/ALUhw/MULT/mux_out[4][10] ,
         \DataPath/ALUhw/MULT/mux_out[4][11] ,
         \DataPath/ALUhw/MULT/mux_out[4][12] ,
         \DataPath/ALUhw/MULT/mux_out[4][13] ,
         \DataPath/ALUhw/MULT/mux_out[4][14] ,
         \DataPath/ALUhw/MULT/mux_out[4][15] ,
         \DataPath/ALUhw/MULT/mux_out[4][16] ,
         \DataPath/ALUhw/MULT/mux_out[4][17] ,
         \DataPath/ALUhw/MULT/mux_out[4][18] ,
         \DataPath/ALUhw/MULT/mux_out[4][19] ,
         \DataPath/ALUhw/MULT/mux_out[4][20] ,
         \DataPath/ALUhw/MULT/mux_out[4][21] ,
         \DataPath/ALUhw/MULT/mux_out[4][22] ,
         \DataPath/ALUhw/MULT/mux_out[4][23] ,
         \DataPath/ALUhw/MULT/mux_out[4][24] ,
         \DataPath/ALUhw/MULT/mux_out[4][25] ,
         \DataPath/ALUhw/MULT/mux_out[4][26] ,
         \DataPath/ALUhw/MULT/mux_out[4][27] ,
         \DataPath/ALUhw/MULT/mux_out[4][28] ,
         \DataPath/ALUhw/MULT/mux_out[4][29] ,
         \DataPath/ALUhw/MULT/mux_out[4][30] ,
         \DataPath/ALUhw/MULT/mux_out[4][31] ,
         \DataPath/ALUhw/MULT/mux_out[3][6] ,
         \DataPath/ALUhw/MULT/mux_out[3][7] ,
         \DataPath/ALUhw/MULT/mux_out[3][8] ,
         \DataPath/ALUhw/MULT/mux_out[3][9] ,
         \DataPath/ALUhw/MULT/mux_out[3][10] ,
         \DataPath/ALUhw/MULT/mux_out[3][11] ,
         \DataPath/ALUhw/MULT/mux_out[3][12] ,
         \DataPath/ALUhw/MULT/mux_out[3][13] ,
         \DataPath/ALUhw/MULT/mux_out[3][14] ,
         \DataPath/ALUhw/MULT/mux_out[3][15] ,
         \DataPath/ALUhw/MULT/mux_out[3][16] ,
         \DataPath/ALUhw/MULT/mux_out[3][17] ,
         \DataPath/ALUhw/MULT/mux_out[3][18] ,
         \DataPath/ALUhw/MULT/mux_out[3][19] ,
         \DataPath/ALUhw/MULT/mux_out[3][20] ,
         \DataPath/ALUhw/MULT/mux_out[3][21] ,
         \DataPath/ALUhw/MULT/mux_out[3][22] ,
         \DataPath/ALUhw/MULT/mux_out[3][23] ,
         \DataPath/ALUhw/MULT/mux_out[3][24] ,
         \DataPath/ALUhw/MULT/mux_out[3][25] ,
         \DataPath/ALUhw/MULT/mux_out[3][26] ,
         \DataPath/ALUhw/MULT/mux_out[3][27] ,
         \DataPath/ALUhw/MULT/mux_out[3][28] ,
         \DataPath/ALUhw/MULT/mux_out[3][29] ,
         \DataPath/ALUhw/MULT/mux_out[3][30] ,
         \DataPath/ALUhw/MULT/mux_out[3][31] ,
         \DataPath/ALUhw/MULT/mux_out[2][5] ,
         \DataPath/ALUhw/MULT/mux_out[2][6] ,
         \DataPath/ALUhw/MULT/mux_out[2][7] ,
         \DataPath/ALUhw/MULT/mux_out[2][8] ,
         \DataPath/ALUhw/MULT/mux_out[2][9] ,
         \DataPath/ALUhw/MULT/mux_out[2][10] ,
         \DataPath/ALUhw/MULT/mux_out[2][11] ,
         \DataPath/ALUhw/MULT/mux_out[2][12] ,
         \DataPath/ALUhw/MULT/mux_out[2][13] ,
         \DataPath/ALUhw/MULT/mux_out[2][14] ,
         \DataPath/ALUhw/MULT/mux_out[2][15] ,
         \DataPath/ALUhw/MULT/mux_out[2][16] ,
         \DataPath/ALUhw/MULT/mux_out[2][17] ,
         \DataPath/ALUhw/MULT/mux_out[2][18] ,
         \DataPath/ALUhw/MULT/mux_out[2][19] ,
         \DataPath/ALUhw/MULT/mux_out[2][20] ,
         \DataPath/ALUhw/MULT/mux_out[2][21] ,
         \DataPath/ALUhw/MULT/mux_out[2][22] ,
         \DataPath/ALUhw/MULT/mux_out[2][23] ,
         \DataPath/ALUhw/MULT/mux_out[2][24] ,
         \DataPath/ALUhw/MULT/mux_out[2][25] ,
         \DataPath/ALUhw/MULT/mux_out[2][26] ,
         \DataPath/ALUhw/MULT/mux_out[2][27] ,
         \DataPath/ALUhw/MULT/mux_out[2][28] ,
         \DataPath/ALUhw/MULT/mux_out[2][29] ,
         \DataPath/ALUhw/MULT/mux_out[2][30] ,
         \DataPath/ALUhw/MULT/mux_out[2][31] ,
         \DataPath/ALUhw/MULT/mux_out[1][2] ,
         \DataPath/ALUhw/MULT/mux_out[1][3] ,
         \DataPath/ALUhw/MULT/mux_out[1][6] ,
         \DataPath/ALUhw/MULT/mux_out[1][7] ,
         \DataPath/ALUhw/MULT/mux_out[1][8] ,
         \DataPath/ALUhw/MULT/mux_out[1][9] ,
         \DataPath/ALUhw/MULT/mux_out[1][10] ,
         \DataPath/ALUhw/MULT/mux_out[1][11] ,
         \DataPath/ALUhw/MULT/mux_out[1][12] ,
         \DataPath/ALUhw/MULT/mux_out[1][15] ,
         \DataPath/ALUhw/MULT/mux_out[1][16] ,
         \DataPath/ALUhw/MULT/mux_out[1][17] ,
         \DataPath/ALUhw/MULT/mux_out[1][18] ,
         \DataPath/ALUhw/MULT/mux_out[1][19] ,
         \DataPath/ALUhw/MULT/mux_out[1][20] ,
         \DataPath/ALUhw/MULT/mux_out[1][21] ,
         \DataPath/ALUhw/MULT/mux_out[1][22] ,
         \DataPath/ALUhw/MULT/mux_out[1][23] ,
         \DataPath/ALUhw/MULT/mux_out[1][24] ,
         \DataPath/ALUhw/MULT/mux_out[1][25] ,
         \DataPath/ALUhw/MULT/mux_out[1][26] ,
         \DataPath/ALUhw/MULT/mux_out[1][29] ,
         \DataPath/ALUhw/MULT/mux_out[1][30] ,
         \DataPath/ALUhw/MULT/mux_out[1][31] ,
         \DataPath/ALUhw/MULT/mux_out[0][0] ,
         \DataPath/ALUhw/MULT/mux_out[0][4] ,
         \DataPath/ALUhw/MULT/mux_out[0][5] ,
         \DataPath/ALUhw/MULT/mux_out[0][6] ,
         \DataPath/ALUhw/MULT/mux_out[0][7] ,
         \DataPath/ALUhw/MULT/mux_out[0][8] ,
         \DataPath/ALUhw/MULT/mux_out[0][9] ,
         \DataPath/ALUhw/MULT/mux_out[0][10] ,
         \DataPath/ALUhw/MULT/mux_out[0][11] ,
         \DataPath/ALUhw/MULT/mux_out[0][12] ,
         \DataPath/ALUhw/MULT/mux_out[0][13] ,
         \DataPath/ALUhw/MULT/mux_out[0][15] ,
         \DataPath/ALUhw/MULT/mux_out[0][16] ,
         \DataPath/ALUhw/MULT/mux_out[0][24] ,
         \DataPath/ALUhw/MULT/mux_out[0][25] ,
         \DataPath/ALUhw/MULT/mux_out[0][26] ,
         \DataPath/ALUhw/MULT/mux_out[0][31] , \C620/DATA2_2 , \C620/DATA2_3 ,
         \C620/DATA2_4 , \C620/DATA2_5 , \C620/DATA2_6 , \C620/DATA2_7 ,
         \C620/DATA2_8 , \C620/DATA2_9 , \C620/DATA2_10 , \C620/DATA2_11 ,
         \C620/DATA2_12 , \C620/DATA2_13 , \C620/DATA2_14 , \C620/DATA2_15 ,
         \C620/DATA2_16 , \C620/DATA2_23 , \C620/DATA2_24 , \C620/DATA2_25 ,
         \C620/DATA2_26 , \C620/DATA2_27 , \C620/DATA2_29 , \C620/DATA2_31 ,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n90, n99, n102,
         n165, n166, n167, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n208, n210, n217, n218,
         n222, n223, n359, n360, n361, n362, n363, n366, n367, n368, n369,
         n370, n380, n381, n406, n465, n466, n470, n471, n481, n497, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n537, n539, n555, n556, n558, n560, n562, n564, n566, n568, n570,
         n572, n574, n576, n578, n580, n582, n583, n584, n589, n590, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n835, n836, n849, n877, n892, n896, n898, n900,
         n902, n904, n906, n908, n910, n912, n914, n916, n918, n920, n922,
         n924, n926, n928, n930, n934, n936, n938, n940, n942, n944, n946,
         n948, n950, n952, n954, n956, n958, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n982, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1019, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1056, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1093, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1130, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n2011, n2133, n2165, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2346, n2348, n2350, n2352, n2354,
         n2356, n2358, n2360, n2362, n2364, n2366, n2371, n2373, n2375, n2377,
         n2383, n2386, n2389, n2392, n2396, n2398, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2775, n2776, n2777, n2778, n2779, n2780, n2846, n2847,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2861, n2866,
         n2867, n2868, n2869, n2870, n2872, n2886, n2889, n2890, n3147, n3153,
         n3197, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3307, n3309,
         n3311, n3313, n3315, n3317, n3319, n3321, n3323, n3325, n3327, n3329,
         n3331, n3333, n3335, n3337, n3339, n3341, n3343, n3345, n3347, n3349,
         n3351, n3353, n3355, n3357, n3359, n3361, n3363, n3365, n3367, n3374,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3412, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3450, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3488, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3526, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3564,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3602, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3640, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3677, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3714, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3751,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3786, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3821, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3856, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3891, n3895, n3897,
         n3899, n3901, n3903, n3905, n3907, n3909, n3911, n3913, n3915, n3917,
         n3919, n3921, n3923, n3925, n3927, n3929, n3931, n3933, n3935, n3937,
         n3939, n3941, n3943, n3945, n3947, n3949, n3951, n3953, n3955, n3959,
         n3963, n3965, n3967, n3969, n3971, n3973, n3975, n3977, n3979, n3981,
         n3983, n3985, n3987, n3989, n3991, n3993, n3995, n3997, n3999, n4001,
         n4003, n4005, n4007, n4009, n4011, n4013, n4015, n4017, n4019, n4021,
         n4023, n4027, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4062, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4097, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4132, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4167,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4202, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4237, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4272, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4307, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4342,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4377, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4412, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4447, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4482, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4517,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4552, n4556, n4558, n4560, n4562, n4564, n4566, n4568, n4570,
         n4572, n4574, n4576, n4578, n4580, n4582, n4584, n4586, n4588, n4590,
         n4592, n4594, n4596, n4598, n4600, n4602, n4604, n4606, n4608, n4610,
         n4612, n4614, n4616, n4620, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4655, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4690, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4725,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4760, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4795, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4830, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4865, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4900,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4935, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4970, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5005, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5040, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5075,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5110, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5145, n5149, n5151, n5153, n5155, n5157, n5159,
         n5161, n5163, n5165, n5167, n5169, n5171, n5173, n5175, n5177, n5179,
         n5181, n5183, n5185, n5187, n5189, n5191, n5193, n5195, n5197, n5199,
         n5201, n5203, n5205, n5207, n5209, n5212, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5248, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5283,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5318, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5353, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5388, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5423, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5458,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5493, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5528, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5563, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5602, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5639,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5676, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5713, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5750, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5789, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5825,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5861, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5897, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5933, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5969, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6005,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6042, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6078, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6723,
         n6724, n6725, n6726, n6727, n6728, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7124, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7166, n7168, n7169, n7170, \intadd_2/B[3] , \intadd_2/B[2] ,
         \intadd_2/B[1] , \intadd_2/B[0] , \intadd_2/SUM[3] ,
         \intadd_2/SUM[1] , \intadd_2/SUM[0] , \intadd_2/CO , \intadd_2/n33 ,
         \intadd_2/n32 , \intadd_2/n30 , \intadd_2/n28 , \intadd_2/n27 ,
         \intadd_2/n25 , \intadd_2/n23 , \intadd_2/n22 , \intadd_2/n18 ,
         \intadd_2/n17 , \intadd_2/n16 , \intadd_2/n15 , \intadd_2/n14 ,
         \intadd_2/n13 , \intadd_2/n11 , \intadd_2/n9 , \intadd_2/n4 ,
         \intadd_2/n3 , \intadd_2/n1 , \intadd_0/A[0] , \intadd_0/B[4] ,
         \intadd_0/B[3] , \intadd_0/B[2] , \intadd_0/B[1] , \intadd_0/B[0] ,
         \intadd_0/SUM[4] , \intadd_0/SUM[3] , \intadd_0/SUM[2] ,
         \intadd_0/SUM[1] , \intadd_0/SUM[0] , \intadd_0/n45 , \intadd_0/n44 ,
         \intadd_0/n41 , \intadd_0/n40 , \intadd_0/n38 , \intadd_0/n36 ,
         \intadd_0/n35 , \intadd_0/n33 , \intadd_0/n31 , \intadd_0/n30 ,
         \intadd_0/n29 , \intadd_0/n28 , \intadd_0/n27 , \intadd_0/n26 ,
         \intadd_0/n25 , \intadd_0/n24 , \intadd_0/n23 , \intadd_0/n22 ,
         \intadd_0/n21 , \intadd_0/n19 , \intadd_0/n17 , \intadd_0/n16 ,
         \intadd_0/n15 , \intadd_0/n14 , \intadd_0/n5 , \intadd_0/n4 ,
         \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 , \intadd_1/A[4] ,
         \intadd_1/A[3] , \intadd_1/A[1] , \intadd_1/A[0] , \intadd_1/B[4] ,
         \intadd_1/B[2] , \intadd_1/B[1] , \intadd_1/B[0] , \intadd_1/CI ,
         \intadd_1/SUM[4] , \intadd_1/SUM[3] , \intadd_1/SUM[2] ,
         \intadd_1/SUM[1] , \intadd_1/SUM[0] , \intadd_1/CO , \intadd_1/n36 ,
         \intadd_1/n35 , \intadd_1/n34 , \intadd_1/n33 , \intadd_1/n32 ,
         \intadd_1/n31 , \intadd_1/n30 , \intadd_1/n29 , \intadd_1/n28 ,
         \intadd_1/n27 , \intadd_1/n26 , \intadd_1/n25 , \intadd_1/n24 ,
         \intadd_1/n23 , \intadd_1/n22 , \intadd_1/n21 , \intadd_1/n20 ,
         \intadd_1/n19 , \intadd_1/n18 , \intadd_1/n17 , \intadd_1/n16 ,
         \intadd_1/n15 , \intadd_1/n13 , \intadd_1/n12 , \intadd_1/n11 ,
         \intadd_1/n10 , \intadd_1/n8 , \intadd_1/n5 , \intadd_1/n4 ,
         \intadd_1/n3 , \intadd_1/n2 , \intadd_1/n1 ,
         \DP_OP_1091J1_126_6973/n72 , \DP_OP_1091J1_126_6973/n37 ,
         \DP_OP_1091J1_126_6973/n30 , \DP_OP_1091J1_126_6973/n29 ,
         \DP_OP_1091J1_126_6973/n28 , \DP_OP_1091J1_126_6973/n27 ,
         \DP_OP_1091J1_126_6973/n26 , \DP_OP_1091J1_126_6973/n25 ,
         \DP_OP_1091J1_126_6973/n24 , \DP_OP_1091J1_126_6973/n23 ,
         \DP_OP_1091J1_126_6973/n22 , \DP_OP_1091J1_126_6973/n21 ,
         \DP_OP_1091J1_126_6973/n20 , \DP_OP_1091J1_126_6973/n19 ,
         \DP_OP_1091J1_126_6973/n18 , \DP_OP_1091J1_126_6973/n17 ,
         \DP_OP_1091J1_126_6973/n16 , \DP_OP_1091J1_126_6973/n15 ,
         \DP_OP_1091J1_126_6973/n13 , \DP_OP_1091J1_126_6973/n10 ,
         \DP_OP_1091J1_126_6973/n9 , \DP_OP_1091J1_126_6973/n8 ,
         \DP_OP_1091J1_126_6973/n7 , \DP_OP_1091J1_126_6973/n6 ,
         \DP_OP_1091J1_126_6973/n5 , \DP_OP_751_130_6421/n1781 ,
         \DP_OP_751_130_6421/n1780 , \DP_OP_751_130_6421/n1779 ,
         \DP_OP_751_130_6421/n1778 , \DP_OP_751_130_6421/n1777 ,
         \DP_OP_751_130_6421/n1776 , \DP_OP_751_130_6421/n1775 ,
         \DP_OP_751_130_6421/n1771 , \DP_OP_751_130_6421/n1763 ,
         \DP_OP_751_130_6421/n1762 , \DP_OP_751_130_6421/n1761 ,
         \DP_OP_751_130_6421/n1756 , \DP_OP_751_130_6421/n1753 ,
         \DP_OP_751_130_6421/n1752 , \DP_OP_751_130_6421/n1744 ,
         \DP_OP_751_130_6421/n1743 , \DP_OP_751_130_6421/n1742 ,
         \DP_OP_751_130_6421/n1741 , \DP_OP_751_130_6421/n1740 ,
         \DP_OP_751_130_6421/n1736 , \DP_OP_751_130_6421/n1735 ,
         \DP_OP_751_130_6421/n1734 , \DP_OP_751_130_6421/n1733 ,
         \DP_OP_751_130_6421/n1732 , \DP_OP_751_130_6421/n1731 ,
         \DP_OP_751_130_6421/n1730 , \DP_OP_751_130_6421/n1729 ,
         \DP_OP_751_130_6421/n1728 , \DP_OP_751_130_6421/n1727 ,
         \DP_OP_751_130_6421/n1726 , \DP_OP_751_130_6421/n1725 ,
         \DP_OP_751_130_6421/n1724 , \DP_OP_751_130_6421/n1721 ,
         \DP_OP_751_130_6421/n1719 , \DP_OP_751_130_6421/n1714 ,
         \DP_OP_751_130_6421/n1713 , \DP_OP_751_130_6421/n1712 ,
         \DP_OP_751_130_6421/n1711 , \DP_OP_751_130_6421/n1710 ,
         \DP_OP_751_130_6421/n1706 , \DP_OP_751_130_6421/n1705 ,
         \DP_OP_751_130_6421/n1704 , \DP_OP_751_130_6421/n1703 ,
         \DP_OP_751_130_6421/n1702 , \DP_OP_751_130_6421/n1701 ,
         \DP_OP_751_130_6421/n1700 , \DP_OP_751_130_6421/n1699 ,
         \DP_OP_751_130_6421/n1698 , \DP_OP_751_130_6421/n1697 ,
         \DP_OP_751_130_6421/n1696 , \DP_OP_751_130_6421/n1693 ,
         \DP_OP_751_130_6421/n1692 , \DP_OP_751_130_6421/n1691 ,
         \DP_OP_751_130_6421/n1686 , \DP_OP_751_130_6421/n1685 ,
         \DP_OP_751_130_6421/n1684 , \DP_OP_751_130_6421/n1683 ,
         \DP_OP_751_130_6421/n1682 , \DP_OP_751_130_6421/n1681 ,
         \DP_OP_751_130_6421/n1680 , \DP_OP_751_130_6421/n1679 ,
         \DP_OP_751_130_6421/n1678 , \DP_OP_751_130_6421/n1677 ,
         \DP_OP_751_130_6421/n1676 , \DP_OP_751_130_6421/n1675 ,
         \DP_OP_751_130_6421/n1674 , \DP_OP_751_130_6421/n1673 ,
         \DP_OP_751_130_6421/n1672 , \DP_OP_751_130_6421/n1671 ,
         \DP_OP_751_130_6421/n1670 , \DP_OP_751_130_6421/n1669 ,
         \DP_OP_751_130_6421/n1668 , \DP_OP_751_130_6421/n1667 ,
         \DP_OP_751_130_6421/n1666 , \DP_OP_751_130_6421/n1665 ,
         \DP_OP_751_130_6421/n1664 , \DP_OP_751_130_6421/n1663 ,
         \DP_OP_751_130_6421/n1662 , \DP_OP_751_130_6421/n1661 ,
         \DP_OP_751_130_6421/n1660 , \DP_OP_751_130_6421/n1659 ,
         \DP_OP_751_130_6421/n1658 , \DP_OP_751_130_6421/n1657 ,
         \DP_OP_751_130_6421/n1656 , \DP_OP_751_130_6421/n1655 ,
         \DP_OP_751_130_6421/n1654 , \DP_OP_751_130_6421/n1653 ,
         \DP_OP_751_130_6421/n1652 , \DP_OP_751_130_6421/n1651 ,
         \DP_OP_751_130_6421/n1650 , \DP_OP_751_130_6421/n1649 ,
         \DP_OP_751_130_6421/n1648 , \DP_OP_751_130_6421/n1647 ,
         \DP_OP_751_130_6421/n1646 , \DP_OP_751_130_6421/n1645 ,
         \DP_OP_751_130_6421/n1644 , \DP_OP_751_130_6421/n1643 ,
         \DP_OP_751_130_6421/n1642 , \DP_OP_751_130_6421/n1641 ,
         \DP_OP_751_130_6421/n1640 , \DP_OP_751_130_6421/n1639 ,
         \DP_OP_751_130_6421/n1638 , \DP_OP_751_130_6421/n1637 ,
         \DP_OP_751_130_6421/n1636 , \DP_OP_751_130_6421/n1635 ,
         \DP_OP_751_130_6421/n1634 , \DP_OP_751_130_6421/n1633 ,
         \DP_OP_751_130_6421/n1632 , \DP_OP_751_130_6421/n1631 ,
         \DP_OP_751_130_6421/n1630 , \DP_OP_751_130_6421/n1629 ,
         \DP_OP_751_130_6421/n1628 , \DP_OP_751_130_6421/n1626 ,
         \DP_OP_751_130_6421/n1617 , \DP_OP_751_130_6421/n1615 ,
         \DP_OP_751_130_6421/n1614 , \DP_OP_751_130_6421/n1613 ,
         \DP_OP_751_130_6421/n1612 , \DP_OP_751_130_6421/n1611 ,
         \DP_OP_751_130_6421/n1610 , \DP_OP_751_130_6421/n1609 ,
         \DP_OP_751_130_6421/n1608 , \DP_OP_751_130_6421/n1607 ,
         \DP_OP_751_130_6421/n1606 , \DP_OP_751_130_6421/n1605 ,
         \DP_OP_751_130_6421/n1604 , \DP_OP_751_130_6421/n1603 ,
         \DP_OP_751_130_6421/n1602 , \DP_OP_751_130_6421/n1601 ,
         \DP_OP_751_130_6421/n1600 , \DP_OP_751_130_6421/n1599 ,
         \DP_OP_751_130_6421/n1598 , \DP_OP_751_130_6421/n1597 ,
         \DP_OP_751_130_6421/n1596 , \DP_OP_751_130_6421/n1595 ,
         \DP_OP_751_130_6421/n1594 , \DP_OP_751_130_6421/n1593 ,
         \DP_OP_751_130_6421/n1592 , \DP_OP_751_130_6421/n1591 ,
         \DP_OP_751_130_6421/n1590 , \DP_OP_751_130_6421/n1582 ,
         \DP_OP_751_130_6421/n1581 , \DP_OP_751_130_6421/n1580 ,
         \DP_OP_751_130_6421/n1579 , \DP_OP_751_130_6421/n1578 ,
         \DP_OP_751_130_6421/n1577 , \DP_OP_751_130_6421/n1576 ,
         \DP_OP_751_130_6421/n1575 , \DP_OP_751_130_6421/n1574 ,
         \DP_OP_751_130_6421/n1573 , \DP_OP_751_130_6421/n1572 ,
         \DP_OP_751_130_6421/n1571 , \DP_OP_751_130_6421/n1570 ,
         \DP_OP_751_130_6421/n1569 , \DP_OP_751_130_6421/n1568 ,
         \DP_OP_751_130_6421/n1567 , \DP_OP_751_130_6421/n1566 ,
         \DP_OP_751_130_6421/n1565 , \DP_OP_751_130_6421/n1564 ,
         \DP_OP_751_130_6421/n1563 , \DP_OP_751_130_6421/n1562 ,
         \DP_OP_751_130_6421/n1561 , \DP_OP_751_130_6421/n1560 ,
         \DP_OP_751_130_6421/n1559 , \DP_OP_751_130_6421/n1558 ,
         \DP_OP_751_130_6421/n1557 , \DP_OP_751_130_6421/n1556 ,
         \DP_OP_751_130_6421/n1555 , \DP_OP_751_130_6421/n1554 ,
         \DP_OP_751_130_6421/n1553 , \DP_OP_751_130_6421/n1552 ,
         \DP_OP_751_130_6421/n1551 , \DP_OP_751_130_6421/n1550 ,
         \DP_OP_751_130_6421/n1549 , \DP_OP_751_130_6421/n1548 ,
         \DP_OP_751_130_6421/n1547 , \DP_OP_751_130_6421/n1546 ,
         \DP_OP_751_130_6421/n1545 , \DP_OP_751_130_6421/n1544 ,
         \DP_OP_751_130_6421/n1543 , \DP_OP_751_130_6421/n1542 ,
         \DP_OP_751_130_6421/n1541 , \DP_OP_751_130_6421/n1540 ,
         \DP_OP_751_130_6421/n1539 , \DP_OP_751_130_6421/n1538 ,
         \DP_OP_751_130_6421/n1537 , \DP_OP_751_130_6421/n1536 ,
         \DP_OP_751_130_6421/n1535 , \DP_OP_751_130_6421/n1534 ,
         \DP_OP_751_130_6421/n1533 , \DP_OP_751_130_6421/n1532 ,
         \DP_OP_751_130_6421/n1531 , \DP_OP_751_130_6421/n1530 ,
         \DP_OP_751_130_6421/n1529 , \DP_OP_751_130_6421/n1528 ,
         \DP_OP_751_130_6421/n1515 , \DP_OP_751_130_6421/n1514 ,
         \DP_OP_751_130_6421/n1513 , \DP_OP_751_130_6421/n1512 ,
         \DP_OP_751_130_6421/n1511 , \DP_OP_751_130_6421/n1510 ,
         \DP_OP_751_130_6421/n1509 , \DP_OP_751_130_6421/n1508 ,
         \DP_OP_751_130_6421/n1507 , \DP_OP_751_130_6421/n1506 ,
         \DP_OP_751_130_6421/n1505 , \DP_OP_751_130_6421/n1504 ,
         \DP_OP_751_130_6421/n1503 , \DP_OP_751_130_6421/n1502 ,
         \DP_OP_751_130_6421/n1501 , \DP_OP_751_130_6421/n1500 ,
         \DP_OP_751_130_6421/n1499 , \DP_OP_751_130_6421/n1498 ,
         \DP_OP_751_130_6421/n1497 , \DP_OP_751_130_6421/n1496 ,
         \DP_OP_751_130_6421/n1495 , \DP_OP_751_130_6421/n1494 ,
         \DP_OP_751_130_6421/n1493 , \DP_OP_751_130_6421/n1492 ,
         \DP_OP_751_130_6421/n1491 , \DP_OP_751_130_6421/n1490 ,
         \DP_OP_751_130_6421/n1489 , \DP_OP_751_130_6421/n1480 ,
         \DP_OP_751_130_6421/n1479 , \DP_OP_751_130_6421/n1478 ,
         \DP_OP_751_130_6421/n1477 , \DP_OP_751_130_6421/n1476 ,
         \DP_OP_751_130_6421/n1475 , \DP_OP_751_130_6421/n1474 ,
         \DP_OP_751_130_6421/n1473 , \DP_OP_751_130_6421/n1472 ,
         \DP_OP_751_130_6421/n1471 , \DP_OP_751_130_6421/n1470 ,
         \DP_OP_751_130_6421/n1469 , \DP_OP_751_130_6421/n1468 ,
         \DP_OP_751_130_6421/n1467 , \DP_OP_751_130_6421/n1466 ,
         \DP_OP_751_130_6421/n1465 , \DP_OP_751_130_6421/n1464 ,
         \DP_OP_751_130_6421/n1463 , \DP_OP_751_130_6421/n1462 ,
         \DP_OP_751_130_6421/n1461 , \DP_OP_751_130_6421/n1460 ,
         \DP_OP_751_130_6421/n1459 , \DP_OP_751_130_6421/n1458 ,
         \DP_OP_751_130_6421/n1457 , \DP_OP_751_130_6421/n1456 ,
         \DP_OP_751_130_6421/n1455 , \DP_OP_751_130_6421/n1454 ,
         \DP_OP_751_130_6421/n1453 , \DP_OP_751_130_6421/n1452 ,
         \DP_OP_751_130_6421/n1451 , \DP_OP_751_130_6421/n1450 ,
         \DP_OP_751_130_6421/n1449 , \DP_OP_751_130_6421/n1448 ,
         \DP_OP_751_130_6421/n1447 , \DP_OP_751_130_6421/n1446 ,
         \DP_OP_751_130_6421/n1445 , \DP_OP_751_130_6421/n1444 ,
         \DP_OP_751_130_6421/n1443 , \DP_OP_751_130_6421/n1442 ,
         \DP_OP_751_130_6421/n1441 , \DP_OP_751_130_6421/n1440 ,
         \DP_OP_751_130_6421/n1439 , \DP_OP_751_130_6421/n1438 ,
         \DP_OP_751_130_6421/n1437 , \DP_OP_751_130_6421/n1436 ,
         \DP_OP_751_130_6421/n1435 , \DP_OP_751_130_6421/n1434 ,
         \DP_OP_751_130_6421/n1433 , \DP_OP_751_130_6421/n1431 ,
         \DP_OP_751_130_6421/n1430 , \DP_OP_751_130_6421/n1413 ,
         \DP_OP_751_130_6421/n1411 , \DP_OP_751_130_6421/n1410 ,
         \DP_OP_751_130_6421/n1409 , \DP_OP_751_130_6421/n1408 ,
         \DP_OP_751_130_6421/n1407 , \DP_OP_751_130_6421/n1406 ,
         \DP_OP_751_130_6421/n1405 , \DP_OP_751_130_6421/n1404 ,
         \DP_OP_751_130_6421/n1403 , \DP_OP_751_130_6421/n1402 ,
         \DP_OP_751_130_6421/n1401 , \DP_OP_751_130_6421/n1400 ,
         \DP_OP_751_130_6421/n1399 , \DP_OP_751_130_6421/n1398 ,
         \DP_OP_751_130_6421/n1397 , \DP_OP_751_130_6421/n1396 ,
         \DP_OP_751_130_6421/n1395 , \DP_OP_751_130_6421/n1394 ,
         \DP_OP_751_130_6421/n1393 , \DP_OP_751_130_6421/n1392 ,
         \DP_OP_751_130_6421/n1391 , \DP_OP_751_130_6421/n1390 ,
         \DP_OP_751_130_6421/n1389 , \DP_OP_751_130_6421/n1378 ,
         \DP_OP_751_130_6421/n1377 , \DP_OP_751_130_6421/n1376 ,
         \DP_OP_751_130_6421/n1375 , \DP_OP_751_130_6421/n1374 ,
         \DP_OP_751_130_6421/n1373 , \DP_OP_751_130_6421/n1372 ,
         \DP_OP_751_130_6421/n1371 , \DP_OP_751_130_6421/n1370 ,
         \DP_OP_751_130_6421/n1369 , \DP_OP_751_130_6421/n1368 ,
         \DP_OP_751_130_6421/n1367 , \DP_OP_751_130_6421/n1366 ,
         \DP_OP_751_130_6421/n1365 , \DP_OP_751_130_6421/n1364 ,
         \DP_OP_751_130_6421/n1363 , \DP_OP_751_130_6421/n1362 ,
         \DP_OP_751_130_6421/n1361 , \DP_OP_751_130_6421/n1360 ,
         \DP_OP_751_130_6421/n1359 , \DP_OP_751_130_6421/n1358 ,
         \DP_OP_751_130_6421/n1357 , \DP_OP_751_130_6421/n1356 ,
         \DP_OP_751_130_6421/n1355 , \DP_OP_751_130_6421/n1354 ,
         \DP_OP_751_130_6421/n1353 , \DP_OP_751_130_6421/n1352 ,
         \DP_OP_751_130_6421/n1351 , \DP_OP_751_130_6421/n1350 ,
         \DP_OP_751_130_6421/n1349 , \DP_OP_751_130_6421/n1348 ,
         \DP_OP_751_130_6421/n1347 , \DP_OP_751_130_6421/n1346 ,
         \DP_OP_751_130_6421/n1345 , \DP_OP_751_130_6421/n1344 ,
         \DP_OP_751_130_6421/n1343 , \DP_OP_751_130_6421/n1342 ,
         \DP_OP_751_130_6421/n1341 , \DP_OP_751_130_6421/n1340 ,
         \DP_OP_751_130_6421/n1339 , \DP_OP_751_130_6421/n1338 ,
         \DP_OP_751_130_6421/n1337 , \DP_OP_751_130_6421/n1336 ,
         \DP_OP_751_130_6421/n1335 , \DP_OP_751_130_6421/n1334 ,
         \DP_OP_751_130_6421/n1333 , \DP_OP_751_130_6421/n1332 ,
         \DP_OP_751_130_6421/n1311 , \DP_OP_751_130_6421/n1310 ,
         \DP_OP_751_130_6421/n1309 , \DP_OP_751_130_6421/n1308 ,
         \DP_OP_751_130_6421/n1307 , \DP_OP_751_130_6421/n1306 ,
         \DP_OP_751_130_6421/n1305 , \DP_OP_751_130_6421/n1304 ,
         \DP_OP_751_130_6421/n1303 , \DP_OP_751_130_6421/n1302 ,
         \DP_OP_751_130_6421/n1301 , \DP_OP_751_130_6421/n1300 ,
         \DP_OP_751_130_6421/n1299 , \DP_OP_751_130_6421/n1298 ,
         \DP_OP_751_130_6421/n1297 , \DP_OP_751_130_6421/n1296 ,
         \DP_OP_751_130_6421/n1295 , \DP_OP_751_130_6421/n1294 ,
         \DP_OP_751_130_6421/n1293 , \DP_OP_751_130_6421/n1292 ,
         \DP_OP_751_130_6421/n1291 , \DP_OP_751_130_6421/n1290 ,
         \DP_OP_751_130_6421/n1289 , \DP_OP_751_130_6421/n1276 ,
         \DP_OP_751_130_6421/n1275 , \DP_OP_751_130_6421/n1274 ,
         \DP_OP_751_130_6421/n1273 , \DP_OP_751_130_6421/n1272 ,
         \DP_OP_751_130_6421/n1271 , \DP_OP_751_130_6421/n1270 ,
         \DP_OP_751_130_6421/n1269 , \DP_OP_751_130_6421/n1268 ,
         \DP_OP_751_130_6421/n1267 , \DP_OP_751_130_6421/n1266 ,
         \DP_OP_751_130_6421/n1265 , \DP_OP_751_130_6421/n1264 ,
         \DP_OP_751_130_6421/n1263 , \DP_OP_751_130_6421/n1262 ,
         \DP_OP_751_130_6421/n1261 , \DP_OP_751_130_6421/n1260 ,
         \DP_OP_751_130_6421/n1259 , \DP_OP_751_130_6421/n1258 ,
         \DP_OP_751_130_6421/n1257 , \DP_OP_751_130_6421/n1256 ,
         \DP_OP_751_130_6421/n1255 , \DP_OP_751_130_6421/n1254 ,
         \DP_OP_751_130_6421/n1253 , \DP_OP_751_130_6421/n1252 ,
         \DP_OP_751_130_6421/n1251 , \DP_OP_751_130_6421/n1250 ,
         \DP_OP_751_130_6421/n1249 , \DP_OP_751_130_6421/n1248 ,
         \DP_OP_751_130_6421/n1247 , \DP_OP_751_130_6421/n1246 ,
         \DP_OP_751_130_6421/n1245 , \DP_OP_751_130_6421/n1244 ,
         \DP_OP_751_130_6421/n1243 , \DP_OP_751_130_6421/n1242 ,
         \DP_OP_751_130_6421/n1241 , \DP_OP_751_130_6421/n1240 ,
         \DP_OP_751_130_6421/n1239 , \DP_OP_751_130_6421/n1238 ,
         \DP_OP_751_130_6421/n1237 , \DP_OP_751_130_6421/n1236 ,
         \DP_OP_751_130_6421/n1235 , \DP_OP_751_130_6421/n1234 ,
         \DP_OP_751_130_6421/n1209 , \DP_OP_751_130_6421/n1208 ,
         \DP_OP_751_130_6421/n1207 , \DP_OP_751_130_6421/n1206 ,
         \DP_OP_751_130_6421/n1205 , \DP_OP_751_130_6421/n1204 ,
         \DP_OP_751_130_6421/n1203 , \DP_OP_751_130_6421/n1202 ,
         \DP_OP_751_130_6421/n1201 , \DP_OP_751_130_6421/n1200 ,
         \DP_OP_751_130_6421/n1199 , \DP_OP_751_130_6421/n1198 ,
         \DP_OP_751_130_6421/n1197 , \DP_OP_751_130_6421/n1196 ,
         \DP_OP_751_130_6421/n1195 , \DP_OP_751_130_6421/n1194 ,
         \DP_OP_751_130_6421/n1193 , \DP_OP_751_130_6421/n1192 ,
         \DP_OP_751_130_6421/n1191 , \DP_OP_751_130_6421/n1190 ,
         \DP_OP_751_130_6421/n1189 , \DP_OP_751_130_6421/n1174 ,
         \DP_OP_751_130_6421/n1173 , \DP_OP_751_130_6421/n1172 ,
         \DP_OP_751_130_6421/n1171 , \DP_OP_751_130_6421/n1170 ,
         \DP_OP_751_130_6421/n1169 , \DP_OP_751_130_6421/n1168 ,
         \DP_OP_751_130_6421/n1167 , \DP_OP_751_130_6421/n1166 ,
         \DP_OP_751_130_6421/n1165 , \DP_OP_751_130_6421/n1164 ,
         \DP_OP_751_130_6421/n1163 , \DP_OP_751_130_6421/n1162 ,
         \DP_OP_751_130_6421/n1161 , \DP_OP_751_130_6421/n1160 ,
         \DP_OP_751_130_6421/n1159 , \DP_OP_751_130_6421/n1158 ,
         \DP_OP_751_130_6421/n1157 , \DP_OP_751_130_6421/n1156 ,
         \DP_OP_751_130_6421/n1155 , \DP_OP_751_130_6421/n1154 ,
         \DP_OP_751_130_6421/n1153 , \DP_OP_751_130_6421/n1152 ,
         \DP_OP_751_130_6421/n1151 , \DP_OP_751_130_6421/n1150 ,
         \DP_OP_751_130_6421/n1149 , \DP_OP_751_130_6421/n1148 ,
         \DP_OP_751_130_6421/n1147 , \DP_OP_751_130_6421/n1146 ,
         \DP_OP_751_130_6421/n1145 , \DP_OP_751_130_6421/n1144 ,
         \DP_OP_751_130_6421/n1143 , \DP_OP_751_130_6421/n1142 ,
         \DP_OP_751_130_6421/n1141 , \DP_OP_751_130_6421/n1140 ,
         \DP_OP_751_130_6421/n1139 , \DP_OP_751_130_6421/n1138 ,
         \DP_OP_751_130_6421/n1137 , \DP_OP_751_130_6421/n1136 ,
         \DP_OP_751_130_6421/n1107 , \DP_OP_751_130_6421/n1106 ,
         \DP_OP_751_130_6421/n1105 , \DP_OP_751_130_6421/n1104 ,
         \DP_OP_751_130_6421/n1103 , \DP_OP_751_130_6421/n1102 ,
         \DP_OP_751_130_6421/n1101 , \DP_OP_751_130_6421/n1100 ,
         \DP_OP_751_130_6421/n1099 , \DP_OP_751_130_6421/n1098 ,
         \DP_OP_751_130_6421/n1097 , \DP_OP_751_130_6421/n1096 ,
         \DP_OP_751_130_6421/n1095 , \DP_OP_751_130_6421/n1094 ,
         \DP_OP_751_130_6421/n1093 , \DP_OP_751_130_6421/n1092 ,
         \DP_OP_751_130_6421/n1091 , \DP_OP_751_130_6421/n1090 ,
         \DP_OP_751_130_6421/n1089 , \DP_OP_751_130_6421/n1072 ,
         \DP_OP_751_130_6421/n1071 , \DP_OP_751_130_6421/n1070 ,
         \DP_OP_751_130_6421/n1069 , \DP_OP_751_130_6421/n1068 ,
         \DP_OP_751_130_6421/n1067 , \DP_OP_751_130_6421/n1066 ,
         \DP_OP_751_130_6421/n1065 , \DP_OP_751_130_6421/n1064 ,
         \DP_OP_751_130_6421/n1063 , \DP_OP_751_130_6421/n1062 ,
         \DP_OP_751_130_6421/n1061 , \DP_OP_751_130_6421/n1060 ,
         \DP_OP_751_130_6421/n1059 , \DP_OP_751_130_6421/n1058 ,
         \DP_OP_751_130_6421/n1057 , \DP_OP_751_130_6421/n1056 ,
         \DP_OP_751_130_6421/n1055 , \DP_OP_751_130_6421/n1054 ,
         \DP_OP_751_130_6421/n1053 , \DP_OP_751_130_6421/n1052 ,
         \DP_OP_751_130_6421/n1051 , \DP_OP_751_130_6421/n1050 ,
         \DP_OP_751_130_6421/n1049 , \DP_OP_751_130_6421/n1048 ,
         \DP_OP_751_130_6421/n1047 , \DP_OP_751_130_6421/n1046 ,
         \DP_OP_751_130_6421/n1045 , \DP_OP_751_130_6421/n1044 ,
         \DP_OP_751_130_6421/n1043 , \DP_OP_751_130_6421/n1042 ,
         \DP_OP_751_130_6421/n1041 , \DP_OP_751_130_6421/n1040 ,
         \DP_OP_751_130_6421/n1039 , \DP_OP_751_130_6421/n1038 ,
         \DP_OP_751_130_6421/n1005 , \DP_OP_751_130_6421/n1004 ,
         \DP_OP_751_130_6421/n1003 , \DP_OP_751_130_6421/n1002 ,
         \DP_OP_751_130_6421/n1001 , \DP_OP_751_130_6421/n1000 ,
         \DP_OP_751_130_6421/n999 , \DP_OP_751_130_6421/n998 ,
         \DP_OP_751_130_6421/n997 , \DP_OP_751_130_6421/n996 ,
         \DP_OP_751_130_6421/n995 , \DP_OP_751_130_6421/n994 ,
         \DP_OP_751_130_6421/n993 , \DP_OP_751_130_6421/n992 ,
         \DP_OP_751_130_6421/n991 , \DP_OP_751_130_6421/n990 ,
         \DP_OP_751_130_6421/n989 , \DP_OP_751_130_6421/n970 ,
         \DP_OP_751_130_6421/n969 , \DP_OP_751_130_6421/n968 ,
         \DP_OP_751_130_6421/n967 , \DP_OP_751_130_6421/n966 ,
         \DP_OP_751_130_6421/n965 , \DP_OP_751_130_6421/n964 ,
         \DP_OP_751_130_6421/n963 , \DP_OP_751_130_6421/n962 ,
         \DP_OP_751_130_6421/n961 , \DP_OP_751_130_6421/n960 ,
         \DP_OP_751_130_6421/n959 , \DP_OP_751_130_6421/n958 ,
         \DP_OP_751_130_6421/n957 , \DP_OP_751_130_6421/n956 ,
         \DP_OP_751_130_6421/n955 , \DP_OP_751_130_6421/n954 ,
         \DP_OP_751_130_6421/n953 , \DP_OP_751_130_6421/n952 ,
         \DP_OP_751_130_6421/n951 , \DP_OP_751_130_6421/n950 ,
         \DP_OP_751_130_6421/n949 , \DP_OP_751_130_6421/n948 ,
         \DP_OP_751_130_6421/n947 , \DP_OP_751_130_6421/n946 ,
         \DP_OP_751_130_6421/n945 , \DP_OP_751_130_6421/n944 ,
         \DP_OP_751_130_6421/n943 , \DP_OP_751_130_6421/n942 ,
         \DP_OP_751_130_6421/n941 , \DP_OP_751_130_6421/n940 ,
         \DP_OP_751_130_6421/n903 , \DP_OP_751_130_6421/n902 ,
         \DP_OP_751_130_6421/n901 , \DP_OP_751_130_6421/n900 ,
         \DP_OP_751_130_6421/n899 , \DP_OP_751_130_6421/n898 ,
         \DP_OP_751_130_6421/n897 , \DP_OP_751_130_6421/n896 ,
         \DP_OP_751_130_6421/n895 , \DP_OP_751_130_6421/n894 ,
         \DP_OP_751_130_6421/n893 , \DP_OP_751_130_6421/n892 ,
         \DP_OP_751_130_6421/n891 , \DP_OP_751_130_6421/n890 ,
         \DP_OP_751_130_6421/n889 , \DP_OP_751_130_6421/n868 ,
         \DP_OP_751_130_6421/n867 , \DP_OP_751_130_6421/n866 ,
         \DP_OP_751_130_6421/n865 , \DP_OP_751_130_6421/n864 ,
         \DP_OP_751_130_6421/n863 , \DP_OP_751_130_6421/n862 ,
         \DP_OP_751_130_6421/n861 , \DP_OP_751_130_6421/n860 ,
         \DP_OP_751_130_6421/n859 , \DP_OP_751_130_6421/n858 ,
         \DP_OP_751_130_6421/n857 , \DP_OP_751_130_6421/n856 ,
         \DP_OP_751_130_6421/n855 , \DP_OP_751_130_6421/n854 ,
         \DP_OP_751_130_6421/n853 , \DP_OP_751_130_6421/n852 ,
         \DP_OP_751_130_6421/n851 , \DP_OP_751_130_6421/n850 ,
         \DP_OP_751_130_6421/n849 , \DP_OP_751_130_6421/n848 ,
         \DP_OP_751_130_6421/n847 , \DP_OP_751_130_6421/n846 ,
         \DP_OP_751_130_6421/n845 , \DP_OP_751_130_6421/n844 ,
         \DP_OP_751_130_6421/n843 , \DP_OP_751_130_6421/n842 ,
         \DP_OP_751_130_6421/n801 , \DP_OP_751_130_6421/n800 ,
         \DP_OP_751_130_6421/n799 , \DP_OP_751_130_6421/n798 ,
         \DP_OP_751_130_6421/n797 , \DP_OP_751_130_6421/n796 ,
         \DP_OP_751_130_6421/n795 , \DP_OP_751_130_6421/n794 ,
         \DP_OP_751_130_6421/n793 , \DP_OP_751_130_6421/n792 ,
         \DP_OP_751_130_6421/n791 , \DP_OP_751_130_6421/n790 ,
         \DP_OP_751_130_6421/n789 , \DP_OP_751_130_6421/n766 ,
         \DP_OP_751_130_6421/n765 , \DP_OP_751_130_6421/n764 ,
         \DP_OP_751_130_6421/n763 , \DP_OP_751_130_6421/n762 ,
         \DP_OP_751_130_6421/n761 , \DP_OP_751_130_6421/n760 ,
         \DP_OP_751_130_6421/n759 , \DP_OP_751_130_6421/n758 ,
         \DP_OP_751_130_6421/n757 , \DP_OP_751_130_6421/n756 ,
         \DP_OP_751_130_6421/n755 , \DP_OP_751_130_6421/n754 ,
         \DP_OP_751_130_6421/n753 , \DP_OP_751_130_6421/n752 ,
         \DP_OP_751_130_6421/n751 , \DP_OP_751_130_6421/n750 ,
         \DP_OP_751_130_6421/n749 , \DP_OP_751_130_6421/n748 ,
         \DP_OP_751_130_6421/n747 , \DP_OP_751_130_6421/n746 ,
         \DP_OP_751_130_6421/n745 , \DP_OP_751_130_6421/n744 ,
         \DP_OP_751_130_6421/n699 , \DP_OP_751_130_6421/n698 ,
         \DP_OP_751_130_6421/n697 , \DP_OP_751_130_6421/n696 ,
         \DP_OP_751_130_6421/n695 , \DP_OP_751_130_6421/n694 ,
         \DP_OP_751_130_6421/n693 , \DP_OP_751_130_6421/n692 ,
         \DP_OP_751_130_6421/n691 , \DP_OP_751_130_6421/n690 ,
         \DP_OP_751_130_6421/n689 , \DP_OP_751_130_6421/n664 ,
         \DP_OP_751_130_6421/n663 , \DP_OP_751_130_6421/n662 ,
         \DP_OP_751_130_6421/n661 , \DP_OP_751_130_6421/n660 ,
         \DP_OP_751_130_6421/n659 , \DP_OP_751_130_6421/n658 ,
         \DP_OP_751_130_6421/n657 , \DP_OP_751_130_6421/n656 ,
         \DP_OP_751_130_6421/n655 , \DP_OP_751_130_6421/n654 ,
         \DP_OP_751_130_6421/n653 , \DP_OP_751_130_6421/n652 ,
         \DP_OP_751_130_6421/n651 , \DP_OP_751_130_6421/n650 ,
         \DP_OP_751_130_6421/n649 , \DP_OP_751_130_6421/n648 ,
         \DP_OP_751_130_6421/n647 , \DP_OP_751_130_6421/n646 ,
         \DP_OP_751_130_6421/n597 , \DP_OP_751_130_6421/n596 ,
         \DP_OP_751_130_6421/n595 , \DP_OP_751_130_6421/n594 ,
         \DP_OP_751_130_6421/n593 , \DP_OP_751_130_6421/n592 ,
         \DP_OP_751_130_6421/n591 , \DP_OP_751_130_6421/n590 ,
         \DP_OP_751_130_6421/n589 , \DP_OP_751_130_6421/n562 ,
         \DP_OP_751_130_6421/n561 , \DP_OP_751_130_6421/n560 ,
         \DP_OP_751_130_6421/n559 , \DP_OP_751_130_6421/n558 ,
         \DP_OP_751_130_6421/n557 , \DP_OP_751_130_6421/n556 ,
         \DP_OP_751_130_6421/n555 , \DP_OP_751_130_6421/n554 ,
         \DP_OP_751_130_6421/n553 , \DP_OP_751_130_6421/n552 ,
         \DP_OP_751_130_6421/n551 , \DP_OP_751_130_6421/n550 ,
         \DP_OP_751_130_6421/n549 , \DP_OP_751_130_6421/n548 ,
         \DP_OP_751_130_6421/n495 , \DP_OP_751_130_6421/n494 ,
         \DP_OP_751_130_6421/n493 , \DP_OP_751_130_6421/n492 ,
         \DP_OP_751_130_6421/n491 , \DP_OP_751_130_6421/n490 ,
         \DP_OP_751_130_6421/n489 , \DP_OP_751_130_6421/n460 ,
         \DP_OP_751_130_6421/n459 , \DP_OP_751_130_6421/n458 ,
         \DP_OP_751_130_6421/n457 , \DP_OP_751_130_6421/n456 ,
         \DP_OP_751_130_6421/n455 , \DP_OP_751_130_6421/n454 ,
         \DP_OP_751_130_6421/n453 , \DP_OP_751_130_6421/n452 ,
         \DP_OP_751_130_6421/n451 , \DP_OP_751_130_6421/n450 ,
         \DP_OP_751_130_6421/n393 , \DP_OP_751_130_6421/n392 ,
         \DP_OP_751_130_6421/n391 , \DP_OP_751_130_6421/n390 ,
         \DP_OP_751_130_6421/n389 , \DP_OP_751_130_6421/n358 ,
         \DP_OP_751_130_6421/n357 , \DP_OP_751_130_6421/n356 ,
         \DP_OP_751_130_6421/n355 , \DP_OP_751_130_6421/n354 ,
         \DP_OP_751_130_6421/n353 , \DP_OP_751_130_6421/n352 ,
         \DP_OP_751_130_6421/n291 , \DP_OP_751_130_6421/n290 ,
         \DP_OP_751_130_6421/n185 , \DP_OP_751_130_6421/n183 ,
         \DP_OP_751_130_6421/n181 , \DP_OP_751_130_6421/n176 ,
         \DP_OP_751_130_6421/n173 , \DP_OP_751_130_6421/n171 ,
         \DP_OP_751_130_6421/n169 , \DP_OP_751_130_6421/n165 ,
         \DP_OP_751_130_6421/n164 , \DP_OP_751_130_6421/n163 ,
         \DP_OP_751_130_6421/n161 , \DP_OP_751_130_6421/n159 ,
         \DP_OP_751_130_6421/n158 , \DP_OP_751_130_6421/n155 ,
         \DP_OP_751_130_6421/n154 , \DP_OP_751_130_6421/n153 ,
         \DP_OP_751_130_6421/n152 , \DP_OP_751_130_6421/n151 ,
         \DP_OP_751_130_6421/n150 , \DP_OP_751_130_6421/n148 ,
         \DP_OP_751_130_6421/n147 , \DP_OP_751_130_6421/n146 ,
         \DP_OP_751_130_6421/n145 , \DP_OP_751_130_6421/n144 ,
         \DP_OP_751_130_6421/n142 , \DP_OP_751_130_6421/n140 ,
         \DP_OP_751_130_6421/n139 , \DP_OP_751_130_6421/n138 ,
         \DP_OP_751_130_6421/n137 , \DP_OP_751_130_6421/n136 ,
         \DP_OP_751_130_6421/n134 , \DP_OP_751_130_6421/n132 ,
         \DP_OP_751_130_6421/n131 , \DP_OP_751_130_6421/n130 ,
         \DP_OP_751_130_6421/n129 , \DP_OP_751_130_6421/n128 ,
         \DP_OP_751_130_6421/n126 , \DP_OP_751_130_6421/n124 ,
         \DP_OP_751_130_6421/n123 , \DP_OP_751_130_6421/n122 ,
         \DP_OP_751_130_6421/n120 , \DP_OP_751_130_6421/n118 ,
         \DP_OP_751_130_6421/n117 , \DP_OP_751_130_6421/n116 ,
         \DP_OP_751_130_6421/n115 , \DP_OP_751_130_6421/n114 ,
         \DP_OP_751_130_6421/n112 , \DP_OP_751_130_6421/n110 ,
         \DP_OP_751_130_6421/n109 , \DP_OP_751_130_6421/n108 ,
         \DP_OP_751_130_6421/n107 , \DP_OP_751_130_6421/n106 ,
         \DP_OP_751_130_6421/n104 , \DP_OP_751_130_6421/n102 ,
         \DP_OP_751_130_6421/n101 , \DP_OP_751_130_6421/n100 ,
         \DP_OP_751_130_6421/n99 , \DP_OP_751_130_6421/n98 ,
         \DP_OP_751_130_6421/n97 , \DP_OP_751_130_6421/n96 ,
         \DP_OP_751_130_6421/n95 , \DP_OP_751_130_6421/n94 ,
         \DP_OP_751_130_6421/n92 , \DP_OP_751_130_6421/n90 ,
         \DP_OP_751_130_6421/n89 , \DP_OP_751_130_6421/n88 ,
         \DP_OP_751_130_6421/n87 , \DP_OP_751_130_6421/n86 ,
         \DP_OP_751_130_6421/n84 , \DP_OP_751_130_6421/n82 ,
         \DP_OP_751_130_6421/n81 , \DP_OP_751_130_6421/n80 ,
         \DP_OP_751_130_6421/n79 , \DP_OP_751_130_6421/n78 ,
         \DP_OP_751_130_6421/n74 , \DP_OP_751_130_6421/n73 ,
         \DP_OP_751_130_6421/n72 , \DP_OP_751_130_6421/n71 ,
         \DP_OP_751_130_6421/n66 , \DP_OP_751_130_6421/n64 ,
         \DP_OP_751_130_6421/n62 , \DP_OP_751_130_6421/n61 ,
         \DP_OP_751_130_6421/n60 , \DP_OP_751_130_6421/n22 ,
         \DP_OP_751_130_6421/n20 , \DP_OP_751_130_6421/n18 ,
         \DP_OP_751_130_6421/n17 , \DP_OP_751_130_6421/n16 ,
         \DP_OP_751_130_6421/n13 , \DP_OP_751_130_6421/n10 ,
         \DP_OP_751_130_6421/n9 , \DP_OP_751_130_6421/n8 ,
         \DP_OP_751_130_6421/n7 , \DP_OP_751_130_6421/n6 ,
         \DP_OP_751_130_6421/n5 , \DP_OP_751_130_6421/n4 , n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852;
  wire   [31:0] IR;
  wire   [4:0] i_ALU_OP;
  wire   [4:0] i_ADD_WB;
  wire   [31:0] i_RD1;
  wire   [31:0] i_RD2;
  wire   [4:0] i_ADD_RS1;
  wire   [4:0] i_ADD_RS2;
  wire   [4:0] i_ADD_WS1;
  assign IRAM_ISSUE = 1'b1;
  assign DRAMRF_ADDRESS[1] = 1'b0;
  assign DATA_SIZE_RF[1] = 1'b0;
  assign DATA_SIZE_RF[0] = 1'b0;
  assign DRAMRF_ADDRESS[0] = 1'b0;

  hazard_table_N_REGS_LOG5 \DECODEhw/HAZARD_CTRL  ( .CLK(CLK), .RST(RST), 
        .WR1(\DECODEhw/i_WR1 ), .WR2(i_WF), .ADD_WR1(i_ADD_WS1), .ADD_WR2(
        i_ADD_WB), .ADD_CHECK1(i_ADD_RS1), .ADD_CHECK2(i_ADD_RS2), .BUSY(
        i_HAZARD_SIG_CU), .BUSY_WINDOW(i_BUSY_WINDOW) );
  in_loc_selblock_NBIT_DATA32_N8_F5 \DataPath/RF/SELBLOCK_INLOC  ( .regs({
        \DataPath/RF/bus_reg_dataout[2559] , 
        \DataPath/RF/bus_reg_dataout[2558] , 
        \DataPath/RF/bus_reg_dataout[2557] , 
        \DataPath/RF/bus_reg_dataout[2556] , 
        \DataPath/RF/bus_reg_dataout[2555] , 
        \DataPath/RF/bus_reg_dataout[2554] , 
        \DataPath/RF/bus_reg_dataout[2553] , 
        \DataPath/RF/bus_reg_dataout[2552] , 
        \DataPath/RF/bus_reg_dataout[2551] , 
        \DataPath/RF/bus_reg_dataout[2550] , 
        \DataPath/RF/bus_reg_dataout[2549] , 
        \DataPath/RF/bus_reg_dataout[2548] , 
        \DataPath/RF/bus_reg_dataout[2547] , 
        \DataPath/RF/bus_reg_dataout[2546] , 
        \DataPath/RF/bus_reg_dataout[2545] , 
        \DataPath/RF/bus_reg_dataout[2544] , 
        \DataPath/RF/bus_reg_dataout[2543] , 
        \DataPath/RF/bus_reg_dataout[2542] , 
        \DataPath/RF/bus_reg_dataout[2541] , 
        \DataPath/RF/bus_reg_dataout[2540] , 
        \DataPath/RF/bus_reg_dataout[2539] , 
        \DataPath/RF/bus_reg_dataout[2538] , 
        \DataPath/RF/bus_reg_dataout[2537] , 
        \DataPath/RF/bus_reg_dataout[2536] , 
        \DataPath/RF/bus_reg_dataout[2535] , 
        \DataPath/RF/bus_reg_dataout[2534] , 
        \DataPath/RF/bus_reg_dataout[2533] , 
        \DataPath/RF/bus_reg_dataout[2532] , 
        \DataPath/RF/bus_reg_dataout[2531] , 
        \DataPath/RF/bus_reg_dataout[2530] , 
        \DataPath/RF/bus_reg_dataout[2529] , 
        \DataPath/RF/bus_reg_dataout[2528] , 
        \DataPath/RF/bus_reg_dataout[2527] , 
        \DataPath/RF/bus_reg_dataout[2526] , 
        \DataPath/RF/bus_reg_dataout[2525] , 
        \DataPath/RF/bus_reg_dataout[2524] , 
        \DataPath/RF/bus_reg_dataout[2523] , 
        \DataPath/RF/bus_reg_dataout[2522] , 
        \DataPath/RF/bus_reg_dataout[2521] , 
        \DataPath/RF/bus_reg_dataout[2520] , 
        \DataPath/RF/bus_reg_dataout[2519] , 
        \DataPath/RF/bus_reg_dataout[2518] , 
        \DataPath/RF/bus_reg_dataout[2517] , 
        \DataPath/RF/bus_reg_dataout[2516] , 
        \DataPath/RF/bus_reg_dataout[2515] , 
        \DataPath/RF/bus_reg_dataout[2514] , 
        \DataPath/RF/bus_reg_dataout[2513] , 
        \DataPath/RF/bus_reg_dataout[2512] , 
        \DataPath/RF/bus_reg_dataout[2511] , 
        \DataPath/RF/bus_reg_dataout[2510] , 
        \DataPath/RF/bus_reg_dataout[2509] , 
        \DataPath/RF/bus_reg_dataout[2508] , 
        \DataPath/RF/bus_reg_dataout[2507] , 
        \DataPath/RF/bus_reg_dataout[2506] , 
        \DataPath/RF/bus_reg_dataout[2505] , 
        \DataPath/RF/bus_reg_dataout[2504] , 
        \DataPath/RF/bus_reg_dataout[2503] , 
        \DataPath/RF/bus_reg_dataout[2502] , 
        \DataPath/RF/bus_reg_dataout[2501] , 
        \DataPath/RF/bus_reg_dataout[2500] , 
        \DataPath/RF/bus_reg_dataout[2499] , 
        \DataPath/RF/bus_reg_dataout[2498] , 
        \DataPath/RF/bus_reg_dataout[2497] , 
        \DataPath/RF/bus_reg_dataout[2496] , 
        \DataPath/RF/bus_reg_dataout[2495] , 
        \DataPath/RF/bus_reg_dataout[2494] , 
        \DataPath/RF/bus_reg_dataout[2493] , 
        \DataPath/RF/bus_reg_dataout[2492] , 
        \DataPath/RF/bus_reg_dataout[2491] , 
        \DataPath/RF/bus_reg_dataout[2490] , 
        \DataPath/RF/bus_reg_dataout[2489] , 
        \DataPath/RF/bus_reg_dataout[2488] , 
        \DataPath/RF/bus_reg_dataout[2487] , 
        \DataPath/RF/bus_reg_dataout[2486] , 
        \DataPath/RF/bus_reg_dataout[2485] , 
        \DataPath/RF/bus_reg_dataout[2484] , 
        \DataPath/RF/bus_reg_dataout[2483] , 
        \DataPath/RF/bus_reg_dataout[2482] , 
        \DataPath/RF/bus_reg_dataout[2481] , 
        \DataPath/RF/bus_reg_dataout[2480] , 
        \DataPath/RF/bus_reg_dataout[2479] , 
        \DataPath/RF/bus_reg_dataout[2478] , 
        \DataPath/RF/bus_reg_dataout[2477] , 
        \DataPath/RF/bus_reg_dataout[2476] , 
        \DataPath/RF/bus_reg_dataout[2475] , 
        \DataPath/RF/bus_reg_dataout[2474] , 
        \DataPath/RF/bus_reg_dataout[2473] , 
        \DataPath/RF/bus_reg_dataout[2472] , 
        \DataPath/RF/bus_reg_dataout[2471] , 
        \DataPath/RF/bus_reg_dataout[2470] , 
        \DataPath/RF/bus_reg_dataout[2469] , 
        \DataPath/RF/bus_reg_dataout[2468] , 
        \DataPath/RF/bus_reg_dataout[2467] , 
        \DataPath/RF/bus_reg_dataout[2466] , 
        \DataPath/RF/bus_reg_dataout[2465] , 
        \DataPath/RF/bus_reg_dataout[2464] , 
        \DataPath/RF/bus_reg_dataout[2463] , 
        \DataPath/RF/bus_reg_dataout[2462] , 
        \DataPath/RF/bus_reg_dataout[2461] , 
        \DataPath/RF/bus_reg_dataout[2460] , 
        \DataPath/RF/bus_reg_dataout[2459] , 
        \DataPath/RF/bus_reg_dataout[2458] , 
        \DataPath/RF/bus_reg_dataout[2457] , 
        \DataPath/RF/bus_reg_dataout[2456] , 
        \DataPath/RF/bus_reg_dataout[2455] , 
        \DataPath/RF/bus_reg_dataout[2454] , 
        \DataPath/RF/bus_reg_dataout[2453] , 
        \DataPath/RF/bus_reg_dataout[2452] , 
        \DataPath/RF/bus_reg_dataout[2451] , 
        \DataPath/RF/bus_reg_dataout[2450] , 
        \DataPath/RF/bus_reg_dataout[2449] , 
        \DataPath/RF/bus_reg_dataout[2448] , 
        \DataPath/RF/bus_reg_dataout[2447] , 
        \DataPath/RF/bus_reg_dataout[2446] , 
        \DataPath/RF/bus_reg_dataout[2445] , 
        \DataPath/RF/bus_reg_dataout[2444] , 
        \DataPath/RF/bus_reg_dataout[2443] , 
        \DataPath/RF/bus_reg_dataout[2442] , 
        \DataPath/RF/bus_reg_dataout[2441] , 
        \DataPath/RF/bus_reg_dataout[2440] , 
        \DataPath/RF/bus_reg_dataout[2439] , 
        \DataPath/RF/bus_reg_dataout[2438] , 
        \DataPath/RF/bus_reg_dataout[2437] , 
        \DataPath/RF/bus_reg_dataout[2436] , 
        \DataPath/RF/bus_reg_dataout[2435] , 
        \DataPath/RF/bus_reg_dataout[2434] , 
        \DataPath/RF/bus_reg_dataout[2433] , 
        \DataPath/RF/bus_reg_dataout[2432] , 
        \DataPath/RF/bus_reg_dataout[2431] , 
        \DataPath/RF/bus_reg_dataout[2430] , 
        \DataPath/RF/bus_reg_dataout[2429] , 
        \DataPath/RF/bus_reg_dataout[2428] , 
        \DataPath/RF/bus_reg_dataout[2427] , 
        \DataPath/RF/bus_reg_dataout[2426] , 
        \DataPath/RF/bus_reg_dataout[2425] , 
        \DataPath/RF/bus_reg_dataout[2424] , 
        \DataPath/RF/bus_reg_dataout[2423] , 
        \DataPath/RF/bus_reg_dataout[2422] , 
        \DataPath/RF/bus_reg_dataout[2421] , 
        \DataPath/RF/bus_reg_dataout[2420] , 
        \DataPath/RF/bus_reg_dataout[2419] , 
        \DataPath/RF/bus_reg_dataout[2418] , 
        \DataPath/RF/bus_reg_dataout[2417] , 
        \DataPath/RF/bus_reg_dataout[2416] , 
        \DataPath/RF/bus_reg_dataout[2415] , 
        \DataPath/RF/bus_reg_dataout[2414] , 
        \DataPath/RF/bus_reg_dataout[2413] , 
        \DataPath/RF/bus_reg_dataout[2412] , 
        \DataPath/RF/bus_reg_dataout[2411] , 
        \DataPath/RF/bus_reg_dataout[2410] , 
        \DataPath/RF/bus_reg_dataout[2409] , 
        \DataPath/RF/bus_reg_dataout[2408] , 
        \DataPath/RF/bus_reg_dataout[2407] , 
        \DataPath/RF/bus_reg_dataout[2406] , 
        \DataPath/RF/bus_reg_dataout[2405] , 
        \DataPath/RF/bus_reg_dataout[2404] , 
        \DataPath/RF/bus_reg_dataout[2403] , 
        \DataPath/RF/bus_reg_dataout[2402] , 
        \DataPath/RF/bus_reg_dataout[2401] , 
        \DataPath/RF/bus_reg_dataout[2400] , 
        \DataPath/RF/bus_reg_dataout[2399] , 
        \DataPath/RF/bus_reg_dataout[2398] , 
        \DataPath/RF/bus_reg_dataout[2397] , 
        \DataPath/RF/bus_reg_dataout[2396] , 
        \DataPath/RF/bus_reg_dataout[2395] , 
        \DataPath/RF/bus_reg_dataout[2394] , 
        \DataPath/RF/bus_reg_dataout[2393] , 
        \DataPath/RF/bus_reg_dataout[2392] , 
        \DataPath/RF/bus_reg_dataout[2391] , 
        \DataPath/RF/bus_reg_dataout[2390] , 
        \DataPath/RF/bus_reg_dataout[2389] , 
        \DataPath/RF/bus_reg_dataout[2388] , 
        \DataPath/RF/bus_reg_dataout[2387] , 
        \DataPath/RF/bus_reg_dataout[2386] , 
        \DataPath/RF/bus_reg_dataout[2385] , 
        \DataPath/RF/bus_reg_dataout[2384] , 
        \DataPath/RF/bus_reg_dataout[2383] , 
        \DataPath/RF/bus_reg_dataout[2382] , 
        \DataPath/RF/bus_reg_dataout[2381] , 
        \DataPath/RF/bus_reg_dataout[2380] , 
        \DataPath/RF/bus_reg_dataout[2379] , 
        \DataPath/RF/bus_reg_dataout[2378] , 
        \DataPath/RF/bus_reg_dataout[2377] , 
        \DataPath/RF/bus_reg_dataout[2376] , 
        \DataPath/RF/bus_reg_dataout[2375] , 
        \DataPath/RF/bus_reg_dataout[2374] , 
        \DataPath/RF/bus_reg_dataout[2373] , 
        \DataPath/RF/bus_reg_dataout[2372] , 
        \DataPath/RF/bus_reg_dataout[2371] , 
        \DataPath/RF/bus_reg_dataout[2370] , 
        \DataPath/RF/bus_reg_dataout[2369] , 
        \DataPath/RF/bus_reg_dataout[2368] , 
        \DataPath/RF/bus_reg_dataout[2367] , 
        \DataPath/RF/bus_reg_dataout[2366] , 
        \DataPath/RF/bus_reg_dataout[2365] , 
        \DataPath/RF/bus_reg_dataout[2364] , 
        \DataPath/RF/bus_reg_dataout[2363] , 
        \DataPath/RF/bus_reg_dataout[2362] , 
        \DataPath/RF/bus_reg_dataout[2361] , 
        \DataPath/RF/bus_reg_dataout[2360] , 
        \DataPath/RF/bus_reg_dataout[2359] , 
        \DataPath/RF/bus_reg_dataout[2358] , 
        \DataPath/RF/bus_reg_dataout[2357] , 
        \DataPath/RF/bus_reg_dataout[2356] , 
        \DataPath/RF/bus_reg_dataout[2355] , 
        \DataPath/RF/bus_reg_dataout[2354] , 
        \DataPath/RF/bus_reg_dataout[2353] , 
        \DataPath/RF/bus_reg_dataout[2352] , 
        \DataPath/RF/bus_reg_dataout[2351] , 
        \DataPath/RF/bus_reg_dataout[2350] , 
        \DataPath/RF/bus_reg_dataout[2349] , 
        \DataPath/RF/bus_reg_dataout[2348] , 
        \DataPath/RF/bus_reg_dataout[2347] , 
        \DataPath/RF/bus_reg_dataout[2346] , 
        \DataPath/RF/bus_reg_dataout[2345] , 
        \DataPath/RF/bus_reg_dataout[2344] , 
        \DataPath/RF/bus_reg_dataout[2343] , 
        \DataPath/RF/bus_reg_dataout[2342] , 
        \DataPath/RF/bus_reg_dataout[2341] , 
        \DataPath/RF/bus_reg_dataout[2340] , 
        \DataPath/RF/bus_reg_dataout[2339] , 
        \DataPath/RF/bus_reg_dataout[2338] , 
        \DataPath/RF/bus_reg_dataout[2337] , 
        \DataPath/RF/bus_reg_dataout[2336] , 
        \DataPath/RF/bus_reg_dataout[2335] , 
        \DataPath/RF/bus_reg_dataout[2334] , 
        \DataPath/RF/bus_reg_dataout[2333] , 
        \DataPath/RF/bus_reg_dataout[2332] , 
        \DataPath/RF/bus_reg_dataout[2331] , 
        \DataPath/RF/bus_reg_dataout[2330] , 
        \DataPath/RF/bus_reg_dataout[2329] , 
        \DataPath/RF/bus_reg_dataout[2328] , 
        \DataPath/RF/bus_reg_dataout[2327] , 
        \DataPath/RF/bus_reg_dataout[2326] , 
        \DataPath/RF/bus_reg_dataout[2325] , 
        \DataPath/RF/bus_reg_dataout[2324] , 
        \DataPath/RF/bus_reg_dataout[2323] , 
        \DataPath/RF/bus_reg_dataout[2322] , 
        \DataPath/RF/bus_reg_dataout[2321] , 
        \DataPath/RF/bus_reg_dataout[2320] , 
        \DataPath/RF/bus_reg_dataout[2319] , 
        \DataPath/RF/bus_reg_dataout[2318] , 
        \DataPath/RF/bus_reg_dataout[2317] , 
        \DataPath/RF/bus_reg_dataout[2316] , 
        \DataPath/RF/bus_reg_dataout[2315] , 
        \DataPath/RF/bus_reg_dataout[2314] , 
        \DataPath/RF/bus_reg_dataout[2313] , 
        \DataPath/RF/bus_reg_dataout[2312] , 
        \DataPath/RF/bus_reg_dataout[2311] , 
        \DataPath/RF/bus_reg_dataout[2310] , 
        \DataPath/RF/bus_reg_dataout[2309] , 
        \DataPath/RF/bus_reg_dataout[2308] , 
        \DataPath/RF/bus_reg_dataout[2307] , 
        \DataPath/RF/bus_reg_dataout[2306] , 
        \DataPath/RF/bus_reg_dataout[2305] , 
        \DataPath/RF/bus_reg_dataout[2304] , 
        \DataPath/RF/bus_reg_dataout[2303] , 
        \DataPath/RF/bus_reg_dataout[2302] , 
        \DataPath/RF/bus_reg_dataout[2301] , 
        \DataPath/RF/bus_reg_dataout[2300] , 
        \DataPath/RF/bus_reg_dataout[2299] , 
        \DataPath/RF/bus_reg_dataout[2298] , 
        \DataPath/RF/bus_reg_dataout[2297] , 
        \DataPath/RF/bus_reg_dataout[2296] , 
        \DataPath/RF/bus_reg_dataout[2295] , 
        \DataPath/RF/bus_reg_dataout[2294] , 
        \DataPath/RF/bus_reg_dataout[2293] , 
        \DataPath/RF/bus_reg_dataout[2292] , 
        \DataPath/RF/bus_reg_dataout[2291] , 
        \DataPath/RF/bus_reg_dataout[2290] , 
        \DataPath/RF/bus_reg_dataout[2289] , 
        \DataPath/RF/bus_reg_dataout[2288] , 
        \DataPath/RF/bus_reg_dataout[2287] , 
        \DataPath/RF/bus_reg_dataout[2286] , 
        \DataPath/RF/bus_reg_dataout[2285] , 
        \DataPath/RF/bus_reg_dataout[2284] , 
        \DataPath/RF/bus_reg_dataout[2283] , 
        \DataPath/RF/bus_reg_dataout[2282] , 
        \DataPath/RF/bus_reg_dataout[2281] , 
        \DataPath/RF/bus_reg_dataout[2280] , 
        \DataPath/RF/bus_reg_dataout[2279] , 
        \DataPath/RF/bus_reg_dataout[2278] , 
        \DataPath/RF/bus_reg_dataout[2277] , 
        \DataPath/RF/bus_reg_dataout[2276] , 
        \DataPath/RF/bus_reg_dataout[2275] , 
        \DataPath/RF/bus_reg_dataout[2274] , 
        \DataPath/RF/bus_reg_dataout[2273] , 
        \DataPath/RF/bus_reg_dataout[2272] , 
        \DataPath/RF/bus_reg_dataout[2271] , 
        \DataPath/RF/bus_reg_dataout[2270] , 
        \DataPath/RF/bus_reg_dataout[2269] , 
        \DataPath/RF/bus_reg_dataout[2268] , 
        \DataPath/RF/bus_reg_dataout[2267] , 
        \DataPath/RF/bus_reg_dataout[2266] , 
        \DataPath/RF/bus_reg_dataout[2265] , 
        \DataPath/RF/bus_reg_dataout[2264] , 
        \DataPath/RF/bus_reg_dataout[2263] , 
        \DataPath/RF/bus_reg_dataout[2262] , 
        \DataPath/RF/bus_reg_dataout[2261] , 
        \DataPath/RF/bus_reg_dataout[2260] , 
        \DataPath/RF/bus_reg_dataout[2259] , 
        \DataPath/RF/bus_reg_dataout[2258] , 
        \DataPath/RF/bus_reg_dataout[2257] , 
        \DataPath/RF/bus_reg_dataout[2256] , 
        \DataPath/RF/bus_reg_dataout[2255] , 
        \DataPath/RF/bus_reg_dataout[2254] , 
        \DataPath/RF/bus_reg_dataout[2253] , 
        \DataPath/RF/bus_reg_dataout[2252] , 
        \DataPath/RF/bus_reg_dataout[2251] , 
        \DataPath/RF/bus_reg_dataout[2250] , 
        \DataPath/RF/bus_reg_dataout[2249] , 
        \DataPath/RF/bus_reg_dataout[2248] , 
        \DataPath/RF/bus_reg_dataout[2247] , 
        \DataPath/RF/bus_reg_dataout[2246] , 
        \DataPath/RF/bus_reg_dataout[2245] , 
        \DataPath/RF/bus_reg_dataout[2244] , 
        \DataPath/RF/bus_reg_dataout[2243] , 
        \DataPath/RF/bus_reg_dataout[2242] , 
        \DataPath/RF/bus_reg_dataout[2241] , 
        \DataPath/RF/bus_reg_dataout[2240] , 
        \DataPath/RF/bus_reg_dataout[2239] , 
        \DataPath/RF/bus_reg_dataout[2238] , 
        \DataPath/RF/bus_reg_dataout[2237] , 
        \DataPath/RF/bus_reg_dataout[2236] , 
        \DataPath/RF/bus_reg_dataout[2235] , 
        \DataPath/RF/bus_reg_dataout[2234] , 
        \DataPath/RF/bus_reg_dataout[2233] , 
        \DataPath/RF/bus_reg_dataout[2232] , 
        \DataPath/RF/bus_reg_dataout[2231] , 
        \DataPath/RF/bus_reg_dataout[2230] , 
        \DataPath/RF/bus_reg_dataout[2229] , 
        \DataPath/RF/bus_reg_dataout[2228] , 
        \DataPath/RF/bus_reg_dataout[2227] , 
        \DataPath/RF/bus_reg_dataout[2226] , 
        \DataPath/RF/bus_reg_dataout[2225] , 
        \DataPath/RF/bus_reg_dataout[2224] , 
        \DataPath/RF/bus_reg_dataout[2223] , 
        \DataPath/RF/bus_reg_dataout[2222] , 
        \DataPath/RF/bus_reg_dataout[2221] , 
        \DataPath/RF/bus_reg_dataout[2220] , 
        \DataPath/RF/bus_reg_dataout[2219] , 
        \DataPath/RF/bus_reg_dataout[2218] , 
        \DataPath/RF/bus_reg_dataout[2217] , 
        \DataPath/RF/bus_reg_dataout[2216] , 
        \DataPath/RF/bus_reg_dataout[2215] , 
        \DataPath/RF/bus_reg_dataout[2214] , 
        \DataPath/RF/bus_reg_dataout[2213] , 
        \DataPath/RF/bus_reg_dataout[2212] , 
        \DataPath/RF/bus_reg_dataout[2211] , 
        \DataPath/RF/bus_reg_dataout[2210] , 
        \DataPath/RF/bus_reg_dataout[2209] , 
        \DataPath/RF/bus_reg_dataout[2208] , 
        \DataPath/RF/bus_reg_dataout[2207] , 
        \DataPath/RF/bus_reg_dataout[2206] , 
        \DataPath/RF/bus_reg_dataout[2205] , 
        \DataPath/RF/bus_reg_dataout[2204] , 
        \DataPath/RF/bus_reg_dataout[2203] , 
        \DataPath/RF/bus_reg_dataout[2202] , 
        \DataPath/RF/bus_reg_dataout[2201] , 
        \DataPath/RF/bus_reg_dataout[2200] , 
        \DataPath/RF/bus_reg_dataout[2199] , 
        \DataPath/RF/bus_reg_dataout[2198] , 
        \DataPath/RF/bus_reg_dataout[2197] , 
        \DataPath/RF/bus_reg_dataout[2196] , 
        \DataPath/RF/bus_reg_dataout[2195] , 
        \DataPath/RF/bus_reg_dataout[2194] , 
        \DataPath/RF/bus_reg_dataout[2193] , 
        \DataPath/RF/bus_reg_dataout[2192] , 
        \DataPath/RF/bus_reg_dataout[2191] , 
        \DataPath/RF/bus_reg_dataout[2190] , 
        \DataPath/RF/bus_reg_dataout[2189] , 
        \DataPath/RF/bus_reg_dataout[2188] , 
        \DataPath/RF/bus_reg_dataout[2187] , 
        \DataPath/RF/bus_reg_dataout[2186] , 
        \DataPath/RF/bus_reg_dataout[2185] , 
        \DataPath/RF/bus_reg_dataout[2184] , 
        \DataPath/RF/bus_reg_dataout[2183] , 
        \DataPath/RF/bus_reg_dataout[2182] , 
        \DataPath/RF/bus_reg_dataout[2181] , 
        \DataPath/RF/bus_reg_dataout[2180] , 
        \DataPath/RF/bus_reg_dataout[2179] , 
        \DataPath/RF/bus_reg_dataout[2178] , 
        \DataPath/RF/bus_reg_dataout[2177] , 
        \DataPath/RF/bus_reg_dataout[2176] , 
        \DataPath/RF/bus_reg_dataout[2175] , 
        \DataPath/RF/bus_reg_dataout[2174] , 
        \DataPath/RF/bus_reg_dataout[2173] , 
        \DataPath/RF/bus_reg_dataout[2172] , 
        \DataPath/RF/bus_reg_dataout[2171] , 
        \DataPath/RF/bus_reg_dataout[2170] , 
        \DataPath/RF/bus_reg_dataout[2169] , 
        \DataPath/RF/bus_reg_dataout[2168] , 
        \DataPath/RF/bus_reg_dataout[2167] , 
        \DataPath/RF/bus_reg_dataout[2166] , 
        \DataPath/RF/bus_reg_dataout[2165] , 
        \DataPath/RF/bus_reg_dataout[2164] , 
        \DataPath/RF/bus_reg_dataout[2163] , 
        \DataPath/RF/bus_reg_dataout[2162] , 
        \DataPath/RF/bus_reg_dataout[2161] , 
        \DataPath/RF/bus_reg_dataout[2160] , 
        \DataPath/RF/bus_reg_dataout[2159] , 
        \DataPath/RF/bus_reg_dataout[2158] , 
        \DataPath/RF/bus_reg_dataout[2157] , 
        \DataPath/RF/bus_reg_dataout[2156] , 
        \DataPath/RF/bus_reg_dataout[2155] , 
        \DataPath/RF/bus_reg_dataout[2154] , 
        \DataPath/RF/bus_reg_dataout[2153] , 
        \DataPath/RF/bus_reg_dataout[2152] , 
        \DataPath/RF/bus_reg_dataout[2151] , 
        \DataPath/RF/bus_reg_dataout[2150] , 
        \DataPath/RF/bus_reg_dataout[2149] , 
        \DataPath/RF/bus_reg_dataout[2148] , 
        \DataPath/RF/bus_reg_dataout[2147] , 
        \DataPath/RF/bus_reg_dataout[2146] , 
        \DataPath/RF/bus_reg_dataout[2145] , 
        \DataPath/RF/bus_reg_dataout[2144] , 
        \DataPath/RF/bus_reg_dataout[2143] , 
        \DataPath/RF/bus_reg_dataout[2142] , 
        \DataPath/RF/bus_reg_dataout[2141] , 
        \DataPath/RF/bus_reg_dataout[2140] , 
        \DataPath/RF/bus_reg_dataout[2139] , 
        \DataPath/RF/bus_reg_dataout[2138] , 
        \DataPath/RF/bus_reg_dataout[2137] , 
        \DataPath/RF/bus_reg_dataout[2136] , 
        \DataPath/RF/bus_reg_dataout[2135] , 
        \DataPath/RF/bus_reg_dataout[2134] , 
        \DataPath/RF/bus_reg_dataout[2133] , 
        \DataPath/RF/bus_reg_dataout[2132] , 
        \DataPath/RF/bus_reg_dataout[2131] , 
        \DataPath/RF/bus_reg_dataout[2130] , 
        \DataPath/RF/bus_reg_dataout[2129] , 
        \DataPath/RF/bus_reg_dataout[2128] , 
        \DataPath/RF/bus_reg_dataout[2127] , 
        \DataPath/RF/bus_reg_dataout[2126] , 
        \DataPath/RF/bus_reg_dataout[2125] , 
        \DataPath/RF/bus_reg_dataout[2124] , 
        \DataPath/RF/bus_reg_dataout[2123] , 
        \DataPath/RF/bus_reg_dataout[2122] , 
        \DataPath/RF/bus_reg_dataout[2121] , 
        \DataPath/RF/bus_reg_dataout[2120] , 
        \DataPath/RF/bus_reg_dataout[2119] , 
        \DataPath/RF/bus_reg_dataout[2118] , 
        \DataPath/RF/bus_reg_dataout[2117] , 
        \DataPath/RF/bus_reg_dataout[2116] , 
        \DataPath/RF/bus_reg_dataout[2115] , 
        \DataPath/RF/bus_reg_dataout[2114] , 
        \DataPath/RF/bus_reg_dataout[2113] , 
        \DataPath/RF/bus_reg_dataout[2112] , 
        \DataPath/RF/bus_reg_dataout[2111] , 
        \DataPath/RF/bus_reg_dataout[2110] , 
        \DataPath/RF/bus_reg_dataout[2109] , 
        \DataPath/RF/bus_reg_dataout[2108] , 
        \DataPath/RF/bus_reg_dataout[2107] , 
        \DataPath/RF/bus_reg_dataout[2106] , 
        \DataPath/RF/bus_reg_dataout[2105] , 
        \DataPath/RF/bus_reg_dataout[2104] , 
        \DataPath/RF/bus_reg_dataout[2103] , 
        \DataPath/RF/bus_reg_dataout[2102] , 
        \DataPath/RF/bus_reg_dataout[2101] , 
        \DataPath/RF/bus_reg_dataout[2100] , 
        \DataPath/RF/bus_reg_dataout[2099] , 
        \DataPath/RF/bus_reg_dataout[2098] , 
        \DataPath/RF/bus_reg_dataout[2097] , 
        \DataPath/RF/bus_reg_dataout[2096] , 
        \DataPath/RF/bus_reg_dataout[2095] , 
        \DataPath/RF/bus_reg_dataout[2094] , 
        \DataPath/RF/bus_reg_dataout[2093] , 
        \DataPath/RF/bus_reg_dataout[2092] , 
        \DataPath/RF/bus_reg_dataout[2091] , 
        \DataPath/RF/bus_reg_dataout[2090] , 
        \DataPath/RF/bus_reg_dataout[2089] , 
        \DataPath/RF/bus_reg_dataout[2088] , 
        \DataPath/RF/bus_reg_dataout[2087] , 
        \DataPath/RF/bus_reg_dataout[2086] , 
        \DataPath/RF/bus_reg_dataout[2085] , 
        \DataPath/RF/bus_reg_dataout[2084] , 
        \DataPath/RF/bus_reg_dataout[2083] , 
        \DataPath/RF/bus_reg_dataout[2082] , 
        \DataPath/RF/bus_reg_dataout[2081] , 
        \DataPath/RF/bus_reg_dataout[2080] , 
        \DataPath/RF/bus_reg_dataout[2079] , 
        \DataPath/RF/bus_reg_dataout[2078] , 
        \DataPath/RF/bus_reg_dataout[2077] , 
        \DataPath/RF/bus_reg_dataout[2076] , 
        \DataPath/RF/bus_reg_dataout[2075] , 
        \DataPath/RF/bus_reg_dataout[2074] , 
        \DataPath/RF/bus_reg_dataout[2073] , 
        \DataPath/RF/bus_reg_dataout[2072] , 
        \DataPath/RF/bus_reg_dataout[2071] , 
        \DataPath/RF/bus_reg_dataout[2070] , 
        \DataPath/RF/bus_reg_dataout[2069] , 
        \DataPath/RF/bus_reg_dataout[2068] , 
        \DataPath/RF/bus_reg_dataout[2067] , 
        \DataPath/RF/bus_reg_dataout[2066] , 
        \DataPath/RF/bus_reg_dataout[2065] , 
        \DataPath/RF/bus_reg_dataout[2064] , 
        \DataPath/RF/bus_reg_dataout[2063] , 
        \DataPath/RF/bus_reg_dataout[2062] , 
        \DataPath/RF/bus_reg_dataout[2061] , 
        \DataPath/RF/bus_reg_dataout[2060] , 
        \DataPath/RF/bus_reg_dataout[2059] , 
        \DataPath/RF/bus_reg_dataout[2058] , 
        \DataPath/RF/bus_reg_dataout[2057] , 
        \DataPath/RF/bus_reg_dataout[2056] , 
        \DataPath/RF/bus_reg_dataout[2055] , 
        \DataPath/RF/bus_reg_dataout[2054] , 
        \DataPath/RF/bus_reg_dataout[2053] , 
        \DataPath/RF/bus_reg_dataout[2052] , 
        \DataPath/RF/bus_reg_dataout[2051] , 
        \DataPath/RF/bus_reg_dataout[2050] , 
        \DataPath/RF/bus_reg_dataout[2049] , 
        \DataPath/RF/bus_reg_dataout[2048] , 
        \DataPath/RF/bus_reg_dataout[2047] , 
        \DataPath/RF/bus_reg_dataout[2046] , 
        \DataPath/RF/bus_reg_dataout[2045] , 
        \DataPath/RF/bus_reg_dataout[2044] , 
        \DataPath/RF/bus_reg_dataout[2043] , 
        \DataPath/RF/bus_reg_dataout[2042] , 
        \DataPath/RF/bus_reg_dataout[2041] , 
        \DataPath/RF/bus_reg_dataout[2040] , 
        \DataPath/RF/bus_reg_dataout[2039] , 
        \DataPath/RF/bus_reg_dataout[2038] , 
        \DataPath/RF/bus_reg_dataout[2037] , 
        \DataPath/RF/bus_reg_dataout[2036] , 
        \DataPath/RF/bus_reg_dataout[2035] , 
        \DataPath/RF/bus_reg_dataout[2034] , 
        \DataPath/RF/bus_reg_dataout[2033] , 
        \DataPath/RF/bus_reg_dataout[2032] , 
        \DataPath/RF/bus_reg_dataout[2031] , 
        \DataPath/RF/bus_reg_dataout[2030] , 
        \DataPath/RF/bus_reg_dataout[2029] , 
        \DataPath/RF/bus_reg_dataout[2028] , 
        \DataPath/RF/bus_reg_dataout[2027] , 
        \DataPath/RF/bus_reg_dataout[2026] , 
        \DataPath/RF/bus_reg_dataout[2025] , 
        \DataPath/RF/bus_reg_dataout[2024] , 
        \DataPath/RF/bus_reg_dataout[2023] , 
        \DataPath/RF/bus_reg_dataout[2022] , 
        \DataPath/RF/bus_reg_dataout[2021] , 
        \DataPath/RF/bus_reg_dataout[2020] , 
        \DataPath/RF/bus_reg_dataout[2019] , 
        \DataPath/RF/bus_reg_dataout[2018] , 
        \DataPath/RF/bus_reg_dataout[2017] , 
        \DataPath/RF/bus_reg_dataout[2016] , 
        \DataPath/RF/bus_reg_dataout[2015] , 
        \DataPath/RF/bus_reg_dataout[2014] , 
        \DataPath/RF/bus_reg_dataout[2013] , 
        \DataPath/RF/bus_reg_dataout[2012] , 
        \DataPath/RF/bus_reg_dataout[2011] , 
        \DataPath/RF/bus_reg_dataout[2010] , 
        \DataPath/RF/bus_reg_dataout[2009] , 
        \DataPath/RF/bus_reg_dataout[2008] , 
        \DataPath/RF/bus_reg_dataout[2007] , 
        \DataPath/RF/bus_reg_dataout[2006] , 
        \DataPath/RF/bus_reg_dataout[2005] , 
        \DataPath/RF/bus_reg_dataout[2004] , 
        \DataPath/RF/bus_reg_dataout[2003] , 
        \DataPath/RF/bus_reg_dataout[2002] , 
        \DataPath/RF/bus_reg_dataout[2001] , 
        \DataPath/RF/bus_reg_dataout[2000] , 
        \DataPath/RF/bus_reg_dataout[1999] , 
        \DataPath/RF/bus_reg_dataout[1998] , 
        \DataPath/RF/bus_reg_dataout[1997] , 
        \DataPath/RF/bus_reg_dataout[1996] , 
        \DataPath/RF/bus_reg_dataout[1995] , 
        \DataPath/RF/bus_reg_dataout[1994] , 
        \DataPath/RF/bus_reg_dataout[1993] , 
        \DataPath/RF/bus_reg_dataout[1992] , 
        \DataPath/RF/bus_reg_dataout[1991] , 
        \DataPath/RF/bus_reg_dataout[1990] , 
        \DataPath/RF/bus_reg_dataout[1989] , 
        \DataPath/RF/bus_reg_dataout[1988] , 
        \DataPath/RF/bus_reg_dataout[1987] , 
        \DataPath/RF/bus_reg_dataout[1986] , 
        \DataPath/RF/bus_reg_dataout[1985] , 
        \DataPath/RF/bus_reg_dataout[1984] , 
        \DataPath/RF/bus_reg_dataout[1983] , 
        \DataPath/RF/bus_reg_dataout[1982] , 
        \DataPath/RF/bus_reg_dataout[1981] , 
        \DataPath/RF/bus_reg_dataout[1980] , 
        \DataPath/RF/bus_reg_dataout[1979] , 
        \DataPath/RF/bus_reg_dataout[1978] , 
        \DataPath/RF/bus_reg_dataout[1977] , 
        \DataPath/RF/bus_reg_dataout[1976] , 
        \DataPath/RF/bus_reg_dataout[1975] , 
        \DataPath/RF/bus_reg_dataout[1974] , 
        \DataPath/RF/bus_reg_dataout[1973] , 
        \DataPath/RF/bus_reg_dataout[1972] , 
        \DataPath/RF/bus_reg_dataout[1971] , 
        \DataPath/RF/bus_reg_dataout[1970] , 
        \DataPath/RF/bus_reg_dataout[1969] , 
        \DataPath/RF/bus_reg_dataout[1968] , 
        \DataPath/RF/bus_reg_dataout[1967] , 
        \DataPath/RF/bus_reg_dataout[1966] , 
        \DataPath/RF/bus_reg_dataout[1965] , 
        \DataPath/RF/bus_reg_dataout[1964] , 
        \DataPath/RF/bus_reg_dataout[1963] , 
        \DataPath/RF/bus_reg_dataout[1962] , 
        \DataPath/RF/bus_reg_dataout[1961] , 
        \DataPath/RF/bus_reg_dataout[1960] , 
        \DataPath/RF/bus_reg_dataout[1959] , 
        \DataPath/RF/bus_reg_dataout[1958] , 
        \DataPath/RF/bus_reg_dataout[1957] , 
        \DataPath/RF/bus_reg_dataout[1956] , 
        \DataPath/RF/bus_reg_dataout[1955] , 
        \DataPath/RF/bus_reg_dataout[1954] , 
        \DataPath/RF/bus_reg_dataout[1953] , 
        \DataPath/RF/bus_reg_dataout[1952] , 
        \DataPath/RF/bus_reg_dataout[1951] , 
        \DataPath/RF/bus_reg_dataout[1950] , 
        \DataPath/RF/bus_reg_dataout[1949] , 
        \DataPath/RF/bus_reg_dataout[1948] , 
        \DataPath/RF/bus_reg_dataout[1947] , 
        \DataPath/RF/bus_reg_dataout[1946] , 
        \DataPath/RF/bus_reg_dataout[1945] , 
        \DataPath/RF/bus_reg_dataout[1944] , 
        \DataPath/RF/bus_reg_dataout[1943] , 
        \DataPath/RF/bus_reg_dataout[1942] , 
        \DataPath/RF/bus_reg_dataout[1941] , 
        \DataPath/RF/bus_reg_dataout[1940] , 
        \DataPath/RF/bus_reg_dataout[1939] , 
        \DataPath/RF/bus_reg_dataout[1938] , 
        \DataPath/RF/bus_reg_dataout[1937] , 
        \DataPath/RF/bus_reg_dataout[1936] , 
        \DataPath/RF/bus_reg_dataout[1935] , 
        \DataPath/RF/bus_reg_dataout[1934] , 
        \DataPath/RF/bus_reg_dataout[1933] , 
        \DataPath/RF/bus_reg_dataout[1932] , 
        \DataPath/RF/bus_reg_dataout[1931] , 
        \DataPath/RF/bus_reg_dataout[1930] , 
        \DataPath/RF/bus_reg_dataout[1929] , 
        \DataPath/RF/bus_reg_dataout[1928] , 
        \DataPath/RF/bus_reg_dataout[1927] , 
        \DataPath/RF/bus_reg_dataout[1926] , 
        \DataPath/RF/bus_reg_dataout[1925] , 
        \DataPath/RF/bus_reg_dataout[1924] , 
        \DataPath/RF/bus_reg_dataout[1923] , 
        \DataPath/RF/bus_reg_dataout[1922] , 
        \DataPath/RF/bus_reg_dataout[1921] , 
        \DataPath/RF/bus_reg_dataout[1920] , 
        \DataPath/RF/bus_reg_dataout[1919] , 
        \DataPath/RF/bus_reg_dataout[1918] , 
        \DataPath/RF/bus_reg_dataout[1917] , 
        \DataPath/RF/bus_reg_dataout[1916] , 
        \DataPath/RF/bus_reg_dataout[1915] , 
        \DataPath/RF/bus_reg_dataout[1914] , 
        \DataPath/RF/bus_reg_dataout[1913] , 
        \DataPath/RF/bus_reg_dataout[1912] , 
        \DataPath/RF/bus_reg_dataout[1911] , 
        \DataPath/RF/bus_reg_dataout[1910] , 
        \DataPath/RF/bus_reg_dataout[1909] , 
        \DataPath/RF/bus_reg_dataout[1908] , 
        \DataPath/RF/bus_reg_dataout[1907] , 
        \DataPath/RF/bus_reg_dataout[1906] , 
        \DataPath/RF/bus_reg_dataout[1905] , 
        \DataPath/RF/bus_reg_dataout[1904] , 
        \DataPath/RF/bus_reg_dataout[1903] , 
        \DataPath/RF/bus_reg_dataout[1902] , 
        \DataPath/RF/bus_reg_dataout[1901] , 
        \DataPath/RF/bus_reg_dataout[1900] , 
        \DataPath/RF/bus_reg_dataout[1899] , 
        \DataPath/RF/bus_reg_dataout[1898] , 
        \DataPath/RF/bus_reg_dataout[1897] , 
        \DataPath/RF/bus_reg_dataout[1896] , 
        \DataPath/RF/bus_reg_dataout[1895] , 
        \DataPath/RF/bus_reg_dataout[1894] , 
        \DataPath/RF/bus_reg_dataout[1893] , 
        \DataPath/RF/bus_reg_dataout[1892] , 
        \DataPath/RF/bus_reg_dataout[1891] , 
        \DataPath/RF/bus_reg_dataout[1890] , 
        \DataPath/RF/bus_reg_dataout[1889] , 
        \DataPath/RF/bus_reg_dataout[1888] , 
        \DataPath/RF/bus_reg_dataout[1887] , 
        \DataPath/RF/bus_reg_dataout[1886] , 
        \DataPath/RF/bus_reg_dataout[1885] , 
        \DataPath/RF/bus_reg_dataout[1884] , 
        \DataPath/RF/bus_reg_dataout[1883] , 
        \DataPath/RF/bus_reg_dataout[1882] , 
        \DataPath/RF/bus_reg_dataout[1881] , 
        \DataPath/RF/bus_reg_dataout[1880] , 
        \DataPath/RF/bus_reg_dataout[1879] , 
        \DataPath/RF/bus_reg_dataout[1878] , 
        \DataPath/RF/bus_reg_dataout[1877] , 
        \DataPath/RF/bus_reg_dataout[1876] , 
        \DataPath/RF/bus_reg_dataout[1875] , 
        \DataPath/RF/bus_reg_dataout[1874] , 
        \DataPath/RF/bus_reg_dataout[1873] , 
        \DataPath/RF/bus_reg_dataout[1872] , 
        \DataPath/RF/bus_reg_dataout[1871] , 
        \DataPath/RF/bus_reg_dataout[1870] , 
        \DataPath/RF/bus_reg_dataout[1869] , 
        \DataPath/RF/bus_reg_dataout[1868] , 
        \DataPath/RF/bus_reg_dataout[1867] , 
        \DataPath/RF/bus_reg_dataout[1866] , 
        \DataPath/RF/bus_reg_dataout[1865] , 
        \DataPath/RF/bus_reg_dataout[1864] , 
        \DataPath/RF/bus_reg_dataout[1863] , 
        \DataPath/RF/bus_reg_dataout[1862] , 
        \DataPath/RF/bus_reg_dataout[1861] , 
        \DataPath/RF/bus_reg_dataout[1860] , 
        \DataPath/RF/bus_reg_dataout[1859] , 
        \DataPath/RF/bus_reg_dataout[1858] , 
        \DataPath/RF/bus_reg_dataout[1857] , 
        \DataPath/RF/bus_reg_dataout[1856] , 
        \DataPath/RF/bus_reg_dataout[1855] , 
        \DataPath/RF/bus_reg_dataout[1854] , 
        \DataPath/RF/bus_reg_dataout[1853] , 
        \DataPath/RF/bus_reg_dataout[1852] , 
        \DataPath/RF/bus_reg_dataout[1851] , 
        \DataPath/RF/bus_reg_dataout[1850] , 
        \DataPath/RF/bus_reg_dataout[1849] , 
        \DataPath/RF/bus_reg_dataout[1848] , 
        \DataPath/RF/bus_reg_dataout[1847] , 
        \DataPath/RF/bus_reg_dataout[1846] , 
        \DataPath/RF/bus_reg_dataout[1845] , 
        \DataPath/RF/bus_reg_dataout[1844] , 
        \DataPath/RF/bus_reg_dataout[1843] , 
        \DataPath/RF/bus_reg_dataout[1842] , 
        \DataPath/RF/bus_reg_dataout[1841] , 
        \DataPath/RF/bus_reg_dataout[1840] , 
        \DataPath/RF/bus_reg_dataout[1839] , 
        \DataPath/RF/bus_reg_dataout[1838] , 
        \DataPath/RF/bus_reg_dataout[1837] , 
        \DataPath/RF/bus_reg_dataout[1836] , 
        \DataPath/RF/bus_reg_dataout[1835] , 
        \DataPath/RF/bus_reg_dataout[1834] , 
        \DataPath/RF/bus_reg_dataout[1833] , 
        \DataPath/RF/bus_reg_dataout[1832] , 
        \DataPath/RF/bus_reg_dataout[1831] , 
        \DataPath/RF/bus_reg_dataout[1830] , 
        \DataPath/RF/bus_reg_dataout[1829] , 
        \DataPath/RF/bus_reg_dataout[1828] , 
        \DataPath/RF/bus_reg_dataout[1827] , 
        \DataPath/RF/bus_reg_dataout[1826] , 
        \DataPath/RF/bus_reg_dataout[1825] , 
        \DataPath/RF/bus_reg_dataout[1824] , 
        \DataPath/RF/bus_reg_dataout[1823] , 
        \DataPath/RF/bus_reg_dataout[1822] , 
        \DataPath/RF/bus_reg_dataout[1821] , 
        \DataPath/RF/bus_reg_dataout[1820] , 
        \DataPath/RF/bus_reg_dataout[1819] , 
        \DataPath/RF/bus_reg_dataout[1818] , 
        \DataPath/RF/bus_reg_dataout[1817] , 
        \DataPath/RF/bus_reg_dataout[1816] , 
        \DataPath/RF/bus_reg_dataout[1815] , 
        \DataPath/RF/bus_reg_dataout[1814] , 
        \DataPath/RF/bus_reg_dataout[1813] , 
        \DataPath/RF/bus_reg_dataout[1812] , 
        \DataPath/RF/bus_reg_dataout[1811] , 
        \DataPath/RF/bus_reg_dataout[1810] , 
        \DataPath/RF/bus_reg_dataout[1809] , 
        \DataPath/RF/bus_reg_dataout[1808] , 
        \DataPath/RF/bus_reg_dataout[1807] , 
        \DataPath/RF/bus_reg_dataout[1806] , 
        \DataPath/RF/bus_reg_dataout[1805] , 
        \DataPath/RF/bus_reg_dataout[1804] , 
        \DataPath/RF/bus_reg_dataout[1803] , 
        \DataPath/RF/bus_reg_dataout[1802] , 
        \DataPath/RF/bus_reg_dataout[1801] , 
        \DataPath/RF/bus_reg_dataout[1800] , 
        \DataPath/RF/bus_reg_dataout[1799] , 
        \DataPath/RF/bus_reg_dataout[1798] , 
        \DataPath/RF/bus_reg_dataout[1797] , 
        \DataPath/RF/bus_reg_dataout[1796] , 
        \DataPath/RF/bus_reg_dataout[1795] , 
        \DataPath/RF/bus_reg_dataout[1794] , 
        \DataPath/RF/bus_reg_dataout[1793] , 
        \DataPath/RF/bus_reg_dataout[1792] , 
        \DataPath/RF/bus_reg_dataout[1791] , 
        \DataPath/RF/bus_reg_dataout[1790] , 
        \DataPath/RF/bus_reg_dataout[1789] , 
        \DataPath/RF/bus_reg_dataout[1788] , 
        \DataPath/RF/bus_reg_dataout[1787] , 
        \DataPath/RF/bus_reg_dataout[1786] , 
        \DataPath/RF/bus_reg_dataout[1785] , 
        \DataPath/RF/bus_reg_dataout[1784] , 
        \DataPath/RF/bus_reg_dataout[1783] , 
        \DataPath/RF/bus_reg_dataout[1782] , 
        \DataPath/RF/bus_reg_dataout[1781] , 
        \DataPath/RF/bus_reg_dataout[1780] , 
        \DataPath/RF/bus_reg_dataout[1779] , 
        \DataPath/RF/bus_reg_dataout[1778] , 
        \DataPath/RF/bus_reg_dataout[1777] , 
        \DataPath/RF/bus_reg_dataout[1776] , 
        \DataPath/RF/bus_reg_dataout[1775] , 
        \DataPath/RF/bus_reg_dataout[1774] , 
        \DataPath/RF/bus_reg_dataout[1773] , 
        \DataPath/RF/bus_reg_dataout[1772] , 
        \DataPath/RF/bus_reg_dataout[1771] , 
        \DataPath/RF/bus_reg_dataout[1770] , 
        \DataPath/RF/bus_reg_dataout[1769] , 
        \DataPath/RF/bus_reg_dataout[1768] , 
        \DataPath/RF/bus_reg_dataout[1767] , 
        \DataPath/RF/bus_reg_dataout[1766] , 
        \DataPath/RF/bus_reg_dataout[1765] , 
        \DataPath/RF/bus_reg_dataout[1764] , 
        \DataPath/RF/bus_reg_dataout[1763] , 
        \DataPath/RF/bus_reg_dataout[1762] , 
        \DataPath/RF/bus_reg_dataout[1761] , 
        \DataPath/RF/bus_reg_dataout[1760] , 
        \DataPath/RF/bus_reg_dataout[1759] , 
        \DataPath/RF/bus_reg_dataout[1758] , 
        \DataPath/RF/bus_reg_dataout[1757] , 
        \DataPath/RF/bus_reg_dataout[1756] , 
        \DataPath/RF/bus_reg_dataout[1755] , 
        \DataPath/RF/bus_reg_dataout[1754] , 
        \DataPath/RF/bus_reg_dataout[1753] , 
        \DataPath/RF/bus_reg_dataout[1752] , 
        \DataPath/RF/bus_reg_dataout[1751] , 
        \DataPath/RF/bus_reg_dataout[1750] , 
        \DataPath/RF/bus_reg_dataout[1749] , 
        \DataPath/RF/bus_reg_dataout[1748] , 
        \DataPath/RF/bus_reg_dataout[1747] , 
        \DataPath/RF/bus_reg_dataout[1746] , 
        \DataPath/RF/bus_reg_dataout[1745] , 
        \DataPath/RF/bus_reg_dataout[1744] , 
        \DataPath/RF/bus_reg_dataout[1743] , 
        \DataPath/RF/bus_reg_dataout[1742] , 
        \DataPath/RF/bus_reg_dataout[1741] , 
        \DataPath/RF/bus_reg_dataout[1740] , 
        \DataPath/RF/bus_reg_dataout[1739] , 
        \DataPath/RF/bus_reg_dataout[1738] , 
        \DataPath/RF/bus_reg_dataout[1737] , 
        \DataPath/RF/bus_reg_dataout[1736] , 
        \DataPath/RF/bus_reg_dataout[1735] , 
        \DataPath/RF/bus_reg_dataout[1734] , 
        \DataPath/RF/bus_reg_dataout[1733] , 
        \DataPath/RF/bus_reg_dataout[1732] , 
        \DataPath/RF/bus_reg_dataout[1731] , 
        \DataPath/RF/bus_reg_dataout[1730] , 
        \DataPath/RF/bus_reg_dataout[1729] , 
        \DataPath/RF/bus_reg_dataout[1728] , 
        \DataPath/RF/bus_reg_dataout[1727] , 
        \DataPath/RF/bus_reg_dataout[1726] , 
        \DataPath/RF/bus_reg_dataout[1725] , 
        \DataPath/RF/bus_reg_dataout[1724] , 
        \DataPath/RF/bus_reg_dataout[1723] , 
        \DataPath/RF/bus_reg_dataout[1722] , 
        \DataPath/RF/bus_reg_dataout[1721] , 
        \DataPath/RF/bus_reg_dataout[1720] , 
        \DataPath/RF/bus_reg_dataout[1719] , 
        \DataPath/RF/bus_reg_dataout[1718] , 
        \DataPath/RF/bus_reg_dataout[1717] , 
        \DataPath/RF/bus_reg_dataout[1716] , 
        \DataPath/RF/bus_reg_dataout[1715] , 
        \DataPath/RF/bus_reg_dataout[1714] , 
        \DataPath/RF/bus_reg_dataout[1713] , 
        \DataPath/RF/bus_reg_dataout[1712] , 
        \DataPath/RF/bus_reg_dataout[1711] , 
        \DataPath/RF/bus_reg_dataout[1710] , 
        \DataPath/RF/bus_reg_dataout[1709] , 
        \DataPath/RF/bus_reg_dataout[1708] , 
        \DataPath/RF/bus_reg_dataout[1707] , 
        \DataPath/RF/bus_reg_dataout[1706] , 
        \DataPath/RF/bus_reg_dataout[1705] , 
        \DataPath/RF/bus_reg_dataout[1704] , 
        \DataPath/RF/bus_reg_dataout[1703] , 
        \DataPath/RF/bus_reg_dataout[1702] , 
        \DataPath/RF/bus_reg_dataout[1701] , 
        \DataPath/RF/bus_reg_dataout[1700] , 
        \DataPath/RF/bus_reg_dataout[1699] , 
        \DataPath/RF/bus_reg_dataout[1698] , 
        \DataPath/RF/bus_reg_dataout[1697] , 
        \DataPath/RF/bus_reg_dataout[1696] , 
        \DataPath/RF/bus_reg_dataout[1695] , 
        \DataPath/RF/bus_reg_dataout[1694] , 
        \DataPath/RF/bus_reg_dataout[1693] , 
        \DataPath/RF/bus_reg_dataout[1692] , 
        \DataPath/RF/bus_reg_dataout[1691] , 
        \DataPath/RF/bus_reg_dataout[1690] , 
        \DataPath/RF/bus_reg_dataout[1689] , 
        \DataPath/RF/bus_reg_dataout[1688] , 
        \DataPath/RF/bus_reg_dataout[1687] , 
        \DataPath/RF/bus_reg_dataout[1686] , 
        \DataPath/RF/bus_reg_dataout[1685] , 
        \DataPath/RF/bus_reg_dataout[1684] , 
        \DataPath/RF/bus_reg_dataout[1683] , 
        \DataPath/RF/bus_reg_dataout[1682] , 
        \DataPath/RF/bus_reg_dataout[1681] , 
        \DataPath/RF/bus_reg_dataout[1680] , 
        \DataPath/RF/bus_reg_dataout[1679] , 
        \DataPath/RF/bus_reg_dataout[1678] , 
        \DataPath/RF/bus_reg_dataout[1677] , 
        \DataPath/RF/bus_reg_dataout[1676] , 
        \DataPath/RF/bus_reg_dataout[1675] , 
        \DataPath/RF/bus_reg_dataout[1674] , 
        \DataPath/RF/bus_reg_dataout[1673] , 
        \DataPath/RF/bus_reg_dataout[1672] , 
        \DataPath/RF/bus_reg_dataout[1671] , 
        \DataPath/RF/bus_reg_dataout[1670] , 
        \DataPath/RF/bus_reg_dataout[1669] , 
        \DataPath/RF/bus_reg_dataout[1668] , 
        \DataPath/RF/bus_reg_dataout[1667] , 
        \DataPath/RF/bus_reg_dataout[1666] , 
        \DataPath/RF/bus_reg_dataout[1665] , 
        \DataPath/RF/bus_reg_dataout[1664] , 
        \DataPath/RF/bus_reg_dataout[1663] , 
        \DataPath/RF/bus_reg_dataout[1662] , 
        \DataPath/RF/bus_reg_dataout[1661] , 
        \DataPath/RF/bus_reg_dataout[1660] , 
        \DataPath/RF/bus_reg_dataout[1659] , 
        \DataPath/RF/bus_reg_dataout[1658] , 
        \DataPath/RF/bus_reg_dataout[1657] , 
        \DataPath/RF/bus_reg_dataout[1656] , 
        \DataPath/RF/bus_reg_dataout[1655] , 
        \DataPath/RF/bus_reg_dataout[1654] , 
        \DataPath/RF/bus_reg_dataout[1653] , 
        \DataPath/RF/bus_reg_dataout[1652] , 
        \DataPath/RF/bus_reg_dataout[1651] , 
        \DataPath/RF/bus_reg_dataout[1650] , 
        \DataPath/RF/bus_reg_dataout[1649] , 
        \DataPath/RF/bus_reg_dataout[1648] , 
        \DataPath/RF/bus_reg_dataout[1647] , 
        \DataPath/RF/bus_reg_dataout[1646] , 
        \DataPath/RF/bus_reg_dataout[1645] , 
        \DataPath/RF/bus_reg_dataout[1644] , 
        \DataPath/RF/bus_reg_dataout[1643] , 
        \DataPath/RF/bus_reg_dataout[1642] , 
        \DataPath/RF/bus_reg_dataout[1641] , 
        \DataPath/RF/bus_reg_dataout[1640] , 
        \DataPath/RF/bus_reg_dataout[1639] , 
        \DataPath/RF/bus_reg_dataout[1638] , 
        \DataPath/RF/bus_reg_dataout[1637] , 
        \DataPath/RF/bus_reg_dataout[1636] , 
        \DataPath/RF/bus_reg_dataout[1635] , 
        \DataPath/RF/bus_reg_dataout[1634] , 
        \DataPath/RF/bus_reg_dataout[1633] , 
        \DataPath/RF/bus_reg_dataout[1632] , 
        \DataPath/RF/bus_reg_dataout[1631] , 
        \DataPath/RF/bus_reg_dataout[1630] , 
        \DataPath/RF/bus_reg_dataout[1629] , 
        \DataPath/RF/bus_reg_dataout[1628] , 
        \DataPath/RF/bus_reg_dataout[1627] , 
        \DataPath/RF/bus_reg_dataout[1626] , 
        \DataPath/RF/bus_reg_dataout[1625] , 
        \DataPath/RF/bus_reg_dataout[1624] , 
        \DataPath/RF/bus_reg_dataout[1623] , 
        \DataPath/RF/bus_reg_dataout[1622] , 
        \DataPath/RF/bus_reg_dataout[1621] , 
        \DataPath/RF/bus_reg_dataout[1620] , 
        \DataPath/RF/bus_reg_dataout[1619] , 
        \DataPath/RF/bus_reg_dataout[1618] , 
        \DataPath/RF/bus_reg_dataout[1617] , 
        \DataPath/RF/bus_reg_dataout[1616] , 
        \DataPath/RF/bus_reg_dataout[1615] , 
        \DataPath/RF/bus_reg_dataout[1614] , 
        \DataPath/RF/bus_reg_dataout[1613] , 
        \DataPath/RF/bus_reg_dataout[1612] , 
        \DataPath/RF/bus_reg_dataout[1611] , 
        \DataPath/RF/bus_reg_dataout[1610] , 
        \DataPath/RF/bus_reg_dataout[1609] , 
        \DataPath/RF/bus_reg_dataout[1608] , 
        \DataPath/RF/bus_reg_dataout[1607] , 
        \DataPath/RF/bus_reg_dataout[1606] , 
        \DataPath/RF/bus_reg_dataout[1605] , 
        \DataPath/RF/bus_reg_dataout[1604] , 
        \DataPath/RF/bus_reg_dataout[1603] , 
        \DataPath/RF/bus_reg_dataout[1602] , 
        \DataPath/RF/bus_reg_dataout[1601] , 
        \DataPath/RF/bus_reg_dataout[1600] , 
        \DataPath/RF/bus_reg_dataout[1599] , 
        \DataPath/RF/bus_reg_dataout[1598] , 
        \DataPath/RF/bus_reg_dataout[1597] , 
        \DataPath/RF/bus_reg_dataout[1596] , 
        \DataPath/RF/bus_reg_dataout[1595] , 
        \DataPath/RF/bus_reg_dataout[1594] , 
        \DataPath/RF/bus_reg_dataout[1593] , 
        \DataPath/RF/bus_reg_dataout[1592] , 
        \DataPath/RF/bus_reg_dataout[1591] , 
        \DataPath/RF/bus_reg_dataout[1590] , 
        \DataPath/RF/bus_reg_dataout[1589] , 
        \DataPath/RF/bus_reg_dataout[1588] , 
        \DataPath/RF/bus_reg_dataout[1587] , 
        \DataPath/RF/bus_reg_dataout[1586] , 
        \DataPath/RF/bus_reg_dataout[1585] , 
        \DataPath/RF/bus_reg_dataout[1584] , 
        \DataPath/RF/bus_reg_dataout[1583] , 
        \DataPath/RF/bus_reg_dataout[1582] , 
        \DataPath/RF/bus_reg_dataout[1581] , 
        \DataPath/RF/bus_reg_dataout[1580] , 
        \DataPath/RF/bus_reg_dataout[1579] , 
        \DataPath/RF/bus_reg_dataout[1578] , 
        \DataPath/RF/bus_reg_dataout[1577] , 
        \DataPath/RF/bus_reg_dataout[1576] , 
        \DataPath/RF/bus_reg_dataout[1575] , 
        \DataPath/RF/bus_reg_dataout[1574] , 
        \DataPath/RF/bus_reg_dataout[1573] , 
        \DataPath/RF/bus_reg_dataout[1572] , 
        \DataPath/RF/bus_reg_dataout[1571] , 
        \DataPath/RF/bus_reg_dataout[1570] , 
        \DataPath/RF/bus_reg_dataout[1569] , 
        \DataPath/RF/bus_reg_dataout[1568] , 
        \DataPath/RF/bus_reg_dataout[1567] , 
        \DataPath/RF/bus_reg_dataout[1566] , 
        \DataPath/RF/bus_reg_dataout[1565] , 
        \DataPath/RF/bus_reg_dataout[1564] , 
        \DataPath/RF/bus_reg_dataout[1563] , 
        \DataPath/RF/bus_reg_dataout[1562] , 
        \DataPath/RF/bus_reg_dataout[1561] , 
        \DataPath/RF/bus_reg_dataout[1560] , 
        \DataPath/RF/bus_reg_dataout[1559] , 
        \DataPath/RF/bus_reg_dataout[1558] , 
        \DataPath/RF/bus_reg_dataout[1557] , 
        \DataPath/RF/bus_reg_dataout[1556] , 
        \DataPath/RF/bus_reg_dataout[1555] , 
        \DataPath/RF/bus_reg_dataout[1554] , 
        \DataPath/RF/bus_reg_dataout[1553] , 
        \DataPath/RF/bus_reg_dataout[1552] , 
        \DataPath/RF/bus_reg_dataout[1551] , 
        \DataPath/RF/bus_reg_dataout[1550] , 
        \DataPath/RF/bus_reg_dataout[1549] , 
        \DataPath/RF/bus_reg_dataout[1548] , 
        \DataPath/RF/bus_reg_dataout[1547] , 
        \DataPath/RF/bus_reg_dataout[1546] , 
        \DataPath/RF/bus_reg_dataout[1545] , 
        \DataPath/RF/bus_reg_dataout[1544] , 
        \DataPath/RF/bus_reg_dataout[1543] , 
        \DataPath/RF/bus_reg_dataout[1542] , 
        \DataPath/RF/bus_reg_dataout[1541] , 
        \DataPath/RF/bus_reg_dataout[1540] , 
        \DataPath/RF/bus_reg_dataout[1539] , 
        \DataPath/RF/bus_reg_dataout[1538] , 
        \DataPath/RF/bus_reg_dataout[1537] , 
        \DataPath/RF/bus_reg_dataout[1536] , 
        \DataPath/RF/bus_reg_dataout[1535] , 
        \DataPath/RF/bus_reg_dataout[1534] , 
        \DataPath/RF/bus_reg_dataout[1533] , 
        \DataPath/RF/bus_reg_dataout[1532] , 
        \DataPath/RF/bus_reg_dataout[1531] , 
        \DataPath/RF/bus_reg_dataout[1530] , 
        \DataPath/RF/bus_reg_dataout[1529] , 
        \DataPath/RF/bus_reg_dataout[1528] , 
        \DataPath/RF/bus_reg_dataout[1527] , 
        \DataPath/RF/bus_reg_dataout[1526] , 
        \DataPath/RF/bus_reg_dataout[1525] , 
        \DataPath/RF/bus_reg_dataout[1524] , 
        \DataPath/RF/bus_reg_dataout[1523] , 
        \DataPath/RF/bus_reg_dataout[1522] , 
        \DataPath/RF/bus_reg_dataout[1521] , 
        \DataPath/RF/bus_reg_dataout[1520] , 
        \DataPath/RF/bus_reg_dataout[1519] , 
        \DataPath/RF/bus_reg_dataout[1518] , 
        \DataPath/RF/bus_reg_dataout[1517] , 
        \DataPath/RF/bus_reg_dataout[1516] , 
        \DataPath/RF/bus_reg_dataout[1515] , 
        \DataPath/RF/bus_reg_dataout[1514] , 
        \DataPath/RF/bus_reg_dataout[1513] , 
        \DataPath/RF/bus_reg_dataout[1512] , 
        \DataPath/RF/bus_reg_dataout[1511] , 
        \DataPath/RF/bus_reg_dataout[1510] , 
        \DataPath/RF/bus_reg_dataout[1509] , 
        \DataPath/RF/bus_reg_dataout[1508] , 
        \DataPath/RF/bus_reg_dataout[1507] , 
        \DataPath/RF/bus_reg_dataout[1506] , 
        \DataPath/RF/bus_reg_dataout[1505] , 
        \DataPath/RF/bus_reg_dataout[1504] , 
        \DataPath/RF/bus_reg_dataout[1503] , 
        \DataPath/RF/bus_reg_dataout[1502] , 
        \DataPath/RF/bus_reg_dataout[1501] , 
        \DataPath/RF/bus_reg_dataout[1500] , 
        \DataPath/RF/bus_reg_dataout[1499] , 
        \DataPath/RF/bus_reg_dataout[1498] , 
        \DataPath/RF/bus_reg_dataout[1497] , 
        \DataPath/RF/bus_reg_dataout[1496] , 
        \DataPath/RF/bus_reg_dataout[1495] , 
        \DataPath/RF/bus_reg_dataout[1494] , 
        \DataPath/RF/bus_reg_dataout[1493] , 
        \DataPath/RF/bus_reg_dataout[1492] , 
        \DataPath/RF/bus_reg_dataout[1491] , 
        \DataPath/RF/bus_reg_dataout[1490] , 
        \DataPath/RF/bus_reg_dataout[1489] , 
        \DataPath/RF/bus_reg_dataout[1488] , 
        \DataPath/RF/bus_reg_dataout[1487] , 
        \DataPath/RF/bus_reg_dataout[1486] , 
        \DataPath/RF/bus_reg_dataout[1485] , 
        \DataPath/RF/bus_reg_dataout[1484] , 
        \DataPath/RF/bus_reg_dataout[1483] , 
        \DataPath/RF/bus_reg_dataout[1482] , 
        \DataPath/RF/bus_reg_dataout[1481] , 
        \DataPath/RF/bus_reg_dataout[1480] , 
        \DataPath/RF/bus_reg_dataout[1479] , 
        \DataPath/RF/bus_reg_dataout[1478] , 
        \DataPath/RF/bus_reg_dataout[1477] , 
        \DataPath/RF/bus_reg_dataout[1476] , 
        \DataPath/RF/bus_reg_dataout[1475] , 
        \DataPath/RF/bus_reg_dataout[1474] , 
        \DataPath/RF/bus_reg_dataout[1473] , 
        \DataPath/RF/bus_reg_dataout[1472] , 
        \DataPath/RF/bus_reg_dataout[1471] , 
        \DataPath/RF/bus_reg_dataout[1470] , 
        \DataPath/RF/bus_reg_dataout[1469] , 
        \DataPath/RF/bus_reg_dataout[1468] , 
        \DataPath/RF/bus_reg_dataout[1467] , 
        \DataPath/RF/bus_reg_dataout[1466] , 
        \DataPath/RF/bus_reg_dataout[1465] , 
        \DataPath/RF/bus_reg_dataout[1464] , 
        \DataPath/RF/bus_reg_dataout[1463] , 
        \DataPath/RF/bus_reg_dataout[1462] , 
        \DataPath/RF/bus_reg_dataout[1461] , 
        \DataPath/RF/bus_reg_dataout[1460] , 
        \DataPath/RF/bus_reg_dataout[1459] , 
        \DataPath/RF/bus_reg_dataout[1458] , 
        \DataPath/RF/bus_reg_dataout[1457] , 
        \DataPath/RF/bus_reg_dataout[1456] , 
        \DataPath/RF/bus_reg_dataout[1455] , 
        \DataPath/RF/bus_reg_dataout[1454] , 
        \DataPath/RF/bus_reg_dataout[1453] , 
        \DataPath/RF/bus_reg_dataout[1452] , 
        \DataPath/RF/bus_reg_dataout[1451] , 
        \DataPath/RF/bus_reg_dataout[1450] , 
        \DataPath/RF/bus_reg_dataout[1449] , 
        \DataPath/RF/bus_reg_dataout[1448] , 
        \DataPath/RF/bus_reg_dataout[1447] , 
        \DataPath/RF/bus_reg_dataout[1446] , 
        \DataPath/RF/bus_reg_dataout[1445] , 
        \DataPath/RF/bus_reg_dataout[1444] , 
        \DataPath/RF/bus_reg_dataout[1443] , 
        \DataPath/RF/bus_reg_dataout[1442] , 
        \DataPath/RF/bus_reg_dataout[1441] , 
        \DataPath/RF/bus_reg_dataout[1440] , 
        \DataPath/RF/bus_reg_dataout[1439] , 
        \DataPath/RF/bus_reg_dataout[1438] , 
        \DataPath/RF/bus_reg_dataout[1437] , 
        \DataPath/RF/bus_reg_dataout[1436] , 
        \DataPath/RF/bus_reg_dataout[1435] , 
        \DataPath/RF/bus_reg_dataout[1434] , 
        \DataPath/RF/bus_reg_dataout[1433] , 
        \DataPath/RF/bus_reg_dataout[1432] , 
        \DataPath/RF/bus_reg_dataout[1431] , 
        \DataPath/RF/bus_reg_dataout[1430] , 
        \DataPath/RF/bus_reg_dataout[1429] , 
        \DataPath/RF/bus_reg_dataout[1428] , 
        \DataPath/RF/bus_reg_dataout[1427] , 
        \DataPath/RF/bus_reg_dataout[1426] , 
        \DataPath/RF/bus_reg_dataout[1425] , 
        \DataPath/RF/bus_reg_dataout[1424] , 
        \DataPath/RF/bus_reg_dataout[1423] , 
        \DataPath/RF/bus_reg_dataout[1422] , 
        \DataPath/RF/bus_reg_dataout[1421] , 
        \DataPath/RF/bus_reg_dataout[1420] , 
        \DataPath/RF/bus_reg_dataout[1419] , 
        \DataPath/RF/bus_reg_dataout[1418] , 
        \DataPath/RF/bus_reg_dataout[1417] , 
        \DataPath/RF/bus_reg_dataout[1416] , 
        \DataPath/RF/bus_reg_dataout[1415] , 
        \DataPath/RF/bus_reg_dataout[1414] , 
        \DataPath/RF/bus_reg_dataout[1413] , 
        \DataPath/RF/bus_reg_dataout[1412] , 
        \DataPath/RF/bus_reg_dataout[1411] , 
        \DataPath/RF/bus_reg_dataout[1410] , 
        \DataPath/RF/bus_reg_dataout[1409] , 
        \DataPath/RF/bus_reg_dataout[1408] , 
        \DataPath/RF/bus_reg_dataout[1407] , 
        \DataPath/RF/bus_reg_dataout[1406] , 
        \DataPath/RF/bus_reg_dataout[1405] , 
        \DataPath/RF/bus_reg_dataout[1404] , 
        \DataPath/RF/bus_reg_dataout[1403] , 
        \DataPath/RF/bus_reg_dataout[1402] , 
        \DataPath/RF/bus_reg_dataout[1401] , 
        \DataPath/RF/bus_reg_dataout[1400] , 
        \DataPath/RF/bus_reg_dataout[1399] , 
        \DataPath/RF/bus_reg_dataout[1398] , 
        \DataPath/RF/bus_reg_dataout[1397] , 
        \DataPath/RF/bus_reg_dataout[1396] , 
        \DataPath/RF/bus_reg_dataout[1395] , 
        \DataPath/RF/bus_reg_dataout[1394] , 
        \DataPath/RF/bus_reg_dataout[1393] , 
        \DataPath/RF/bus_reg_dataout[1392] , 
        \DataPath/RF/bus_reg_dataout[1391] , 
        \DataPath/RF/bus_reg_dataout[1390] , 
        \DataPath/RF/bus_reg_dataout[1389] , 
        \DataPath/RF/bus_reg_dataout[1388] , 
        \DataPath/RF/bus_reg_dataout[1387] , 
        \DataPath/RF/bus_reg_dataout[1386] , 
        \DataPath/RF/bus_reg_dataout[1385] , 
        \DataPath/RF/bus_reg_dataout[1384] , 
        \DataPath/RF/bus_reg_dataout[1383] , 
        \DataPath/RF/bus_reg_dataout[1382] , 
        \DataPath/RF/bus_reg_dataout[1381] , 
        \DataPath/RF/bus_reg_dataout[1380] , 
        \DataPath/RF/bus_reg_dataout[1379] , 
        \DataPath/RF/bus_reg_dataout[1378] , 
        \DataPath/RF/bus_reg_dataout[1377] , 
        \DataPath/RF/bus_reg_dataout[1376] , 
        \DataPath/RF/bus_reg_dataout[1375] , 
        \DataPath/RF/bus_reg_dataout[1374] , 
        \DataPath/RF/bus_reg_dataout[1373] , 
        \DataPath/RF/bus_reg_dataout[1372] , 
        \DataPath/RF/bus_reg_dataout[1371] , 
        \DataPath/RF/bus_reg_dataout[1370] , 
        \DataPath/RF/bus_reg_dataout[1369] , 
        \DataPath/RF/bus_reg_dataout[1368] , 
        \DataPath/RF/bus_reg_dataout[1367] , 
        \DataPath/RF/bus_reg_dataout[1366] , 
        \DataPath/RF/bus_reg_dataout[1365] , 
        \DataPath/RF/bus_reg_dataout[1364] , 
        \DataPath/RF/bus_reg_dataout[1363] , 
        \DataPath/RF/bus_reg_dataout[1362] , 
        \DataPath/RF/bus_reg_dataout[1361] , 
        \DataPath/RF/bus_reg_dataout[1360] , 
        \DataPath/RF/bus_reg_dataout[1359] , 
        \DataPath/RF/bus_reg_dataout[1358] , 
        \DataPath/RF/bus_reg_dataout[1357] , 
        \DataPath/RF/bus_reg_dataout[1356] , 
        \DataPath/RF/bus_reg_dataout[1355] , 
        \DataPath/RF/bus_reg_dataout[1354] , 
        \DataPath/RF/bus_reg_dataout[1353] , 
        \DataPath/RF/bus_reg_dataout[1352] , 
        \DataPath/RF/bus_reg_dataout[1351] , 
        \DataPath/RF/bus_reg_dataout[1350] , 
        \DataPath/RF/bus_reg_dataout[1349] , 
        \DataPath/RF/bus_reg_dataout[1348] , 
        \DataPath/RF/bus_reg_dataout[1347] , 
        \DataPath/RF/bus_reg_dataout[1346] , 
        \DataPath/RF/bus_reg_dataout[1345] , 
        \DataPath/RF/bus_reg_dataout[1344] , 
        \DataPath/RF/bus_reg_dataout[1343] , 
        \DataPath/RF/bus_reg_dataout[1342] , 
        \DataPath/RF/bus_reg_dataout[1341] , 
        \DataPath/RF/bus_reg_dataout[1340] , 
        \DataPath/RF/bus_reg_dataout[1339] , 
        \DataPath/RF/bus_reg_dataout[1338] , 
        \DataPath/RF/bus_reg_dataout[1337] , 
        \DataPath/RF/bus_reg_dataout[1336] , 
        \DataPath/RF/bus_reg_dataout[1335] , 
        \DataPath/RF/bus_reg_dataout[1334] , 
        \DataPath/RF/bus_reg_dataout[1333] , 
        \DataPath/RF/bus_reg_dataout[1332] , 
        \DataPath/RF/bus_reg_dataout[1331] , 
        \DataPath/RF/bus_reg_dataout[1330] , 
        \DataPath/RF/bus_reg_dataout[1329] , 
        \DataPath/RF/bus_reg_dataout[1328] , 
        \DataPath/RF/bus_reg_dataout[1327] , 
        \DataPath/RF/bus_reg_dataout[1326] , 
        \DataPath/RF/bus_reg_dataout[1325] , 
        \DataPath/RF/bus_reg_dataout[1324] , 
        \DataPath/RF/bus_reg_dataout[1323] , 
        \DataPath/RF/bus_reg_dataout[1322] , 
        \DataPath/RF/bus_reg_dataout[1321] , 
        \DataPath/RF/bus_reg_dataout[1320] , 
        \DataPath/RF/bus_reg_dataout[1319] , 
        \DataPath/RF/bus_reg_dataout[1318] , 
        \DataPath/RF/bus_reg_dataout[1317] , 
        \DataPath/RF/bus_reg_dataout[1316] , 
        \DataPath/RF/bus_reg_dataout[1315] , 
        \DataPath/RF/bus_reg_dataout[1314] , 
        \DataPath/RF/bus_reg_dataout[1313] , 
        \DataPath/RF/bus_reg_dataout[1312] , 
        \DataPath/RF/bus_reg_dataout[1311] , 
        \DataPath/RF/bus_reg_dataout[1310] , 
        \DataPath/RF/bus_reg_dataout[1309] , 
        \DataPath/RF/bus_reg_dataout[1308] , 
        \DataPath/RF/bus_reg_dataout[1307] , 
        \DataPath/RF/bus_reg_dataout[1306] , 
        \DataPath/RF/bus_reg_dataout[1305] , 
        \DataPath/RF/bus_reg_dataout[1304] , 
        \DataPath/RF/bus_reg_dataout[1303] , 
        \DataPath/RF/bus_reg_dataout[1302] , 
        \DataPath/RF/bus_reg_dataout[1301] , 
        \DataPath/RF/bus_reg_dataout[1300] , 
        \DataPath/RF/bus_reg_dataout[1299] , 
        \DataPath/RF/bus_reg_dataout[1298] , 
        \DataPath/RF/bus_reg_dataout[1297] , 
        \DataPath/RF/bus_reg_dataout[1296] , 
        \DataPath/RF/bus_reg_dataout[1295] , 
        \DataPath/RF/bus_reg_dataout[1294] , 
        \DataPath/RF/bus_reg_dataout[1293] , 
        \DataPath/RF/bus_reg_dataout[1292] , 
        \DataPath/RF/bus_reg_dataout[1291] , 
        \DataPath/RF/bus_reg_dataout[1290] , 
        \DataPath/RF/bus_reg_dataout[1289] , 
        \DataPath/RF/bus_reg_dataout[1288] , 
        \DataPath/RF/bus_reg_dataout[1287] , 
        \DataPath/RF/bus_reg_dataout[1286] , 
        \DataPath/RF/bus_reg_dataout[1285] , 
        \DataPath/RF/bus_reg_dataout[1284] , 
        \DataPath/RF/bus_reg_dataout[1283] , 
        \DataPath/RF/bus_reg_dataout[1282] , 
        \DataPath/RF/bus_reg_dataout[1281] , 
        \DataPath/RF/bus_reg_dataout[1280] , 
        \DataPath/RF/bus_reg_dataout[1279] , 
        \DataPath/RF/bus_reg_dataout[1278] , 
        \DataPath/RF/bus_reg_dataout[1277] , 
        \DataPath/RF/bus_reg_dataout[1276] , 
        \DataPath/RF/bus_reg_dataout[1275] , 
        \DataPath/RF/bus_reg_dataout[1274] , 
        \DataPath/RF/bus_reg_dataout[1273] , 
        \DataPath/RF/bus_reg_dataout[1272] , 
        \DataPath/RF/bus_reg_dataout[1271] , 
        \DataPath/RF/bus_reg_dataout[1270] , 
        \DataPath/RF/bus_reg_dataout[1269] , 
        \DataPath/RF/bus_reg_dataout[1268] , 
        \DataPath/RF/bus_reg_dataout[1267] , 
        \DataPath/RF/bus_reg_dataout[1266] , 
        \DataPath/RF/bus_reg_dataout[1265] , 
        \DataPath/RF/bus_reg_dataout[1264] , 
        \DataPath/RF/bus_reg_dataout[1263] , 
        \DataPath/RF/bus_reg_dataout[1262] , 
        \DataPath/RF/bus_reg_dataout[1261] , 
        \DataPath/RF/bus_reg_dataout[1260] , 
        \DataPath/RF/bus_reg_dataout[1259] , 
        \DataPath/RF/bus_reg_dataout[1258] , 
        \DataPath/RF/bus_reg_dataout[1257] , 
        \DataPath/RF/bus_reg_dataout[1256] , 
        \DataPath/RF/bus_reg_dataout[1255] , 
        \DataPath/RF/bus_reg_dataout[1254] , 
        \DataPath/RF/bus_reg_dataout[1253] , 
        \DataPath/RF/bus_reg_dataout[1252] , 
        \DataPath/RF/bus_reg_dataout[1251] , 
        \DataPath/RF/bus_reg_dataout[1250] , 
        \DataPath/RF/bus_reg_dataout[1249] , 
        \DataPath/RF/bus_reg_dataout[1248] , 
        \DataPath/RF/bus_reg_dataout[1247] , 
        \DataPath/RF/bus_reg_dataout[1246] , 
        \DataPath/RF/bus_reg_dataout[1245] , 
        \DataPath/RF/bus_reg_dataout[1244] , 
        \DataPath/RF/bus_reg_dataout[1243] , 
        \DataPath/RF/bus_reg_dataout[1242] , 
        \DataPath/RF/bus_reg_dataout[1241] , 
        \DataPath/RF/bus_reg_dataout[1240] , 
        \DataPath/RF/bus_reg_dataout[1239] , 
        \DataPath/RF/bus_reg_dataout[1238] , 
        \DataPath/RF/bus_reg_dataout[1237] , 
        \DataPath/RF/bus_reg_dataout[1236] , 
        \DataPath/RF/bus_reg_dataout[1235] , 
        \DataPath/RF/bus_reg_dataout[1234] , 
        \DataPath/RF/bus_reg_dataout[1233] , 
        \DataPath/RF/bus_reg_dataout[1232] , 
        \DataPath/RF/bus_reg_dataout[1231] , 
        \DataPath/RF/bus_reg_dataout[1230] , 
        \DataPath/RF/bus_reg_dataout[1229] , 
        \DataPath/RF/bus_reg_dataout[1228] , 
        \DataPath/RF/bus_reg_dataout[1227] , 
        \DataPath/RF/bus_reg_dataout[1226] , 
        \DataPath/RF/bus_reg_dataout[1225] , 
        \DataPath/RF/bus_reg_dataout[1224] , 
        \DataPath/RF/bus_reg_dataout[1223] , 
        \DataPath/RF/bus_reg_dataout[1222] , 
        \DataPath/RF/bus_reg_dataout[1221] , 
        \DataPath/RF/bus_reg_dataout[1220] , 
        \DataPath/RF/bus_reg_dataout[1219] , 
        \DataPath/RF/bus_reg_dataout[1218] , 
        \DataPath/RF/bus_reg_dataout[1217] , 
        \DataPath/RF/bus_reg_dataout[1216] , 
        \DataPath/RF/bus_reg_dataout[1215] , 
        \DataPath/RF/bus_reg_dataout[1214] , 
        \DataPath/RF/bus_reg_dataout[1213] , 
        \DataPath/RF/bus_reg_dataout[1212] , 
        \DataPath/RF/bus_reg_dataout[1211] , 
        \DataPath/RF/bus_reg_dataout[1210] , 
        \DataPath/RF/bus_reg_dataout[1209] , 
        \DataPath/RF/bus_reg_dataout[1208] , 
        \DataPath/RF/bus_reg_dataout[1207] , 
        \DataPath/RF/bus_reg_dataout[1206] , 
        \DataPath/RF/bus_reg_dataout[1205] , 
        \DataPath/RF/bus_reg_dataout[1204] , 
        \DataPath/RF/bus_reg_dataout[1203] , 
        \DataPath/RF/bus_reg_dataout[1202] , 
        \DataPath/RF/bus_reg_dataout[1201] , 
        \DataPath/RF/bus_reg_dataout[1200] , 
        \DataPath/RF/bus_reg_dataout[1199] , 
        \DataPath/RF/bus_reg_dataout[1198] , 
        \DataPath/RF/bus_reg_dataout[1197] , 
        \DataPath/RF/bus_reg_dataout[1196] , 
        \DataPath/RF/bus_reg_dataout[1195] , 
        \DataPath/RF/bus_reg_dataout[1194] , 
        \DataPath/RF/bus_reg_dataout[1193] , 
        \DataPath/RF/bus_reg_dataout[1192] , 
        \DataPath/RF/bus_reg_dataout[1191] , 
        \DataPath/RF/bus_reg_dataout[1190] , 
        \DataPath/RF/bus_reg_dataout[1189] , 
        \DataPath/RF/bus_reg_dataout[1188] , 
        \DataPath/RF/bus_reg_dataout[1187] , 
        \DataPath/RF/bus_reg_dataout[1186] , 
        \DataPath/RF/bus_reg_dataout[1185] , 
        \DataPath/RF/bus_reg_dataout[1184] , 
        \DataPath/RF/bus_reg_dataout[1183] , 
        \DataPath/RF/bus_reg_dataout[1182] , 
        \DataPath/RF/bus_reg_dataout[1181] , 
        \DataPath/RF/bus_reg_dataout[1180] , 
        \DataPath/RF/bus_reg_dataout[1179] , 
        \DataPath/RF/bus_reg_dataout[1178] , 
        \DataPath/RF/bus_reg_dataout[1177] , 
        \DataPath/RF/bus_reg_dataout[1176] , 
        \DataPath/RF/bus_reg_dataout[1175] , 
        \DataPath/RF/bus_reg_dataout[1174] , 
        \DataPath/RF/bus_reg_dataout[1173] , 
        \DataPath/RF/bus_reg_dataout[1172] , 
        \DataPath/RF/bus_reg_dataout[1171] , 
        \DataPath/RF/bus_reg_dataout[1170] , 
        \DataPath/RF/bus_reg_dataout[1169] , 
        \DataPath/RF/bus_reg_dataout[1168] , 
        \DataPath/RF/bus_reg_dataout[1167] , 
        \DataPath/RF/bus_reg_dataout[1166] , 
        \DataPath/RF/bus_reg_dataout[1165] , 
        \DataPath/RF/bus_reg_dataout[1164] , 
        \DataPath/RF/bus_reg_dataout[1163] , 
        \DataPath/RF/bus_reg_dataout[1162] , 
        \DataPath/RF/bus_reg_dataout[1161] , 
        \DataPath/RF/bus_reg_dataout[1160] , 
        \DataPath/RF/bus_reg_dataout[1159] , 
        \DataPath/RF/bus_reg_dataout[1158] , 
        \DataPath/RF/bus_reg_dataout[1157] , 
        \DataPath/RF/bus_reg_dataout[1156] , 
        \DataPath/RF/bus_reg_dataout[1155] , 
        \DataPath/RF/bus_reg_dataout[1154] , 
        \DataPath/RF/bus_reg_dataout[1153] , 
        \DataPath/RF/bus_reg_dataout[1152] , 
        \DataPath/RF/bus_reg_dataout[1151] , 
        \DataPath/RF/bus_reg_dataout[1150] , 
        \DataPath/RF/bus_reg_dataout[1149] , 
        \DataPath/RF/bus_reg_dataout[1148] , 
        \DataPath/RF/bus_reg_dataout[1147] , 
        \DataPath/RF/bus_reg_dataout[1146] , 
        \DataPath/RF/bus_reg_dataout[1145] , 
        \DataPath/RF/bus_reg_dataout[1144] , 
        \DataPath/RF/bus_reg_dataout[1143] , 
        \DataPath/RF/bus_reg_dataout[1142] , 
        \DataPath/RF/bus_reg_dataout[1141] , 
        \DataPath/RF/bus_reg_dataout[1140] , 
        \DataPath/RF/bus_reg_dataout[1139] , 
        \DataPath/RF/bus_reg_dataout[1138] , 
        \DataPath/RF/bus_reg_dataout[1137] , 
        \DataPath/RF/bus_reg_dataout[1136] , 
        \DataPath/RF/bus_reg_dataout[1135] , 
        \DataPath/RF/bus_reg_dataout[1134] , 
        \DataPath/RF/bus_reg_dataout[1133] , 
        \DataPath/RF/bus_reg_dataout[1132] , 
        \DataPath/RF/bus_reg_dataout[1131] , 
        \DataPath/RF/bus_reg_dataout[1130] , 
        \DataPath/RF/bus_reg_dataout[1129] , 
        \DataPath/RF/bus_reg_dataout[1128] , 
        \DataPath/RF/bus_reg_dataout[1127] , 
        \DataPath/RF/bus_reg_dataout[1126] , 
        \DataPath/RF/bus_reg_dataout[1125] , 
        \DataPath/RF/bus_reg_dataout[1124] , 
        \DataPath/RF/bus_reg_dataout[1123] , 
        \DataPath/RF/bus_reg_dataout[1122] , 
        \DataPath/RF/bus_reg_dataout[1121] , 
        \DataPath/RF/bus_reg_dataout[1120] , 
        \DataPath/RF/bus_reg_dataout[1119] , 
        \DataPath/RF/bus_reg_dataout[1118] , 
        \DataPath/RF/bus_reg_dataout[1117] , 
        \DataPath/RF/bus_reg_dataout[1116] , 
        \DataPath/RF/bus_reg_dataout[1115] , 
        \DataPath/RF/bus_reg_dataout[1114] , 
        \DataPath/RF/bus_reg_dataout[1113] , 
        \DataPath/RF/bus_reg_dataout[1112] , 
        \DataPath/RF/bus_reg_dataout[1111] , 
        \DataPath/RF/bus_reg_dataout[1110] , 
        \DataPath/RF/bus_reg_dataout[1109] , 
        \DataPath/RF/bus_reg_dataout[1108] , 
        \DataPath/RF/bus_reg_dataout[1107] , 
        \DataPath/RF/bus_reg_dataout[1106] , 
        \DataPath/RF/bus_reg_dataout[1105] , 
        \DataPath/RF/bus_reg_dataout[1104] , 
        \DataPath/RF/bus_reg_dataout[1103] , 
        \DataPath/RF/bus_reg_dataout[1102] , 
        \DataPath/RF/bus_reg_dataout[1101] , 
        \DataPath/RF/bus_reg_dataout[1100] , 
        \DataPath/RF/bus_reg_dataout[1099] , 
        \DataPath/RF/bus_reg_dataout[1098] , 
        \DataPath/RF/bus_reg_dataout[1097] , 
        \DataPath/RF/bus_reg_dataout[1096] , 
        \DataPath/RF/bus_reg_dataout[1095] , 
        \DataPath/RF/bus_reg_dataout[1094] , 
        \DataPath/RF/bus_reg_dataout[1093] , 
        \DataPath/RF/bus_reg_dataout[1092] , 
        \DataPath/RF/bus_reg_dataout[1091] , 
        \DataPath/RF/bus_reg_dataout[1090] , 
        \DataPath/RF/bus_reg_dataout[1089] , 
        \DataPath/RF/bus_reg_dataout[1088] , 
        \DataPath/RF/bus_reg_dataout[1087] , 
        \DataPath/RF/bus_reg_dataout[1086] , 
        \DataPath/RF/bus_reg_dataout[1085] , 
        \DataPath/RF/bus_reg_dataout[1084] , 
        \DataPath/RF/bus_reg_dataout[1083] , 
        \DataPath/RF/bus_reg_dataout[1082] , 
        \DataPath/RF/bus_reg_dataout[1081] , 
        \DataPath/RF/bus_reg_dataout[1080] , 
        \DataPath/RF/bus_reg_dataout[1079] , 
        \DataPath/RF/bus_reg_dataout[1078] , 
        \DataPath/RF/bus_reg_dataout[1077] , 
        \DataPath/RF/bus_reg_dataout[1076] , 
        \DataPath/RF/bus_reg_dataout[1075] , 
        \DataPath/RF/bus_reg_dataout[1074] , 
        \DataPath/RF/bus_reg_dataout[1073] , 
        \DataPath/RF/bus_reg_dataout[1072] , 
        \DataPath/RF/bus_reg_dataout[1071] , 
        \DataPath/RF/bus_reg_dataout[1070] , 
        \DataPath/RF/bus_reg_dataout[1069] , 
        \DataPath/RF/bus_reg_dataout[1068] , 
        \DataPath/RF/bus_reg_dataout[1067] , 
        \DataPath/RF/bus_reg_dataout[1066] , 
        \DataPath/RF/bus_reg_dataout[1065] , 
        \DataPath/RF/bus_reg_dataout[1064] , 
        \DataPath/RF/bus_reg_dataout[1063] , 
        \DataPath/RF/bus_reg_dataout[1062] , 
        \DataPath/RF/bus_reg_dataout[1061] , 
        \DataPath/RF/bus_reg_dataout[1060] , 
        \DataPath/RF/bus_reg_dataout[1059] , 
        \DataPath/RF/bus_reg_dataout[1058] , 
        \DataPath/RF/bus_reg_dataout[1057] , 
        \DataPath/RF/bus_reg_dataout[1056] , 
        \DataPath/RF/bus_reg_dataout[1055] , 
        \DataPath/RF/bus_reg_dataout[1054] , 
        \DataPath/RF/bus_reg_dataout[1053] , 
        \DataPath/RF/bus_reg_dataout[1052] , 
        \DataPath/RF/bus_reg_dataout[1051] , 
        \DataPath/RF/bus_reg_dataout[1050] , 
        \DataPath/RF/bus_reg_dataout[1049] , 
        \DataPath/RF/bus_reg_dataout[1048] , 
        \DataPath/RF/bus_reg_dataout[1047] , 
        \DataPath/RF/bus_reg_dataout[1046] , 
        \DataPath/RF/bus_reg_dataout[1045] , 
        \DataPath/RF/bus_reg_dataout[1044] , 
        \DataPath/RF/bus_reg_dataout[1043] , 
        \DataPath/RF/bus_reg_dataout[1042] , 
        \DataPath/RF/bus_reg_dataout[1041] , 
        \DataPath/RF/bus_reg_dataout[1040] , 
        \DataPath/RF/bus_reg_dataout[1039] , 
        \DataPath/RF/bus_reg_dataout[1038] , 
        \DataPath/RF/bus_reg_dataout[1037] , 
        \DataPath/RF/bus_reg_dataout[1036] , 
        \DataPath/RF/bus_reg_dataout[1035] , 
        \DataPath/RF/bus_reg_dataout[1034] , 
        \DataPath/RF/bus_reg_dataout[1033] , 
        \DataPath/RF/bus_reg_dataout[1032] , 
        \DataPath/RF/bus_reg_dataout[1031] , 
        \DataPath/RF/bus_reg_dataout[1030] , 
        \DataPath/RF/bus_reg_dataout[1029] , 
        \DataPath/RF/bus_reg_dataout[1028] , 
        \DataPath/RF/bus_reg_dataout[1027] , 
        \DataPath/RF/bus_reg_dataout[1026] , 
        \DataPath/RF/bus_reg_dataout[1025] , 
        \DataPath/RF/bus_reg_dataout[1024] , 
        \DataPath/RF/bus_reg_dataout[1023] , 
        \DataPath/RF/bus_reg_dataout[1022] , 
        \DataPath/RF/bus_reg_dataout[1021] , 
        \DataPath/RF/bus_reg_dataout[1020] , 
        \DataPath/RF/bus_reg_dataout[1019] , 
        \DataPath/RF/bus_reg_dataout[1018] , 
        \DataPath/RF/bus_reg_dataout[1017] , 
        \DataPath/RF/bus_reg_dataout[1016] , 
        \DataPath/RF/bus_reg_dataout[1015] , 
        \DataPath/RF/bus_reg_dataout[1014] , 
        \DataPath/RF/bus_reg_dataout[1013] , 
        \DataPath/RF/bus_reg_dataout[1012] , 
        \DataPath/RF/bus_reg_dataout[1011] , 
        \DataPath/RF/bus_reg_dataout[1010] , 
        \DataPath/RF/bus_reg_dataout[1009] , 
        \DataPath/RF/bus_reg_dataout[1008] , 
        \DataPath/RF/bus_reg_dataout[1007] , 
        \DataPath/RF/bus_reg_dataout[1006] , 
        \DataPath/RF/bus_reg_dataout[1005] , 
        \DataPath/RF/bus_reg_dataout[1004] , 
        \DataPath/RF/bus_reg_dataout[1003] , 
        \DataPath/RF/bus_reg_dataout[1002] , 
        \DataPath/RF/bus_reg_dataout[1001] , 
        \DataPath/RF/bus_reg_dataout[1000] , 
        \DataPath/RF/bus_reg_dataout[999] , \DataPath/RF/bus_reg_dataout[998] , 
        \DataPath/RF/bus_reg_dataout[997] , \DataPath/RF/bus_reg_dataout[996] , 
        \DataPath/RF/bus_reg_dataout[995] , \DataPath/RF/bus_reg_dataout[994] , 
        \DataPath/RF/bus_reg_dataout[993] , \DataPath/RF/bus_reg_dataout[992] , 
        \DataPath/RF/bus_reg_dataout[991] , \DataPath/RF/bus_reg_dataout[990] , 
        \DataPath/RF/bus_reg_dataout[989] , \DataPath/RF/bus_reg_dataout[988] , 
        \DataPath/RF/bus_reg_dataout[987] , \DataPath/RF/bus_reg_dataout[986] , 
        \DataPath/RF/bus_reg_dataout[985] , \DataPath/RF/bus_reg_dataout[984] , 
        \DataPath/RF/bus_reg_dataout[983] , \DataPath/RF/bus_reg_dataout[982] , 
        \DataPath/RF/bus_reg_dataout[981] , \DataPath/RF/bus_reg_dataout[980] , 
        \DataPath/RF/bus_reg_dataout[979] , \DataPath/RF/bus_reg_dataout[978] , 
        \DataPath/RF/bus_reg_dataout[977] , \DataPath/RF/bus_reg_dataout[976] , 
        \DataPath/RF/bus_reg_dataout[975] , \DataPath/RF/bus_reg_dataout[974] , 
        \DataPath/RF/bus_reg_dataout[973] , \DataPath/RF/bus_reg_dataout[972] , 
        \DataPath/RF/bus_reg_dataout[971] , \DataPath/RF/bus_reg_dataout[970] , 
        \DataPath/RF/bus_reg_dataout[969] , \DataPath/RF/bus_reg_dataout[968] , 
        \DataPath/RF/bus_reg_dataout[967] , \DataPath/RF/bus_reg_dataout[966] , 
        \DataPath/RF/bus_reg_dataout[965] , \DataPath/RF/bus_reg_dataout[964] , 
        \DataPath/RF/bus_reg_dataout[963] , \DataPath/RF/bus_reg_dataout[962] , 
        \DataPath/RF/bus_reg_dataout[961] , \DataPath/RF/bus_reg_dataout[960] , 
        \DataPath/RF/bus_reg_dataout[959] , \DataPath/RF/bus_reg_dataout[958] , 
        \DataPath/RF/bus_reg_dataout[957] , \DataPath/RF/bus_reg_dataout[956] , 
        \DataPath/RF/bus_reg_dataout[955] , \DataPath/RF/bus_reg_dataout[954] , 
        \DataPath/RF/bus_reg_dataout[953] , \DataPath/RF/bus_reg_dataout[952] , 
        \DataPath/RF/bus_reg_dataout[951] , \DataPath/RF/bus_reg_dataout[950] , 
        \DataPath/RF/bus_reg_dataout[949] , \DataPath/RF/bus_reg_dataout[948] , 
        \DataPath/RF/bus_reg_dataout[947] , \DataPath/RF/bus_reg_dataout[946] , 
        \DataPath/RF/bus_reg_dataout[945] , \DataPath/RF/bus_reg_dataout[944] , 
        \DataPath/RF/bus_reg_dataout[943] , \DataPath/RF/bus_reg_dataout[942] , 
        \DataPath/RF/bus_reg_dataout[941] , \DataPath/RF/bus_reg_dataout[940] , 
        \DataPath/RF/bus_reg_dataout[939] , \DataPath/RF/bus_reg_dataout[938] , 
        \DataPath/RF/bus_reg_dataout[937] , \DataPath/RF/bus_reg_dataout[936] , 
        \DataPath/RF/bus_reg_dataout[935] , \DataPath/RF/bus_reg_dataout[934] , 
        \DataPath/RF/bus_reg_dataout[933] , \DataPath/RF/bus_reg_dataout[932] , 
        \DataPath/RF/bus_reg_dataout[931] , \DataPath/RF/bus_reg_dataout[930] , 
        \DataPath/RF/bus_reg_dataout[929] , \DataPath/RF/bus_reg_dataout[928] , 
        \DataPath/RF/bus_reg_dataout[927] , \DataPath/RF/bus_reg_dataout[926] , 
        \DataPath/RF/bus_reg_dataout[925] , \DataPath/RF/bus_reg_dataout[924] , 
        \DataPath/RF/bus_reg_dataout[923] , \DataPath/RF/bus_reg_dataout[922] , 
        \DataPath/RF/bus_reg_dataout[921] , \DataPath/RF/bus_reg_dataout[920] , 
        \DataPath/RF/bus_reg_dataout[919] , \DataPath/RF/bus_reg_dataout[918] , 
        \DataPath/RF/bus_reg_dataout[917] , \DataPath/RF/bus_reg_dataout[916] , 
        \DataPath/RF/bus_reg_dataout[915] , \DataPath/RF/bus_reg_dataout[914] , 
        \DataPath/RF/bus_reg_dataout[913] , \DataPath/RF/bus_reg_dataout[912] , 
        \DataPath/RF/bus_reg_dataout[911] , \DataPath/RF/bus_reg_dataout[910] , 
        \DataPath/RF/bus_reg_dataout[909] , \DataPath/RF/bus_reg_dataout[908] , 
        \DataPath/RF/bus_reg_dataout[907] , \DataPath/RF/bus_reg_dataout[906] , 
        \DataPath/RF/bus_reg_dataout[905] , \DataPath/RF/bus_reg_dataout[904] , 
        \DataPath/RF/bus_reg_dataout[903] , \DataPath/RF/bus_reg_dataout[902] , 
        \DataPath/RF/bus_reg_dataout[901] , \DataPath/RF/bus_reg_dataout[900] , 
        \DataPath/RF/bus_reg_dataout[899] , \DataPath/RF/bus_reg_dataout[898] , 
        \DataPath/RF/bus_reg_dataout[897] , \DataPath/RF/bus_reg_dataout[896] , 
        \DataPath/RF/bus_reg_dataout[895] , \DataPath/RF/bus_reg_dataout[894] , 
        \DataPath/RF/bus_reg_dataout[893] , \DataPath/RF/bus_reg_dataout[892] , 
        \DataPath/RF/bus_reg_dataout[891] , \DataPath/RF/bus_reg_dataout[890] , 
        \DataPath/RF/bus_reg_dataout[889] , \DataPath/RF/bus_reg_dataout[888] , 
        \DataPath/RF/bus_reg_dataout[887] , \DataPath/RF/bus_reg_dataout[886] , 
        \DataPath/RF/bus_reg_dataout[885] , \DataPath/RF/bus_reg_dataout[884] , 
        \DataPath/RF/bus_reg_dataout[883] , \DataPath/RF/bus_reg_dataout[882] , 
        \DataPath/RF/bus_reg_dataout[881] , \DataPath/RF/bus_reg_dataout[880] , 
        \DataPath/RF/bus_reg_dataout[879] , \DataPath/RF/bus_reg_dataout[878] , 
        \DataPath/RF/bus_reg_dataout[877] , \DataPath/RF/bus_reg_dataout[876] , 
        \DataPath/RF/bus_reg_dataout[875] , \DataPath/RF/bus_reg_dataout[874] , 
        \DataPath/RF/bus_reg_dataout[873] , \DataPath/RF/bus_reg_dataout[872] , 
        \DataPath/RF/bus_reg_dataout[871] , \DataPath/RF/bus_reg_dataout[870] , 
        \DataPath/RF/bus_reg_dataout[869] , \DataPath/RF/bus_reg_dataout[868] , 
        \DataPath/RF/bus_reg_dataout[867] , \DataPath/RF/bus_reg_dataout[866] , 
        \DataPath/RF/bus_reg_dataout[865] , \DataPath/RF/bus_reg_dataout[864] , 
        \DataPath/RF/bus_reg_dataout[863] , \DataPath/RF/bus_reg_dataout[862] , 
        \DataPath/RF/bus_reg_dataout[861] , \DataPath/RF/bus_reg_dataout[860] , 
        \DataPath/RF/bus_reg_dataout[859] , \DataPath/RF/bus_reg_dataout[858] , 
        \DataPath/RF/bus_reg_dataout[857] , \DataPath/RF/bus_reg_dataout[856] , 
        \DataPath/RF/bus_reg_dataout[855] , \DataPath/RF/bus_reg_dataout[854] , 
        \DataPath/RF/bus_reg_dataout[853] , \DataPath/RF/bus_reg_dataout[852] , 
        \DataPath/RF/bus_reg_dataout[851] , \DataPath/RF/bus_reg_dataout[850] , 
        \DataPath/RF/bus_reg_dataout[849] , \DataPath/RF/bus_reg_dataout[848] , 
        \DataPath/RF/bus_reg_dataout[847] , \DataPath/RF/bus_reg_dataout[846] , 
        \DataPath/RF/bus_reg_dataout[845] , \DataPath/RF/bus_reg_dataout[844] , 
        \DataPath/RF/bus_reg_dataout[843] , \DataPath/RF/bus_reg_dataout[842] , 
        \DataPath/RF/bus_reg_dataout[841] , \DataPath/RF/bus_reg_dataout[840] , 
        \DataPath/RF/bus_reg_dataout[839] , \DataPath/RF/bus_reg_dataout[838] , 
        \DataPath/RF/bus_reg_dataout[837] , \DataPath/RF/bus_reg_dataout[836] , 
        \DataPath/RF/bus_reg_dataout[835] , \DataPath/RF/bus_reg_dataout[834] , 
        \DataPath/RF/bus_reg_dataout[833] , \DataPath/RF/bus_reg_dataout[832] , 
        \DataPath/RF/bus_reg_dataout[831] , \DataPath/RF/bus_reg_dataout[830] , 
        \DataPath/RF/bus_reg_dataout[829] , \DataPath/RF/bus_reg_dataout[828] , 
        \DataPath/RF/bus_reg_dataout[827] , \DataPath/RF/bus_reg_dataout[826] , 
        \DataPath/RF/bus_reg_dataout[825] , \DataPath/RF/bus_reg_dataout[824] , 
        \DataPath/RF/bus_reg_dataout[823] , \DataPath/RF/bus_reg_dataout[822] , 
        \DataPath/RF/bus_reg_dataout[821] , \DataPath/RF/bus_reg_dataout[820] , 
        \DataPath/RF/bus_reg_dataout[819] , \DataPath/RF/bus_reg_dataout[818] , 
        \DataPath/RF/bus_reg_dataout[817] , \DataPath/RF/bus_reg_dataout[816] , 
        \DataPath/RF/bus_reg_dataout[815] , \DataPath/RF/bus_reg_dataout[814] , 
        \DataPath/RF/bus_reg_dataout[813] , \DataPath/RF/bus_reg_dataout[812] , 
        \DataPath/RF/bus_reg_dataout[811] , \DataPath/RF/bus_reg_dataout[810] , 
        \DataPath/RF/bus_reg_dataout[809] , \DataPath/RF/bus_reg_dataout[808] , 
        \DataPath/RF/bus_reg_dataout[807] , \DataPath/RF/bus_reg_dataout[806] , 
        \DataPath/RF/bus_reg_dataout[805] , \DataPath/RF/bus_reg_dataout[804] , 
        \DataPath/RF/bus_reg_dataout[803] , \DataPath/RF/bus_reg_dataout[802] , 
        \DataPath/RF/bus_reg_dataout[801] , \DataPath/RF/bus_reg_dataout[800] , 
        \DataPath/RF/bus_reg_dataout[799] , \DataPath/RF/bus_reg_dataout[798] , 
        \DataPath/RF/bus_reg_dataout[797] , \DataPath/RF/bus_reg_dataout[796] , 
        \DataPath/RF/bus_reg_dataout[795] , \DataPath/RF/bus_reg_dataout[794] , 
        \DataPath/RF/bus_reg_dataout[793] , \DataPath/RF/bus_reg_dataout[792] , 
        \DataPath/RF/bus_reg_dataout[791] , \DataPath/RF/bus_reg_dataout[790] , 
        \DataPath/RF/bus_reg_dataout[789] , \DataPath/RF/bus_reg_dataout[788] , 
        \DataPath/RF/bus_reg_dataout[787] , \DataPath/RF/bus_reg_dataout[786] , 
        \DataPath/RF/bus_reg_dataout[785] , \DataPath/RF/bus_reg_dataout[784] , 
        \DataPath/RF/bus_reg_dataout[783] , \DataPath/RF/bus_reg_dataout[782] , 
        \DataPath/RF/bus_reg_dataout[781] , \DataPath/RF/bus_reg_dataout[780] , 
        \DataPath/RF/bus_reg_dataout[779] , \DataPath/RF/bus_reg_dataout[778] , 
        \DataPath/RF/bus_reg_dataout[777] , \DataPath/RF/bus_reg_dataout[776] , 
        \DataPath/RF/bus_reg_dataout[775] , \DataPath/RF/bus_reg_dataout[774] , 
        \DataPath/RF/bus_reg_dataout[773] , \DataPath/RF/bus_reg_dataout[772] , 
        \DataPath/RF/bus_reg_dataout[771] , \DataPath/RF/bus_reg_dataout[770] , 
        \DataPath/RF/bus_reg_dataout[769] , \DataPath/RF/bus_reg_dataout[768] , 
        \DataPath/RF/bus_reg_dataout[767] , \DataPath/RF/bus_reg_dataout[766] , 
        \DataPath/RF/bus_reg_dataout[765] , \DataPath/RF/bus_reg_dataout[764] , 
        \DataPath/RF/bus_reg_dataout[763] , \DataPath/RF/bus_reg_dataout[762] , 
        \DataPath/RF/bus_reg_dataout[761] , \DataPath/RF/bus_reg_dataout[760] , 
        \DataPath/RF/bus_reg_dataout[759] , \DataPath/RF/bus_reg_dataout[758] , 
        \DataPath/RF/bus_reg_dataout[757] , \DataPath/RF/bus_reg_dataout[756] , 
        \DataPath/RF/bus_reg_dataout[755] , \DataPath/RF/bus_reg_dataout[754] , 
        \DataPath/RF/bus_reg_dataout[753] , \DataPath/RF/bus_reg_dataout[752] , 
        \DataPath/RF/bus_reg_dataout[751] , \DataPath/RF/bus_reg_dataout[750] , 
        \DataPath/RF/bus_reg_dataout[749] , \DataPath/RF/bus_reg_dataout[748] , 
        \DataPath/RF/bus_reg_dataout[747] , \DataPath/RF/bus_reg_dataout[746] , 
        \DataPath/RF/bus_reg_dataout[745] , \DataPath/RF/bus_reg_dataout[744] , 
        \DataPath/RF/bus_reg_dataout[743] , \DataPath/RF/bus_reg_dataout[742] , 
        \DataPath/RF/bus_reg_dataout[741] , \DataPath/RF/bus_reg_dataout[740] , 
        \DataPath/RF/bus_reg_dataout[739] , \DataPath/RF/bus_reg_dataout[738] , 
        \DataPath/RF/bus_reg_dataout[737] , \DataPath/RF/bus_reg_dataout[736] , 
        \DataPath/RF/bus_reg_dataout[735] , \DataPath/RF/bus_reg_dataout[734] , 
        \DataPath/RF/bus_reg_dataout[733] , \DataPath/RF/bus_reg_dataout[732] , 
        \DataPath/RF/bus_reg_dataout[731] , \DataPath/RF/bus_reg_dataout[730] , 
        \DataPath/RF/bus_reg_dataout[729] , \DataPath/RF/bus_reg_dataout[728] , 
        \DataPath/RF/bus_reg_dataout[727] , \DataPath/RF/bus_reg_dataout[726] , 
        \DataPath/RF/bus_reg_dataout[725] , \DataPath/RF/bus_reg_dataout[724] , 
        \DataPath/RF/bus_reg_dataout[723] , \DataPath/RF/bus_reg_dataout[722] , 
        \DataPath/RF/bus_reg_dataout[721] , \DataPath/RF/bus_reg_dataout[720] , 
        \DataPath/RF/bus_reg_dataout[719] , \DataPath/RF/bus_reg_dataout[718] , 
        \DataPath/RF/bus_reg_dataout[717] , \DataPath/RF/bus_reg_dataout[716] , 
        \DataPath/RF/bus_reg_dataout[715] , \DataPath/RF/bus_reg_dataout[714] , 
        \DataPath/RF/bus_reg_dataout[713] , \DataPath/RF/bus_reg_dataout[712] , 
        \DataPath/RF/bus_reg_dataout[711] , \DataPath/RF/bus_reg_dataout[710] , 
        \DataPath/RF/bus_reg_dataout[709] , \DataPath/RF/bus_reg_dataout[708] , 
        \DataPath/RF/bus_reg_dataout[707] , \DataPath/RF/bus_reg_dataout[706] , 
        \DataPath/RF/bus_reg_dataout[705] , \DataPath/RF/bus_reg_dataout[704] , 
        \DataPath/RF/bus_reg_dataout[703] , \DataPath/RF/bus_reg_dataout[702] , 
        \DataPath/RF/bus_reg_dataout[701] , \DataPath/RF/bus_reg_dataout[700] , 
        \DataPath/RF/bus_reg_dataout[699] , \DataPath/RF/bus_reg_dataout[698] , 
        \DataPath/RF/bus_reg_dataout[697] , \DataPath/RF/bus_reg_dataout[696] , 
        \DataPath/RF/bus_reg_dataout[695] , \DataPath/RF/bus_reg_dataout[694] , 
        \DataPath/RF/bus_reg_dataout[693] , \DataPath/RF/bus_reg_dataout[692] , 
        \DataPath/RF/bus_reg_dataout[691] , \DataPath/RF/bus_reg_dataout[690] , 
        \DataPath/RF/bus_reg_dataout[689] , \DataPath/RF/bus_reg_dataout[688] , 
        \DataPath/RF/bus_reg_dataout[687] , \DataPath/RF/bus_reg_dataout[686] , 
        \DataPath/RF/bus_reg_dataout[685] , \DataPath/RF/bus_reg_dataout[684] , 
        \DataPath/RF/bus_reg_dataout[683] , \DataPath/RF/bus_reg_dataout[682] , 
        \DataPath/RF/bus_reg_dataout[681] , \DataPath/RF/bus_reg_dataout[680] , 
        \DataPath/RF/bus_reg_dataout[679] , \DataPath/RF/bus_reg_dataout[678] , 
        \DataPath/RF/bus_reg_dataout[677] , \DataPath/RF/bus_reg_dataout[676] , 
        \DataPath/RF/bus_reg_dataout[675] , \DataPath/RF/bus_reg_dataout[674] , 
        \DataPath/RF/bus_reg_dataout[673] , \DataPath/RF/bus_reg_dataout[672] , 
        \DataPath/RF/bus_reg_dataout[671] , \DataPath/RF/bus_reg_dataout[670] , 
        \DataPath/RF/bus_reg_dataout[669] , \DataPath/RF/bus_reg_dataout[668] , 
        \DataPath/RF/bus_reg_dataout[667] , \DataPath/RF/bus_reg_dataout[666] , 
        \DataPath/RF/bus_reg_dataout[665] , \DataPath/RF/bus_reg_dataout[664] , 
        \DataPath/RF/bus_reg_dataout[663] , \DataPath/RF/bus_reg_dataout[662] , 
        \DataPath/RF/bus_reg_dataout[661] , \DataPath/RF/bus_reg_dataout[660] , 
        \DataPath/RF/bus_reg_dataout[659] , \DataPath/RF/bus_reg_dataout[658] , 
        \DataPath/RF/bus_reg_dataout[657] , \DataPath/RF/bus_reg_dataout[656] , 
        \DataPath/RF/bus_reg_dataout[655] , \DataPath/RF/bus_reg_dataout[654] , 
        \DataPath/RF/bus_reg_dataout[653] , \DataPath/RF/bus_reg_dataout[652] , 
        \DataPath/RF/bus_reg_dataout[651] , \DataPath/RF/bus_reg_dataout[650] , 
        \DataPath/RF/bus_reg_dataout[649] , \DataPath/RF/bus_reg_dataout[648] , 
        \DataPath/RF/bus_reg_dataout[647] , \DataPath/RF/bus_reg_dataout[646] , 
        \DataPath/RF/bus_reg_dataout[645] , \DataPath/RF/bus_reg_dataout[644] , 
        \DataPath/RF/bus_reg_dataout[643] , \DataPath/RF/bus_reg_dataout[642] , 
        \DataPath/RF/bus_reg_dataout[641] , \DataPath/RF/bus_reg_dataout[640] , 
        \DataPath/RF/bus_reg_dataout[639] , \DataPath/RF/bus_reg_dataout[638] , 
        \DataPath/RF/bus_reg_dataout[637] , \DataPath/RF/bus_reg_dataout[636] , 
        \DataPath/RF/bus_reg_dataout[635] , \DataPath/RF/bus_reg_dataout[634] , 
        \DataPath/RF/bus_reg_dataout[633] , \DataPath/RF/bus_reg_dataout[632] , 
        \DataPath/RF/bus_reg_dataout[631] , \DataPath/RF/bus_reg_dataout[630] , 
        \DataPath/RF/bus_reg_dataout[629] , \DataPath/RF/bus_reg_dataout[628] , 
        \DataPath/RF/bus_reg_dataout[627] , \DataPath/RF/bus_reg_dataout[626] , 
        \DataPath/RF/bus_reg_dataout[625] , \DataPath/RF/bus_reg_dataout[624] , 
        \DataPath/RF/bus_reg_dataout[623] , \DataPath/RF/bus_reg_dataout[622] , 
        \DataPath/RF/bus_reg_dataout[621] , \DataPath/RF/bus_reg_dataout[620] , 
        \DataPath/RF/bus_reg_dataout[619] , \DataPath/RF/bus_reg_dataout[618] , 
        \DataPath/RF/bus_reg_dataout[617] , \DataPath/RF/bus_reg_dataout[616] , 
        \DataPath/RF/bus_reg_dataout[615] , \DataPath/RF/bus_reg_dataout[614] , 
        \DataPath/RF/bus_reg_dataout[613] , \DataPath/RF/bus_reg_dataout[612] , 
        \DataPath/RF/bus_reg_dataout[611] , \DataPath/RF/bus_reg_dataout[610] , 
        \DataPath/RF/bus_reg_dataout[609] , \DataPath/RF/bus_reg_dataout[608] , 
        \DataPath/RF/bus_reg_dataout[607] , \DataPath/RF/bus_reg_dataout[606] , 
        \DataPath/RF/bus_reg_dataout[605] , \DataPath/RF/bus_reg_dataout[604] , 
        \DataPath/RF/bus_reg_dataout[603] , \DataPath/RF/bus_reg_dataout[602] , 
        \DataPath/RF/bus_reg_dataout[601] , \DataPath/RF/bus_reg_dataout[600] , 
        \DataPath/RF/bus_reg_dataout[599] , \DataPath/RF/bus_reg_dataout[598] , 
        \DataPath/RF/bus_reg_dataout[597] , \DataPath/RF/bus_reg_dataout[596] , 
        \DataPath/RF/bus_reg_dataout[595] , \DataPath/RF/bus_reg_dataout[594] , 
        \DataPath/RF/bus_reg_dataout[593] , \DataPath/RF/bus_reg_dataout[592] , 
        \DataPath/RF/bus_reg_dataout[591] , \DataPath/RF/bus_reg_dataout[590] , 
        \DataPath/RF/bus_reg_dataout[589] , \DataPath/RF/bus_reg_dataout[588] , 
        \DataPath/RF/bus_reg_dataout[587] , \DataPath/RF/bus_reg_dataout[586] , 
        \DataPath/RF/bus_reg_dataout[585] , \DataPath/RF/bus_reg_dataout[584] , 
        \DataPath/RF/bus_reg_dataout[583] , \DataPath/RF/bus_reg_dataout[582] , 
        \DataPath/RF/bus_reg_dataout[581] , \DataPath/RF/bus_reg_dataout[580] , 
        \DataPath/RF/bus_reg_dataout[579] , \DataPath/RF/bus_reg_dataout[578] , 
        \DataPath/RF/bus_reg_dataout[577] , \DataPath/RF/bus_reg_dataout[576] , 
        \DataPath/RF/bus_reg_dataout[575] , \DataPath/RF/bus_reg_dataout[574] , 
        \DataPath/RF/bus_reg_dataout[573] , \DataPath/RF/bus_reg_dataout[572] , 
        \DataPath/RF/bus_reg_dataout[571] , \DataPath/RF/bus_reg_dataout[570] , 
        \DataPath/RF/bus_reg_dataout[569] , \DataPath/RF/bus_reg_dataout[568] , 
        \DataPath/RF/bus_reg_dataout[567] , \DataPath/RF/bus_reg_dataout[566] , 
        \DataPath/RF/bus_reg_dataout[565] , \DataPath/RF/bus_reg_dataout[564] , 
        \DataPath/RF/bus_reg_dataout[563] , \DataPath/RF/bus_reg_dataout[562] , 
        \DataPath/RF/bus_reg_dataout[561] , \DataPath/RF/bus_reg_dataout[560] , 
        \DataPath/RF/bus_reg_dataout[559] , \DataPath/RF/bus_reg_dataout[558] , 
        \DataPath/RF/bus_reg_dataout[557] , \DataPath/RF/bus_reg_dataout[556] , 
        \DataPath/RF/bus_reg_dataout[555] , \DataPath/RF/bus_reg_dataout[554] , 
        \DataPath/RF/bus_reg_dataout[553] , \DataPath/RF/bus_reg_dataout[552] , 
        \DataPath/RF/bus_reg_dataout[551] , \DataPath/RF/bus_reg_dataout[550] , 
        \DataPath/RF/bus_reg_dataout[549] , \DataPath/RF/bus_reg_dataout[548] , 
        \DataPath/RF/bus_reg_dataout[547] , \DataPath/RF/bus_reg_dataout[546] , 
        \DataPath/RF/bus_reg_dataout[545] , \DataPath/RF/bus_reg_dataout[544] , 
        \DataPath/RF/bus_reg_dataout[543] , \DataPath/RF/bus_reg_dataout[542] , 
        \DataPath/RF/bus_reg_dataout[541] , \DataPath/RF/bus_reg_dataout[540] , 
        \DataPath/RF/bus_reg_dataout[539] , \DataPath/RF/bus_reg_dataout[538] , 
        \DataPath/RF/bus_reg_dataout[537] , \DataPath/RF/bus_reg_dataout[536] , 
        \DataPath/RF/bus_reg_dataout[535] , \DataPath/RF/bus_reg_dataout[534] , 
        \DataPath/RF/bus_reg_dataout[533] , \DataPath/RF/bus_reg_dataout[532] , 
        \DataPath/RF/bus_reg_dataout[531] , \DataPath/RF/bus_reg_dataout[530] , 
        \DataPath/RF/bus_reg_dataout[529] , \DataPath/RF/bus_reg_dataout[528] , 
        \DataPath/RF/bus_reg_dataout[527] , \DataPath/RF/bus_reg_dataout[526] , 
        \DataPath/RF/bus_reg_dataout[525] , \DataPath/RF/bus_reg_dataout[524] , 
        \DataPath/RF/bus_reg_dataout[523] , \DataPath/RF/bus_reg_dataout[522] , 
        \DataPath/RF/bus_reg_dataout[521] , \DataPath/RF/bus_reg_dataout[520] , 
        \DataPath/RF/bus_reg_dataout[519] , \DataPath/RF/bus_reg_dataout[518] , 
        \DataPath/RF/bus_reg_dataout[517] , \DataPath/RF/bus_reg_dataout[516] , 
        \DataPath/RF/bus_reg_dataout[515] , \DataPath/RF/bus_reg_dataout[514] , 
        \DataPath/RF/bus_reg_dataout[513] , \DataPath/RF/bus_reg_dataout[512] , 
        \DataPath/RF/bus_reg_dataout[511] , \DataPath/RF/bus_reg_dataout[510] , 
        \DataPath/RF/bus_reg_dataout[509] , \DataPath/RF/bus_reg_dataout[508] , 
        \DataPath/RF/bus_reg_dataout[507] , \DataPath/RF/bus_reg_dataout[506] , 
        \DataPath/RF/bus_reg_dataout[505] , \DataPath/RF/bus_reg_dataout[504] , 
        \DataPath/RF/bus_reg_dataout[503] , \DataPath/RF/bus_reg_dataout[502] , 
        \DataPath/RF/bus_reg_dataout[501] , \DataPath/RF/bus_reg_dataout[500] , 
        \DataPath/RF/bus_reg_dataout[499] , \DataPath/RF/bus_reg_dataout[498] , 
        \DataPath/RF/bus_reg_dataout[497] , \DataPath/RF/bus_reg_dataout[496] , 
        \DataPath/RF/bus_reg_dataout[495] , \DataPath/RF/bus_reg_dataout[494] , 
        \DataPath/RF/bus_reg_dataout[493] , \DataPath/RF/bus_reg_dataout[492] , 
        \DataPath/RF/bus_reg_dataout[491] , \DataPath/RF/bus_reg_dataout[490] , 
        \DataPath/RF/bus_reg_dataout[489] , \DataPath/RF/bus_reg_dataout[488] , 
        \DataPath/RF/bus_reg_dataout[487] , \DataPath/RF/bus_reg_dataout[486] , 
        \DataPath/RF/bus_reg_dataout[485] , \DataPath/RF/bus_reg_dataout[484] , 
        \DataPath/RF/bus_reg_dataout[483] , \DataPath/RF/bus_reg_dataout[482] , 
        \DataPath/RF/bus_reg_dataout[481] , \DataPath/RF/bus_reg_dataout[480] , 
        \DataPath/RF/bus_reg_dataout[479] , \DataPath/RF/bus_reg_dataout[478] , 
        \DataPath/RF/bus_reg_dataout[477] , \DataPath/RF/bus_reg_dataout[476] , 
        \DataPath/RF/bus_reg_dataout[475] , \DataPath/RF/bus_reg_dataout[474] , 
        \DataPath/RF/bus_reg_dataout[473] , \DataPath/RF/bus_reg_dataout[472] , 
        \DataPath/RF/bus_reg_dataout[471] , \DataPath/RF/bus_reg_dataout[470] , 
        \DataPath/RF/bus_reg_dataout[469] , \DataPath/RF/bus_reg_dataout[468] , 
        \DataPath/RF/bus_reg_dataout[467] , \DataPath/RF/bus_reg_dataout[466] , 
        \DataPath/RF/bus_reg_dataout[465] , \DataPath/RF/bus_reg_dataout[464] , 
        \DataPath/RF/bus_reg_dataout[463] , \DataPath/RF/bus_reg_dataout[462] , 
        \DataPath/RF/bus_reg_dataout[461] , \DataPath/RF/bus_reg_dataout[460] , 
        \DataPath/RF/bus_reg_dataout[459] , \DataPath/RF/bus_reg_dataout[458] , 
        \DataPath/RF/bus_reg_dataout[457] , \DataPath/RF/bus_reg_dataout[456] , 
        \DataPath/RF/bus_reg_dataout[455] , \DataPath/RF/bus_reg_dataout[454] , 
        \DataPath/RF/bus_reg_dataout[453] , \DataPath/RF/bus_reg_dataout[452] , 
        \DataPath/RF/bus_reg_dataout[451] , \DataPath/RF/bus_reg_dataout[450] , 
        \DataPath/RF/bus_reg_dataout[449] , \DataPath/RF/bus_reg_dataout[448] , 
        \DataPath/RF/bus_reg_dataout[447] , \DataPath/RF/bus_reg_dataout[446] , 
        \DataPath/RF/bus_reg_dataout[445] , \DataPath/RF/bus_reg_dataout[444] , 
        \DataPath/RF/bus_reg_dataout[443] , \DataPath/RF/bus_reg_dataout[442] , 
        \DataPath/RF/bus_reg_dataout[441] , \DataPath/RF/bus_reg_dataout[440] , 
        \DataPath/RF/bus_reg_dataout[439] , \DataPath/RF/bus_reg_dataout[438] , 
        \DataPath/RF/bus_reg_dataout[437] , \DataPath/RF/bus_reg_dataout[436] , 
        \DataPath/RF/bus_reg_dataout[435] , \DataPath/RF/bus_reg_dataout[434] , 
        \DataPath/RF/bus_reg_dataout[433] , \DataPath/RF/bus_reg_dataout[432] , 
        \DataPath/RF/bus_reg_dataout[431] , \DataPath/RF/bus_reg_dataout[430] , 
        \DataPath/RF/bus_reg_dataout[429] , \DataPath/RF/bus_reg_dataout[428] , 
        \DataPath/RF/bus_reg_dataout[427] , \DataPath/RF/bus_reg_dataout[426] , 
        \DataPath/RF/bus_reg_dataout[425] , \DataPath/RF/bus_reg_dataout[424] , 
        \DataPath/RF/bus_reg_dataout[423] , \DataPath/RF/bus_reg_dataout[422] , 
        \DataPath/RF/bus_reg_dataout[421] , \DataPath/RF/bus_reg_dataout[420] , 
        \DataPath/RF/bus_reg_dataout[419] , \DataPath/RF/bus_reg_dataout[418] , 
        \DataPath/RF/bus_reg_dataout[417] , \DataPath/RF/bus_reg_dataout[416] , 
        \DataPath/RF/bus_reg_dataout[415] , \DataPath/RF/bus_reg_dataout[414] , 
        \DataPath/RF/bus_reg_dataout[413] , \DataPath/RF/bus_reg_dataout[412] , 
        \DataPath/RF/bus_reg_dataout[411] , \DataPath/RF/bus_reg_dataout[410] , 
        \DataPath/RF/bus_reg_dataout[409] , \DataPath/RF/bus_reg_dataout[408] , 
        \DataPath/RF/bus_reg_dataout[407] , \DataPath/RF/bus_reg_dataout[406] , 
        \DataPath/RF/bus_reg_dataout[405] , \DataPath/RF/bus_reg_dataout[404] , 
        \DataPath/RF/bus_reg_dataout[403] , \DataPath/RF/bus_reg_dataout[402] , 
        \DataPath/RF/bus_reg_dataout[401] , \DataPath/RF/bus_reg_dataout[400] , 
        \DataPath/RF/bus_reg_dataout[399] , \DataPath/RF/bus_reg_dataout[398] , 
        \DataPath/RF/bus_reg_dataout[397] , \DataPath/RF/bus_reg_dataout[396] , 
        \DataPath/RF/bus_reg_dataout[395] , \DataPath/RF/bus_reg_dataout[394] , 
        \DataPath/RF/bus_reg_dataout[393] , \DataPath/RF/bus_reg_dataout[392] , 
        \DataPath/RF/bus_reg_dataout[391] , \DataPath/RF/bus_reg_dataout[390] , 
        \DataPath/RF/bus_reg_dataout[389] , \DataPath/RF/bus_reg_dataout[388] , 
        \DataPath/RF/bus_reg_dataout[387] , \DataPath/RF/bus_reg_dataout[386] , 
        \DataPath/RF/bus_reg_dataout[385] , \DataPath/RF/bus_reg_dataout[384] , 
        \DataPath/RF/bus_reg_dataout[383] , \DataPath/RF/bus_reg_dataout[382] , 
        \DataPath/RF/bus_reg_dataout[381] , \DataPath/RF/bus_reg_dataout[380] , 
        \DataPath/RF/bus_reg_dataout[379] , \DataPath/RF/bus_reg_dataout[378] , 
        \DataPath/RF/bus_reg_dataout[377] , \DataPath/RF/bus_reg_dataout[376] , 
        \DataPath/RF/bus_reg_dataout[375] , \DataPath/RF/bus_reg_dataout[374] , 
        \DataPath/RF/bus_reg_dataout[373] , \DataPath/RF/bus_reg_dataout[372] , 
        \DataPath/RF/bus_reg_dataout[371] , \DataPath/RF/bus_reg_dataout[370] , 
        \DataPath/RF/bus_reg_dataout[369] , \DataPath/RF/bus_reg_dataout[368] , 
        \DataPath/RF/bus_reg_dataout[367] , \DataPath/RF/bus_reg_dataout[366] , 
        \DataPath/RF/bus_reg_dataout[365] , \DataPath/RF/bus_reg_dataout[364] , 
        \DataPath/RF/bus_reg_dataout[363] , \DataPath/RF/bus_reg_dataout[362] , 
        \DataPath/RF/bus_reg_dataout[361] , \DataPath/RF/bus_reg_dataout[360] , 
        \DataPath/RF/bus_reg_dataout[359] , \DataPath/RF/bus_reg_dataout[358] , 
        \DataPath/RF/bus_reg_dataout[357] , \DataPath/RF/bus_reg_dataout[356] , 
        \DataPath/RF/bus_reg_dataout[355] , \DataPath/RF/bus_reg_dataout[354] , 
        \DataPath/RF/bus_reg_dataout[353] , \DataPath/RF/bus_reg_dataout[352] , 
        \DataPath/RF/bus_reg_dataout[351] , \DataPath/RF/bus_reg_dataout[350] , 
        \DataPath/RF/bus_reg_dataout[349] , \DataPath/RF/bus_reg_dataout[348] , 
        \DataPath/RF/bus_reg_dataout[347] , \DataPath/RF/bus_reg_dataout[346] , 
        \DataPath/RF/bus_reg_dataout[345] , \DataPath/RF/bus_reg_dataout[344] , 
        \DataPath/RF/bus_reg_dataout[343] , \DataPath/RF/bus_reg_dataout[342] , 
        \DataPath/RF/bus_reg_dataout[341] , \DataPath/RF/bus_reg_dataout[340] , 
        \DataPath/RF/bus_reg_dataout[339] , \DataPath/RF/bus_reg_dataout[338] , 
        \DataPath/RF/bus_reg_dataout[337] , \DataPath/RF/bus_reg_dataout[336] , 
        \DataPath/RF/bus_reg_dataout[335] , \DataPath/RF/bus_reg_dataout[334] , 
        \DataPath/RF/bus_reg_dataout[333] , \DataPath/RF/bus_reg_dataout[332] , 
        \DataPath/RF/bus_reg_dataout[331] , \DataPath/RF/bus_reg_dataout[330] , 
        \DataPath/RF/bus_reg_dataout[329] , \DataPath/RF/bus_reg_dataout[328] , 
        \DataPath/RF/bus_reg_dataout[327] , \DataPath/RF/bus_reg_dataout[326] , 
        \DataPath/RF/bus_reg_dataout[325] , \DataPath/RF/bus_reg_dataout[324] , 
        \DataPath/RF/bus_reg_dataout[323] , \DataPath/RF/bus_reg_dataout[322] , 
        \DataPath/RF/bus_reg_dataout[321] , \DataPath/RF/bus_reg_dataout[320] , 
        \DataPath/RF/bus_reg_dataout[319] , \DataPath/RF/bus_reg_dataout[318] , 
        \DataPath/RF/bus_reg_dataout[317] , \DataPath/RF/bus_reg_dataout[316] , 
        \DataPath/RF/bus_reg_dataout[315] , \DataPath/RF/bus_reg_dataout[314] , 
        \DataPath/RF/bus_reg_dataout[313] , \DataPath/RF/bus_reg_dataout[312] , 
        \DataPath/RF/bus_reg_dataout[311] , \DataPath/RF/bus_reg_dataout[310] , 
        \DataPath/RF/bus_reg_dataout[309] , \DataPath/RF/bus_reg_dataout[308] , 
        \DataPath/RF/bus_reg_dataout[307] , \DataPath/RF/bus_reg_dataout[306] , 
        \DataPath/RF/bus_reg_dataout[305] , \DataPath/RF/bus_reg_dataout[304] , 
        \DataPath/RF/bus_reg_dataout[303] , \DataPath/RF/bus_reg_dataout[302] , 
        \DataPath/RF/bus_reg_dataout[301] , \DataPath/RF/bus_reg_dataout[300] , 
        \DataPath/RF/bus_reg_dataout[299] , \DataPath/RF/bus_reg_dataout[298] , 
        \DataPath/RF/bus_reg_dataout[297] , \DataPath/RF/bus_reg_dataout[296] , 
        \DataPath/RF/bus_reg_dataout[295] , \DataPath/RF/bus_reg_dataout[294] , 
        \DataPath/RF/bus_reg_dataout[293] , \DataPath/RF/bus_reg_dataout[292] , 
        \DataPath/RF/bus_reg_dataout[291] , \DataPath/RF/bus_reg_dataout[290] , 
        \DataPath/RF/bus_reg_dataout[289] , \DataPath/RF/bus_reg_dataout[288] , 
        \DataPath/RF/bus_reg_dataout[287] , \DataPath/RF/bus_reg_dataout[286] , 
        \DataPath/RF/bus_reg_dataout[285] , \DataPath/RF/bus_reg_dataout[284] , 
        \DataPath/RF/bus_reg_dataout[283] , \DataPath/RF/bus_reg_dataout[282] , 
        \DataPath/RF/bus_reg_dataout[281] , \DataPath/RF/bus_reg_dataout[280] , 
        \DataPath/RF/bus_reg_dataout[279] , \DataPath/RF/bus_reg_dataout[278] , 
        \DataPath/RF/bus_reg_dataout[277] , \DataPath/RF/bus_reg_dataout[276] , 
        \DataPath/RF/bus_reg_dataout[275] , \DataPath/RF/bus_reg_dataout[274] , 
        \DataPath/RF/bus_reg_dataout[273] , \DataPath/RF/bus_reg_dataout[272] , 
        \DataPath/RF/bus_reg_dataout[271] , \DataPath/RF/bus_reg_dataout[270] , 
        \DataPath/RF/bus_reg_dataout[269] , \DataPath/RF/bus_reg_dataout[268] , 
        \DataPath/RF/bus_reg_dataout[267] , \DataPath/RF/bus_reg_dataout[266] , 
        \DataPath/RF/bus_reg_dataout[265] , \DataPath/RF/bus_reg_dataout[264] , 
        \DataPath/RF/bus_reg_dataout[263] , \DataPath/RF/bus_reg_dataout[262] , 
        \DataPath/RF/bus_reg_dataout[261] , \DataPath/RF/bus_reg_dataout[260] , 
        \DataPath/RF/bus_reg_dataout[259] , \DataPath/RF/bus_reg_dataout[258] , 
        \DataPath/RF/bus_reg_dataout[257] , \DataPath/RF/bus_reg_dataout[256] , 
        \DataPath/RF/bus_reg_dataout[255] , \DataPath/RF/bus_reg_dataout[254] , 
        \DataPath/RF/bus_reg_dataout[253] , \DataPath/RF/bus_reg_dataout[252] , 
        \DataPath/RF/bus_reg_dataout[251] , \DataPath/RF/bus_reg_dataout[250] , 
        \DataPath/RF/bus_reg_dataout[249] , \DataPath/RF/bus_reg_dataout[248] , 
        \DataPath/RF/bus_reg_dataout[247] , \DataPath/RF/bus_reg_dataout[246] , 
        \DataPath/RF/bus_reg_dataout[245] , \DataPath/RF/bus_reg_dataout[244] , 
        \DataPath/RF/bus_reg_dataout[243] , \DataPath/RF/bus_reg_dataout[242] , 
        \DataPath/RF/bus_reg_dataout[241] , \DataPath/RF/bus_reg_dataout[240] , 
        \DataPath/RF/bus_reg_dataout[239] , \DataPath/RF/bus_reg_dataout[238] , 
        \DataPath/RF/bus_reg_dataout[237] , \DataPath/RF/bus_reg_dataout[236] , 
        \DataPath/RF/bus_reg_dataout[235] , \DataPath/RF/bus_reg_dataout[234] , 
        \DataPath/RF/bus_reg_dataout[233] , \DataPath/RF/bus_reg_dataout[232] , 
        \DataPath/RF/bus_reg_dataout[231] , \DataPath/RF/bus_reg_dataout[230] , 
        \DataPath/RF/bus_reg_dataout[229] , \DataPath/RF/bus_reg_dataout[228] , 
        \DataPath/RF/bus_reg_dataout[227] , \DataPath/RF/bus_reg_dataout[226] , 
        \DataPath/RF/bus_reg_dataout[225] , \DataPath/RF/bus_reg_dataout[224] , 
        \DataPath/RF/bus_reg_dataout[223] , \DataPath/RF/bus_reg_dataout[222] , 
        \DataPath/RF/bus_reg_dataout[221] , \DataPath/RF/bus_reg_dataout[220] , 
        \DataPath/RF/bus_reg_dataout[219] , \DataPath/RF/bus_reg_dataout[218] , 
        \DataPath/RF/bus_reg_dataout[217] , \DataPath/RF/bus_reg_dataout[216] , 
        \DataPath/RF/bus_reg_dataout[215] , \DataPath/RF/bus_reg_dataout[214] , 
        \DataPath/RF/bus_reg_dataout[213] , \DataPath/RF/bus_reg_dataout[212] , 
        \DataPath/RF/bus_reg_dataout[211] , \DataPath/RF/bus_reg_dataout[210] , 
        \DataPath/RF/bus_reg_dataout[209] , \DataPath/RF/bus_reg_dataout[208] , 
        \DataPath/RF/bus_reg_dataout[207] , \DataPath/RF/bus_reg_dataout[206] , 
        \DataPath/RF/bus_reg_dataout[205] , \DataPath/RF/bus_reg_dataout[204] , 
        \DataPath/RF/bus_reg_dataout[203] , \DataPath/RF/bus_reg_dataout[202] , 
        \DataPath/RF/bus_reg_dataout[201] , \DataPath/RF/bus_reg_dataout[200] , 
        \DataPath/RF/bus_reg_dataout[199] , \DataPath/RF/bus_reg_dataout[198] , 
        \DataPath/RF/bus_reg_dataout[197] , \DataPath/RF/bus_reg_dataout[196] , 
        \DataPath/RF/bus_reg_dataout[195] , \DataPath/RF/bus_reg_dataout[194] , 
        \DataPath/RF/bus_reg_dataout[193] , \DataPath/RF/bus_reg_dataout[192] , 
        \DataPath/RF/bus_reg_dataout[191] , \DataPath/RF/bus_reg_dataout[190] , 
        \DataPath/RF/bus_reg_dataout[189] , \DataPath/RF/bus_reg_dataout[188] , 
        \DataPath/RF/bus_reg_dataout[187] , \DataPath/RF/bus_reg_dataout[186] , 
        \DataPath/RF/bus_reg_dataout[185] , \DataPath/RF/bus_reg_dataout[184] , 
        \DataPath/RF/bus_reg_dataout[183] , \DataPath/RF/bus_reg_dataout[182] , 
        \DataPath/RF/bus_reg_dataout[181] , \DataPath/RF/bus_reg_dataout[180] , 
        \DataPath/RF/bus_reg_dataout[179] , \DataPath/RF/bus_reg_dataout[178] , 
        \DataPath/RF/bus_reg_dataout[177] , \DataPath/RF/bus_reg_dataout[176] , 
        \DataPath/RF/bus_reg_dataout[175] , \DataPath/RF/bus_reg_dataout[174] , 
        \DataPath/RF/bus_reg_dataout[173] , \DataPath/RF/bus_reg_dataout[172] , 
        \DataPath/RF/bus_reg_dataout[171] , \DataPath/RF/bus_reg_dataout[170] , 
        \DataPath/RF/bus_reg_dataout[169] , \DataPath/RF/bus_reg_dataout[168] , 
        \DataPath/RF/bus_reg_dataout[167] , \DataPath/RF/bus_reg_dataout[166] , 
        \DataPath/RF/bus_reg_dataout[165] , \DataPath/RF/bus_reg_dataout[164] , 
        \DataPath/RF/bus_reg_dataout[163] , \DataPath/RF/bus_reg_dataout[162] , 
        \DataPath/RF/bus_reg_dataout[161] , \DataPath/RF/bus_reg_dataout[160] , 
        \DataPath/RF/bus_reg_dataout[159] , \DataPath/RF/bus_reg_dataout[158] , 
        \DataPath/RF/bus_reg_dataout[157] , \DataPath/RF/bus_reg_dataout[156] , 
        \DataPath/RF/bus_reg_dataout[155] , \DataPath/RF/bus_reg_dataout[154] , 
        \DataPath/RF/bus_reg_dataout[153] , \DataPath/RF/bus_reg_dataout[152] , 
        \DataPath/RF/bus_reg_dataout[151] , \DataPath/RF/bus_reg_dataout[150] , 
        \DataPath/RF/bus_reg_dataout[149] , \DataPath/RF/bus_reg_dataout[148] , 
        \DataPath/RF/bus_reg_dataout[147] , \DataPath/RF/bus_reg_dataout[146] , 
        \DataPath/RF/bus_reg_dataout[145] , \DataPath/RF/bus_reg_dataout[144] , 
        \DataPath/RF/bus_reg_dataout[143] , \DataPath/RF/bus_reg_dataout[142] , 
        \DataPath/RF/bus_reg_dataout[141] , \DataPath/RF/bus_reg_dataout[140] , 
        \DataPath/RF/bus_reg_dataout[139] , \DataPath/RF/bus_reg_dataout[138] , 
        \DataPath/RF/bus_reg_dataout[137] , \DataPath/RF/bus_reg_dataout[136] , 
        \DataPath/RF/bus_reg_dataout[135] , \DataPath/RF/bus_reg_dataout[134] , 
        \DataPath/RF/bus_reg_dataout[133] , \DataPath/RF/bus_reg_dataout[132] , 
        \DataPath/RF/bus_reg_dataout[131] , \DataPath/RF/bus_reg_dataout[130] , 
        \DataPath/RF/bus_reg_dataout[129] , \DataPath/RF/bus_reg_dataout[128] , 
        \DataPath/RF/bus_reg_dataout[127] , \DataPath/RF/bus_reg_dataout[126] , 
        \DataPath/RF/bus_reg_dataout[125] , \DataPath/RF/bus_reg_dataout[124] , 
        \DataPath/RF/bus_reg_dataout[123] , \DataPath/RF/bus_reg_dataout[122] , 
        \DataPath/RF/bus_reg_dataout[121] , \DataPath/RF/bus_reg_dataout[120] , 
        \DataPath/RF/bus_reg_dataout[119] , \DataPath/RF/bus_reg_dataout[118] , 
        \DataPath/RF/bus_reg_dataout[117] , \DataPath/RF/bus_reg_dataout[116] , 
        \DataPath/RF/bus_reg_dataout[115] , \DataPath/RF/bus_reg_dataout[114] , 
        \DataPath/RF/bus_reg_dataout[113] , \DataPath/RF/bus_reg_dataout[112] , 
        \DataPath/RF/bus_reg_dataout[111] , \DataPath/RF/bus_reg_dataout[110] , 
        \DataPath/RF/bus_reg_dataout[109] , \DataPath/RF/bus_reg_dataout[108] , 
        \DataPath/RF/bus_reg_dataout[107] , \DataPath/RF/bus_reg_dataout[106] , 
        \DataPath/RF/bus_reg_dataout[105] , \DataPath/RF/bus_reg_dataout[104] , 
        \DataPath/RF/bus_reg_dataout[103] , \DataPath/RF/bus_reg_dataout[102] , 
        \DataPath/RF/bus_reg_dataout[101] , \DataPath/RF/bus_reg_dataout[100] , 
        \DataPath/RF/bus_reg_dataout[99] , \DataPath/RF/bus_reg_dataout[98] , 
        \DataPath/RF/bus_reg_dataout[97] , \DataPath/RF/bus_reg_dataout[96] , 
        \DataPath/RF/bus_reg_dataout[95] , \DataPath/RF/bus_reg_dataout[94] , 
        \DataPath/RF/bus_reg_dataout[93] , \DataPath/RF/bus_reg_dataout[92] , 
        \DataPath/RF/bus_reg_dataout[91] , \DataPath/RF/bus_reg_dataout[90] , 
        \DataPath/RF/bus_reg_dataout[89] , \DataPath/RF/bus_reg_dataout[88] , 
        \DataPath/RF/bus_reg_dataout[87] , \DataPath/RF/bus_reg_dataout[86] , 
        \DataPath/RF/bus_reg_dataout[85] , \DataPath/RF/bus_reg_dataout[84] , 
        \DataPath/RF/bus_reg_dataout[83] , \DataPath/RF/bus_reg_dataout[82] , 
        \DataPath/RF/bus_reg_dataout[81] , \DataPath/RF/bus_reg_dataout[80] , 
        \DataPath/RF/bus_reg_dataout[79] , \DataPath/RF/bus_reg_dataout[78] , 
        \DataPath/RF/bus_reg_dataout[77] , \DataPath/RF/bus_reg_dataout[76] , 
        \DataPath/RF/bus_reg_dataout[75] , \DataPath/RF/bus_reg_dataout[74] , 
        \DataPath/RF/bus_reg_dataout[73] , \DataPath/RF/bus_reg_dataout[72] , 
        \DataPath/RF/bus_reg_dataout[71] , \DataPath/RF/bus_reg_dataout[70] , 
        \DataPath/RF/bus_reg_dataout[69] , \DataPath/RF/bus_reg_dataout[68] , 
        \DataPath/RF/bus_reg_dataout[67] , \DataPath/RF/bus_reg_dataout[66] , 
        \DataPath/RF/bus_reg_dataout[65] , \DataPath/RF/bus_reg_dataout[64] , 
        \DataPath/RF/bus_reg_dataout[63] , \DataPath/RF/bus_reg_dataout[62] , 
        \DataPath/RF/bus_reg_dataout[61] , \DataPath/RF/bus_reg_dataout[60] , 
        \DataPath/RF/bus_reg_dataout[59] , \DataPath/RF/bus_reg_dataout[58] , 
        \DataPath/RF/bus_reg_dataout[57] , \DataPath/RF/bus_reg_dataout[56] , 
        \DataPath/RF/bus_reg_dataout[55] , \DataPath/RF/bus_reg_dataout[54] , 
        \DataPath/RF/bus_reg_dataout[53] , \DataPath/RF/bus_reg_dataout[52] , 
        \DataPath/RF/bus_reg_dataout[51] , \DataPath/RF/bus_reg_dataout[50] , 
        \DataPath/RF/bus_reg_dataout[49] , \DataPath/RF/bus_reg_dataout[48] , 
        \DataPath/RF/bus_reg_dataout[47] , \DataPath/RF/bus_reg_dataout[46] , 
        \DataPath/RF/bus_reg_dataout[45] , \DataPath/RF/bus_reg_dataout[44] , 
        \DataPath/RF/bus_reg_dataout[43] , \DataPath/RF/bus_reg_dataout[42] , 
        \DataPath/RF/bus_reg_dataout[41] , \DataPath/RF/bus_reg_dataout[40] , 
        \DataPath/RF/bus_reg_dataout[39] , \DataPath/RF/bus_reg_dataout[38] , 
        \DataPath/RF/bus_reg_dataout[37] , \DataPath/RF/bus_reg_dataout[36] , 
        \DataPath/RF/bus_reg_dataout[35] , \DataPath/RF/bus_reg_dataout[34] , 
        \DataPath/RF/bus_reg_dataout[33] , \DataPath/RF/bus_reg_dataout[32] , 
        \DataPath/RF/bus_reg_dataout[31] , \DataPath/RF/bus_reg_dataout[30] , 
        \DataPath/RF/bus_reg_dataout[29] , \DataPath/RF/bus_reg_dataout[28] , 
        \DataPath/RF/bus_reg_dataout[27] , \DataPath/RF/bus_reg_dataout[26] , 
        \DataPath/RF/bus_reg_dataout[25] , \DataPath/RF/bus_reg_dataout[24] , 
        \DataPath/RF/bus_reg_dataout[23] , \DataPath/RF/bus_reg_dataout[22] , 
        \DataPath/RF/bus_reg_dataout[21] , \DataPath/RF/bus_reg_dataout[20] , 
        \DataPath/RF/bus_reg_dataout[19] , \DataPath/RF/bus_reg_dataout[18] , 
        \DataPath/RF/bus_reg_dataout[17] , \DataPath/RF/bus_reg_dataout[16] , 
        \DataPath/RF/bus_reg_dataout[15] , \DataPath/RF/bus_reg_dataout[14] , 
        \DataPath/RF/bus_reg_dataout[13] , \DataPath/RF/bus_reg_dataout[12] , 
        \DataPath/RF/bus_reg_dataout[11] , \DataPath/RF/bus_reg_dataout[10] , 
        \DataPath/RF/bus_reg_dataout[9] , \DataPath/RF/bus_reg_dataout[8] , 
        \DataPath/RF/bus_reg_dataout[7] , \DataPath/RF/bus_reg_dataout[6] , 
        \DataPath/RF/bus_reg_dataout[5] , \DataPath/RF/bus_reg_dataout[4] , 
        \DataPath/RF/bus_reg_dataout[3] , \DataPath/RF/bus_reg_dataout[2] , 
        \DataPath/RF/bus_reg_dataout[1] , \DataPath/RF/bus_reg_dataout[0] }), 
        .win({n8281, \DataPath/RF/c_swin[3] , \DataPath/RF/c_swin[2] , 
        \DataPath/RF/c_swin[1] , \DataPath/RF/c_swin[0] }), .curr_proc_regs({
        \DataPath/RF/bus_sel_savedwin_data[511] , 
        \DataPath/RF/bus_sel_savedwin_data[510] , 
        \DataPath/RF/bus_sel_savedwin_data[509] , 
        \DataPath/RF/bus_sel_savedwin_data[508] , 
        \DataPath/RF/bus_sel_savedwin_data[507] , 
        \DataPath/RF/bus_sel_savedwin_data[506] , 
        \DataPath/RF/bus_sel_savedwin_data[505] , 
        \DataPath/RF/bus_sel_savedwin_data[504] , 
        \DataPath/RF/bus_sel_savedwin_data[503] , 
        \DataPath/RF/bus_sel_savedwin_data[502] , 
        \DataPath/RF/bus_sel_savedwin_data[501] , 
        \DataPath/RF/bus_sel_savedwin_data[500] , 
        \DataPath/RF/bus_sel_savedwin_data[499] , 
        \DataPath/RF/bus_sel_savedwin_data[498] , 
        \DataPath/RF/bus_sel_savedwin_data[497] , 
        \DataPath/RF/bus_sel_savedwin_data[496] , 
        \DataPath/RF/bus_sel_savedwin_data[495] , 
        \DataPath/RF/bus_sel_savedwin_data[494] , 
        \DataPath/RF/bus_sel_savedwin_data[493] , 
        \DataPath/RF/bus_sel_savedwin_data[492] , 
        \DataPath/RF/bus_sel_savedwin_data[491] , 
        \DataPath/RF/bus_sel_savedwin_data[490] , 
        \DataPath/RF/bus_sel_savedwin_data[489] , 
        \DataPath/RF/bus_sel_savedwin_data[488] , 
        \DataPath/RF/bus_sel_savedwin_data[487] , 
        \DataPath/RF/bus_sel_savedwin_data[486] , 
        \DataPath/RF/bus_sel_savedwin_data[485] , 
        \DataPath/RF/bus_sel_savedwin_data[484] , 
        \DataPath/RF/bus_sel_savedwin_data[483] , 
        \DataPath/RF/bus_sel_savedwin_data[482] , 
        \DataPath/RF/bus_sel_savedwin_data[481] , 
        \DataPath/RF/bus_sel_savedwin_data[480] , 
        \DataPath/RF/bus_sel_savedwin_data[479] , 
        \DataPath/RF/bus_sel_savedwin_data[478] , 
        \DataPath/RF/bus_sel_savedwin_data[477] , 
        \DataPath/RF/bus_sel_savedwin_data[476] , 
        \DataPath/RF/bus_sel_savedwin_data[475] , 
        \DataPath/RF/bus_sel_savedwin_data[474] , 
        \DataPath/RF/bus_sel_savedwin_data[473] , 
        \DataPath/RF/bus_sel_savedwin_data[472] , 
        \DataPath/RF/bus_sel_savedwin_data[471] , 
        \DataPath/RF/bus_sel_savedwin_data[470] , 
        \DataPath/RF/bus_sel_savedwin_data[469] , 
        \DataPath/RF/bus_sel_savedwin_data[468] , 
        \DataPath/RF/bus_sel_savedwin_data[467] , 
        \DataPath/RF/bus_sel_savedwin_data[466] , 
        \DataPath/RF/bus_sel_savedwin_data[465] , 
        \DataPath/RF/bus_sel_savedwin_data[464] , 
        \DataPath/RF/bus_sel_savedwin_data[463] , 
        \DataPath/RF/bus_sel_savedwin_data[462] , 
        \DataPath/RF/bus_sel_savedwin_data[461] , 
        \DataPath/RF/bus_sel_savedwin_data[460] , 
        \DataPath/RF/bus_sel_savedwin_data[459] , 
        \DataPath/RF/bus_sel_savedwin_data[458] , 
        \DataPath/RF/bus_sel_savedwin_data[457] , 
        \DataPath/RF/bus_sel_savedwin_data[456] , 
        \DataPath/RF/bus_sel_savedwin_data[455] , 
        \DataPath/RF/bus_sel_savedwin_data[454] , 
        \DataPath/RF/bus_sel_savedwin_data[453] , 
        \DataPath/RF/bus_sel_savedwin_data[452] , 
        \DataPath/RF/bus_sel_savedwin_data[451] , 
        \DataPath/RF/bus_sel_savedwin_data[450] , 
        \DataPath/RF/bus_sel_savedwin_data[449] , 
        \DataPath/RF/bus_sel_savedwin_data[448] , 
        \DataPath/RF/bus_sel_savedwin_data[447] , 
        \DataPath/RF/bus_sel_savedwin_data[446] , 
        \DataPath/RF/bus_sel_savedwin_data[445] , 
        \DataPath/RF/bus_sel_savedwin_data[444] , 
        \DataPath/RF/bus_sel_savedwin_data[443] , 
        \DataPath/RF/bus_sel_savedwin_data[442] , 
        \DataPath/RF/bus_sel_savedwin_data[441] , 
        \DataPath/RF/bus_sel_savedwin_data[440] , 
        \DataPath/RF/bus_sel_savedwin_data[439] , 
        \DataPath/RF/bus_sel_savedwin_data[438] , 
        \DataPath/RF/bus_sel_savedwin_data[437] , 
        \DataPath/RF/bus_sel_savedwin_data[436] , 
        \DataPath/RF/bus_sel_savedwin_data[435] , 
        \DataPath/RF/bus_sel_savedwin_data[434] , 
        \DataPath/RF/bus_sel_savedwin_data[433] , 
        \DataPath/RF/bus_sel_savedwin_data[432] , 
        \DataPath/RF/bus_sel_savedwin_data[431] , 
        \DataPath/RF/bus_sel_savedwin_data[430] , 
        \DataPath/RF/bus_sel_savedwin_data[429] , 
        \DataPath/RF/bus_sel_savedwin_data[428] , 
        \DataPath/RF/bus_sel_savedwin_data[427] , 
        \DataPath/RF/bus_sel_savedwin_data[426] , 
        \DataPath/RF/bus_sel_savedwin_data[425] , 
        \DataPath/RF/bus_sel_savedwin_data[424] , 
        \DataPath/RF/bus_sel_savedwin_data[423] , 
        \DataPath/RF/bus_sel_savedwin_data[422] , 
        \DataPath/RF/bus_sel_savedwin_data[421] , 
        \DataPath/RF/bus_sel_savedwin_data[420] , 
        \DataPath/RF/bus_sel_savedwin_data[419] , 
        \DataPath/RF/bus_sel_savedwin_data[418] , 
        \DataPath/RF/bus_sel_savedwin_data[417] , 
        \DataPath/RF/bus_sel_savedwin_data[416] , 
        \DataPath/RF/bus_sel_savedwin_data[415] , 
        \DataPath/RF/bus_sel_savedwin_data[414] , 
        \DataPath/RF/bus_sel_savedwin_data[413] , 
        \DataPath/RF/bus_sel_savedwin_data[412] , 
        \DataPath/RF/bus_sel_savedwin_data[411] , 
        \DataPath/RF/bus_sel_savedwin_data[410] , 
        \DataPath/RF/bus_sel_savedwin_data[409] , 
        \DataPath/RF/bus_sel_savedwin_data[408] , 
        \DataPath/RF/bus_sel_savedwin_data[407] , 
        \DataPath/RF/bus_sel_savedwin_data[406] , 
        \DataPath/RF/bus_sel_savedwin_data[405] , 
        \DataPath/RF/bus_sel_savedwin_data[404] , 
        \DataPath/RF/bus_sel_savedwin_data[403] , 
        \DataPath/RF/bus_sel_savedwin_data[402] , 
        \DataPath/RF/bus_sel_savedwin_data[401] , 
        \DataPath/RF/bus_sel_savedwin_data[400] , 
        \DataPath/RF/bus_sel_savedwin_data[399] , 
        \DataPath/RF/bus_sel_savedwin_data[398] , 
        \DataPath/RF/bus_sel_savedwin_data[397] , 
        \DataPath/RF/bus_sel_savedwin_data[396] , 
        \DataPath/RF/bus_sel_savedwin_data[395] , 
        \DataPath/RF/bus_sel_savedwin_data[394] , 
        \DataPath/RF/bus_sel_savedwin_data[393] , 
        \DataPath/RF/bus_sel_savedwin_data[392] , 
        \DataPath/RF/bus_sel_savedwin_data[391] , 
        \DataPath/RF/bus_sel_savedwin_data[390] , 
        \DataPath/RF/bus_sel_savedwin_data[389] , 
        \DataPath/RF/bus_sel_savedwin_data[388] , 
        \DataPath/RF/bus_sel_savedwin_data[387] , 
        \DataPath/RF/bus_sel_savedwin_data[386] , 
        \DataPath/RF/bus_sel_savedwin_data[385] , 
        \DataPath/RF/bus_sel_savedwin_data[384] , 
        \DataPath/RF/bus_sel_savedwin_data[383] , 
        \DataPath/RF/bus_sel_savedwin_data[382] , 
        \DataPath/RF/bus_sel_savedwin_data[381] , 
        \DataPath/RF/bus_sel_savedwin_data[380] , 
        \DataPath/RF/bus_sel_savedwin_data[379] , 
        \DataPath/RF/bus_sel_savedwin_data[378] , 
        \DataPath/RF/bus_sel_savedwin_data[377] , 
        \DataPath/RF/bus_sel_savedwin_data[376] , 
        \DataPath/RF/bus_sel_savedwin_data[375] , 
        \DataPath/RF/bus_sel_savedwin_data[374] , 
        \DataPath/RF/bus_sel_savedwin_data[373] , 
        \DataPath/RF/bus_sel_savedwin_data[372] , 
        \DataPath/RF/bus_sel_savedwin_data[371] , 
        \DataPath/RF/bus_sel_savedwin_data[370] , 
        \DataPath/RF/bus_sel_savedwin_data[369] , 
        \DataPath/RF/bus_sel_savedwin_data[368] , 
        \DataPath/RF/bus_sel_savedwin_data[367] , 
        \DataPath/RF/bus_sel_savedwin_data[366] , 
        \DataPath/RF/bus_sel_savedwin_data[365] , 
        \DataPath/RF/bus_sel_savedwin_data[364] , 
        \DataPath/RF/bus_sel_savedwin_data[363] , 
        \DataPath/RF/bus_sel_savedwin_data[362] , 
        \DataPath/RF/bus_sel_savedwin_data[361] , 
        \DataPath/RF/bus_sel_savedwin_data[360] , 
        \DataPath/RF/bus_sel_savedwin_data[359] , 
        \DataPath/RF/bus_sel_savedwin_data[358] , 
        \DataPath/RF/bus_sel_savedwin_data[357] , 
        \DataPath/RF/bus_sel_savedwin_data[356] , 
        \DataPath/RF/bus_sel_savedwin_data[355] , 
        \DataPath/RF/bus_sel_savedwin_data[354] , 
        \DataPath/RF/bus_sel_savedwin_data[353] , 
        \DataPath/RF/bus_sel_savedwin_data[352] , 
        \DataPath/RF/bus_sel_savedwin_data[351] , 
        \DataPath/RF/bus_sel_savedwin_data[350] , 
        \DataPath/RF/bus_sel_savedwin_data[349] , 
        \DataPath/RF/bus_sel_savedwin_data[348] , 
        \DataPath/RF/bus_sel_savedwin_data[347] , 
        \DataPath/RF/bus_sel_savedwin_data[346] , 
        \DataPath/RF/bus_sel_savedwin_data[345] , 
        \DataPath/RF/bus_sel_savedwin_data[344] , 
        \DataPath/RF/bus_sel_savedwin_data[343] , 
        \DataPath/RF/bus_sel_savedwin_data[342] , 
        \DataPath/RF/bus_sel_savedwin_data[341] , 
        \DataPath/RF/bus_sel_savedwin_data[340] , 
        \DataPath/RF/bus_sel_savedwin_data[339] , 
        \DataPath/RF/bus_sel_savedwin_data[338] , 
        \DataPath/RF/bus_sel_savedwin_data[337] , 
        \DataPath/RF/bus_sel_savedwin_data[336] , 
        \DataPath/RF/bus_sel_savedwin_data[335] , 
        \DataPath/RF/bus_sel_savedwin_data[334] , 
        \DataPath/RF/bus_sel_savedwin_data[333] , 
        \DataPath/RF/bus_sel_savedwin_data[332] , 
        \DataPath/RF/bus_sel_savedwin_data[331] , 
        \DataPath/RF/bus_sel_savedwin_data[330] , 
        \DataPath/RF/bus_sel_savedwin_data[329] , 
        \DataPath/RF/bus_sel_savedwin_data[328] , 
        \DataPath/RF/bus_sel_savedwin_data[327] , 
        \DataPath/RF/bus_sel_savedwin_data[326] , 
        \DataPath/RF/bus_sel_savedwin_data[325] , 
        \DataPath/RF/bus_sel_savedwin_data[324] , 
        \DataPath/RF/bus_sel_savedwin_data[323] , 
        \DataPath/RF/bus_sel_savedwin_data[322] , 
        \DataPath/RF/bus_sel_savedwin_data[321] , 
        \DataPath/RF/bus_sel_savedwin_data[320] , 
        \DataPath/RF/bus_sel_savedwin_data[319] , 
        \DataPath/RF/bus_sel_savedwin_data[318] , 
        \DataPath/RF/bus_sel_savedwin_data[317] , 
        \DataPath/RF/bus_sel_savedwin_data[316] , 
        \DataPath/RF/bus_sel_savedwin_data[315] , 
        \DataPath/RF/bus_sel_savedwin_data[314] , 
        \DataPath/RF/bus_sel_savedwin_data[313] , 
        \DataPath/RF/bus_sel_savedwin_data[312] , 
        \DataPath/RF/bus_sel_savedwin_data[311] , 
        \DataPath/RF/bus_sel_savedwin_data[310] , 
        \DataPath/RF/bus_sel_savedwin_data[309] , 
        \DataPath/RF/bus_sel_savedwin_data[308] , 
        \DataPath/RF/bus_sel_savedwin_data[307] , 
        \DataPath/RF/bus_sel_savedwin_data[306] , 
        \DataPath/RF/bus_sel_savedwin_data[305] , 
        \DataPath/RF/bus_sel_savedwin_data[304] , 
        \DataPath/RF/bus_sel_savedwin_data[303] , 
        \DataPath/RF/bus_sel_savedwin_data[302] , 
        \DataPath/RF/bus_sel_savedwin_data[301] , 
        \DataPath/RF/bus_sel_savedwin_data[300] , 
        \DataPath/RF/bus_sel_savedwin_data[299] , 
        \DataPath/RF/bus_sel_savedwin_data[298] , 
        \DataPath/RF/bus_sel_savedwin_data[297] , 
        \DataPath/RF/bus_sel_savedwin_data[296] , 
        \DataPath/RF/bus_sel_savedwin_data[295] , 
        \DataPath/RF/bus_sel_savedwin_data[294] , 
        \DataPath/RF/bus_sel_savedwin_data[293] , 
        \DataPath/RF/bus_sel_savedwin_data[292] , 
        \DataPath/RF/bus_sel_savedwin_data[291] , 
        \DataPath/RF/bus_sel_savedwin_data[290] , 
        \DataPath/RF/bus_sel_savedwin_data[289] , 
        \DataPath/RF/bus_sel_savedwin_data[288] , 
        \DataPath/RF/bus_sel_savedwin_data[287] , 
        \DataPath/RF/bus_sel_savedwin_data[286] , 
        \DataPath/RF/bus_sel_savedwin_data[285] , 
        \DataPath/RF/bus_sel_savedwin_data[284] , 
        \DataPath/RF/bus_sel_savedwin_data[283] , 
        \DataPath/RF/bus_sel_savedwin_data[282] , 
        \DataPath/RF/bus_sel_savedwin_data[281] , 
        \DataPath/RF/bus_sel_savedwin_data[280] , 
        \DataPath/RF/bus_sel_savedwin_data[279] , 
        \DataPath/RF/bus_sel_savedwin_data[278] , 
        \DataPath/RF/bus_sel_savedwin_data[277] , 
        \DataPath/RF/bus_sel_savedwin_data[276] , 
        \DataPath/RF/bus_sel_savedwin_data[275] , 
        \DataPath/RF/bus_sel_savedwin_data[274] , 
        \DataPath/RF/bus_sel_savedwin_data[273] , 
        \DataPath/RF/bus_sel_savedwin_data[272] , 
        \DataPath/RF/bus_sel_savedwin_data[271] , 
        \DataPath/RF/bus_sel_savedwin_data[270] , 
        \DataPath/RF/bus_sel_savedwin_data[269] , 
        \DataPath/RF/bus_sel_savedwin_data[268] , 
        \DataPath/RF/bus_sel_savedwin_data[267] , 
        \DataPath/RF/bus_sel_savedwin_data[266] , 
        \DataPath/RF/bus_sel_savedwin_data[265] , 
        \DataPath/RF/bus_sel_savedwin_data[264] , 
        \DataPath/RF/bus_sel_savedwin_data[263] , 
        \DataPath/RF/bus_sel_savedwin_data[262] , 
        \DataPath/RF/bus_sel_savedwin_data[261] , 
        \DataPath/RF/bus_sel_savedwin_data[260] , 
        \DataPath/RF/bus_sel_savedwin_data[259] , 
        \DataPath/RF/bus_sel_savedwin_data[258] , 
        \DataPath/RF/bus_sel_savedwin_data[257] , 
        \DataPath/RF/bus_sel_savedwin_data[256] , 
        \DataPath/RF/bus_sel_savedwin_data[255] , 
        \DataPath/RF/bus_sel_savedwin_data[254] , 
        \DataPath/RF/bus_sel_savedwin_data[253] , 
        \DataPath/RF/bus_sel_savedwin_data[252] , 
        \DataPath/RF/bus_sel_savedwin_data[251] , 
        \DataPath/RF/bus_sel_savedwin_data[250] , 
        \DataPath/RF/bus_sel_savedwin_data[249] , 
        \DataPath/RF/bus_sel_savedwin_data[248] , 
        \DataPath/RF/bus_sel_savedwin_data[247] , 
        \DataPath/RF/bus_sel_savedwin_data[246] , 
        \DataPath/RF/bus_sel_savedwin_data[245] , 
        \DataPath/RF/bus_sel_savedwin_data[244] , 
        \DataPath/RF/bus_sel_savedwin_data[243] , 
        \DataPath/RF/bus_sel_savedwin_data[242] , 
        \DataPath/RF/bus_sel_savedwin_data[241] , 
        \DataPath/RF/bus_sel_savedwin_data[240] , 
        \DataPath/RF/bus_sel_savedwin_data[239] , 
        \DataPath/RF/bus_sel_savedwin_data[238] , 
        \DataPath/RF/bus_sel_savedwin_data[237] , 
        \DataPath/RF/bus_sel_savedwin_data[236] , 
        \DataPath/RF/bus_sel_savedwin_data[235] , 
        \DataPath/RF/bus_sel_savedwin_data[234] , 
        \DataPath/RF/bus_sel_savedwin_data[233] , 
        \DataPath/RF/bus_sel_savedwin_data[232] , 
        \DataPath/RF/bus_sel_savedwin_data[231] , 
        \DataPath/RF/bus_sel_savedwin_data[230] , 
        \DataPath/RF/bus_sel_savedwin_data[229] , 
        \DataPath/RF/bus_sel_savedwin_data[228] , 
        \DataPath/RF/bus_sel_savedwin_data[227] , 
        \DataPath/RF/bus_sel_savedwin_data[226] , 
        \DataPath/RF/bus_sel_savedwin_data[225] , 
        \DataPath/RF/bus_sel_savedwin_data[224] , 
        \DataPath/RF/bus_sel_savedwin_data[223] , 
        \DataPath/RF/bus_sel_savedwin_data[222] , 
        \DataPath/RF/bus_sel_savedwin_data[221] , 
        \DataPath/RF/bus_sel_savedwin_data[220] , 
        \DataPath/RF/bus_sel_savedwin_data[219] , 
        \DataPath/RF/bus_sel_savedwin_data[218] , 
        \DataPath/RF/bus_sel_savedwin_data[217] , 
        \DataPath/RF/bus_sel_savedwin_data[216] , 
        \DataPath/RF/bus_sel_savedwin_data[215] , 
        \DataPath/RF/bus_sel_savedwin_data[214] , 
        \DataPath/RF/bus_sel_savedwin_data[213] , 
        \DataPath/RF/bus_sel_savedwin_data[212] , 
        \DataPath/RF/bus_sel_savedwin_data[211] , 
        \DataPath/RF/bus_sel_savedwin_data[210] , 
        \DataPath/RF/bus_sel_savedwin_data[209] , 
        \DataPath/RF/bus_sel_savedwin_data[208] , 
        \DataPath/RF/bus_sel_savedwin_data[207] , 
        \DataPath/RF/bus_sel_savedwin_data[206] , 
        \DataPath/RF/bus_sel_savedwin_data[205] , 
        \DataPath/RF/bus_sel_savedwin_data[204] , 
        \DataPath/RF/bus_sel_savedwin_data[203] , 
        \DataPath/RF/bus_sel_savedwin_data[202] , 
        \DataPath/RF/bus_sel_savedwin_data[201] , 
        \DataPath/RF/bus_sel_savedwin_data[200] , 
        \DataPath/RF/bus_sel_savedwin_data[199] , 
        \DataPath/RF/bus_sel_savedwin_data[198] , 
        \DataPath/RF/bus_sel_savedwin_data[197] , 
        \DataPath/RF/bus_sel_savedwin_data[196] , 
        \DataPath/RF/bus_sel_savedwin_data[195] , 
        \DataPath/RF/bus_sel_savedwin_data[194] , 
        \DataPath/RF/bus_sel_savedwin_data[193] , 
        \DataPath/RF/bus_sel_savedwin_data[192] , 
        \DataPath/RF/bus_sel_savedwin_data[191] , 
        \DataPath/RF/bus_sel_savedwin_data[190] , 
        \DataPath/RF/bus_sel_savedwin_data[189] , 
        \DataPath/RF/bus_sel_savedwin_data[188] , 
        \DataPath/RF/bus_sel_savedwin_data[187] , 
        \DataPath/RF/bus_sel_savedwin_data[186] , 
        \DataPath/RF/bus_sel_savedwin_data[185] , 
        \DataPath/RF/bus_sel_savedwin_data[184] , 
        \DataPath/RF/bus_sel_savedwin_data[183] , 
        \DataPath/RF/bus_sel_savedwin_data[182] , 
        \DataPath/RF/bus_sel_savedwin_data[181] , 
        \DataPath/RF/bus_sel_savedwin_data[180] , 
        \DataPath/RF/bus_sel_savedwin_data[179] , 
        \DataPath/RF/bus_sel_savedwin_data[178] , 
        \DataPath/RF/bus_sel_savedwin_data[177] , 
        \DataPath/RF/bus_sel_savedwin_data[176] , 
        \DataPath/RF/bus_sel_savedwin_data[175] , 
        \DataPath/RF/bus_sel_savedwin_data[174] , 
        \DataPath/RF/bus_sel_savedwin_data[173] , 
        \DataPath/RF/bus_sel_savedwin_data[172] , 
        \DataPath/RF/bus_sel_savedwin_data[171] , 
        \DataPath/RF/bus_sel_savedwin_data[170] , 
        \DataPath/RF/bus_sel_savedwin_data[169] , 
        \DataPath/RF/bus_sel_savedwin_data[168] , 
        \DataPath/RF/bus_sel_savedwin_data[167] , 
        \DataPath/RF/bus_sel_savedwin_data[166] , 
        \DataPath/RF/bus_sel_savedwin_data[165] , 
        \DataPath/RF/bus_sel_savedwin_data[164] , 
        \DataPath/RF/bus_sel_savedwin_data[163] , 
        \DataPath/RF/bus_sel_savedwin_data[162] , 
        \DataPath/RF/bus_sel_savedwin_data[161] , 
        \DataPath/RF/bus_sel_savedwin_data[160] , 
        \DataPath/RF/bus_sel_savedwin_data[159] , 
        \DataPath/RF/bus_sel_savedwin_data[158] , 
        \DataPath/RF/bus_sel_savedwin_data[157] , 
        \DataPath/RF/bus_sel_savedwin_data[156] , 
        \DataPath/RF/bus_sel_savedwin_data[155] , 
        \DataPath/RF/bus_sel_savedwin_data[154] , 
        \DataPath/RF/bus_sel_savedwin_data[153] , 
        \DataPath/RF/bus_sel_savedwin_data[152] , 
        \DataPath/RF/bus_sel_savedwin_data[151] , 
        \DataPath/RF/bus_sel_savedwin_data[150] , 
        \DataPath/RF/bus_sel_savedwin_data[149] , 
        \DataPath/RF/bus_sel_savedwin_data[148] , 
        \DataPath/RF/bus_sel_savedwin_data[147] , 
        \DataPath/RF/bus_sel_savedwin_data[146] , 
        \DataPath/RF/bus_sel_savedwin_data[145] , 
        \DataPath/RF/bus_sel_savedwin_data[144] , 
        \DataPath/RF/bus_sel_savedwin_data[143] , 
        \DataPath/RF/bus_sel_savedwin_data[142] , 
        \DataPath/RF/bus_sel_savedwin_data[141] , 
        \DataPath/RF/bus_sel_savedwin_data[140] , 
        \DataPath/RF/bus_sel_savedwin_data[139] , 
        \DataPath/RF/bus_sel_savedwin_data[138] , 
        \DataPath/RF/bus_sel_savedwin_data[137] , 
        \DataPath/RF/bus_sel_savedwin_data[136] , 
        \DataPath/RF/bus_sel_savedwin_data[135] , 
        \DataPath/RF/bus_sel_savedwin_data[134] , 
        \DataPath/RF/bus_sel_savedwin_data[133] , 
        \DataPath/RF/bus_sel_savedwin_data[132] , 
        \DataPath/RF/bus_sel_savedwin_data[131] , 
        \DataPath/RF/bus_sel_savedwin_data[130] , 
        \DataPath/RF/bus_sel_savedwin_data[129] , 
        \DataPath/RF/bus_sel_savedwin_data[128] , 
        \DataPath/RF/bus_sel_savedwin_data[127] , 
        \DataPath/RF/bus_sel_savedwin_data[126] , 
        \DataPath/RF/bus_sel_savedwin_data[125] , 
        \DataPath/RF/bus_sel_savedwin_data[124] , 
        \DataPath/RF/bus_sel_savedwin_data[123] , 
        \DataPath/RF/bus_sel_savedwin_data[122] , 
        \DataPath/RF/bus_sel_savedwin_data[121] , 
        \DataPath/RF/bus_sel_savedwin_data[120] , 
        \DataPath/RF/bus_sel_savedwin_data[119] , 
        \DataPath/RF/bus_sel_savedwin_data[118] , 
        \DataPath/RF/bus_sel_savedwin_data[117] , 
        \DataPath/RF/bus_sel_savedwin_data[116] , 
        \DataPath/RF/bus_sel_savedwin_data[115] , 
        \DataPath/RF/bus_sel_savedwin_data[114] , 
        \DataPath/RF/bus_sel_savedwin_data[113] , 
        \DataPath/RF/bus_sel_savedwin_data[112] , 
        \DataPath/RF/bus_sel_savedwin_data[111] , 
        \DataPath/RF/bus_sel_savedwin_data[110] , 
        \DataPath/RF/bus_sel_savedwin_data[109] , 
        \DataPath/RF/bus_sel_savedwin_data[108] , 
        \DataPath/RF/bus_sel_savedwin_data[107] , 
        \DataPath/RF/bus_sel_savedwin_data[106] , 
        \DataPath/RF/bus_sel_savedwin_data[105] , 
        \DataPath/RF/bus_sel_savedwin_data[104] , 
        \DataPath/RF/bus_sel_savedwin_data[103] , 
        \DataPath/RF/bus_sel_savedwin_data[102] , 
        \DataPath/RF/bus_sel_savedwin_data[101] , 
        \DataPath/RF/bus_sel_savedwin_data[100] , 
        \DataPath/RF/bus_sel_savedwin_data[99] , 
        \DataPath/RF/bus_sel_savedwin_data[98] , 
        \DataPath/RF/bus_sel_savedwin_data[97] , 
        \DataPath/RF/bus_sel_savedwin_data[96] , 
        \DataPath/RF/bus_sel_savedwin_data[95] , 
        \DataPath/RF/bus_sel_savedwin_data[94] , 
        \DataPath/RF/bus_sel_savedwin_data[93] , 
        \DataPath/RF/bus_sel_savedwin_data[92] , 
        \DataPath/RF/bus_sel_savedwin_data[91] , 
        \DataPath/RF/bus_sel_savedwin_data[90] , 
        \DataPath/RF/bus_sel_savedwin_data[89] , 
        \DataPath/RF/bus_sel_savedwin_data[88] , 
        \DataPath/RF/bus_sel_savedwin_data[87] , 
        \DataPath/RF/bus_sel_savedwin_data[86] , 
        \DataPath/RF/bus_sel_savedwin_data[85] , 
        \DataPath/RF/bus_sel_savedwin_data[84] , 
        \DataPath/RF/bus_sel_savedwin_data[83] , 
        \DataPath/RF/bus_sel_savedwin_data[82] , 
        \DataPath/RF/bus_sel_savedwin_data[81] , 
        \DataPath/RF/bus_sel_savedwin_data[80] , 
        \DataPath/RF/bus_sel_savedwin_data[79] , 
        \DataPath/RF/bus_sel_savedwin_data[78] , 
        \DataPath/RF/bus_sel_savedwin_data[77] , 
        \DataPath/RF/bus_sel_savedwin_data[76] , 
        \DataPath/RF/bus_sel_savedwin_data[75] , 
        \DataPath/RF/bus_sel_savedwin_data[74] , 
        \DataPath/RF/bus_sel_savedwin_data[73] , 
        \DataPath/RF/bus_sel_savedwin_data[72] , 
        \DataPath/RF/bus_sel_savedwin_data[71] , 
        \DataPath/RF/bus_sel_savedwin_data[70] , 
        \DataPath/RF/bus_sel_savedwin_data[69] , 
        \DataPath/RF/bus_sel_savedwin_data[68] , 
        \DataPath/RF/bus_sel_savedwin_data[67] , 
        \DataPath/RF/bus_sel_savedwin_data[66] , 
        \DataPath/RF/bus_sel_savedwin_data[65] , 
        \DataPath/RF/bus_sel_savedwin_data[64] , 
        \DataPath/RF/bus_sel_savedwin_data[63] , 
        \DataPath/RF/bus_sel_savedwin_data[62] , 
        \DataPath/RF/bus_sel_savedwin_data[61] , 
        \DataPath/RF/bus_sel_savedwin_data[60] , 
        \DataPath/RF/bus_sel_savedwin_data[59] , 
        \DataPath/RF/bus_sel_savedwin_data[58] , 
        \DataPath/RF/bus_sel_savedwin_data[57] , 
        \DataPath/RF/bus_sel_savedwin_data[56] , 
        \DataPath/RF/bus_sel_savedwin_data[55] , 
        \DataPath/RF/bus_sel_savedwin_data[54] , 
        \DataPath/RF/bus_sel_savedwin_data[53] , 
        \DataPath/RF/bus_sel_savedwin_data[52] , 
        \DataPath/RF/bus_sel_savedwin_data[51] , 
        \DataPath/RF/bus_sel_savedwin_data[50] , 
        \DataPath/RF/bus_sel_savedwin_data[49] , 
        \DataPath/RF/bus_sel_savedwin_data[48] , 
        \DataPath/RF/bus_sel_savedwin_data[47] , 
        \DataPath/RF/bus_sel_savedwin_data[46] , 
        \DataPath/RF/bus_sel_savedwin_data[45] , 
        \DataPath/RF/bus_sel_savedwin_data[44] , 
        \DataPath/RF/bus_sel_savedwin_data[43] , 
        \DataPath/RF/bus_sel_savedwin_data[42] , 
        \DataPath/RF/bus_sel_savedwin_data[41] , 
        \DataPath/RF/bus_sel_savedwin_data[40] , 
        \DataPath/RF/bus_sel_savedwin_data[39] , 
        \DataPath/RF/bus_sel_savedwin_data[38] , 
        \DataPath/RF/bus_sel_savedwin_data[37] , 
        \DataPath/RF/bus_sel_savedwin_data[36] , 
        \DataPath/RF/bus_sel_savedwin_data[35] , 
        \DataPath/RF/bus_sel_savedwin_data[34] , 
        \DataPath/RF/bus_sel_savedwin_data[33] , 
        \DataPath/RF/bus_sel_savedwin_data[32] , 
        \DataPath/RF/bus_sel_savedwin_data[31] , 
        \DataPath/RF/bus_sel_savedwin_data[30] , 
        \DataPath/RF/bus_sel_savedwin_data[29] , 
        \DataPath/RF/bus_sel_savedwin_data[28] , 
        \DataPath/RF/bus_sel_savedwin_data[27] , 
        \DataPath/RF/bus_sel_savedwin_data[26] , 
        \DataPath/RF/bus_sel_savedwin_data[25] , 
        \DataPath/RF/bus_sel_savedwin_data[24] , 
        \DataPath/RF/bus_sel_savedwin_data[23] , 
        \DataPath/RF/bus_sel_savedwin_data[22] , 
        \DataPath/RF/bus_sel_savedwin_data[21] , 
        \DataPath/RF/bus_sel_savedwin_data[20] , 
        \DataPath/RF/bus_sel_savedwin_data[19] , 
        \DataPath/RF/bus_sel_savedwin_data[18] , 
        \DataPath/RF/bus_sel_savedwin_data[17] , 
        \DataPath/RF/bus_sel_savedwin_data[16] , 
        \DataPath/RF/bus_sel_savedwin_data[15] , 
        \DataPath/RF/bus_sel_savedwin_data[14] , 
        \DataPath/RF/bus_sel_savedwin_data[13] , 
        \DataPath/RF/bus_sel_savedwin_data[12] , 
        \DataPath/RF/bus_sel_savedwin_data[11] , 
        \DataPath/RF/bus_sel_savedwin_data[10] , 
        \DataPath/RF/bus_sel_savedwin_data[9] , 
        \DataPath/RF/bus_sel_savedwin_data[8] , 
        \DataPath/RF/bus_sel_savedwin_data[7] , 
        \DataPath/RF/bus_sel_savedwin_data[6] , 
        \DataPath/RF/bus_sel_savedwin_data[5] , 
        \DataPath/RF/bus_sel_savedwin_data[4] , 
        \DataPath/RF/bus_sel_savedwin_data[3] , 
        \DataPath/RF/bus_sel_savedwin_data[2] , 
        \DataPath/RF/bus_sel_savedwin_data[1] , 
        \DataPath/RF/bus_sel_savedwin_data[0] }) );
  mux_N32_M5_1 \DataPath/RF/RDPORT1  ( .S(i_ADD_RS2), .Q({
        \DataPath/RF/bus_selected_win_data[767] , 
        \DataPath/RF/bus_selected_win_data[766] , 
        \DataPath/RF/bus_selected_win_data[765] , 
        \DataPath/RF/bus_selected_win_data[764] , 
        \DataPath/RF/bus_selected_win_data[763] , 
        \DataPath/RF/bus_selected_win_data[762] , 
        \DataPath/RF/bus_selected_win_data[761] , 
        \DataPath/RF/bus_selected_win_data[760] , 
        \DataPath/RF/bus_selected_win_data[759] , 
        \DataPath/RF/bus_selected_win_data[758] , 
        \DataPath/RF/bus_selected_win_data[757] , 
        \DataPath/RF/bus_selected_win_data[756] , 
        \DataPath/RF/bus_selected_win_data[755] , 
        \DataPath/RF/bus_selected_win_data[754] , 
        \DataPath/RF/bus_selected_win_data[753] , 
        \DataPath/RF/bus_selected_win_data[752] , 
        \DataPath/RF/bus_selected_win_data[751] , 
        \DataPath/RF/bus_selected_win_data[750] , 
        \DataPath/RF/bus_selected_win_data[749] , 
        \DataPath/RF/bus_selected_win_data[748] , 
        \DataPath/RF/bus_selected_win_data[747] , 
        \DataPath/RF/bus_selected_win_data[746] , 
        \DataPath/RF/bus_selected_win_data[745] , 
        \DataPath/RF/bus_selected_win_data[744] , 
        \DataPath/RF/bus_selected_win_data[743] , 
        \DataPath/RF/bus_selected_win_data[742] , 
        \DataPath/RF/bus_selected_win_data[741] , 
        \DataPath/RF/bus_selected_win_data[740] , 
        \DataPath/RF/bus_selected_win_data[739] , 
        \DataPath/RF/bus_selected_win_data[738] , 
        \DataPath/RF/bus_selected_win_data[737] , 
        \DataPath/RF/bus_selected_win_data[736] , 
        \DataPath/RF/bus_selected_win_data[735] , 
        \DataPath/RF/bus_selected_win_data[734] , 
        \DataPath/RF/bus_selected_win_data[733] , 
        \DataPath/RF/bus_selected_win_data[732] , 
        \DataPath/RF/bus_selected_win_data[731] , 
        \DataPath/RF/bus_selected_win_data[730] , 
        \DataPath/RF/bus_selected_win_data[729] , 
        \DataPath/RF/bus_selected_win_data[728] , 
        \DataPath/RF/bus_selected_win_data[727] , 
        \DataPath/RF/bus_selected_win_data[726] , 
        \DataPath/RF/bus_selected_win_data[725] , 
        \DataPath/RF/bus_selected_win_data[724] , 
        \DataPath/RF/bus_selected_win_data[723] , 
        \DataPath/RF/bus_selected_win_data[722] , 
        \DataPath/RF/bus_selected_win_data[721] , 
        \DataPath/RF/bus_selected_win_data[720] , 
        \DataPath/RF/bus_selected_win_data[719] , 
        \DataPath/RF/bus_selected_win_data[718] , 
        \DataPath/RF/bus_selected_win_data[717] , 
        \DataPath/RF/bus_selected_win_data[716] , 
        \DataPath/RF/bus_selected_win_data[715] , 
        \DataPath/RF/bus_selected_win_data[714] , 
        \DataPath/RF/bus_selected_win_data[713] , 
        \DataPath/RF/bus_selected_win_data[712] , 
        \DataPath/RF/bus_selected_win_data[711] , 
        \DataPath/RF/bus_selected_win_data[710] , 
        \DataPath/RF/bus_selected_win_data[709] , 
        \DataPath/RF/bus_selected_win_data[708] , 
        \DataPath/RF/bus_selected_win_data[707] , 
        \DataPath/RF/bus_selected_win_data[706] , 
        \DataPath/RF/bus_selected_win_data[705] , 
        \DataPath/RF/bus_selected_win_data[704] , 
        \DataPath/RF/bus_selected_win_data[703] , 
        \DataPath/RF/bus_selected_win_data[702] , 
        \DataPath/RF/bus_selected_win_data[701] , 
        \DataPath/RF/bus_selected_win_data[700] , 
        \DataPath/RF/bus_selected_win_data[699] , 
        \DataPath/RF/bus_selected_win_data[698] , 
        \DataPath/RF/bus_selected_win_data[697] , 
        \DataPath/RF/bus_selected_win_data[696] , 
        \DataPath/RF/bus_selected_win_data[695] , 
        \DataPath/RF/bus_selected_win_data[694] , 
        \DataPath/RF/bus_selected_win_data[693] , 
        \DataPath/RF/bus_selected_win_data[692] , 
        \DataPath/RF/bus_selected_win_data[691] , 
        \DataPath/RF/bus_selected_win_data[690] , 
        \DataPath/RF/bus_selected_win_data[689] , 
        \DataPath/RF/bus_selected_win_data[688] , 
        \DataPath/RF/bus_selected_win_data[687] , 
        \DataPath/RF/bus_selected_win_data[686] , 
        \DataPath/RF/bus_selected_win_data[685] , 
        \DataPath/RF/bus_selected_win_data[684] , 
        \DataPath/RF/bus_selected_win_data[683] , 
        \DataPath/RF/bus_selected_win_data[682] , 
        \DataPath/RF/bus_selected_win_data[681] , 
        \DataPath/RF/bus_selected_win_data[680] , 
        \DataPath/RF/bus_selected_win_data[679] , 
        \DataPath/RF/bus_selected_win_data[678] , 
        \DataPath/RF/bus_selected_win_data[677] , 
        \DataPath/RF/bus_selected_win_data[676] , 
        \DataPath/RF/bus_selected_win_data[675] , 
        \DataPath/RF/bus_selected_win_data[674] , 
        \DataPath/RF/bus_selected_win_data[673] , 
        \DataPath/RF/bus_selected_win_data[672] , 
        \DataPath/RF/bus_selected_win_data[671] , 
        \DataPath/RF/bus_selected_win_data[670] , 
        \DataPath/RF/bus_selected_win_data[669] , 
        \DataPath/RF/bus_selected_win_data[668] , 
        \DataPath/RF/bus_selected_win_data[667] , 
        \DataPath/RF/bus_selected_win_data[666] , 
        \DataPath/RF/bus_selected_win_data[665] , 
        \DataPath/RF/bus_selected_win_data[664] , 
        \DataPath/RF/bus_selected_win_data[663] , 
        \DataPath/RF/bus_selected_win_data[662] , 
        \DataPath/RF/bus_selected_win_data[661] , 
        \DataPath/RF/bus_selected_win_data[660] , 
        \DataPath/RF/bus_selected_win_data[659] , 
        \DataPath/RF/bus_selected_win_data[658] , 
        \DataPath/RF/bus_selected_win_data[657] , 
        \DataPath/RF/bus_selected_win_data[656] , 
        \DataPath/RF/bus_selected_win_data[655] , 
        \DataPath/RF/bus_selected_win_data[654] , 
        \DataPath/RF/bus_selected_win_data[653] , 
        \DataPath/RF/bus_selected_win_data[652] , 
        \DataPath/RF/bus_selected_win_data[651] , 
        \DataPath/RF/bus_selected_win_data[650] , 
        \DataPath/RF/bus_selected_win_data[649] , 
        \DataPath/RF/bus_selected_win_data[648] , 
        \DataPath/RF/bus_selected_win_data[647] , 
        \DataPath/RF/bus_selected_win_data[646] , 
        \DataPath/RF/bus_selected_win_data[645] , 
        \DataPath/RF/bus_selected_win_data[644] , 
        \DataPath/RF/bus_selected_win_data[643] , 
        \DataPath/RF/bus_selected_win_data[642] , 
        \DataPath/RF/bus_selected_win_data[641] , 
        \DataPath/RF/bus_selected_win_data[640] , 
        \DataPath/RF/bus_selected_win_data[639] , 
        \DataPath/RF/bus_selected_win_data[638] , 
        \DataPath/RF/bus_selected_win_data[637] , 
        \DataPath/RF/bus_selected_win_data[636] , 
        \DataPath/RF/bus_selected_win_data[635] , 
        \DataPath/RF/bus_selected_win_data[634] , 
        \DataPath/RF/bus_selected_win_data[633] , 
        \DataPath/RF/bus_selected_win_data[632] , 
        \DataPath/RF/bus_selected_win_data[631] , 
        \DataPath/RF/bus_selected_win_data[630] , 
        \DataPath/RF/bus_selected_win_data[629] , 
        \DataPath/RF/bus_selected_win_data[628] , 
        \DataPath/RF/bus_selected_win_data[627] , 
        \DataPath/RF/bus_selected_win_data[626] , 
        \DataPath/RF/bus_selected_win_data[625] , 
        \DataPath/RF/bus_selected_win_data[624] , 
        \DataPath/RF/bus_selected_win_data[623] , 
        \DataPath/RF/bus_selected_win_data[622] , 
        \DataPath/RF/bus_selected_win_data[621] , 
        \DataPath/RF/bus_selected_win_data[620] , 
        \DataPath/RF/bus_selected_win_data[619] , 
        \DataPath/RF/bus_selected_win_data[618] , 
        \DataPath/RF/bus_selected_win_data[617] , 
        \DataPath/RF/bus_selected_win_data[616] , 
        \DataPath/RF/bus_selected_win_data[615] , 
        \DataPath/RF/bus_selected_win_data[614] , 
        \DataPath/RF/bus_selected_win_data[613] , 
        \DataPath/RF/bus_selected_win_data[612] , 
        \DataPath/RF/bus_selected_win_data[611] , 
        \DataPath/RF/bus_selected_win_data[610] , 
        \DataPath/RF/bus_selected_win_data[609] , 
        \DataPath/RF/bus_selected_win_data[608] , 
        \DataPath/RF/bus_selected_win_data[607] , 
        \DataPath/RF/bus_selected_win_data[606] , 
        \DataPath/RF/bus_selected_win_data[605] , 
        \DataPath/RF/bus_selected_win_data[604] , 
        \DataPath/RF/bus_selected_win_data[603] , 
        \DataPath/RF/bus_selected_win_data[602] , 
        \DataPath/RF/bus_selected_win_data[601] , 
        \DataPath/RF/bus_selected_win_data[600] , 
        \DataPath/RF/bus_selected_win_data[599] , 
        \DataPath/RF/bus_selected_win_data[598] , 
        \DataPath/RF/bus_selected_win_data[597] , 
        \DataPath/RF/bus_selected_win_data[596] , 
        \DataPath/RF/bus_selected_win_data[595] , 
        \DataPath/RF/bus_selected_win_data[594] , 
        \DataPath/RF/bus_selected_win_data[593] , 
        \DataPath/RF/bus_selected_win_data[592] , 
        \DataPath/RF/bus_selected_win_data[591] , 
        \DataPath/RF/bus_selected_win_data[590] , 
        \DataPath/RF/bus_selected_win_data[589] , 
        \DataPath/RF/bus_selected_win_data[588] , 
        \DataPath/RF/bus_selected_win_data[587] , 
        \DataPath/RF/bus_selected_win_data[586] , 
        \DataPath/RF/bus_selected_win_data[585] , 
        \DataPath/RF/bus_selected_win_data[584] , 
        \DataPath/RF/bus_selected_win_data[583] , 
        \DataPath/RF/bus_selected_win_data[582] , 
        \DataPath/RF/bus_selected_win_data[581] , 
        \DataPath/RF/bus_selected_win_data[580] , 
        \DataPath/RF/bus_selected_win_data[579] , 
        \DataPath/RF/bus_selected_win_data[578] , 
        \DataPath/RF/bus_selected_win_data[577] , 
        \DataPath/RF/bus_selected_win_data[576] , 
        \DataPath/RF/bus_selected_win_data[575] , 
        \DataPath/RF/bus_selected_win_data[574] , 
        \DataPath/RF/bus_selected_win_data[573] , 
        \DataPath/RF/bus_selected_win_data[572] , 
        \DataPath/RF/bus_selected_win_data[571] , 
        \DataPath/RF/bus_selected_win_data[570] , 
        \DataPath/RF/bus_selected_win_data[569] , 
        \DataPath/RF/bus_selected_win_data[568] , 
        \DataPath/RF/bus_selected_win_data[567] , 
        \DataPath/RF/bus_selected_win_data[566] , 
        \DataPath/RF/bus_selected_win_data[565] , 
        \DataPath/RF/bus_selected_win_data[564] , 
        \DataPath/RF/bus_selected_win_data[563] , 
        \DataPath/RF/bus_selected_win_data[562] , 
        \DataPath/RF/bus_selected_win_data[561] , 
        \DataPath/RF/bus_selected_win_data[560] , 
        \DataPath/RF/bus_selected_win_data[559] , 
        \DataPath/RF/bus_selected_win_data[558] , 
        \DataPath/RF/bus_selected_win_data[557] , 
        \DataPath/RF/bus_selected_win_data[556] , 
        \DataPath/RF/bus_selected_win_data[555] , 
        \DataPath/RF/bus_selected_win_data[554] , 
        \DataPath/RF/bus_selected_win_data[553] , 
        \DataPath/RF/bus_selected_win_data[552] , 
        \DataPath/RF/bus_selected_win_data[551] , 
        \DataPath/RF/bus_selected_win_data[550] , 
        \DataPath/RF/bus_selected_win_data[549] , 
        \DataPath/RF/bus_selected_win_data[548] , 
        \DataPath/RF/bus_selected_win_data[547] , 
        \DataPath/RF/bus_selected_win_data[546] , 
        \DataPath/RF/bus_selected_win_data[545] , 
        \DataPath/RF/bus_selected_win_data[544] , 
        \DataPath/RF/bus_selected_win_data[543] , 
        \DataPath/RF/bus_selected_win_data[542] , 
        \DataPath/RF/bus_selected_win_data[541] , 
        \DataPath/RF/bus_selected_win_data[540] , 
        \DataPath/RF/bus_selected_win_data[539] , 
        \DataPath/RF/bus_selected_win_data[538] , 
        \DataPath/RF/bus_selected_win_data[537] , 
        \DataPath/RF/bus_selected_win_data[536] , 
        \DataPath/RF/bus_selected_win_data[535] , 
        \DataPath/RF/bus_selected_win_data[534] , 
        \DataPath/RF/bus_selected_win_data[533] , 
        \DataPath/RF/bus_selected_win_data[532] , 
        \DataPath/RF/bus_selected_win_data[531] , 
        \DataPath/RF/bus_selected_win_data[530] , 
        \DataPath/RF/bus_selected_win_data[529] , 
        \DataPath/RF/bus_selected_win_data[528] , 
        \DataPath/RF/bus_selected_win_data[527] , 
        \DataPath/RF/bus_selected_win_data[526] , 
        \DataPath/RF/bus_selected_win_data[525] , 
        \DataPath/RF/bus_selected_win_data[524] , 
        \DataPath/RF/bus_selected_win_data[523] , 
        \DataPath/RF/bus_selected_win_data[522] , 
        \DataPath/RF/bus_selected_win_data[521] , 
        \DataPath/RF/bus_selected_win_data[520] , 
        \DataPath/RF/bus_selected_win_data[519] , 
        \DataPath/RF/bus_selected_win_data[518] , 
        \DataPath/RF/bus_selected_win_data[517] , 
        \DataPath/RF/bus_selected_win_data[516] , 
        \DataPath/RF/bus_selected_win_data[515] , 
        \DataPath/RF/bus_selected_win_data[514] , 
        \DataPath/RF/bus_selected_win_data[513] , 
        \DataPath/RF/bus_selected_win_data[512] , 
        \DataPath/RF/bus_selected_win_data[511] , 
        \DataPath/RF/bus_selected_win_data[510] , 
        \DataPath/RF/bus_selected_win_data[509] , 
        \DataPath/RF/bus_selected_win_data[508] , 
        \DataPath/RF/bus_selected_win_data[507] , 
        \DataPath/RF/bus_selected_win_data[506] , 
        \DataPath/RF/bus_selected_win_data[505] , 
        \DataPath/RF/bus_selected_win_data[504] , 
        \DataPath/RF/bus_selected_win_data[503] , 
        \DataPath/RF/bus_selected_win_data[502] , 
        \DataPath/RF/bus_selected_win_data[501] , 
        \DataPath/RF/bus_selected_win_data[500] , 
        \DataPath/RF/bus_selected_win_data[499] , 
        \DataPath/RF/bus_selected_win_data[498] , 
        \DataPath/RF/bus_selected_win_data[497] , 
        \DataPath/RF/bus_selected_win_data[496] , 
        \DataPath/RF/bus_selected_win_data[495] , 
        \DataPath/RF/bus_selected_win_data[494] , 
        \DataPath/RF/bus_selected_win_data[493] , 
        \DataPath/RF/bus_selected_win_data[492] , 
        \DataPath/RF/bus_selected_win_data[491] , 
        \DataPath/RF/bus_selected_win_data[490] , 
        \DataPath/RF/bus_selected_win_data[489] , 
        \DataPath/RF/bus_selected_win_data[488] , 
        \DataPath/RF/bus_selected_win_data[487] , 
        \DataPath/RF/bus_selected_win_data[486] , 
        \DataPath/RF/bus_selected_win_data[485] , 
        \DataPath/RF/bus_selected_win_data[484] , 
        \DataPath/RF/bus_selected_win_data[483] , 
        \DataPath/RF/bus_selected_win_data[482] , 
        \DataPath/RF/bus_selected_win_data[481] , 
        \DataPath/RF/bus_selected_win_data[480] , 
        \DataPath/RF/bus_selected_win_data[479] , 
        \DataPath/RF/bus_selected_win_data[478] , 
        \DataPath/RF/bus_selected_win_data[477] , 
        \DataPath/RF/bus_selected_win_data[476] , 
        \DataPath/RF/bus_selected_win_data[475] , 
        \DataPath/RF/bus_selected_win_data[474] , 
        \DataPath/RF/bus_selected_win_data[473] , 
        \DataPath/RF/bus_selected_win_data[472] , 
        \DataPath/RF/bus_selected_win_data[471] , 
        \DataPath/RF/bus_selected_win_data[470] , 
        \DataPath/RF/bus_selected_win_data[469] , 
        \DataPath/RF/bus_selected_win_data[468] , 
        \DataPath/RF/bus_selected_win_data[467] , 
        \DataPath/RF/bus_selected_win_data[466] , 
        \DataPath/RF/bus_selected_win_data[465] , 
        \DataPath/RF/bus_selected_win_data[464] , 
        \DataPath/RF/bus_selected_win_data[463] , 
        \DataPath/RF/bus_selected_win_data[462] , 
        \DataPath/RF/bus_selected_win_data[461] , 
        \DataPath/RF/bus_selected_win_data[460] , 
        \DataPath/RF/bus_selected_win_data[459] , 
        \DataPath/RF/bus_selected_win_data[458] , 
        \DataPath/RF/bus_selected_win_data[457] , 
        \DataPath/RF/bus_selected_win_data[456] , 
        \DataPath/RF/bus_selected_win_data[455] , 
        \DataPath/RF/bus_selected_win_data[454] , 
        \DataPath/RF/bus_selected_win_data[453] , 
        \DataPath/RF/bus_selected_win_data[452] , 
        \DataPath/RF/bus_selected_win_data[451] , 
        \DataPath/RF/bus_selected_win_data[450] , 
        \DataPath/RF/bus_selected_win_data[449] , 
        \DataPath/RF/bus_selected_win_data[448] , 
        \DataPath/RF/bus_selected_win_data[447] , 
        \DataPath/RF/bus_selected_win_data[446] , 
        \DataPath/RF/bus_selected_win_data[445] , 
        \DataPath/RF/bus_selected_win_data[444] , 
        \DataPath/RF/bus_selected_win_data[443] , 
        \DataPath/RF/bus_selected_win_data[442] , 
        \DataPath/RF/bus_selected_win_data[441] , 
        \DataPath/RF/bus_selected_win_data[440] , 
        \DataPath/RF/bus_selected_win_data[439] , 
        \DataPath/RF/bus_selected_win_data[438] , 
        \DataPath/RF/bus_selected_win_data[437] , 
        \DataPath/RF/bus_selected_win_data[436] , 
        \DataPath/RF/bus_selected_win_data[435] , 
        \DataPath/RF/bus_selected_win_data[434] , 
        \DataPath/RF/bus_selected_win_data[433] , 
        \DataPath/RF/bus_selected_win_data[432] , 
        \DataPath/RF/bus_selected_win_data[431] , 
        \DataPath/RF/bus_selected_win_data[430] , 
        \DataPath/RF/bus_selected_win_data[429] , 
        \DataPath/RF/bus_selected_win_data[428] , 
        \DataPath/RF/bus_selected_win_data[427] , 
        \DataPath/RF/bus_selected_win_data[426] , 
        \DataPath/RF/bus_selected_win_data[425] , 
        \DataPath/RF/bus_selected_win_data[424] , 
        \DataPath/RF/bus_selected_win_data[423] , 
        \DataPath/RF/bus_selected_win_data[422] , 
        \DataPath/RF/bus_selected_win_data[421] , 
        \DataPath/RF/bus_selected_win_data[420] , 
        \DataPath/RF/bus_selected_win_data[419] , 
        \DataPath/RF/bus_selected_win_data[418] , 
        \DataPath/RF/bus_selected_win_data[417] , 
        \DataPath/RF/bus_selected_win_data[416] , 
        \DataPath/RF/bus_selected_win_data[415] , 
        \DataPath/RF/bus_selected_win_data[414] , 
        \DataPath/RF/bus_selected_win_data[413] , 
        \DataPath/RF/bus_selected_win_data[412] , 
        \DataPath/RF/bus_selected_win_data[411] , 
        \DataPath/RF/bus_selected_win_data[410] , 
        \DataPath/RF/bus_selected_win_data[409] , 
        \DataPath/RF/bus_selected_win_data[408] , 
        \DataPath/RF/bus_selected_win_data[407] , 
        \DataPath/RF/bus_selected_win_data[406] , 
        \DataPath/RF/bus_selected_win_data[405] , 
        \DataPath/RF/bus_selected_win_data[404] , 
        \DataPath/RF/bus_selected_win_data[403] , 
        \DataPath/RF/bus_selected_win_data[402] , 
        \DataPath/RF/bus_selected_win_data[401] , 
        \DataPath/RF/bus_selected_win_data[400] , 
        \DataPath/RF/bus_selected_win_data[399] , 
        \DataPath/RF/bus_selected_win_data[398] , 
        \DataPath/RF/bus_selected_win_data[397] , 
        \DataPath/RF/bus_selected_win_data[396] , 
        \DataPath/RF/bus_selected_win_data[395] , 
        \DataPath/RF/bus_selected_win_data[394] , 
        \DataPath/RF/bus_selected_win_data[393] , 
        \DataPath/RF/bus_selected_win_data[392] , 
        \DataPath/RF/bus_selected_win_data[391] , 
        \DataPath/RF/bus_selected_win_data[390] , 
        \DataPath/RF/bus_selected_win_data[389] , 
        \DataPath/RF/bus_selected_win_data[388] , 
        \DataPath/RF/bus_selected_win_data[387] , 
        \DataPath/RF/bus_selected_win_data[386] , 
        \DataPath/RF/bus_selected_win_data[385] , 
        \DataPath/RF/bus_selected_win_data[384] , 
        \DataPath/RF/bus_selected_win_data[383] , 
        \DataPath/RF/bus_selected_win_data[382] , 
        \DataPath/RF/bus_selected_win_data[381] , 
        \DataPath/RF/bus_selected_win_data[380] , 
        \DataPath/RF/bus_selected_win_data[379] , 
        \DataPath/RF/bus_selected_win_data[378] , 
        \DataPath/RF/bus_selected_win_data[377] , 
        \DataPath/RF/bus_selected_win_data[376] , 
        \DataPath/RF/bus_selected_win_data[375] , 
        \DataPath/RF/bus_selected_win_data[374] , 
        \DataPath/RF/bus_selected_win_data[373] , 
        \DataPath/RF/bus_selected_win_data[372] , 
        \DataPath/RF/bus_selected_win_data[371] , 
        \DataPath/RF/bus_selected_win_data[370] , 
        \DataPath/RF/bus_selected_win_data[369] , 
        \DataPath/RF/bus_selected_win_data[368] , 
        \DataPath/RF/bus_selected_win_data[367] , 
        \DataPath/RF/bus_selected_win_data[366] , 
        \DataPath/RF/bus_selected_win_data[365] , 
        \DataPath/RF/bus_selected_win_data[364] , 
        \DataPath/RF/bus_selected_win_data[363] , 
        \DataPath/RF/bus_selected_win_data[362] , 
        \DataPath/RF/bus_selected_win_data[361] , 
        \DataPath/RF/bus_selected_win_data[360] , 
        \DataPath/RF/bus_selected_win_data[359] , 
        \DataPath/RF/bus_selected_win_data[358] , 
        \DataPath/RF/bus_selected_win_data[357] , 
        \DataPath/RF/bus_selected_win_data[356] , 
        \DataPath/RF/bus_selected_win_data[355] , 
        \DataPath/RF/bus_selected_win_data[354] , 
        \DataPath/RF/bus_selected_win_data[353] , 
        \DataPath/RF/bus_selected_win_data[352] , 
        \DataPath/RF/bus_selected_win_data[351] , 
        \DataPath/RF/bus_selected_win_data[350] , 
        \DataPath/RF/bus_selected_win_data[349] , 
        \DataPath/RF/bus_selected_win_data[348] , 
        \DataPath/RF/bus_selected_win_data[347] , 
        \DataPath/RF/bus_selected_win_data[346] , 
        \DataPath/RF/bus_selected_win_data[345] , 
        \DataPath/RF/bus_selected_win_data[344] , 
        \DataPath/RF/bus_selected_win_data[343] , 
        \DataPath/RF/bus_selected_win_data[342] , 
        \DataPath/RF/bus_selected_win_data[341] , 
        \DataPath/RF/bus_selected_win_data[340] , 
        \DataPath/RF/bus_selected_win_data[339] , 
        \DataPath/RF/bus_selected_win_data[338] , 
        \DataPath/RF/bus_selected_win_data[337] , 
        \DataPath/RF/bus_selected_win_data[336] , 
        \DataPath/RF/bus_selected_win_data[335] , 
        \DataPath/RF/bus_selected_win_data[334] , 
        \DataPath/RF/bus_selected_win_data[333] , 
        \DataPath/RF/bus_selected_win_data[332] , 
        \DataPath/RF/bus_selected_win_data[331] , 
        \DataPath/RF/bus_selected_win_data[330] , 
        \DataPath/RF/bus_selected_win_data[329] , 
        \DataPath/RF/bus_selected_win_data[328] , 
        \DataPath/RF/bus_selected_win_data[327] , 
        \DataPath/RF/bus_selected_win_data[326] , 
        \DataPath/RF/bus_selected_win_data[325] , 
        \DataPath/RF/bus_selected_win_data[324] , 
        \DataPath/RF/bus_selected_win_data[323] , 
        \DataPath/RF/bus_selected_win_data[322] , 
        \DataPath/RF/bus_selected_win_data[321] , 
        \DataPath/RF/bus_selected_win_data[320] , 
        \DataPath/RF/bus_selected_win_data[319] , 
        \DataPath/RF/bus_selected_win_data[318] , 
        \DataPath/RF/bus_selected_win_data[317] , 
        \DataPath/RF/bus_selected_win_data[316] , 
        \DataPath/RF/bus_selected_win_data[315] , 
        \DataPath/RF/bus_selected_win_data[314] , 
        \DataPath/RF/bus_selected_win_data[313] , 
        \DataPath/RF/bus_selected_win_data[312] , 
        \DataPath/RF/bus_selected_win_data[311] , 
        \DataPath/RF/bus_selected_win_data[310] , 
        \DataPath/RF/bus_selected_win_data[309] , 
        \DataPath/RF/bus_selected_win_data[308] , 
        \DataPath/RF/bus_selected_win_data[307] , 
        \DataPath/RF/bus_selected_win_data[306] , 
        \DataPath/RF/bus_selected_win_data[305] , 
        \DataPath/RF/bus_selected_win_data[304] , 
        \DataPath/RF/bus_selected_win_data[303] , 
        \DataPath/RF/bus_selected_win_data[302] , 
        \DataPath/RF/bus_selected_win_data[301] , 
        \DataPath/RF/bus_selected_win_data[300] , 
        \DataPath/RF/bus_selected_win_data[299] , 
        \DataPath/RF/bus_selected_win_data[298] , 
        \DataPath/RF/bus_selected_win_data[297] , 
        \DataPath/RF/bus_selected_win_data[296] , 
        \DataPath/RF/bus_selected_win_data[295] , 
        \DataPath/RF/bus_selected_win_data[294] , 
        \DataPath/RF/bus_selected_win_data[293] , 
        \DataPath/RF/bus_selected_win_data[292] , 
        \DataPath/RF/bus_selected_win_data[291] , 
        \DataPath/RF/bus_selected_win_data[290] , 
        \DataPath/RF/bus_selected_win_data[289] , 
        \DataPath/RF/bus_selected_win_data[288] , 
        \DataPath/RF/bus_selected_win_data[287] , 
        \DataPath/RF/bus_selected_win_data[286] , 
        \DataPath/RF/bus_selected_win_data[285] , 
        \DataPath/RF/bus_selected_win_data[284] , 
        \DataPath/RF/bus_selected_win_data[283] , 
        \DataPath/RF/bus_selected_win_data[282] , 
        \DataPath/RF/bus_selected_win_data[281] , 
        \DataPath/RF/bus_selected_win_data[280] , 
        \DataPath/RF/bus_selected_win_data[279] , 
        \DataPath/RF/bus_selected_win_data[278] , 
        \DataPath/RF/bus_selected_win_data[277] , 
        \DataPath/RF/bus_selected_win_data[276] , 
        \DataPath/RF/bus_selected_win_data[275] , 
        \DataPath/RF/bus_selected_win_data[274] , 
        \DataPath/RF/bus_selected_win_data[273] , 
        \DataPath/RF/bus_selected_win_data[272] , 
        \DataPath/RF/bus_selected_win_data[271] , 
        \DataPath/RF/bus_selected_win_data[270] , 
        \DataPath/RF/bus_selected_win_data[269] , 
        \DataPath/RF/bus_selected_win_data[268] , 
        \DataPath/RF/bus_selected_win_data[267] , 
        \DataPath/RF/bus_selected_win_data[266] , 
        \DataPath/RF/bus_selected_win_data[265] , 
        \DataPath/RF/bus_selected_win_data[264] , 
        \DataPath/RF/bus_selected_win_data[263] , 
        \DataPath/RF/bus_selected_win_data[262] , 
        \DataPath/RF/bus_selected_win_data[261] , 
        \DataPath/RF/bus_selected_win_data[260] , 
        \DataPath/RF/bus_selected_win_data[259] , 
        \DataPath/RF/bus_selected_win_data[258] , 
        \DataPath/RF/bus_selected_win_data[257] , 
        \DataPath/RF/bus_selected_win_data[256] , 
        \DataPath/RF/bus_selected_win_data[255] , 
        \DataPath/RF/bus_selected_win_data[254] , 
        \DataPath/RF/bus_selected_win_data[253] , 
        \DataPath/RF/bus_selected_win_data[252] , 
        \DataPath/RF/bus_selected_win_data[251] , 
        \DataPath/RF/bus_selected_win_data[250] , 
        \DataPath/RF/bus_selected_win_data[249] , 
        \DataPath/RF/bus_selected_win_data[248] , 
        \DataPath/RF/bus_selected_win_data[247] , 
        \DataPath/RF/bus_selected_win_data[246] , 
        \DataPath/RF/bus_selected_win_data[245] , 
        \DataPath/RF/bus_selected_win_data[244] , 
        \DataPath/RF/bus_selected_win_data[243] , 
        \DataPath/RF/bus_selected_win_data[242] , 
        \DataPath/RF/bus_selected_win_data[241] , 
        \DataPath/RF/bus_selected_win_data[240] , 
        \DataPath/RF/bus_selected_win_data[239] , 
        \DataPath/RF/bus_selected_win_data[238] , 
        \DataPath/RF/bus_selected_win_data[237] , 
        \DataPath/RF/bus_selected_win_data[236] , 
        \DataPath/RF/bus_selected_win_data[235] , 
        \DataPath/RF/bus_selected_win_data[234] , 
        \DataPath/RF/bus_selected_win_data[233] , 
        \DataPath/RF/bus_selected_win_data[232] , 
        \DataPath/RF/bus_selected_win_data[231] , 
        \DataPath/RF/bus_selected_win_data[230] , 
        \DataPath/RF/bus_selected_win_data[229] , 
        \DataPath/RF/bus_selected_win_data[228] , 
        \DataPath/RF/bus_selected_win_data[227] , 
        \DataPath/RF/bus_selected_win_data[226] , 
        \DataPath/RF/bus_selected_win_data[225] , 
        \DataPath/RF/bus_selected_win_data[224] , 
        \DataPath/RF/bus_selected_win_data[223] , 
        \DataPath/RF/bus_selected_win_data[222] , 
        \DataPath/RF/bus_selected_win_data[221] , 
        \DataPath/RF/bus_selected_win_data[220] , 
        \DataPath/RF/bus_selected_win_data[219] , 
        \DataPath/RF/bus_selected_win_data[218] , 
        \DataPath/RF/bus_selected_win_data[217] , 
        \DataPath/RF/bus_selected_win_data[216] , 
        \DataPath/RF/bus_selected_win_data[215] , 
        \DataPath/RF/bus_selected_win_data[214] , 
        \DataPath/RF/bus_selected_win_data[213] , 
        \DataPath/RF/bus_selected_win_data[212] , 
        \DataPath/RF/bus_selected_win_data[211] , 
        \DataPath/RF/bus_selected_win_data[210] , 
        \DataPath/RF/bus_selected_win_data[209] , 
        \DataPath/RF/bus_selected_win_data[208] , 
        \DataPath/RF/bus_selected_win_data[207] , 
        \DataPath/RF/bus_selected_win_data[206] , 
        \DataPath/RF/bus_selected_win_data[205] , 
        \DataPath/RF/bus_selected_win_data[204] , 
        \DataPath/RF/bus_selected_win_data[203] , 
        \DataPath/RF/bus_selected_win_data[202] , 
        \DataPath/RF/bus_selected_win_data[201] , 
        \DataPath/RF/bus_selected_win_data[200] , 
        \DataPath/RF/bus_selected_win_data[199] , 
        \DataPath/RF/bus_selected_win_data[198] , 
        \DataPath/RF/bus_selected_win_data[197] , 
        \DataPath/RF/bus_selected_win_data[196] , 
        \DataPath/RF/bus_selected_win_data[195] , 
        \DataPath/RF/bus_selected_win_data[194] , 
        \DataPath/RF/bus_selected_win_data[193] , 
        \DataPath/RF/bus_selected_win_data[192] , 
        \DataPath/RF/bus_selected_win_data[191] , 
        \DataPath/RF/bus_selected_win_data[190] , 
        \DataPath/RF/bus_selected_win_data[189] , 
        \DataPath/RF/bus_selected_win_data[188] , 
        \DataPath/RF/bus_selected_win_data[187] , 
        \DataPath/RF/bus_selected_win_data[186] , 
        \DataPath/RF/bus_selected_win_data[185] , 
        \DataPath/RF/bus_selected_win_data[184] , 
        \DataPath/RF/bus_selected_win_data[183] , 
        \DataPath/RF/bus_selected_win_data[182] , 
        \DataPath/RF/bus_selected_win_data[181] , 
        \DataPath/RF/bus_selected_win_data[180] , 
        \DataPath/RF/bus_selected_win_data[179] , 
        \DataPath/RF/bus_selected_win_data[178] , 
        \DataPath/RF/bus_selected_win_data[177] , 
        \DataPath/RF/bus_selected_win_data[176] , 
        \DataPath/RF/bus_selected_win_data[175] , 
        \DataPath/RF/bus_selected_win_data[174] , 
        \DataPath/RF/bus_selected_win_data[173] , 
        \DataPath/RF/bus_selected_win_data[172] , 
        \DataPath/RF/bus_selected_win_data[171] , 
        \DataPath/RF/bus_selected_win_data[170] , 
        \DataPath/RF/bus_selected_win_data[169] , 
        \DataPath/RF/bus_selected_win_data[168] , 
        \DataPath/RF/bus_selected_win_data[167] , 
        \DataPath/RF/bus_selected_win_data[166] , 
        \DataPath/RF/bus_selected_win_data[165] , 
        \DataPath/RF/bus_selected_win_data[164] , 
        \DataPath/RF/bus_selected_win_data[163] , 
        \DataPath/RF/bus_selected_win_data[162] , 
        \DataPath/RF/bus_selected_win_data[161] , 
        \DataPath/RF/bus_selected_win_data[160] , 
        \DataPath/RF/bus_selected_win_data[159] , 
        \DataPath/RF/bus_selected_win_data[158] , 
        \DataPath/RF/bus_selected_win_data[157] , 
        \DataPath/RF/bus_selected_win_data[156] , 
        \DataPath/RF/bus_selected_win_data[155] , 
        \DataPath/RF/bus_selected_win_data[154] , 
        \DataPath/RF/bus_selected_win_data[153] , 
        \DataPath/RF/bus_selected_win_data[152] , 
        \DataPath/RF/bus_selected_win_data[151] , 
        \DataPath/RF/bus_selected_win_data[150] , 
        \DataPath/RF/bus_selected_win_data[149] , 
        \DataPath/RF/bus_selected_win_data[148] , 
        \DataPath/RF/bus_selected_win_data[147] , 
        \DataPath/RF/bus_selected_win_data[146] , 
        \DataPath/RF/bus_selected_win_data[145] , 
        \DataPath/RF/bus_selected_win_data[144] , 
        \DataPath/RF/bus_selected_win_data[143] , 
        \DataPath/RF/bus_selected_win_data[142] , 
        \DataPath/RF/bus_selected_win_data[141] , 
        \DataPath/RF/bus_selected_win_data[140] , 
        \DataPath/RF/bus_selected_win_data[139] , 
        \DataPath/RF/bus_selected_win_data[138] , 
        \DataPath/RF/bus_selected_win_data[137] , 
        \DataPath/RF/bus_selected_win_data[136] , 
        \DataPath/RF/bus_selected_win_data[135] , 
        \DataPath/RF/bus_selected_win_data[134] , 
        \DataPath/RF/bus_selected_win_data[133] , 
        \DataPath/RF/bus_selected_win_data[132] , 
        \DataPath/RF/bus_selected_win_data[131] , 
        \DataPath/RF/bus_selected_win_data[130] , 
        \DataPath/RF/bus_selected_win_data[129] , 
        \DataPath/RF/bus_selected_win_data[128] , 
        \DataPath/RF/bus_selected_win_data[127] , 
        \DataPath/RF/bus_selected_win_data[126] , 
        \DataPath/RF/bus_selected_win_data[125] , 
        \DataPath/RF/bus_selected_win_data[124] , 
        \DataPath/RF/bus_selected_win_data[123] , 
        \DataPath/RF/bus_selected_win_data[122] , 
        \DataPath/RF/bus_selected_win_data[121] , 
        \DataPath/RF/bus_selected_win_data[120] , 
        \DataPath/RF/bus_selected_win_data[119] , 
        \DataPath/RF/bus_selected_win_data[118] , 
        \DataPath/RF/bus_selected_win_data[117] , 
        \DataPath/RF/bus_selected_win_data[116] , 
        \DataPath/RF/bus_selected_win_data[115] , 
        \DataPath/RF/bus_selected_win_data[114] , 
        \DataPath/RF/bus_selected_win_data[113] , 
        \DataPath/RF/bus_selected_win_data[112] , 
        \DataPath/RF/bus_selected_win_data[111] , 
        \DataPath/RF/bus_selected_win_data[110] , 
        \DataPath/RF/bus_selected_win_data[109] , 
        \DataPath/RF/bus_selected_win_data[108] , 
        \DataPath/RF/bus_selected_win_data[107] , 
        \DataPath/RF/bus_selected_win_data[106] , 
        \DataPath/RF/bus_selected_win_data[105] , 
        \DataPath/RF/bus_selected_win_data[104] , 
        \DataPath/RF/bus_selected_win_data[103] , 
        \DataPath/RF/bus_selected_win_data[102] , 
        \DataPath/RF/bus_selected_win_data[101] , 
        \DataPath/RF/bus_selected_win_data[100] , 
        \DataPath/RF/bus_selected_win_data[99] , 
        \DataPath/RF/bus_selected_win_data[98] , 
        \DataPath/RF/bus_selected_win_data[97] , 
        \DataPath/RF/bus_selected_win_data[96] , 
        \DataPath/RF/bus_selected_win_data[95] , 
        \DataPath/RF/bus_selected_win_data[94] , 
        \DataPath/RF/bus_selected_win_data[93] , 
        \DataPath/RF/bus_selected_win_data[92] , 
        \DataPath/RF/bus_selected_win_data[91] , 
        \DataPath/RF/bus_selected_win_data[90] , 
        \DataPath/RF/bus_selected_win_data[89] , 
        \DataPath/RF/bus_selected_win_data[88] , 
        \DataPath/RF/bus_selected_win_data[87] , 
        \DataPath/RF/bus_selected_win_data[86] , 
        \DataPath/RF/bus_selected_win_data[85] , 
        \DataPath/RF/bus_selected_win_data[84] , 
        \DataPath/RF/bus_selected_win_data[83] , 
        \DataPath/RF/bus_selected_win_data[82] , 
        \DataPath/RF/bus_selected_win_data[81] , 
        \DataPath/RF/bus_selected_win_data[80] , 
        \DataPath/RF/bus_selected_win_data[79] , 
        \DataPath/RF/bus_selected_win_data[78] , 
        \DataPath/RF/bus_selected_win_data[77] , 
        \DataPath/RF/bus_selected_win_data[76] , 
        \DataPath/RF/bus_selected_win_data[75] , 
        \DataPath/RF/bus_selected_win_data[74] , 
        \DataPath/RF/bus_selected_win_data[73] , 
        \DataPath/RF/bus_selected_win_data[72] , 
        \DataPath/RF/bus_selected_win_data[71] , 
        \DataPath/RF/bus_selected_win_data[70] , 
        \DataPath/RF/bus_selected_win_data[69] , 
        \DataPath/RF/bus_selected_win_data[68] , 
        \DataPath/RF/bus_selected_win_data[67] , 
        \DataPath/RF/bus_selected_win_data[66] , 
        \DataPath/RF/bus_selected_win_data[65] , 
        \DataPath/RF/bus_selected_win_data[64] , 
        \DataPath/RF/bus_selected_win_data[63] , 
        \DataPath/RF/bus_selected_win_data[62] , 
        \DataPath/RF/bus_selected_win_data[61] , 
        \DataPath/RF/bus_selected_win_data[60] , 
        \DataPath/RF/bus_selected_win_data[59] , 
        \DataPath/RF/bus_selected_win_data[58] , 
        \DataPath/RF/bus_selected_win_data[57] , 
        \DataPath/RF/bus_selected_win_data[56] , 
        \DataPath/RF/bus_selected_win_data[55] , 
        \DataPath/RF/bus_selected_win_data[54] , 
        \DataPath/RF/bus_selected_win_data[53] , 
        \DataPath/RF/bus_selected_win_data[52] , 
        \DataPath/RF/bus_selected_win_data[51] , 
        \DataPath/RF/bus_selected_win_data[50] , 
        \DataPath/RF/bus_selected_win_data[49] , 
        \DataPath/RF/bus_selected_win_data[48] , 
        \DataPath/RF/bus_selected_win_data[47] , 
        \DataPath/RF/bus_selected_win_data[46] , 
        \DataPath/RF/bus_selected_win_data[45] , 
        \DataPath/RF/bus_selected_win_data[44] , 
        \DataPath/RF/bus_selected_win_data[43] , 
        \DataPath/RF/bus_selected_win_data[42] , 
        \DataPath/RF/bus_selected_win_data[41] , 
        \DataPath/RF/bus_selected_win_data[40] , 
        \DataPath/RF/bus_selected_win_data[39] , 
        \DataPath/RF/bus_selected_win_data[38] , 
        \DataPath/RF/bus_selected_win_data[37] , 
        \DataPath/RF/bus_selected_win_data[36] , 
        \DataPath/RF/bus_selected_win_data[35] , 
        \DataPath/RF/bus_selected_win_data[34] , 
        \DataPath/RF/bus_selected_win_data[33] , 
        \DataPath/RF/bus_selected_win_data[32] , 
        \DataPath/RF/bus_selected_win_data[31] , 
        \DataPath/RF/bus_selected_win_data[30] , 
        \DataPath/RF/bus_selected_win_data[29] , 
        \DataPath/RF/bus_selected_win_data[28] , 
        \DataPath/RF/bus_selected_win_data[27] , 
        \DataPath/RF/bus_selected_win_data[26] , 
        \DataPath/RF/bus_selected_win_data[25] , 
        \DataPath/RF/bus_selected_win_data[24] , 
        \DataPath/RF/bus_selected_win_data[23] , 
        \DataPath/RF/bus_selected_win_data[22] , 
        \DataPath/RF/bus_selected_win_data[21] , 
        \DataPath/RF/bus_selected_win_data[20] , 
        \DataPath/RF/bus_selected_win_data[19] , 
        \DataPath/RF/bus_selected_win_data[18] , 
        \DataPath/RF/bus_selected_win_data[17] , 
        \DataPath/RF/bus_selected_win_data[16] , 
        \DataPath/RF/bus_selected_win_data[15] , 
        \DataPath/RF/bus_selected_win_data[14] , 
        \DataPath/RF/bus_selected_win_data[13] , 
        \DataPath/RF/bus_selected_win_data[12] , 
        \DataPath/RF/bus_selected_win_data[11] , 
        \DataPath/RF/bus_selected_win_data[10] , 
        \DataPath/RF/bus_selected_win_data[9] , 
        \DataPath/RF/bus_selected_win_data[8] , 
        \DataPath/RF/bus_selected_win_data[7] , 
        \DataPath/RF/bus_selected_win_data[6] , 
        \DataPath/RF/bus_selected_win_data[5] , 
        \DataPath/RF/bus_selected_win_data[4] , 
        \DataPath/RF/bus_selected_win_data[3] , 
        \DataPath/RF/bus_selected_win_data[2] , 
        \DataPath/RF/bus_selected_win_data[1] , 
        \DataPath/RF/bus_selected_win_data[0] , 
        \DataPath/RF/bus_complete_win_data[255] , 
        \DataPath/RF/bus_complete_win_data[254] , 
        \DataPath/RF/bus_complete_win_data[253] , 
        \DataPath/RF/bus_complete_win_data[252] , 
        \DataPath/RF/bus_complete_win_data[251] , 
        \DataPath/RF/bus_complete_win_data[250] , 
        \DataPath/RF/bus_complete_win_data[249] , 
        \DataPath/RF/bus_complete_win_data[248] , 
        \DataPath/RF/bus_complete_win_data[247] , 
        \DataPath/RF/bus_complete_win_data[246] , 
        \DataPath/RF/bus_complete_win_data[245] , 
        \DataPath/RF/bus_complete_win_data[244] , 
        \DataPath/RF/bus_complete_win_data[243] , 
        \DataPath/RF/bus_complete_win_data[242] , 
        \DataPath/RF/bus_complete_win_data[241] , 
        \DataPath/RF/bus_complete_win_data[240] , 
        \DataPath/RF/bus_complete_win_data[239] , 
        \DataPath/RF/bus_complete_win_data[238] , 
        \DataPath/RF/bus_complete_win_data[237] , 
        \DataPath/RF/bus_complete_win_data[236] , 
        \DataPath/RF/bus_complete_win_data[235] , 
        \DataPath/RF/bus_complete_win_data[234] , 
        \DataPath/RF/bus_complete_win_data[233] , 
        \DataPath/RF/bus_complete_win_data[232] , 
        \DataPath/RF/bus_complete_win_data[231] , 
        \DataPath/RF/bus_complete_win_data[230] , 
        \DataPath/RF/bus_complete_win_data[229] , 
        \DataPath/RF/bus_complete_win_data[228] , 
        \DataPath/RF/bus_complete_win_data[227] , 
        \DataPath/RF/bus_complete_win_data[226] , 
        \DataPath/RF/bus_complete_win_data[225] , 
        \DataPath/RF/bus_complete_win_data[224] , 
        \DataPath/RF/bus_complete_win_data[223] , 
        \DataPath/RF/bus_complete_win_data[222] , 
        \DataPath/RF/bus_complete_win_data[221] , 
        \DataPath/RF/bus_complete_win_data[220] , 
        \DataPath/RF/bus_complete_win_data[219] , 
        \DataPath/RF/bus_complete_win_data[218] , 
        \DataPath/RF/bus_complete_win_data[217] , 
        \DataPath/RF/bus_complete_win_data[216] , 
        \DataPath/RF/bus_complete_win_data[215] , 
        \DataPath/RF/bus_complete_win_data[214] , 
        \DataPath/RF/bus_complete_win_data[213] , 
        \DataPath/RF/bus_complete_win_data[212] , 
        \DataPath/RF/bus_complete_win_data[211] , 
        \DataPath/RF/bus_complete_win_data[210] , 
        \DataPath/RF/bus_complete_win_data[209] , 
        \DataPath/RF/bus_complete_win_data[208] , 
        \DataPath/RF/bus_complete_win_data[207] , 
        \DataPath/RF/bus_complete_win_data[206] , 
        \DataPath/RF/bus_complete_win_data[205] , 
        \DataPath/RF/bus_complete_win_data[204] , 
        \DataPath/RF/bus_complete_win_data[203] , 
        \DataPath/RF/bus_complete_win_data[202] , 
        \DataPath/RF/bus_complete_win_data[201] , 
        \DataPath/RF/bus_complete_win_data[200] , 
        \DataPath/RF/bus_complete_win_data[199] , 
        \DataPath/RF/bus_complete_win_data[198] , 
        \DataPath/RF/bus_complete_win_data[197] , 
        \DataPath/RF/bus_complete_win_data[196] , 
        \DataPath/RF/bus_complete_win_data[195] , 
        \DataPath/RF/bus_complete_win_data[194] , 
        \DataPath/RF/bus_complete_win_data[193] , 
        \DataPath/RF/bus_complete_win_data[192] , 
        \DataPath/RF/bus_complete_win_data[191] , 
        \DataPath/RF/bus_complete_win_data[190] , 
        \DataPath/RF/bus_complete_win_data[189] , 
        \DataPath/RF/bus_complete_win_data[188] , 
        \DataPath/RF/bus_complete_win_data[187] , 
        \DataPath/RF/bus_complete_win_data[186] , 
        \DataPath/RF/bus_complete_win_data[185] , 
        \DataPath/RF/bus_complete_win_data[184] , 
        \DataPath/RF/bus_complete_win_data[183] , 
        \DataPath/RF/bus_complete_win_data[182] , 
        \DataPath/RF/bus_complete_win_data[181] , 
        \DataPath/RF/bus_complete_win_data[180] , 
        \DataPath/RF/bus_complete_win_data[179] , 
        \DataPath/RF/bus_complete_win_data[178] , 
        \DataPath/RF/bus_complete_win_data[177] , 
        \DataPath/RF/bus_complete_win_data[176] , 
        \DataPath/RF/bus_complete_win_data[175] , 
        \DataPath/RF/bus_complete_win_data[174] , 
        \DataPath/RF/bus_complete_win_data[173] , 
        \DataPath/RF/bus_complete_win_data[172] , 
        \DataPath/RF/bus_complete_win_data[171] , 
        \DataPath/RF/bus_complete_win_data[170] , 
        \DataPath/RF/bus_complete_win_data[169] , 
        \DataPath/RF/bus_complete_win_data[168] , 
        \DataPath/RF/bus_complete_win_data[167] , 
        \DataPath/RF/bus_complete_win_data[166] , 
        \DataPath/RF/bus_complete_win_data[165] , 
        \DataPath/RF/bus_complete_win_data[164] , 
        \DataPath/RF/bus_complete_win_data[163] , 
        \DataPath/RF/bus_complete_win_data[162] , 
        \DataPath/RF/bus_complete_win_data[161] , 
        \DataPath/RF/bus_complete_win_data[160] , 
        \DataPath/RF/bus_complete_win_data[159] , 
        \DataPath/RF/bus_complete_win_data[158] , 
        \DataPath/RF/bus_complete_win_data[157] , 
        \DataPath/RF/bus_complete_win_data[156] , 
        \DataPath/RF/bus_complete_win_data[155] , 
        \DataPath/RF/bus_complete_win_data[154] , 
        \DataPath/RF/bus_complete_win_data[153] , 
        \DataPath/RF/bus_complete_win_data[152] , 
        \DataPath/RF/bus_complete_win_data[151] , 
        \DataPath/RF/bus_complete_win_data[150] , 
        \DataPath/RF/bus_complete_win_data[149] , 
        \DataPath/RF/bus_complete_win_data[148] , 
        \DataPath/RF/bus_complete_win_data[147] , 
        \DataPath/RF/bus_complete_win_data[146] , 
        \DataPath/RF/bus_complete_win_data[145] , 
        \DataPath/RF/bus_complete_win_data[144] , 
        \DataPath/RF/bus_complete_win_data[143] , 
        \DataPath/RF/bus_complete_win_data[142] , 
        \DataPath/RF/bus_complete_win_data[141] , 
        \DataPath/RF/bus_complete_win_data[140] , 
        \DataPath/RF/bus_complete_win_data[139] , 
        \DataPath/RF/bus_complete_win_data[138] , 
        \DataPath/RF/bus_complete_win_data[137] , 
        \DataPath/RF/bus_complete_win_data[136] , 
        \DataPath/RF/bus_complete_win_data[135] , 
        \DataPath/RF/bus_complete_win_data[134] , 
        \DataPath/RF/bus_complete_win_data[133] , 
        \DataPath/RF/bus_complete_win_data[132] , 
        \DataPath/RF/bus_complete_win_data[131] , 
        \DataPath/RF/bus_complete_win_data[130] , 
        \DataPath/RF/bus_complete_win_data[129] , 
        \DataPath/RF/bus_complete_win_data[128] , 
        \DataPath/RF/bus_complete_win_data[127] , 
        \DataPath/RF/bus_complete_win_data[126] , 
        \DataPath/RF/bus_complete_win_data[125] , 
        \DataPath/RF/bus_complete_win_data[124] , 
        \DataPath/RF/bus_complete_win_data[123] , 
        \DataPath/RF/bus_complete_win_data[122] , 
        \DataPath/RF/bus_complete_win_data[121] , 
        \DataPath/RF/bus_complete_win_data[120] , 
        \DataPath/RF/bus_complete_win_data[119] , 
        \DataPath/RF/bus_complete_win_data[118] , 
        \DataPath/RF/bus_complete_win_data[117] , 
        \DataPath/RF/bus_complete_win_data[116] , 
        \DataPath/RF/bus_complete_win_data[115] , 
        \DataPath/RF/bus_complete_win_data[114] , 
        \DataPath/RF/bus_complete_win_data[113] , 
        \DataPath/RF/bus_complete_win_data[112] , 
        \DataPath/RF/bus_complete_win_data[111] , 
        \DataPath/RF/bus_complete_win_data[110] , 
        \DataPath/RF/bus_complete_win_data[109] , 
        \DataPath/RF/bus_complete_win_data[108] , 
        \DataPath/RF/bus_complete_win_data[107] , 
        \DataPath/RF/bus_complete_win_data[106] , 
        \DataPath/RF/bus_complete_win_data[105] , 
        \DataPath/RF/bus_complete_win_data[104] , 
        \DataPath/RF/bus_complete_win_data[103] , 
        \DataPath/RF/bus_complete_win_data[102] , 
        \DataPath/RF/bus_complete_win_data[101] , 
        \DataPath/RF/bus_complete_win_data[100] , 
        \DataPath/RF/bus_complete_win_data[99] , 
        \DataPath/RF/bus_complete_win_data[98] , 
        \DataPath/RF/bus_complete_win_data[97] , 
        \DataPath/RF/bus_complete_win_data[96] , 
        \DataPath/RF/bus_complete_win_data[95] , 
        \DataPath/RF/bus_complete_win_data[94] , 
        \DataPath/RF/bus_complete_win_data[93] , 
        \DataPath/RF/bus_complete_win_data[92] , 
        \DataPath/RF/bus_complete_win_data[91] , 
        \DataPath/RF/bus_complete_win_data[90] , 
        \DataPath/RF/bus_complete_win_data[89] , 
        \DataPath/RF/bus_complete_win_data[88] , 
        \DataPath/RF/bus_complete_win_data[87] , 
        \DataPath/RF/bus_complete_win_data[86] , 
        \DataPath/RF/bus_complete_win_data[85] , 
        \DataPath/RF/bus_complete_win_data[84] , 
        \DataPath/RF/bus_complete_win_data[83] , 
        \DataPath/RF/bus_complete_win_data[82] , 
        \DataPath/RF/bus_complete_win_data[81] , 
        \DataPath/RF/bus_complete_win_data[80] , 
        \DataPath/RF/bus_complete_win_data[79] , 
        \DataPath/RF/bus_complete_win_data[78] , 
        \DataPath/RF/bus_complete_win_data[77] , 
        \DataPath/RF/bus_complete_win_data[76] , 
        \DataPath/RF/bus_complete_win_data[75] , 
        \DataPath/RF/bus_complete_win_data[74] , 
        \DataPath/RF/bus_complete_win_data[73] , 
        \DataPath/RF/bus_complete_win_data[72] , 
        \DataPath/RF/bus_complete_win_data[71] , 
        \DataPath/RF/bus_complete_win_data[70] , 
        \DataPath/RF/bus_complete_win_data[69] , 
        \DataPath/RF/bus_complete_win_data[68] , 
        \DataPath/RF/bus_complete_win_data[67] , 
        \DataPath/RF/bus_complete_win_data[66] , 
        \DataPath/RF/bus_complete_win_data[65] , 
        \DataPath/RF/bus_complete_win_data[64] , 
        \DataPath/RF/bus_complete_win_data[63] , 
        \DataPath/RF/bus_complete_win_data[62] , 
        \DataPath/RF/bus_complete_win_data[61] , 
        \DataPath/RF/bus_complete_win_data[60] , 
        \DataPath/RF/bus_complete_win_data[59] , 
        \DataPath/RF/bus_complete_win_data[58] , 
        \DataPath/RF/bus_complete_win_data[57] , 
        \DataPath/RF/bus_complete_win_data[56] , 
        \DataPath/RF/bus_complete_win_data[55] , 
        \DataPath/RF/bus_complete_win_data[54] , 
        \DataPath/RF/bus_complete_win_data[53] , 
        \DataPath/RF/bus_complete_win_data[52] , 
        \DataPath/RF/bus_complete_win_data[51] , 
        \DataPath/RF/bus_complete_win_data[50] , 
        \DataPath/RF/bus_complete_win_data[49] , 
        \DataPath/RF/bus_complete_win_data[48] , 
        \DataPath/RF/bus_complete_win_data[47] , 
        \DataPath/RF/bus_complete_win_data[46] , 
        \DataPath/RF/bus_complete_win_data[45] , 
        \DataPath/RF/bus_complete_win_data[44] , 
        \DataPath/RF/bus_complete_win_data[43] , 
        \DataPath/RF/bus_complete_win_data[42] , 
        \DataPath/RF/bus_complete_win_data[41] , 
        \DataPath/RF/bus_complete_win_data[40] , 
        \DataPath/RF/bus_complete_win_data[39] , 
        \DataPath/RF/bus_complete_win_data[38] , 
        \DataPath/RF/bus_complete_win_data[37] , 
        \DataPath/RF/bus_complete_win_data[36] , 
        \DataPath/RF/bus_complete_win_data[35] , 
        \DataPath/RF/bus_complete_win_data[34] , 
        \DataPath/RF/bus_complete_win_data[33] , 
        \DataPath/RF/bus_complete_win_data[32] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .Y({\DataPath/RF/internal_out2[31] , 
        \DataPath/RF/internal_out2[30] , \DataPath/RF/internal_out2[29] , 
        \DataPath/RF/internal_out2[28] , \DataPath/RF/internal_out2[27] , 
        \DataPath/RF/internal_out2[26] , \DataPath/RF/internal_out2[25] , 
        \DataPath/RF/internal_out2[24] , \DataPath/RF/internal_out2[23] , 
        \DataPath/RF/internal_out2[22] , \DataPath/RF/internal_out2[21] , 
        \DataPath/RF/internal_out2[20] , \DataPath/RF/internal_out2[19] , 
        \DataPath/RF/internal_out2[18] , \DataPath/RF/internal_out2[17] , 
        \DataPath/RF/internal_out2[16] , \DataPath/RF/internal_out2[15] , 
        \DataPath/RF/internal_out2[14] , \DataPath/RF/internal_out2[13] , 
        \DataPath/RF/internal_out2[12] , \DataPath/RF/internal_out2[11] , 
        \DataPath/RF/internal_out2[10] , \DataPath/RF/internal_out2[9] , 
        \DataPath/RF/internal_out2[8] , \DataPath/RF/internal_out2[7] , 
        \DataPath/RF/internal_out2[6] , \DataPath/RF/internal_out2[5] , 
        \DataPath/RF/internal_out2[4] , \DataPath/RF/internal_out2[3] , 
        \DataPath/RF/internal_out2[2] , \DataPath/RF/internal_out2[1] , 
        \DataPath/RF/internal_out2[0] }) );
  mux_N32_M5_0 \DataPath/RF/RDPORT0  ( .S(i_ADD_RS1), .Q({
        \DataPath/RF/bus_selected_win_data[767] , 
        \DataPath/RF/bus_selected_win_data[766] , 
        \DataPath/RF/bus_selected_win_data[765] , 
        \DataPath/RF/bus_selected_win_data[764] , 
        \DataPath/RF/bus_selected_win_data[763] , 
        \DataPath/RF/bus_selected_win_data[762] , 
        \DataPath/RF/bus_selected_win_data[761] , 
        \DataPath/RF/bus_selected_win_data[760] , 
        \DataPath/RF/bus_selected_win_data[759] , 
        \DataPath/RF/bus_selected_win_data[758] , 
        \DataPath/RF/bus_selected_win_data[757] , 
        \DataPath/RF/bus_selected_win_data[756] , 
        \DataPath/RF/bus_selected_win_data[755] , 
        \DataPath/RF/bus_selected_win_data[754] , 
        \DataPath/RF/bus_selected_win_data[753] , 
        \DataPath/RF/bus_selected_win_data[752] , 
        \DataPath/RF/bus_selected_win_data[751] , 
        \DataPath/RF/bus_selected_win_data[750] , 
        \DataPath/RF/bus_selected_win_data[749] , 
        \DataPath/RF/bus_selected_win_data[748] , 
        \DataPath/RF/bus_selected_win_data[747] , 
        \DataPath/RF/bus_selected_win_data[746] , 
        \DataPath/RF/bus_selected_win_data[745] , 
        \DataPath/RF/bus_selected_win_data[744] , 
        \DataPath/RF/bus_selected_win_data[743] , 
        \DataPath/RF/bus_selected_win_data[742] , 
        \DataPath/RF/bus_selected_win_data[741] , 
        \DataPath/RF/bus_selected_win_data[740] , 
        \DataPath/RF/bus_selected_win_data[739] , 
        \DataPath/RF/bus_selected_win_data[738] , 
        \DataPath/RF/bus_selected_win_data[737] , 
        \DataPath/RF/bus_selected_win_data[736] , 
        \DataPath/RF/bus_selected_win_data[735] , 
        \DataPath/RF/bus_selected_win_data[734] , 
        \DataPath/RF/bus_selected_win_data[733] , 
        \DataPath/RF/bus_selected_win_data[732] , 
        \DataPath/RF/bus_selected_win_data[731] , 
        \DataPath/RF/bus_selected_win_data[730] , 
        \DataPath/RF/bus_selected_win_data[729] , 
        \DataPath/RF/bus_selected_win_data[728] , 
        \DataPath/RF/bus_selected_win_data[727] , 
        \DataPath/RF/bus_selected_win_data[726] , 
        \DataPath/RF/bus_selected_win_data[725] , 
        \DataPath/RF/bus_selected_win_data[724] , 
        \DataPath/RF/bus_selected_win_data[723] , 
        \DataPath/RF/bus_selected_win_data[722] , 
        \DataPath/RF/bus_selected_win_data[721] , 
        \DataPath/RF/bus_selected_win_data[720] , 
        \DataPath/RF/bus_selected_win_data[719] , 
        \DataPath/RF/bus_selected_win_data[718] , 
        \DataPath/RF/bus_selected_win_data[717] , 
        \DataPath/RF/bus_selected_win_data[716] , 
        \DataPath/RF/bus_selected_win_data[715] , 
        \DataPath/RF/bus_selected_win_data[714] , 
        \DataPath/RF/bus_selected_win_data[713] , 
        \DataPath/RF/bus_selected_win_data[712] , 
        \DataPath/RF/bus_selected_win_data[711] , 
        \DataPath/RF/bus_selected_win_data[710] , 
        \DataPath/RF/bus_selected_win_data[709] , 
        \DataPath/RF/bus_selected_win_data[708] , 
        \DataPath/RF/bus_selected_win_data[707] , 
        \DataPath/RF/bus_selected_win_data[706] , 
        \DataPath/RF/bus_selected_win_data[705] , 
        \DataPath/RF/bus_selected_win_data[704] , 
        \DataPath/RF/bus_selected_win_data[703] , 
        \DataPath/RF/bus_selected_win_data[702] , 
        \DataPath/RF/bus_selected_win_data[701] , 
        \DataPath/RF/bus_selected_win_data[700] , 
        \DataPath/RF/bus_selected_win_data[699] , 
        \DataPath/RF/bus_selected_win_data[698] , 
        \DataPath/RF/bus_selected_win_data[697] , 
        \DataPath/RF/bus_selected_win_data[696] , 
        \DataPath/RF/bus_selected_win_data[695] , 
        \DataPath/RF/bus_selected_win_data[694] , 
        \DataPath/RF/bus_selected_win_data[693] , 
        \DataPath/RF/bus_selected_win_data[692] , 
        \DataPath/RF/bus_selected_win_data[691] , 
        \DataPath/RF/bus_selected_win_data[690] , 
        \DataPath/RF/bus_selected_win_data[689] , 
        \DataPath/RF/bus_selected_win_data[688] , 
        \DataPath/RF/bus_selected_win_data[687] , 
        \DataPath/RF/bus_selected_win_data[686] , 
        \DataPath/RF/bus_selected_win_data[685] , 
        \DataPath/RF/bus_selected_win_data[684] , 
        \DataPath/RF/bus_selected_win_data[683] , 
        \DataPath/RF/bus_selected_win_data[682] , 
        \DataPath/RF/bus_selected_win_data[681] , 
        \DataPath/RF/bus_selected_win_data[680] , 
        \DataPath/RF/bus_selected_win_data[679] , 
        \DataPath/RF/bus_selected_win_data[678] , 
        \DataPath/RF/bus_selected_win_data[677] , 
        \DataPath/RF/bus_selected_win_data[676] , 
        \DataPath/RF/bus_selected_win_data[675] , 
        \DataPath/RF/bus_selected_win_data[674] , 
        \DataPath/RF/bus_selected_win_data[673] , 
        \DataPath/RF/bus_selected_win_data[672] , 
        \DataPath/RF/bus_selected_win_data[671] , 
        \DataPath/RF/bus_selected_win_data[670] , 
        \DataPath/RF/bus_selected_win_data[669] , 
        \DataPath/RF/bus_selected_win_data[668] , 
        \DataPath/RF/bus_selected_win_data[667] , 
        \DataPath/RF/bus_selected_win_data[666] , 
        \DataPath/RF/bus_selected_win_data[665] , 
        \DataPath/RF/bus_selected_win_data[664] , 
        \DataPath/RF/bus_selected_win_data[663] , 
        \DataPath/RF/bus_selected_win_data[662] , 
        \DataPath/RF/bus_selected_win_data[661] , 
        \DataPath/RF/bus_selected_win_data[660] , 
        \DataPath/RF/bus_selected_win_data[659] , 
        \DataPath/RF/bus_selected_win_data[658] , 
        \DataPath/RF/bus_selected_win_data[657] , 
        \DataPath/RF/bus_selected_win_data[656] , 
        \DataPath/RF/bus_selected_win_data[655] , 
        \DataPath/RF/bus_selected_win_data[654] , 
        \DataPath/RF/bus_selected_win_data[653] , 
        \DataPath/RF/bus_selected_win_data[652] , 
        \DataPath/RF/bus_selected_win_data[651] , 
        \DataPath/RF/bus_selected_win_data[650] , 
        \DataPath/RF/bus_selected_win_data[649] , 
        \DataPath/RF/bus_selected_win_data[648] , 
        \DataPath/RF/bus_selected_win_data[647] , 
        \DataPath/RF/bus_selected_win_data[646] , 
        \DataPath/RF/bus_selected_win_data[645] , 
        \DataPath/RF/bus_selected_win_data[644] , 
        \DataPath/RF/bus_selected_win_data[643] , 
        \DataPath/RF/bus_selected_win_data[642] , 
        \DataPath/RF/bus_selected_win_data[641] , 
        \DataPath/RF/bus_selected_win_data[640] , 
        \DataPath/RF/bus_selected_win_data[639] , 
        \DataPath/RF/bus_selected_win_data[638] , 
        \DataPath/RF/bus_selected_win_data[637] , 
        \DataPath/RF/bus_selected_win_data[636] , 
        \DataPath/RF/bus_selected_win_data[635] , 
        \DataPath/RF/bus_selected_win_data[634] , 
        \DataPath/RF/bus_selected_win_data[633] , 
        \DataPath/RF/bus_selected_win_data[632] , 
        \DataPath/RF/bus_selected_win_data[631] , 
        \DataPath/RF/bus_selected_win_data[630] , 
        \DataPath/RF/bus_selected_win_data[629] , 
        \DataPath/RF/bus_selected_win_data[628] , 
        \DataPath/RF/bus_selected_win_data[627] , 
        \DataPath/RF/bus_selected_win_data[626] , 
        \DataPath/RF/bus_selected_win_data[625] , 
        \DataPath/RF/bus_selected_win_data[624] , 
        \DataPath/RF/bus_selected_win_data[623] , 
        \DataPath/RF/bus_selected_win_data[622] , 
        \DataPath/RF/bus_selected_win_data[621] , 
        \DataPath/RF/bus_selected_win_data[620] , 
        \DataPath/RF/bus_selected_win_data[619] , 
        \DataPath/RF/bus_selected_win_data[618] , 
        \DataPath/RF/bus_selected_win_data[617] , 
        \DataPath/RF/bus_selected_win_data[616] , 
        \DataPath/RF/bus_selected_win_data[615] , 
        \DataPath/RF/bus_selected_win_data[614] , 
        \DataPath/RF/bus_selected_win_data[613] , 
        \DataPath/RF/bus_selected_win_data[612] , 
        \DataPath/RF/bus_selected_win_data[611] , 
        \DataPath/RF/bus_selected_win_data[610] , 
        \DataPath/RF/bus_selected_win_data[609] , 
        \DataPath/RF/bus_selected_win_data[608] , 
        \DataPath/RF/bus_selected_win_data[607] , 
        \DataPath/RF/bus_selected_win_data[606] , 
        \DataPath/RF/bus_selected_win_data[605] , 
        \DataPath/RF/bus_selected_win_data[604] , 
        \DataPath/RF/bus_selected_win_data[603] , 
        \DataPath/RF/bus_selected_win_data[602] , 
        \DataPath/RF/bus_selected_win_data[601] , 
        \DataPath/RF/bus_selected_win_data[600] , 
        \DataPath/RF/bus_selected_win_data[599] , 
        \DataPath/RF/bus_selected_win_data[598] , 
        \DataPath/RF/bus_selected_win_data[597] , 
        \DataPath/RF/bus_selected_win_data[596] , 
        \DataPath/RF/bus_selected_win_data[595] , 
        \DataPath/RF/bus_selected_win_data[594] , 
        \DataPath/RF/bus_selected_win_data[593] , 
        \DataPath/RF/bus_selected_win_data[592] , 
        \DataPath/RF/bus_selected_win_data[591] , 
        \DataPath/RF/bus_selected_win_data[590] , 
        \DataPath/RF/bus_selected_win_data[589] , 
        \DataPath/RF/bus_selected_win_data[588] , 
        \DataPath/RF/bus_selected_win_data[587] , 
        \DataPath/RF/bus_selected_win_data[586] , 
        \DataPath/RF/bus_selected_win_data[585] , 
        \DataPath/RF/bus_selected_win_data[584] , 
        \DataPath/RF/bus_selected_win_data[583] , 
        \DataPath/RF/bus_selected_win_data[582] , 
        \DataPath/RF/bus_selected_win_data[581] , 
        \DataPath/RF/bus_selected_win_data[580] , 
        \DataPath/RF/bus_selected_win_data[579] , 
        \DataPath/RF/bus_selected_win_data[578] , 
        \DataPath/RF/bus_selected_win_data[577] , 
        \DataPath/RF/bus_selected_win_data[576] , 
        \DataPath/RF/bus_selected_win_data[575] , 
        \DataPath/RF/bus_selected_win_data[574] , 
        \DataPath/RF/bus_selected_win_data[573] , 
        \DataPath/RF/bus_selected_win_data[572] , 
        \DataPath/RF/bus_selected_win_data[571] , 
        \DataPath/RF/bus_selected_win_data[570] , 
        \DataPath/RF/bus_selected_win_data[569] , 
        \DataPath/RF/bus_selected_win_data[568] , 
        \DataPath/RF/bus_selected_win_data[567] , 
        \DataPath/RF/bus_selected_win_data[566] , 
        \DataPath/RF/bus_selected_win_data[565] , 
        \DataPath/RF/bus_selected_win_data[564] , 
        \DataPath/RF/bus_selected_win_data[563] , 
        \DataPath/RF/bus_selected_win_data[562] , 
        \DataPath/RF/bus_selected_win_data[561] , 
        \DataPath/RF/bus_selected_win_data[560] , 
        \DataPath/RF/bus_selected_win_data[559] , 
        \DataPath/RF/bus_selected_win_data[558] , 
        \DataPath/RF/bus_selected_win_data[557] , 
        \DataPath/RF/bus_selected_win_data[556] , 
        \DataPath/RF/bus_selected_win_data[555] , 
        \DataPath/RF/bus_selected_win_data[554] , 
        \DataPath/RF/bus_selected_win_data[553] , 
        \DataPath/RF/bus_selected_win_data[552] , 
        \DataPath/RF/bus_selected_win_data[551] , 
        \DataPath/RF/bus_selected_win_data[550] , 
        \DataPath/RF/bus_selected_win_data[549] , 
        \DataPath/RF/bus_selected_win_data[548] , 
        \DataPath/RF/bus_selected_win_data[547] , 
        \DataPath/RF/bus_selected_win_data[546] , 
        \DataPath/RF/bus_selected_win_data[545] , 
        \DataPath/RF/bus_selected_win_data[544] , 
        \DataPath/RF/bus_selected_win_data[543] , 
        \DataPath/RF/bus_selected_win_data[542] , 
        \DataPath/RF/bus_selected_win_data[541] , 
        \DataPath/RF/bus_selected_win_data[540] , 
        \DataPath/RF/bus_selected_win_data[539] , 
        \DataPath/RF/bus_selected_win_data[538] , 
        \DataPath/RF/bus_selected_win_data[537] , 
        \DataPath/RF/bus_selected_win_data[536] , 
        \DataPath/RF/bus_selected_win_data[535] , 
        \DataPath/RF/bus_selected_win_data[534] , 
        \DataPath/RF/bus_selected_win_data[533] , 
        \DataPath/RF/bus_selected_win_data[532] , 
        \DataPath/RF/bus_selected_win_data[531] , 
        \DataPath/RF/bus_selected_win_data[530] , 
        \DataPath/RF/bus_selected_win_data[529] , 
        \DataPath/RF/bus_selected_win_data[528] , 
        \DataPath/RF/bus_selected_win_data[527] , 
        \DataPath/RF/bus_selected_win_data[526] , 
        \DataPath/RF/bus_selected_win_data[525] , 
        \DataPath/RF/bus_selected_win_data[524] , 
        \DataPath/RF/bus_selected_win_data[523] , 
        \DataPath/RF/bus_selected_win_data[522] , 
        \DataPath/RF/bus_selected_win_data[521] , 
        \DataPath/RF/bus_selected_win_data[520] , 
        \DataPath/RF/bus_selected_win_data[519] , 
        \DataPath/RF/bus_selected_win_data[518] , 
        \DataPath/RF/bus_selected_win_data[517] , 
        \DataPath/RF/bus_selected_win_data[516] , 
        \DataPath/RF/bus_selected_win_data[515] , 
        \DataPath/RF/bus_selected_win_data[514] , 
        \DataPath/RF/bus_selected_win_data[513] , 
        \DataPath/RF/bus_selected_win_data[512] , 
        \DataPath/RF/bus_selected_win_data[511] , 
        \DataPath/RF/bus_selected_win_data[510] , 
        \DataPath/RF/bus_selected_win_data[509] , 
        \DataPath/RF/bus_selected_win_data[508] , 
        \DataPath/RF/bus_selected_win_data[507] , 
        \DataPath/RF/bus_selected_win_data[506] , 
        \DataPath/RF/bus_selected_win_data[505] , 
        \DataPath/RF/bus_selected_win_data[504] , 
        \DataPath/RF/bus_selected_win_data[503] , 
        \DataPath/RF/bus_selected_win_data[502] , 
        \DataPath/RF/bus_selected_win_data[501] , 
        \DataPath/RF/bus_selected_win_data[500] , 
        \DataPath/RF/bus_selected_win_data[499] , 
        \DataPath/RF/bus_selected_win_data[498] , 
        \DataPath/RF/bus_selected_win_data[497] , 
        \DataPath/RF/bus_selected_win_data[496] , 
        \DataPath/RF/bus_selected_win_data[495] , 
        \DataPath/RF/bus_selected_win_data[494] , 
        \DataPath/RF/bus_selected_win_data[493] , 
        \DataPath/RF/bus_selected_win_data[492] , 
        \DataPath/RF/bus_selected_win_data[491] , 
        \DataPath/RF/bus_selected_win_data[490] , 
        \DataPath/RF/bus_selected_win_data[489] , 
        \DataPath/RF/bus_selected_win_data[488] , 
        \DataPath/RF/bus_selected_win_data[487] , 
        \DataPath/RF/bus_selected_win_data[486] , 
        \DataPath/RF/bus_selected_win_data[485] , 
        \DataPath/RF/bus_selected_win_data[484] , 
        \DataPath/RF/bus_selected_win_data[483] , 
        \DataPath/RF/bus_selected_win_data[482] , 
        \DataPath/RF/bus_selected_win_data[481] , 
        \DataPath/RF/bus_selected_win_data[480] , 
        \DataPath/RF/bus_selected_win_data[479] , 
        \DataPath/RF/bus_selected_win_data[478] , 
        \DataPath/RF/bus_selected_win_data[477] , 
        \DataPath/RF/bus_selected_win_data[476] , 
        \DataPath/RF/bus_selected_win_data[475] , 
        \DataPath/RF/bus_selected_win_data[474] , 
        \DataPath/RF/bus_selected_win_data[473] , 
        \DataPath/RF/bus_selected_win_data[472] , 
        \DataPath/RF/bus_selected_win_data[471] , 
        \DataPath/RF/bus_selected_win_data[470] , 
        \DataPath/RF/bus_selected_win_data[469] , 
        \DataPath/RF/bus_selected_win_data[468] , 
        \DataPath/RF/bus_selected_win_data[467] , 
        \DataPath/RF/bus_selected_win_data[466] , 
        \DataPath/RF/bus_selected_win_data[465] , 
        \DataPath/RF/bus_selected_win_data[464] , 
        \DataPath/RF/bus_selected_win_data[463] , 
        \DataPath/RF/bus_selected_win_data[462] , 
        \DataPath/RF/bus_selected_win_data[461] , 
        \DataPath/RF/bus_selected_win_data[460] , 
        \DataPath/RF/bus_selected_win_data[459] , 
        \DataPath/RF/bus_selected_win_data[458] , 
        \DataPath/RF/bus_selected_win_data[457] , 
        \DataPath/RF/bus_selected_win_data[456] , 
        \DataPath/RF/bus_selected_win_data[455] , 
        \DataPath/RF/bus_selected_win_data[454] , 
        \DataPath/RF/bus_selected_win_data[453] , 
        \DataPath/RF/bus_selected_win_data[452] , 
        \DataPath/RF/bus_selected_win_data[451] , 
        \DataPath/RF/bus_selected_win_data[450] , 
        \DataPath/RF/bus_selected_win_data[449] , 
        \DataPath/RF/bus_selected_win_data[448] , 
        \DataPath/RF/bus_selected_win_data[447] , 
        \DataPath/RF/bus_selected_win_data[446] , 
        \DataPath/RF/bus_selected_win_data[445] , 
        \DataPath/RF/bus_selected_win_data[444] , 
        \DataPath/RF/bus_selected_win_data[443] , 
        \DataPath/RF/bus_selected_win_data[442] , 
        \DataPath/RF/bus_selected_win_data[441] , 
        \DataPath/RF/bus_selected_win_data[440] , 
        \DataPath/RF/bus_selected_win_data[439] , 
        \DataPath/RF/bus_selected_win_data[438] , 
        \DataPath/RF/bus_selected_win_data[437] , 
        \DataPath/RF/bus_selected_win_data[436] , 
        \DataPath/RF/bus_selected_win_data[435] , 
        \DataPath/RF/bus_selected_win_data[434] , 
        \DataPath/RF/bus_selected_win_data[433] , 
        \DataPath/RF/bus_selected_win_data[432] , 
        \DataPath/RF/bus_selected_win_data[431] , 
        \DataPath/RF/bus_selected_win_data[430] , 
        \DataPath/RF/bus_selected_win_data[429] , 
        \DataPath/RF/bus_selected_win_data[428] , 
        \DataPath/RF/bus_selected_win_data[427] , 
        \DataPath/RF/bus_selected_win_data[426] , 
        \DataPath/RF/bus_selected_win_data[425] , 
        \DataPath/RF/bus_selected_win_data[424] , 
        \DataPath/RF/bus_selected_win_data[423] , 
        \DataPath/RF/bus_selected_win_data[422] , 
        \DataPath/RF/bus_selected_win_data[421] , 
        \DataPath/RF/bus_selected_win_data[420] , 
        \DataPath/RF/bus_selected_win_data[419] , 
        \DataPath/RF/bus_selected_win_data[418] , 
        \DataPath/RF/bus_selected_win_data[417] , 
        \DataPath/RF/bus_selected_win_data[416] , 
        \DataPath/RF/bus_selected_win_data[415] , 
        \DataPath/RF/bus_selected_win_data[414] , 
        \DataPath/RF/bus_selected_win_data[413] , 
        \DataPath/RF/bus_selected_win_data[412] , 
        \DataPath/RF/bus_selected_win_data[411] , 
        \DataPath/RF/bus_selected_win_data[410] , 
        \DataPath/RF/bus_selected_win_data[409] , 
        \DataPath/RF/bus_selected_win_data[408] , 
        \DataPath/RF/bus_selected_win_data[407] , 
        \DataPath/RF/bus_selected_win_data[406] , 
        \DataPath/RF/bus_selected_win_data[405] , 
        \DataPath/RF/bus_selected_win_data[404] , 
        \DataPath/RF/bus_selected_win_data[403] , 
        \DataPath/RF/bus_selected_win_data[402] , 
        \DataPath/RF/bus_selected_win_data[401] , 
        \DataPath/RF/bus_selected_win_data[400] , 
        \DataPath/RF/bus_selected_win_data[399] , 
        \DataPath/RF/bus_selected_win_data[398] , 
        \DataPath/RF/bus_selected_win_data[397] , 
        \DataPath/RF/bus_selected_win_data[396] , 
        \DataPath/RF/bus_selected_win_data[395] , 
        \DataPath/RF/bus_selected_win_data[394] , 
        \DataPath/RF/bus_selected_win_data[393] , 
        \DataPath/RF/bus_selected_win_data[392] , 
        \DataPath/RF/bus_selected_win_data[391] , 
        \DataPath/RF/bus_selected_win_data[390] , 
        \DataPath/RF/bus_selected_win_data[389] , 
        \DataPath/RF/bus_selected_win_data[388] , 
        \DataPath/RF/bus_selected_win_data[387] , 
        \DataPath/RF/bus_selected_win_data[386] , 
        \DataPath/RF/bus_selected_win_data[385] , 
        \DataPath/RF/bus_selected_win_data[384] , 
        \DataPath/RF/bus_selected_win_data[383] , 
        \DataPath/RF/bus_selected_win_data[382] , 
        \DataPath/RF/bus_selected_win_data[381] , 
        \DataPath/RF/bus_selected_win_data[380] , 
        \DataPath/RF/bus_selected_win_data[379] , 
        \DataPath/RF/bus_selected_win_data[378] , 
        \DataPath/RF/bus_selected_win_data[377] , 
        \DataPath/RF/bus_selected_win_data[376] , 
        \DataPath/RF/bus_selected_win_data[375] , 
        \DataPath/RF/bus_selected_win_data[374] , 
        \DataPath/RF/bus_selected_win_data[373] , 
        \DataPath/RF/bus_selected_win_data[372] , 
        \DataPath/RF/bus_selected_win_data[371] , 
        \DataPath/RF/bus_selected_win_data[370] , 
        \DataPath/RF/bus_selected_win_data[369] , 
        \DataPath/RF/bus_selected_win_data[368] , 
        \DataPath/RF/bus_selected_win_data[367] , 
        \DataPath/RF/bus_selected_win_data[366] , 
        \DataPath/RF/bus_selected_win_data[365] , 
        \DataPath/RF/bus_selected_win_data[364] , 
        \DataPath/RF/bus_selected_win_data[363] , 
        \DataPath/RF/bus_selected_win_data[362] , 
        \DataPath/RF/bus_selected_win_data[361] , 
        \DataPath/RF/bus_selected_win_data[360] , 
        \DataPath/RF/bus_selected_win_data[359] , 
        \DataPath/RF/bus_selected_win_data[358] , 
        \DataPath/RF/bus_selected_win_data[357] , 
        \DataPath/RF/bus_selected_win_data[356] , 
        \DataPath/RF/bus_selected_win_data[355] , 
        \DataPath/RF/bus_selected_win_data[354] , 
        \DataPath/RF/bus_selected_win_data[353] , 
        \DataPath/RF/bus_selected_win_data[352] , 
        \DataPath/RF/bus_selected_win_data[351] , 
        \DataPath/RF/bus_selected_win_data[350] , 
        \DataPath/RF/bus_selected_win_data[349] , 
        \DataPath/RF/bus_selected_win_data[348] , 
        \DataPath/RF/bus_selected_win_data[347] , 
        \DataPath/RF/bus_selected_win_data[346] , 
        \DataPath/RF/bus_selected_win_data[345] , 
        \DataPath/RF/bus_selected_win_data[344] , 
        \DataPath/RF/bus_selected_win_data[343] , 
        \DataPath/RF/bus_selected_win_data[342] , 
        \DataPath/RF/bus_selected_win_data[341] , 
        \DataPath/RF/bus_selected_win_data[340] , 
        \DataPath/RF/bus_selected_win_data[339] , 
        \DataPath/RF/bus_selected_win_data[338] , 
        \DataPath/RF/bus_selected_win_data[337] , 
        \DataPath/RF/bus_selected_win_data[336] , 
        \DataPath/RF/bus_selected_win_data[335] , 
        \DataPath/RF/bus_selected_win_data[334] , 
        \DataPath/RF/bus_selected_win_data[333] , 
        \DataPath/RF/bus_selected_win_data[332] , 
        \DataPath/RF/bus_selected_win_data[331] , 
        \DataPath/RF/bus_selected_win_data[330] , 
        \DataPath/RF/bus_selected_win_data[329] , 
        \DataPath/RF/bus_selected_win_data[328] , 
        \DataPath/RF/bus_selected_win_data[327] , 
        \DataPath/RF/bus_selected_win_data[326] , 
        \DataPath/RF/bus_selected_win_data[325] , 
        \DataPath/RF/bus_selected_win_data[324] , 
        \DataPath/RF/bus_selected_win_data[323] , 
        \DataPath/RF/bus_selected_win_data[322] , 
        \DataPath/RF/bus_selected_win_data[321] , 
        \DataPath/RF/bus_selected_win_data[320] , 
        \DataPath/RF/bus_selected_win_data[319] , 
        \DataPath/RF/bus_selected_win_data[318] , 
        \DataPath/RF/bus_selected_win_data[317] , 
        \DataPath/RF/bus_selected_win_data[316] , 
        \DataPath/RF/bus_selected_win_data[315] , 
        \DataPath/RF/bus_selected_win_data[314] , 
        \DataPath/RF/bus_selected_win_data[313] , 
        \DataPath/RF/bus_selected_win_data[312] , 
        \DataPath/RF/bus_selected_win_data[311] , 
        \DataPath/RF/bus_selected_win_data[310] , 
        \DataPath/RF/bus_selected_win_data[309] , 
        \DataPath/RF/bus_selected_win_data[308] , 
        \DataPath/RF/bus_selected_win_data[307] , 
        \DataPath/RF/bus_selected_win_data[306] , 
        \DataPath/RF/bus_selected_win_data[305] , 
        \DataPath/RF/bus_selected_win_data[304] , 
        \DataPath/RF/bus_selected_win_data[303] , 
        \DataPath/RF/bus_selected_win_data[302] , 
        \DataPath/RF/bus_selected_win_data[301] , 
        \DataPath/RF/bus_selected_win_data[300] , 
        \DataPath/RF/bus_selected_win_data[299] , 
        \DataPath/RF/bus_selected_win_data[298] , 
        \DataPath/RF/bus_selected_win_data[297] , 
        \DataPath/RF/bus_selected_win_data[296] , 
        \DataPath/RF/bus_selected_win_data[295] , 
        \DataPath/RF/bus_selected_win_data[294] , 
        \DataPath/RF/bus_selected_win_data[293] , 
        \DataPath/RF/bus_selected_win_data[292] , 
        \DataPath/RF/bus_selected_win_data[291] , 
        \DataPath/RF/bus_selected_win_data[290] , 
        \DataPath/RF/bus_selected_win_data[289] , 
        \DataPath/RF/bus_selected_win_data[288] , 
        \DataPath/RF/bus_selected_win_data[287] , 
        \DataPath/RF/bus_selected_win_data[286] , 
        \DataPath/RF/bus_selected_win_data[285] , 
        \DataPath/RF/bus_selected_win_data[284] , 
        \DataPath/RF/bus_selected_win_data[283] , 
        \DataPath/RF/bus_selected_win_data[282] , 
        \DataPath/RF/bus_selected_win_data[281] , 
        \DataPath/RF/bus_selected_win_data[280] , 
        \DataPath/RF/bus_selected_win_data[279] , 
        \DataPath/RF/bus_selected_win_data[278] , 
        \DataPath/RF/bus_selected_win_data[277] , 
        \DataPath/RF/bus_selected_win_data[276] , 
        \DataPath/RF/bus_selected_win_data[275] , 
        \DataPath/RF/bus_selected_win_data[274] , 
        \DataPath/RF/bus_selected_win_data[273] , 
        \DataPath/RF/bus_selected_win_data[272] , 
        \DataPath/RF/bus_selected_win_data[271] , 
        \DataPath/RF/bus_selected_win_data[270] , 
        \DataPath/RF/bus_selected_win_data[269] , 
        \DataPath/RF/bus_selected_win_data[268] , 
        \DataPath/RF/bus_selected_win_data[267] , 
        \DataPath/RF/bus_selected_win_data[266] , 
        \DataPath/RF/bus_selected_win_data[265] , 
        \DataPath/RF/bus_selected_win_data[264] , 
        \DataPath/RF/bus_selected_win_data[263] , 
        \DataPath/RF/bus_selected_win_data[262] , 
        \DataPath/RF/bus_selected_win_data[261] , 
        \DataPath/RF/bus_selected_win_data[260] , 
        \DataPath/RF/bus_selected_win_data[259] , 
        \DataPath/RF/bus_selected_win_data[258] , 
        \DataPath/RF/bus_selected_win_data[257] , 
        \DataPath/RF/bus_selected_win_data[256] , 
        \DataPath/RF/bus_selected_win_data[255] , 
        \DataPath/RF/bus_selected_win_data[254] , 
        \DataPath/RF/bus_selected_win_data[253] , 
        \DataPath/RF/bus_selected_win_data[252] , 
        \DataPath/RF/bus_selected_win_data[251] , 
        \DataPath/RF/bus_selected_win_data[250] , 
        \DataPath/RF/bus_selected_win_data[249] , 
        \DataPath/RF/bus_selected_win_data[248] , 
        \DataPath/RF/bus_selected_win_data[247] , 
        \DataPath/RF/bus_selected_win_data[246] , 
        \DataPath/RF/bus_selected_win_data[245] , 
        \DataPath/RF/bus_selected_win_data[244] , 
        \DataPath/RF/bus_selected_win_data[243] , 
        \DataPath/RF/bus_selected_win_data[242] , 
        \DataPath/RF/bus_selected_win_data[241] , 
        \DataPath/RF/bus_selected_win_data[240] , 
        \DataPath/RF/bus_selected_win_data[239] , 
        \DataPath/RF/bus_selected_win_data[238] , 
        \DataPath/RF/bus_selected_win_data[237] , 
        \DataPath/RF/bus_selected_win_data[236] , 
        \DataPath/RF/bus_selected_win_data[235] , 
        \DataPath/RF/bus_selected_win_data[234] , 
        \DataPath/RF/bus_selected_win_data[233] , 
        \DataPath/RF/bus_selected_win_data[232] , 
        \DataPath/RF/bus_selected_win_data[231] , 
        \DataPath/RF/bus_selected_win_data[230] , 
        \DataPath/RF/bus_selected_win_data[229] , 
        \DataPath/RF/bus_selected_win_data[228] , 
        \DataPath/RF/bus_selected_win_data[227] , 
        \DataPath/RF/bus_selected_win_data[226] , 
        \DataPath/RF/bus_selected_win_data[225] , 
        \DataPath/RF/bus_selected_win_data[224] , 
        \DataPath/RF/bus_selected_win_data[223] , 
        \DataPath/RF/bus_selected_win_data[222] , 
        \DataPath/RF/bus_selected_win_data[221] , 
        \DataPath/RF/bus_selected_win_data[220] , 
        \DataPath/RF/bus_selected_win_data[219] , 
        \DataPath/RF/bus_selected_win_data[218] , 
        \DataPath/RF/bus_selected_win_data[217] , 
        \DataPath/RF/bus_selected_win_data[216] , 
        \DataPath/RF/bus_selected_win_data[215] , 
        \DataPath/RF/bus_selected_win_data[214] , 
        \DataPath/RF/bus_selected_win_data[213] , 
        \DataPath/RF/bus_selected_win_data[212] , 
        \DataPath/RF/bus_selected_win_data[211] , 
        \DataPath/RF/bus_selected_win_data[210] , 
        \DataPath/RF/bus_selected_win_data[209] , 
        \DataPath/RF/bus_selected_win_data[208] , 
        \DataPath/RF/bus_selected_win_data[207] , 
        \DataPath/RF/bus_selected_win_data[206] , 
        \DataPath/RF/bus_selected_win_data[205] , 
        \DataPath/RF/bus_selected_win_data[204] , 
        \DataPath/RF/bus_selected_win_data[203] , 
        \DataPath/RF/bus_selected_win_data[202] , 
        \DataPath/RF/bus_selected_win_data[201] , 
        \DataPath/RF/bus_selected_win_data[200] , 
        \DataPath/RF/bus_selected_win_data[199] , 
        \DataPath/RF/bus_selected_win_data[198] , 
        \DataPath/RF/bus_selected_win_data[197] , 
        \DataPath/RF/bus_selected_win_data[196] , 
        \DataPath/RF/bus_selected_win_data[195] , 
        \DataPath/RF/bus_selected_win_data[194] , 
        \DataPath/RF/bus_selected_win_data[193] , 
        \DataPath/RF/bus_selected_win_data[192] , 
        \DataPath/RF/bus_selected_win_data[191] , 
        \DataPath/RF/bus_selected_win_data[190] , 
        \DataPath/RF/bus_selected_win_data[189] , 
        \DataPath/RF/bus_selected_win_data[188] , 
        \DataPath/RF/bus_selected_win_data[187] , 
        \DataPath/RF/bus_selected_win_data[186] , 
        \DataPath/RF/bus_selected_win_data[185] , 
        \DataPath/RF/bus_selected_win_data[184] , 
        \DataPath/RF/bus_selected_win_data[183] , 
        \DataPath/RF/bus_selected_win_data[182] , 
        \DataPath/RF/bus_selected_win_data[181] , 
        \DataPath/RF/bus_selected_win_data[180] , 
        \DataPath/RF/bus_selected_win_data[179] , 
        \DataPath/RF/bus_selected_win_data[178] , 
        \DataPath/RF/bus_selected_win_data[177] , 
        \DataPath/RF/bus_selected_win_data[176] , 
        \DataPath/RF/bus_selected_win_data[175] , 
        \DataPath/RF/bus_selected_win_data[174] , 
        \DataPath/RF/bus_selected_win_data[173] , 
        \DataPath/RF/bus_selected_win_data[172] , 
        \DataPath/RF/bus_selected_win_data[171] , 
        \DataPath/RF/bus_selected_win_data[170] , 
        \DataPath/RF/bus_selected_win_data[169] , 
        \DataPath/RF/bus_selected_win_data[168] , 
        \DataPath/RF/bus_selected_win_data[167] , 
        \DataPath/RF/bus_selected_win_data[166] , 
        \DataPath/RF/bus_selected_win_data[165] , 
        \DataPath/RF/bus_selected_win_data[164] , 
        \DataPath/RF/bus_selected_win_data[163] , 
        \DataPath/RF/bus_selected_win_data[162] , 
        \DataPath/RF/bus_selected_win_data[161] , 
        \DataPath/RF/bus_selected_win_data[160] , 
        \DataPath/RF/bus_selected_win_data[159] , 
        \DataPath/RF/bus_selected_win_data[158] , 
        \DataPath/RF/bus_selected_win_data[157] , 
        \DataPath/RF/bus_selected_win_data[156] , 
        \DataPath/RF/bus_selected_win_data[155] , 
        \DataPath/RF/bus_selected_win_data[154] , 
        \DataPath/RF/bus_selected_win_data[153] , 
        \DataPath/RF/bus_selected_win_data[152] , 
        \DataPath/RF/bus_selected_win_data[151] , 
        \DataPath/RF/bus_selected_win_data[150] , 
        \DataPath/RF/bus_selected_win_data[149] , 
        \DataPath/RF/bus_selected_win_data[148] , 
        \DataPath/RF/bus_selected_win_data[147] , 
        \DataPath/RF/bus_selected_win_data[146] , 
        \DataPath/RF/bus_selected_win_data[145] , 
        \DataPath/RF/bus_selected_win_data[144] , 
        \DataPath/RF/bus_selected_win_data[143] , 
        \DataPath/RF/bus_selected_win_data[142] , 
        \DataPath/RF/bus_selected_win_data[141] , 
        \DataPath/RF/bus_selected_win_data[140] , 
        \DataPath/RF/bus_selected_win_data[139] , 
        \DataPath/RF/bus_selected_win_data[138] , 
        \DataPath/RF/bus_selected_win_data[137] , 
        \DataPath/RF/bus_selected_win_data[136] , 
        \DataPath/RF/bus_selected_win_data[135] , 
        \DataPath/RF/bus_selected_win_data[134] , 
        \DataPath/RF/bus_selected_win_data[133] , 
        \DataPath/RF/bus_selected_win_data[132] , 
        \DataPath/RF/bus_selected_win_data[131] , 
        \DataPath/RF/bus_selected_win_data[130] , 
        \DataPath/RF/bus_selected_win_data[129] , 
        \DataPath/RF/bus_selected_win_data[128] , 
        \DataPath/RF/bus_selected_win_data[127] , 
        \DataPath/RF/bus_selected_win_data[126] , 
        \DataPath/RF/bus_selected_win_data[125] , 
        \DataPath/RF/bus_selected_win_data[124] , 
        \DataPath/RF/bus_selected_win_data[123] , 
        \DataPath/RF/bus_selected_win_data[122] , 
        \DataPath/RF/bus_selected_win_data[121] , 
        \DataPath/RF/bus_selected_win_data[120] , 
        \DataPath/RF/bus_selected_win_data[119] , 
        \DataPath/RF/bus_selected_win_data[118] , 
        \DataPath/RF/bus_selected_win_data[117] , 
        \DataPath/RF/bus_selected_win_data[116] , 
        \DataPath/RF/bus_selected_win_data[115] , 
        \DataPath/RF/bus_selected_win_data[114] , 
        \DataPath/RF/bus_selected_win_data[113] , 
        \DataPath/RF/bus_selected_win_data[112] , 
        \DataPath/RF/bus_selected_win_data[111] , 
        \DataPath/RF/bus_selected_win_data[110] , 
        \DataPath/RF/bus_selected_win_data[109] , 
        \DataPath/RF/bus_selected_win_data[108] , 
        \DataPath/RF/bus_selected_win_data[107] , 
        \DataPath/RF/bus_selected_win_data[106] , 
        \DataPath/RF/bus_selected_win_data[105] , 
        \DataPath/RF/bus_selected_win_data[104] , 
        \DataPath/RF/bus_selected_win_data[103] , 
        \DataPath/RF/bus_selected_win_data[102] , 
        \DataPath/RF/bus_selected_win_data[101] , 
        \DataPath/RF/bus_selected_win_data[100] , 
        \DataPath/RF/bus_selected_win_data[99] , 
        \DataPath/RF/bus_selected_win_data[98] , 
        \DataPath/RF/bus_selected_win_data[97] , 
        \DataPath/RF/bus_selected_win_data[96] , 
        \DataPath/RF/bus_selected_win_data[95] , 
        \DataPath/RF/bus_selected_win_data[94] , 
        \DataPath/RF/bus_selected_win_data[93] , 
        \DataPath/RF/bus_selected_win_data[92] , 
        \DataPath/RF/bus_selected_win_data[91] , 
        \DataPath/RF/bus_selected_win_data[90] , 
        \DataPath/RF/bus_selected_win_data[89] , 
        \DataPath/RF/bus_selected_win_data[88] , 
        \DataPath/RF/bus_selected_win_data[87] , 
        \DataPath/RF/bus_selected_win_data[86] , 
        \DataPath/RF/bus_selected_win_data[85] , 
        \DataPath/RF/bus_selected_win_data[84] , 
        \DataPath/RF/bus_selected_win_data[83] , 
        \DataPath/RF/bus_selected_win_data[82] , 
        \DataPath/RF/bus_selected_win_data[81] , 
        \DataPath/RF/bus_selected_win_data[80] , 
        \DataPath/RF/bus_selected_win_data[79] , 
        \DataPath/RF/bus_selected_win_data[78] , 
        \DataPath/RF/bus_selected_win_data[77] , 
        \DataPath/RF/bus_selected_win_data[76] , 
        \DataPath/RF/bus_selected_win_data[75] , 
        \DataPath/RF/bus_selected_win_data[74] , 
        \DataPath/RF/bus_selected_win_data[73] , 
        \DataPath/RF/bus_selected_win_data[72] , 
        \DataPath/RF/bus_selected_win_data[71] , 
        \DataPath/RF/bus_selected_win_data[70] , 
        \DataPath/RF/bus_selected_win_data[69] , 
        \DataPath/RF/bus_selected_win_data[68] , 
        \DataPath/RF/bus_selected_win_data[67] , 
        \DataPath/RF/bus_selected_win_data[66] , 
        \DataPath/RF/bus_selected_win_data[65] , 
        \DataPath/RF/bus_selected_win_data[64] , 
        \DataPath/RF/bus_selected_win_data[63] , 
        \DataPath/RF/bus_selected_win_data[62] , 
        \DataPath/RF/bus_selected_win_data[61] , 
        \DataPath/RF/bus_selected_win_data[60] , 
        \DataPath/RF/bus_selected_win_data[59] , 
        \DataPath/RF/bus_selected_win_data[58] , 
        \DataPath/RF/bus_selected_win_data[57] , 
        \DataPath/RF/bus_selected_win_data[56] , 
        \DataPath/RF/bus_selected_win_data[55] , 
        \DataPath/RF/bus_selected_win_data[54] , 
        \DataPath/RF/bus_selected_win_data[53] , 
        \DataPath/RF/bus_selected_win_data[52] , 
        \DataPath/RF/bus_selected_win_data[51] , 
        \DataPath/RF/bus_selected_win_data[50] , 
        \DataPath/RF/bus_selected_win_data[49] , 
        \DataPath/RF/bus_selected_win_data[48] , 
        \DataPath/RF/bus_selected_win_data[47] , 
        \DataPath/RF/bus_selected_win_data[46] , 
        \DataPath/RF/bus_selected_win_data[45] , 
        \DataPath/RF/bus_selected_win_data[44] , 
        \DataPath/RF/bus_selected_win_data[43] , 
        \DataPath/RF/bus_selected_win_data[42] , 
        \DataPath/RF/bus_selected_win_data[41] , 
        \DataPath/RF/bus_selected_win_data[40] , 
        \DataPath/RF/bus_selected_win_data[39] , 
        \DataPath/RF/bus_selected_win_data[38] , 
        \DataPath/RF/bus_selected_win_data[37] , 
        \DataPath/RF/bus_selected_win_data[36] , 
        \DataPath/RF/bus_selected_win_data[35] , 
        \DataPath/RF/bus_selected_win_data[34] , 
        \DataPath/RF/bus_selected_win_data[33] , 
        \DataPath/RF/bus_selected_win_data[32] , 
        \DataPath/RF/bus_selected_win_data[31] , 
        \DataPath/RF/bus_selected_win_data[30] , 
        \DataPath/RF/bus_selected_win_data[29] , 
        \DataPath/RF/bus_selected_win_data[28] , 
        \DataPath/RF/bus_selected_win_data[27] , 
        \DataPath/RF/bus_selected_win_data[26] , 
        \DataPath/RF/bus_selected_win_data[25] , 
        \DataPath/RF/bus_selected_win_data[24] , 
        \DataPath/RF/bus_selected_win_data[23] , 
        \DataPath/RF/bus_selected_win_data[22] , 
        \DataPath/RF/bus_selected_win_data[21] , 
        \DataPath/RF/bus_selected_win_data[20] , 
        \DataPath/RF/bus_selected_win_data[19] , 
        \DataPath/RF/bus_selected_win_data[18] , 
        \DataPath/RF/bus_selected_win_data[17] , 
        \DataPath/RF/bus_selected_win_data[16] , 
        \DataPath/RF/bus_selected_win_data[15] , 
        \DataPath/RF/bus_selected_win_data[14] , 
        \DataPath/RF/bus_selected_win_data[13] , 
        \DataPath/RF/bus_selected_win_data[12] , 
        \DataPath/RF/bus_selected_win_data[11] , 
        \DataPath/RF/bus_selected_win_data[10] , 
        \DataPath/RF/bus_selected_win_data[9] , 
        \DataPath/RF/bus_selected_win_data[8] , 
        \DataPath/RF/bus_selected_win_data[7] , 
        \DataPath/RF/bus_selected_win_data[6] , 
        \DataPath/RF/bus_selected_win_data[5] , 
        \DataPath/RF/bus_selected_win_data[4] , 
        \DataPath/RF/bus_selected_win_data[3] , 
        \DataPath/RF/bus_selected_win_data[2] , 
        \DataPath/RF/bus_selected_win_data[1] , 
        \DataPath/RF/bus_selected_win_data[0] , 
        \DataPath/RF/bus_complete_win_data[255] , 
        \DataPath/RF/bus_complete_win_data[254] , 
        \DataPath/RF/bus_complete_win_data[253] , 
        \DataPath/RF/bus_complete_win_data[252] , 
        \DataPath/RF/bus_complete_win_data[251] , 
        \DataPath/RF/bus_complete_win_data[250] , 
        \DataPath/RF/bus_complete_win_data[249] , 
        \DataPath/RF/bus_complete_win_data[248] , 
        \DataPath/RF/bus_complete_win_data[247] , 
        \DataPath/RF/bus_complete_win_data[246] , 
        \DataPath/RF/bus_complete_win_data[245] , 
        \DataPath/RF/bus_complete_win_data[244] , 
        \DataPath/RF/bus_complete_win_data[243] , 
        \DataPath/RF/bus_complete_win_data[242] , 
        \DataPath/RF/bus_complete_win_data[241] , 
        \DataPath/RF/bus_complete_win_data[240] , 
        \DataPath/RF/bus_complete_win_data[239] , 
        \DataPath/RF/bus_complete_win_data[238] , 
        \DataPath/RF/bus_complete_win_data[237] , 
        \DataPath/RF/bus_complete_win_data[236] , 
        \DataPath/RF/bus_complete_win_data[235] , 
        \DataPath/RF/bus_complete_win_data[234] , 
        \DataPath/RF/bus_complete_win_data[233] , 
        \DataPath/RF/bus_complete_win_data[232] , 
        \DataPath/RF/bus_complete_win_data[231] , 
        \DataPath/RF/bus_complete_win_data[230] , 
        \DataPath/RF/bus_complete_win_data[229] , 
        \DataPath/RF/bus_complete_win_data[228] , 
        \DataPath/RF/bus_complete_win_data[227] , 
        \DataPath/RF/bus_complete_win_data[226] , 
        \DataPath/RF/bus_complete_win_data[225] , 
        \DataPath/RF/bus_complete_win_data[224] , 
        \DataPath/RF/bus_complete_win_data[223] , 
        \DataPath/RF/bus_complete_win_data[222] , 
        \DataPath/RF/bus_complete_win_data[221] , 
        \DataPath/RF/bus_complete_win_data[220] , 
        \DataPath/RF/bus_complete_win_data[219] , 
        \DataPath/RF/bus_complete_win_data[218] , 
        \DataPath/RF/bus_complete_win_data[217] , 
        \DataPath/RF/bus_complete_win_data[216] , 
        \DataPath/RF/bus_complete_win_data[215] , 
        \DataPath/RF/bus_complete_win_data[214] , 
        \DataPath/RF/bus_complete_win_data[213] , 
        \DataPath/RF/bus_complete_win_data[212] , 
        \DataPath/RF/bus_complete_win_data[211] , 
        \DataPath/RF/bus_complete_win_data[210] , 
        \DataPath/RF/bus_complete_win_data[209] , 
        \DataPath/RF/bus_complete_win_data[208] , 
        \DataPath/RF/bus_complete_win_data[207] , 
        \DataPath/RF/bus_complete_win_data[206] , 
        \DataPath/RF/bus_complete_win_data[205] , 
        \DataPath/RF/bus_complete_win_data[204] , 
        \DataPath/RF/bus_complete_win_data[203] , 
        \DataPath/RF/bus_complete_win_data[202] , 
        \DataPath/RF/bus_complete_win_data[201] , 
        \DataPath/RF/bus_complete_win_data[200] , 
        \DataPath/RF/bus_complete_win_data[199] , 
        \DataPath/RF/bus_complete_win_data[198] , 
        \DataPath/RF/bus_complete_win_data[197] , 
        \DataPath/RF/bus_complete_win_data[196] , 
        \DataPath/RF/bus_complete_win_data[195] , 
        \DataPath/RF/bus_complete_win_data[194] , 
        \DataPath/RF/bus_complete_win_data[193] , 
        \DataPath/RF/bus_complete_win_data[192] , 
        \DataPath/RF/bus_complete_win_data[191] , 
        \DataPath/RF/bus_complete_win_data[190] , 
        \DataPath/RF/bus_complete_win_data[189] , 
        \DataPath/RF/bus_complete_win_data[188] , 
        \DataPath/RF/bus_complete_win_data[187] , 
        \DataPath/RF/bus_complete_win_data[186] , 
        \DataPath/RF/bus_complete_win_data[185] , 
        \DataPath/RF/bus_complete_win_data[184] , 
        \DataPath/RF/bus_complete_win_data[183] , 
        \DataPath/RF/bus_complete_win_data[182] , 
        \DataPath/RF/bus_complete_win_data[181] , 
        \DataPath/RF/bus_complete_win_data[180] , 
        \DataPath/RF/bus_complete_win_data[179] , 
        \DataPath/RF/bus_complete_win_data[178] , 
        \DataPath/RF/bus_complete_win_data[177] , 
        \DataPath/RF/bus_complete_win_data[176] , 
        \DataPath/RF/bus_complete_win_data[175] , 
        \DataPath/RF/bus_complete_win_data[174] , 
        \DataPath/RF/bus_complete_win_data[173] , 
        \DataPath/RF/bus_complete_win_data[172] , 
        \DataPath/RF/bus_complete_win_data[171] , 
        \DataPath/RF/bus_complete_win_data[170] , 
        \DataPath/RF/bus_complete_win_data[169] , 
        \DataPath/RF/bus_complete_win_data[168] , 
        \DataPath/RF/bus_complete_win_data[167] , 
        \DataPath/RF/bus_complete_win_data[166] , 
        \DataPath/RF/bus_complete_win_data[165] , 
        \DataPath/RF/bus_complete_win_data[164] , 
        \DataPath/RF/bus_complete_win_data[163] , 
        \DataPath/RF/bus_complete_win_data[162] , 
        \DataPath/RF/bus_complete_win_data[161] , 
        \DataPath/RF/bus_complete_win_data[160] , 
        \DataPath/RF/bus_complete_win_data[159] , 
        \DataPath/RF/bus_complete_win_data[158] , 
        \DataPath/RF/bus_complete_win_data[157] , 
        \DataPath/RF/bus_complete_win_data[156] , 
        \DataPath/RF/bus_complete_win_data[155] , 
        \DataPath/RF/bus_complete_win_data[154] , 
        \DataPath/RF/bus_complete_win_data[153] , 
        \DataPath/RF/bus_complete_win_data[152] , 
        \DataPath/RF/bus_complete_win_data[151] , 
        \DataPath/RF/bus_complete_win_data[150] , 
        \DataPath/RF/bus_complete_win_data[149] , 
        \DataPath/RF/bus_complete_win_data[148] , 
        \DataPath/RF/bus_complete_win_data[147] , 
        \DataPath/RF/bus_complete_win_data[146] , 
        \DataPath/RF/bus_complete_win_data[145] , 
        \DataPath/RF/bus_complete_win_data[144] , 
        \DataPath/RF/bus_complete_win_data[143] , 
        \DataPath/RF/bus_complete_win_data[142] , 
        \DataPath/RF/bus_complete_win_data[141] , 
        \DataPath/RF/bus_complete_win_data[140] , 
        \DataPath/RF/bus_complete_win_data[139] , 
        \DataPath/RF/bus_complete_win_data[138] , 
        \DataPath/RF/bus_complete_win_data[137] , 
        \DataPath/RF/bus_complete_win_data[136] , 
        \DataPath/RF/bus_complete_win_data[135] , 
        \DataPath/RF/bus_complete_win_data[134] , 
        \DataPath/RF/bus_complete_win_data[133] , 
        \DataPath/RF/bus_complete_win_data[132] , 
        \DataPath/RF/bus_complete_win_data[131] , 
        \DataPath/RF/bus_complete_win_data[130] , 
        \DataPath/RF/bus_complete_win_data[129] , 
        \DataPath/RF/bus_complete_win_data[128] , 
        \DataPath/RF/bus_complete_win_data[127] , 
        \DataPath/RF/bus_complete_win_data[126] , 
        \DataPath/RF/bus_complete_win_data[125] , 
        \DataPath/RF/bus_complete_win_data[124] , 
        \DataPath/RF/bus_complete_win_data[123] , 
        \DataPath/RF/bus_complete_win_data[122] , 
        \DataPath/RF/bus_complete_win_data[121] , 
        \DataPath/RF/bus_complete_win_data[120] , 
        \DataPath/RF/bus_complete_win_data[119] , 
        \DataPath/RF/bus_complete_win_data[118] , 
        \DataPath/RF/bus_complete_win_data[117] , 
        \DataPath/RF/bus_complete_win_data[116] , 
        \DataPath/RF/bus_complete_win_data[115] , 
        \DataPath/RF/bus_complete_win_data[114] , 
        \DataPath/RF/bus_complete_win_data[113] , 
        \DataPath/RF/bus_complete_win_data[112] , 
        \DataPath/RF/bus_complete_win_data[111] , 
        \DataPath/RF/bus_complete_win_data[110] , 
        \DataPath/RF/bus_complete_win_data[109] , 
        \DataPath/RF/bus_complete_win_data[108] , 
        \DataPath/RF/bus_complete_win_data[107] , 
        \DataPath/RF/bus_complete_win_data[106] , 
        \DataPath/RF/bus_complete_win_data[105] , 
        \DataPath/RF/bus_complete_win_data[104] , 
        \DataPath/RF/bus_complete_win_data[103] , 
        \DataPath/RF/bus_complete_win_data[102] , 
        \DataPath/RF/bus_complete_win_data[101] , 
        \DataPath/RF/bus_complete_win_data[100] , 
        \DataPath/RF/bus_complete_win_data[99] , 
        \DataPath/RF/bus_complete_win_data[98] , 
        \DataPath/RF/bus_complete_win_data[97] , 
        \DataPath/RF/bus_complete_win_data[96] , 
        \DataPath/RF/bus_complete_win_data[95] , 
        \DataPath/RF/bus_complete_win_data[94] , 
        \DataPath/RF/bus_complete_win_data[93] , 
        \DataPath/RF/bus_complete_win_data[92] , 
        \DataPath/RF/bus_complete_win_data[91] , 
        \DataPath/RF/bus_complete_win_data[90] , 
        \DataPath/RF/bus_complete_win_data[89] , 
        \DataPath/RF/bus_complete_win_data[88] , 
        \DataPath/RF/bus_complete_win_data[87] , 
        \DataPath/RF/bus_complete_win_data[86] , 
        \DataPath/RF/bus_complete_win_data[85] , 
        \DataPath/RF/bus_complete_win_data[84] , 
        \DataPath/RF/bus_complete_win_data[83] , 
        \DataPath/RF/bus_complete_win_data[82] , 
        \DataPath/RF/bus_complete_win_data[81] , 
        \DataPath/RF/bus_complete_win_data[80] , 
        \DataPath/RF/bus_complete_win_data[79] , 
        \DataPath/RF/bus_complete_win_data[78] , 
        \DataPath/RF/bus_complete_win_data[77] , 
        \DataPath/RF/bus_complete_win_data[76] , 
        \DataPath/RF/bus_complete_win_data[75] , 
        \DataPath/RF/bus_complete_win_data[74] , 
        \DataPath/RF/bus_complete_win_data[73] , 
        \DataPath/RF/bus_complete_win_data[72] , 
        \DataPath/RF/bus_complete_win_data[71] , 
        \DataPath/RF/bus_complete_win_data[70] , 
        \DataPath/RF/bus_complete_win_data[69] , 
        \DataPath/RF/bus_complete_win_data[68] , 
        \DataPath/RF/bus_complete_win_data[67] , 
        \DataPath/RF/bus_complete_win_data[66] , 
        \DataPath/RF/bus_complete_win_data[65] , 
        \DataPath/RF/bus_complete_win_data[64] , 
        \DataPath/RF/bus_complete_win_data[63] , 
        \DataPath/RF/bus_complete_win_data[62] , 
        \DataPath/RF/bus_complete_win_data[61] , 
        \DataPath/RF/bus_complete_win_data[60] , 
        \DataPath/RF/bus_complete_win_data[59] , 
        \DataPath/RF/bus_complete_win_data[58] , 
        \DataPath/RF/bus_complete_win_data[57] , 
        \DataPath/RF/bus_complete_win_data[56] , 
        \DataPath/RF/bus_complete_win_data[55] , 
        \DataPath/RF/bus_complete_win_data[54] , 
        \DataPath/RF/bus_complete_win_data[53] , 
        \DataPath/RF/bus_complete_win_data[52] , 
        \DataPath/RF/bus_complete_win_data[51] , 
        \DataPath/RF/bus_complete_win_data[50] , 
        \DataPath/RF/bus_complete_win_data[49] , 
        \DataPath/RF/bus_complete_win_data[48] , 
        \DataPath/RF/bus_complete_win_data[47] , 
        \DataPath/RF/bus_complete_win_data[46] , 
        \DataPath/RF/bus_complete_win_data[45] , 
        \DataPath/RF/bus_complete_win_data[44] , 
        \DataPath/RF/bus_complete_win_data[43] , 
        \DataPath/RF/bus_complete_win_data[42] , 
        \DataPath/RF/bus_complete_win_data[41] , 
        \DataPath/RF/bus_complete_win_data[40] , 
        \DataPath/RF/bus_complete_win_data[39] , 
        \DataPath/RF/bus_complete_win_data[38] , 
        \DataPath/RF/bus_complete_win_data[37] , 
        \DataPath/RF/bus_complete_win_data[36] , 
        \DataPath/RF/bus_complete_win_data[35] , 
        \DataPath/RF/bus_complete_win_data[34] , 
        \DataPath/RF/bus_complete_win_data[33] , 
        \DataPath/RF/bus_complete_win_data[32] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .Y({\DataPath/RF/internal_out1[31] , 
        \DataPath/RF/internal_out1[30] , \DataPath/RF/internal_out1[29] , 
        \DataPath/RF/internal_out1[28] , \DataPath/RF/internal_out1[27] , 
        \DataPath/RF/internal_out1[26] , \DataPath/RF/internal_out1[25] , 
        \DataPath/RF/internal_out1[24] , \DataPath/RF/internal_out1[23] , 
        \DataPath/RF/internal_out1[22] , \DataPath/RF/internal_out1[21] , 
        \DataPath/RF/internal_out1[20] , \DataPath/RF/internal_out1[19] , 
        \DataPath/RF/internal_out1[18] , \DataPath/RF/internal_out1[17] , 
        \DataPath/RF/internal_out1[16] , \DataPath/RF/internal_out1[15] , 
        \DataPath/RF/internal_out1[14] , \DataPath/RF/internal_out1[13] , 
        \DataPath/RF/internal_out1[12] , \DataPath/RF/internal_out1[11] , 
        \DataPath/RF/internal_out1[10] , \DataPath/RF/internal_out1[9] , 
        \DataPath/RF/internal_out1[8] , \DataPath/RF/internal_out1[7] , 
        \DataPath/RF/internal_out1[6] , \DataPath/RF/internal_out1[5] , 
        \DataPath/RF/internal_out1[4] , \DataPath/RF/internal_out1[3] , 
        \DataPath/RF/internal_out1[2] , \DataPath/RF/internal_out1[1] , 
        \DataPath/RF/internal_out1[0] }) );
  select_block_NBIT_DATA32_N8_F5 \DataPath/RF/SEL_BLK  ( .regs({
        \DataPath/RF/bus_reg_dataout[2559] , 
        \DataPath/RF/bus_reg_dataout[2558] , 
        \DataPath/RF/bus_reg_dataout[2557] , 
        \DataPath/RF/bus_reg_dataout[2556] , 
        \DataPath/RF/bus_reg_dataout[2555] , 
        \DataPath/RF/bus_reg_dataout[2554] , 
        \DataPath/RF/bus_reg_dataout[2553] , 
        \DataPath/RF/bus_reg_dataout[2552] , 
        \DataPath/RF/bus_reg_dataout[2551] , 
        \DataPath/RF/bus_reg_dataout[2550] , 
        \DataPath/RF/bus_reg_dataout[2549] , 
        \DataPath/RF/bus_reg_dataout[2548] , 
        \DataPath/RF/bus_reg_dataout[2547] , 
        \DataPath/RF/bus_reg_dataout[2546] , 
        \DataPath/RF/bus_reg_dataout[2545] , 
        \DataPath/RF/bus_reg_dataout[2544] , 
        \DataPath/RF/bus_reg_dataout[2543] , 
        \DataPath/RF/bus_reg_dataout[2542] , 
        \DataPath/RF/bus_reg_dataout[2541] , 
        \DataPath/RF/bus_reg_dataout[2540] , 
        \DataPath/RF/bus_reg_dataout[2539] , 
        \DataPath/RF/bus_reg_dataout[2538] , 
        \DataPath/RF/bus_reg_dataout[2537] , 
        \DataPath/RF/bus_reg_dataout[2536] , 
        \DataPath/RF/bus_reg_dataout[2535] , 
        \DataPath/RF/bus_reg_dataout[2534] , 
        \DataPath/RF/bus_reg_dataout[2533] , 
        \DataPath/RF/bus_reg_dataout[2532] , 
        \DataPath/RF/bus_reg_dataout[2531] , 
        \DataPath/RF/bus_reg_dataout[2530] , 
        \DataPath/RF/bus_reg_dataout[2529] , 
        \DataPath/RF/bus_reg_dataout[2528] , 
        \DataPath/RF/bus_reg_dataout[2527] , 
        \DataPath/RF/bus_reg_dataout[2526] , 
        \DataPath/RF/bus_reg_dataout[2525] , 
        \DataPath/RF/bus_reg_dataout[2524] , 
        \DataPath/RF/bus_reg_dataout[2523] , 
        \DataPath/RF/bus_reg_dataout[2522] , 
        \DataPath/RF/bus_reg_dataout[2521] , 
        \DataPath/RF/bus_reg_dataout[2520] , 
        \DataPath/RF/bus_reg_dataout[2519] , 
        \DataPath/RF/bus_reg_dataout[2518] , 
        \DataPath/RF/bus_reg_dataout[2517] , 
        \DataPath/RF/bus_reg_dataout[2516] , 
        \DataPath/RF/bus_reg_dataout[2515] , 
        \DataPath/RF/bus_reg_dataout[2514] , 
        \DataPath/RF/bus_reg_dataout[2513] , 
        \DataPath/RF/bus_reg_dataout[2512] , 
        \DataPath/RF/bus_reg_dataout[2511] , 
        \DataPath/RF/bus_reg_dataout[2510] , 
        \DataPath/RF/bus_reg_dataout[2509] , 
        \DataPath/RF/bus_reg_dataout[2508] , 
        \DataPath/RF/bus_reg_dataout[2507] , 
        \DataPath/RF/bus_reg_dataout[2506] , 
        \DataPath/RF/bus_reg_dataout[2505] , 
        \DataPath/RF/bus_reg_dataout[2504] , 
        \DataPath/RF/bus_reg_dataout[2503] , 
        \DataPath/RF/bus_reg_dataout[2502] , 
        \DataPath/RF/bus_reg_dataout[2501] , 
        \DataPath/RF/bus_reg_dataout[2500] , 
        \DataPath/RF/bus_reg_dataout[2499] , 
        \DataPath/RF/bus_reg_dataout[2498] , 
        \DataPath/RF/bus_reg_dataout[2497] , 
        \DataPath/RF/bus_reg_dataout[2496] , 
        \DataPath/RF/bus_reg_dataout[2495] , 
        \DataPath/RF/bus_reg_dataout[2494] , 
        \DataPath/RF/bus_reg_dataout[2493] , 
        \DataPath/RF/bus_reg_dataout[2492] , 
        \DataPath/RF/bus_reg_dataout[2491] , 
        \DataPath/RF/bus_reg_dataout[2490] , 
        \DataPath/RF/bus_reg_dataout[2489] , 
        \DataPath/RF/bus_reg_dataout[2488] , 
        \DataPath/RF/bus_reg_dataout[2487] , 
        \DataPath/RF/bus_reg_dataout[2486] , 
        \DataPath/RF/bus_reg_dataout[2485] , 
        \DataPath/RF/bus_reg_dataout[2484] , 
        \DataPath/RF/bus_reg_dataout[2483] , 
        \DataPath/RF/bus_reg_dataout[2482] , 
        \DataPath/RF/bus_reg_dataout[2481] , 
        \DataPath/RF/bus_reg_dataout[2480] , 
        \DataPath/RF/bus_reg_dataout[2479] , 
        \DataPath/RF/bus_reg_dataout[2478] , 
        \DataPath/RF/bus_reg_dataout[2477] , 
        \DataPath/RF/bus_reg_dataout[2476] , 
        \DataPath/RF/bus_reg_dataout[2475] , 
        \DataPath/RF/bus_reg_dataout[2474] , 
        \DataPath/RF/bus_reg_dataout[2473] , 
        \DataPath/RF/bus_reg_dataout[2472] , 
        \DataPath/RF/bus_reg_dataout[2471] , 
        \DataPath/RF/bus_reg_dataout[2470] , 
        \DataPath/RF/bus_reg_dataout[2469] , 
        \DataPath/RF/bus_reg_dataout[2468] , 
        \DataPath/RF/bus_reg_dataout[2467] , 
        \DataPath/RF/bus_reg_dataout[2466] , 
        \DataPath/RF/bus_reg_dataout[2465] , 
        \DataPath/RF/bus_reg_dataout[2464] , 
        \DataPath/RF/bus_reg_dataout[2463] , 
        \DataPath/RF/bus_reg_dataout[2462] , 
        \DataPath/RF/bus_reg_dataout[2461] , 
        \DataPath/RF/bus_reg_dataout[2460] , 
        \DataPath/RF/bus_reg_dataout[2459] , 
        \DataPath/RF/bus_reg_dataout[2458] , 
        \DataPath/RF/bus_reg_dataout[2457] , 
        \DataPath/RF/bus_reg_dataout[2456] , 
        \DataPath/RF/bus_reg_dataout[2455] , 
        \DataPath/RF/bus_reg_dataout[2454] , 
        \DataPath/RF/bus_reg_dataout[2453] , 
        \DataPath/RF/bus_reg_dataout[2452] , 
        \DataPath/RF/bus_reg_dataout[2451] , 
        \DataPath/RF/bus_reg_dataout[2450] , 
        \DataPath/RF/bus_reg_dataout[2449] , 
        \DataPath/RF/bus_reg_dataout[2448] , 
        \DataPath/RF/bus_reg_dataout[2447] , 
        \DataPath/RF/bus_reg_dataout[2446] , 
        \DataPath/RF/bus_reg_dataout[2445] , 
        \DataPath/RF/bus_reg_dataout[2444] , 
        \DataPath/RF/bus_reg_dataout[2443] , 
        \DataPath/RF/bus_reg_dataout[2442] , 
        \DataPath/RF/bus_reg_dataout[2441] , 
        \DataPath/RF/bus_reg_dataout[2440] , 
        \DataPath/RF/bus_reg_dataout[2439] , 
        \DataPath/RF/bus_reg_dataout[2438] , 
        \DataPath/RF/bus_reg_dataout[2437] , 
        \DataPath/RF/bus_reg_dataout[2436] , 
        \DataPath/RF/bus_reg_dataout[2435] , 
        \DataPath/RF/bus_reg_dataout[2434] , 
        \DataPath/RF/bus_reg_dataout[2433] , 
        \DataPath/RF/bus_reg_dataout[2432] , 
        \DataPath/RF/bus_reg_dataout[2431] , 
        \DataPath/RF/bus_reg_dataout[2430] , 
        \DataPath/RF/bus_reg_dataout[2429] , 
        \DataPath/RF/bus_reg_dataout[2428] , 
        \DataPath/RF/bus_reg_dataout[2427] , 
        \DataPath/RF/bus_reg_dataout[2426] , 
        \DataPath/RF/bus_reg_dataout[2425] , 
        \DataPath/RF/bus_reg_dataout[2424] , 
        \DataPath/RF/bus_reg_dataout[2423] , 
        \DataPath/RF/bus_reg_dataout[2422] , 
        \DataPath/RF/bus_reg_dataout[2421] , 
        \DataPath/RF/bus_reg_dataout[2420] , 
        \DataPath/RF/bus_reg_dataout[2419] , 
        \DataPath/RF/bus_reg_dataout[2418] , 
        \DataPath/RF/bus_reg_dataout[2417] , 
        \DataPath/RF/bus_reg_dataout[2416] , 
        \DataPath/RF/bus_reg_dataout[2415] , 
        \DataPath/RF/bus_reg_dataout[2414] , 
        \DataPath/RF/bus_reg_dataout[2413] , 
        \DataPath/RF/bus_reg_dataout[2412] , 
        \DataPath/RF/bus_reg_dataout[2411] , 
        \DataPath/RF/bus_reg_dataout[2410] , 
        \DataPath/RF/bus_reg_dataout[2409] , 
        \DataPath/RF/bus_reg_dataout[2408] , 
        \DataPath/RF/bus_reg_dataout[2407] , 
        \DataPath/RF/bus_reg_dataout[2406] , 
        \DataPath/RF/bus_reg_dataout[2405] , 
        \DataPath/RF/bus_reg_dataout[2404] , 
        \DataPath/RF/bus_reg_dataout[2403] , 
        \DataPath/RF/bus_reg_dataout[2402] , 
        \DataPath/RF/bus_reg_dataout[2401] , 
        \DataPath/RF/bus_reg_dataout[2400] , 
        \DataPath/RF/bus_reg_dataout[2399] , 
        \DataPath/RF/bus_reg_dataout[2398] , 
        \DataPath/RF/bus_reg_dataout[2397] , 
        \DataPath/RF/bus_reg_dataout[2396] , 
        \DataPath/RF/bus_reg_dataout[2395] , 
        \DataPath/RF/bus_reg_dataout[2394] , 
        \DataPath/RF/bus_reg_dataout[2393] , 
        \DataPath/RF/bus_reg_dataout[2392] , 
        \DataPath/RF/bus_reg_dataout[2391] , 
        \DataPath/RF/bus_reg_dataout[2390] , 
        \DataPath/RF/bus_reg_dataout[2389] , 
        \DataPath/RF/bus_reg_dataout[2388] , 
        \DataPath/RF/bus_reg_dataout[2387] , 
        \DataPath/RF/bus_reg_dataout[2386] , 
        \DataPath/RF/bus_reg_dataout[2385] , 
        \DataPath/RF/bus_reg_dataout[2384] , 
        \DataPath/RF/bus_reg_dataout[2383] , 
        \DataPath/RF/bus_reg_dataout[2382] , 
        \DataPath/RF/bus_reg_dataout[2381] , 
        \DataPath/RF/bus_reg_dataout[2380] , 
        \DataPath/RF/bus_reg_dataout[2379] , 
        \DataPath/RF/bus_reg_dataout[2378] , 
        \DataPath/RF/bus_reg_dataout[2377] , 
        \DataPath/RF/bus_reg_dataout[2376] , 
        \DataPath/RF/bus_reg_dataout[2375] , 
        \DataPath/RF/bus_reg_dataout[2374] , 
        \DataPath/RF/bus_reg_dataout[2373] , 
        \DataPath/RF/bus_reg_dataout[2372] , 
        \DataPath/RF/bus_reg_dataout[2371] , 
        \DataPath/RF/bus_reg_dataout[2370] , 
        \DataPath/RF/bus_reg_dataout[2369] , 
        \DataPath/RF/bus_reg_dataout[2368] , 
        \DataPath/RF/bus_reg_dataout[2367] , 
        \DataPath/RF/bus_reg_dataout[2366] , 
        \DataPath/RF/bus_reg_dataout[2365] , 
        \DataPath/RF/bus_reg_dataout[2364] , 
        \DataPath/RF/bus_reg_dataout[2363] , 
        \DataPath/RF/bus_reg_dataout[2362] , 
        \DataPath/RF/bus_reg_dataout[2361] , 
        \DataPath/RF/bus_reg_dataout[2360] , 
        \DataPath/RF/bus_reg_dataout[2359] , 
        \DataPath/RF/bus_reg_dataout[2358] , 
        \DataPath/RF/bus_reg_dataout[2357] , 
        \DataPath/RF/bus_reg_dataout[2356] , 
        \DataPath/RF/bus_reg_dataout[2355] , 
        \DataPath/RF/bus_reg_dataout[2354] , 
        \DataPath/RF/bus_reg_dataout[2353] , 
        \DataPath/RF/bus_reg_dataout[2352] , 
        \DataPath/RF/bus_reg_dataout[2351] , 
        \DataPath/RF/bus_reg_dataout[2350] , 
        \DataPath/RF/bus_reg_dataout[2349] , 
        \DataPath/RF/bus_reg_dataout[2348] , 
        \DataPath/RF/bus_reg_dataout[2347] , 
        \DataPath/RF/bus_reg_dataout[2346] , 
        \DataPath/RF/bus_reg_dataout[2345] , 
        \DataPath/RF/bus_reg_dataout[2344] , 
        \DataPath/RF/bus_reg_dataout[2343] , 
        \DataPath/RF/bus_reg_dataout[2342] , 
        \DataPath/RF/bus_reg_dataout[2341] , 
        \DataPath/RF/bus_reg_dataout[2340] , 
        \DataPath/RF/bus_reg_dataout[2339] , 
        \DataPath/RF/bus_reg_dataout[2338] , 
        \DataPath/RF/bus_reg_dataout[2337] , 
        \DataPath/RF/bus_reg_dataout[2336] , 
        \DataPath/RF/bus_reg_dataout[2335] , 
        \DataPath/RF/bus_reg_dataout[2334] , 
        \DataPath/RF/bus_reg_dataout[2333] , 
        \DataPath/RF/bus_reg_dataout[2332] , 
        \DataPath/RF/bus_reg_dataout[2331] , 
        \DataPath/RF/bus_reg_dataout[2330] , 
        \DataPath/RF/bus_reg_dataout[2329] , 
        \DataPath/RF/bus_reg_dataout[2328] , 
        \DataPath/RF/bus_reg_dataout[2327] , 
        \DataPath/RF/bus_reg_dataout[2326] , 
        \DataPath/RF/bus_reg_dataout[2325] , 
        \DataPath/RF/bus_reg_dataout[2324] , 
        \DataPath/RF/bus_reg_dataout[2323] , 
        \DataPath/RF/bus_reg_dataout[2322] , 
        \DataPath/RF/bus_reg_dataout[2321] , 
        \DataPath/RF/bus_reg_dataout[2320] , 
        \DataPath/RF/bus_reg_dataout[2319] , 
        \DataPath/RF/bus_reg_dataout[2318] , 
        \DataPath/RF/bus_reg_dataout[2317] , 
        \DataPath/RF/bus_reg_dataout[2316] , 
        \DataPath/RF/bus_reg_dataout[2315] , 
        \DataPath/RF/bus_reg_dataout[2314] , 
        \DataPath/RF/bus_reg_dataout[2313] , 
        \DataPath/RF/bus_reg_dataout[2312] , 
        \DataPath/RF/bus_reg_dataout[2311] , 
        \DataPath/RF/bus_reg_dataout[2310] , 
        \DataPath/RF/bus_reg_dataout[2309] , 
        \DataPath/RF/bus_reg_dataout[2308] , 
        \DataPath/RF/bus_reg_dataout[2307] , 
        \DataPath/RF/bus_reg_dataout[2306] , 
        \DataPath/RF/bus_reg_dataout[2305] , 
        \DataPath/RF/bus_reg_dataout[2304] , 
        \DataPath/RF/bus_reg_dataout[2303] , 
        \DataPath/RF/bus_reg_dataout[2302] , 
        \DataPath/RF/bus_reg_dataout[2301] , 
        \DataPath/RF/bus_reg_dataout[2300] , 
        \DataPath/RF/bus_reg_dataout[2299] , 
        \DataPath/RF/bus_reg_dataout[2298] , 
        \DataPath/RF/bus_reg_dataout[2297] , 
        \DataPath/RF/bus_reg_dataout[2296] , 
        \DataPath/RF/bus_reg_dataout[2295] , 
        \DataPath/RF/bus_reg_dataout[2294] , 
        \DataPath/RF/bus_reg_dataout[2293] , 
        \DataPath/RF/bus_reg_dataout[2292] , 
        \DataPath/RF/bus_reg_dataout[2291] , 
        \DataPath/RF/bus_reg_dataout[2290] , 
        \DataPath/RF/bus_reg_dataout[2289] , 
        \DataPath/RF/bus_reg_dataout[2288] , 
        \DataPath/RF/bus_reg_dataout[2287] , 
        \DataPath/RF/bus_reg_dataout[2286] , 
        \DataPath/RF/bus_reg_dataout[2285] , 
        \DataPath/RF/bus_reg_dataout[2284] , 
        \DataPath/RF/bus_reg_dataout[2283] , 
        \DataPath/RF/bus_reg_dataout[2282] , 
        \DataPath/RF/bus_reg_dataout[2281] , 
        \DataPath/RF/bus_reg_dataout[2280] , 
        \DataPath/RF/bus_reg_dataout[2279] , 
        \DataPath/RF/bus_reg_dataout[2278] , 
        \DataPath/RF/bus_reg_dataout[2277] , 
        \DataPath/RF/bus_reg_dataout[2276] , 
        \DataPath/RF/bus_reg_dataout[2275] , 
        \DataPath/RF/bus_reg_dataout[2274] , 
        \DataPath/RF/bus_reg_dataout[2273] , 
        \DataPath/RF/bus_reg_dataout[2272] , 
        \DataPath/RF/bus_reg_dataout[2271] , 
        \DataPath/RF/bus_reg_dataout[2270] , 
        \DataPath/RF/bus_reg_dataout[2269] , 
        \DataPath/RF/bus_reg_dataout[2268] , 
        \DataPath/RF/bus_reg_dataout[2267] , 
        \DataPath/RF/bus_reg_dataout[2266] , 
        \DataPath/RF/bus_reg_dataout[2265] , 
        \DataPath/RF/bus_reg_dataout[2264] , 
        \DataPath/RF/bus_reg_dataout[2263] , 
        \DataPath/RF/bus_reg_dataout[2262] , 
        \DataPath/RF/bus_reg_dataout[2261] , 
        \DataPath/RF/bus_reg_dataout[2260] , 
        \DataPath/RF/bus_reg_dataout[2259] , 
        \DataPath/RF/bus_reg_dataout[2258] , 
        \DataPath/RF/bus_reg_dataout[2257] , 
        \DataPath/RF/bus_reg_dataout[2256] , 
        \DataPath/RF/bus_reg_dataout[2255] , 
        \DataPath/RF/bus_reg_dataout[2254] , 
        \DataPath/RF/bus_reg_dataout[2253] , 
        \DataPath/RF/bus_reg_dataout[2252] , 
        \DataPath/RF/bus_reg_dataout[2251] , 
        \DataPath/RF/bus_reg_dataout[2250] , 
        \DataPath/RF/bus_reg_dataout[2249] , 
        \DataPath/RF/bus_reg_dataout[2248] , 
        \DataPath/RF/bus_reg_dataout[2247] , 
        \DataPath/RF/bus_reg_dataout[2246] , 
        \DataPath/RF/bus_reg_dataout[2245] , 
        \DataPath/RF/bus_reg_dataout[2244] , 
        \DataPath/RF/bus_reg_dataout[2243] , 
        \DataPath/RF/bus_reg_dataout[2242] , 
        \DataPath/RF/bus_reg_dataout[2241] , 
        \DataPath/RF/bus_reg_dataout[2240] , 
        \DataPath/RF/bus_reg_dataout[2239] , 
        \DataPath/RF/bus_reg_dataout[2238] , 
        \DataPath/RF/bus_reg_dataout[2237] , 
        \DataPath/RF/bus_reg_dataout[2236] , 
        \DataPath/RF/bus_reg_dataout[2235] , 
        \DataPath/RF/bus_reg_dataout[2234] , 
        \DataPath/RF/bus_reg_dataout[2233] , 
        \DataPath/RF/bus_reg_dataout[2232] , 
        \DataPath/RF/bus_reg_dataout[2231] , 
        \DataPath/RF/bus_reg_dataout[2230] , 
        \DataPath/RF/bus_reg_dataout[2229] , 
        \DataPath/RF/bus_reg_dataout[2228] , 
        \DataPath/RF/bus_reg_dataout[2227] , 
        \DataPath/RF/bus_reg_dataout[2226] , 
        \DataPath/RF/bus_reg_dataout[2225] , 
        \DataPath/RF/bus_reg_dataout[2224] , 
        \DataPath/RF/bus_reg_dataout[2223] , 
        \DataPath/RF/bus_reg_dataout[2222] , 
        \DataPath/RF/bus_reg_dataout[2221] , 
        \DataPath/RF/bus_reg_dataout[2220] , 
        \DataPath/RF/bus_reg_dataout[2219] , 
        \DataPath/RF/bus_reg_dataout[2218] , 
        \DataPath/RF/bus_reg_dataout[2217] , 
        \DataPath/RF/bus_reg_dataout[2216] , 
        \DataPath/RF/bus_reg_dataout[2215] , 
        \DataPath/RF/bus_reg_dataout[2214] , 
        \DataPath/RF/bus_reg_dataout[2213] , 
        \DataPath/RF/bus_reg_dataout[2212] , 
        \DataPath/RF/bus_reg_dataout[2211] , 
        \DataPath/RF/bus_reg_dataout[2210] , 
        \DataPath/RF/bus_reg_dataout[2209] , 
        \DataPath/RF/bus_reg_dataout[2208] , 
        \DataPath/RF/bus_reg_dataout[2207] , 
        \DataPath/RF/bus_reg_dataout[2206] , 
        \DataPath/RF/bus_reg_dataout[2205] , 
        \DataPath/RF/bus_reg_dataout[2204] , 
        \DataPath/RF/bus_reg_dataout[2203] , 
        \DataPath/RF/bus_reg_dataout[2202] , 
        \DataPath/RF/bus_reg_dataout[2201] , 
        \DataPath/RF/bus_reg_dataout[2200] , 
        \DataPath/RF/bus_reg_dataout[2199] , 
        \DataPath/RF/bus_reg_dataout[2198] , 
        \DataPath/RF/bus_reg_dataout[2197] , 
        \DataPath/RF/bus_reg_dataout[2196] , 
        \DataPath/RF/bus_reg_dataout[2195] , 
        \DataPath/RF/bus_reg_dataout[2194] , 
        \DataPath/RF/bus_reg_dataout[2193] , 
        \DataPath/RF/bus_reg_dataout[2192] , 
        \DataPath/RF/bus_reg_dataout[2191] , 
        \DataPath/RF/bus_reg_dataout[2190] , 
        \DataPath/RF/bus_reg_dataout[2189] , 
        \DataPath/RF/bus_reg_dataout[2188] , 
        \DataPath/RF/bus_reg_dataout[2187] , 
        \DataPath/RF/bus_reg_dataout[2186] , 
        \DataPath/RF/bus_reg_dataout[2185] , 
        \DataPath/RF/bus_reg_dataout[2184] , 
        \DataPath/RF/bus_reg_dataout[2183] , 
        \DataPath/RF/bus_reg_dataout[2182] , 
        \DataPath/RF/bus_reg_dataout[2181] , 
        \DataPath/RF/bus_reg_dataout[2180] , 
        \DataPath/RF/bus_reg_dataout[2179] , 
        \DataPath/RF/bus_reg_dataout[2178] , 
        \DataPath/RF/bus_reg_dataout[2177] , 
        \DataPath/RF/bus_reg_dataout[2176] , 
        \DataPath/RF/bus_reg_dataout[2175] , 
        \DataPath/RF/bus_reg_dataout[2174] , 
        \DataPath/RF/bus_reg_dataout[2173] , 
        \DataPath/RF/bus_reg_dataout[2172] , 
        \DataPath/RF/bus_reg_dataout[2171] , 
        \DataPath/RF/bus_reg_dataout[2170] , 
        \DataPath/RF/bus_reg_dataout[2169] , 
        \DataPath/RF/bus_reg_dataout[2168] , 
        \DataPath/RF/bus_reg_dataout[2167] , 
        \DataPath/RF/bus_reg_dataout[2166] , 
        \DataPath/RF/bus_reg_dataout[2165] , 
        \DataPath/RF/bus_reg_dataout[2164] , 
        \DataPath/RF/bus_reg_dataout[2163] , 
        \DataPath/RF/bus_reg_dataout[2162] , 
        \DataPath/RF/bus_reg_dataout[2161] , 
        \DataPath/RF/bus_reg_dataout[2160] , 
        \DataPath/RF/bus_reg_dataout[2159] , 
        \DataPath/RF/bus_reg_dataout[2158] , 
        \DataPath/RF/bus_reg_dataout[2157] , 
        \DataPath/RF/bus_reg_dataout[2156] , 
        \DataPath/RF/bus_reg_dataout[2155] , 
        \DataPath/RF/bus_reg_dataout[2154] , 
        \DataPath/RF/bus_reg_dataout[2153] , 
        \DataPath/RF/bus_reg_dataout[2152] , 
        \DataPath/RF/bus_reg_dataout[2151] , 
        \DataPath/RF/bus_reg_dataout[2150] , 
        \DataPath/RF/bus_reg_dataout[2149] , 
        \DataPath/RF/bus_reg_dataout[2148] , 
        \DataPath/RF/bus_reg_dataout[2147] , 
        \DataPath/RF/bus_reg_dataout[2146] , 
        \DataPath/RF/bus_reg_dataout[2145] , 
        \DataPath/RF/bus_reg_dataout[2144] , 
        \DataPath/RF/bus_reg_dataout[2143] , 
        \DataPath/RF/bus_reg_dataout[2142] , 
        \DataPath/RF/bus_reg_dataout[2141] , 
        \DataPath/RF/bus_reg_dataout[2140] , 
        \DataPath/RF/bus_reg_dataout[2139] , 
        \DataPath/RF/bus_reg_dataout[2138] , 
        \DataPath/RF/bus_reg_dataout[2137] , 
        \DataPath/RF/bus_reg_dataout[2136] , 
        \DataPath/RF/bus_reg_dataout[2135] , 
        \DataPath/RF/bus_reg_dataout[2134] , 
        \DataPath/RF/bus_reg_dataout[2133] , 
        \DataPath/RF/bus_reg_dataout[2132] , 
        \DataPath/RF/bus_reg_dataout[2131] , 
        \DataPath/RF/bus_reg_dataout[2130] , 
        \DataPath/RF/bus_reg_dataout[2129] , 
        \DataPath/RF/bus_reg_dataout[2128] , 
        \DataPath/RF/bus_reg_dataout[2127] , 
        \DataPath/RF/bus_reg_dataout[2126] , 
        \DataPath/RF/bus_reg_dataout[2125] , 
        \DataPath/RF/bus_reg_dataout[2124] , 
        \DataPath/RF/bus_reg_dataout[2123] , 
        \DataPath/RF/bus_reg_dataout[2122] , 
        \DataPath/RF/bus_reg_dataout[2121] , 
        \DataPath/RF/bus_reg_dataout[2120] , 
        \DataPath/RF/bus_reg_dataout[2119] , 
        \DataPath/RF/bus_reg_dataout[2118] , 
        \DataPath/RF/bus_reg_dataout[2117] , 
        \DataPath/RF/bus_reg_dataout[2116] , 
        \DataPath/RF/bus_reg_dataout[2115] , 
        \DataPath/RF/bus_reg_dataout[2114] , 
        \DataPath/RF/bus_reg_dataout[2113] , 
        \DataPath/RF/bus_reg_dataout[2112] , 
        \DataPath/RF/bus_reg_dataout[2111] , 
        \DataPath/RF/bus_reg_dataout[2110] , 
        \DataPath/RF/bus_reg_dataout[2109] , 
        \DataPath/RF/bus_reg_dataout[2108] , 
        \DataPath/RF/bus_reg_dataout[2107] , 
        \DataPath/RF/bus_reg_dataout[2106] , 
        \DataPath/RF/bus_reg_dataout[2105] , 
        \DataPath/RF/bus_reg_dataout[2104] , 
        \DataPath/RF/bus_reg_dataout[2103] , 
        \DataPath/RF/bus_reg_dataout[2102] , 
        \DataPath/RF/bus_reg_dataout[2101] , 
        \DataPath/RF/bus_reg_dataout[2100] , 
        \DataPath/RF/bus_reg_dataout[2099] , 
        \DataPath/RF/bus_reg_dataout[2098] , 
        \DataPath/RF/bus_reg_dataout[2097] , 
        \DataPath/RF/bus_reg_dataout[2096] , 
        \DataPath/RF/bus_reg_dataout[2095] , 
        \DataPath/RF/bus_reg_dataout[2094] , 
        \DataPath/RF/bus_reg_dataout[2093] , 
        \DataPath/RF/bus_reg_dataout[2092] , 
        \DataPath/RF/bus_reg_dataout[2091] , 
        \DataPath/RF/bus_reg_dataout[2090] , 
        \DataPath/RF/bus_reg_dataout[2089] , 
        \DataPath/RF/bus_reg_dataout[2088] , 
        \DataPath/RF/bus_reg_dataout[2087] , 
        \DataPath/RF/bus_reg_dataout[2086] , 
        \DataPath/RF/bus_reg_dataout[2085] , 
        \DataPath/RF/bus_reg_dataout[2084] , 
        \DataPath/RF/bus_reg_dataout[2083] , 
        \DataPath/RF/bus_reg_dataout[2082] , 
        \DataPath/RF/bus_reg_dataout[2081] , 
        \DataPath/RF/bus_reg_dataout[2080] , 
        \DataPath/RF/bus_reg_dataout[2079] , 
        \DataPath/RF/bus_reg_dataout[2078] , 
        \DataPath/RF/bus_reg_dataout[2077] , 
        \DataPath/RF/bus_reg_dataout[2076] , 
        \DataPath/RF/bus_reg_dataout[2075] , 
        \DataPath/RF/bus_reg_dataout[2074] , 
        \DataPath/RF/bus_reg_dataout[2073] , 
        \DataPath/RF/bus_reg_dataout[2072] , 
        \DataPath/RF/bus_reg_dataout[2071] , 
        \DataPath/RF/bus_reg_dataout[2070] , 
        \DataPath/RF/bus_reg_dataout[2069] , 
        \DataPath/RF/bus_reg_dataout[2068] , 
        \DataPath/RF/bus_reg_dataout[2067] , 
        \DataPath/RF/bus_reg_dataout[2066] , 
        \DataPath/RF/bus_reg_dataout[2065] , 
        \DataPath/RF/bus_reg_dataout[2064] , 
        \DataPath/RF/bus_reg_dataout[2063] , 
        \DataPath/RF/bus_reg_dataout[2062] , 
        \DataPath/RF/bus_reg_dataout[2061] , 
        \DataPath/RF/bus_reg_dataout[2060] , 
        \DataPath/RF/bus_reg_dataout[2059] , 
        \DataPath/RF/bus_reg_dataout[2058] , 
        \DataPath/RF/bus_reg_dataout[2057] , 
        \DataPath/RF/bus_reg_dataout[2056] , 
        \DataPath/RF/bus_reg_dataout[2055] , 
        \DataPath/RF/bus_reg_dataout[2054] , 
        \DataPath/RF/bus_reg_dataout[2053] , 
        \DataPath/RF/bus_reg_dataout[2052] , 
        \DataPath/RF/bus_reg_dataout[2051] , 
        \DataPath/RF/bus_reg_dataout[2050] , 
        \DataPath/RF/bus_reg_dataout[2049] , 
        \DataPath/RF/bus_reg_dataout[2048] , 
        \DataPath/RF/bus_reg_dataout[2047] , 
        \DataPath/RF/bus_reg_dataout[2046] , 
        \DataPath/RF/bus_reg_dataout[2045] , 
        \DataPath/RF/bus_reg_dataout[2044] , 
        \DataPath/RF/bus_reg_dataout[2043] , 
        \DataPath/RF/bus_reg_dataout[2042] , 
        \DataPath/RF/bus_reg_dataout[2041] , 
        \DataPath/RF/bus_reg_dataout[2040] , 
        \DataPath/RF/bus_reg_dataout[2039] , 
        \DataPath/RF/bus_reg_dataout[2038] , 
        \DataPath/RF/bus_reg_dataout[2037] , 
        \DataPath/RF/bus_reg_dataout[2036] , 
        \DataPath/RF/bus_reg_dataout[2035] , 
        \DataPath/RF/bus_reg_dataout[2034] , 
        \DataPath/RF/bus_reg_dataout[2033] , 
        \DataPath/RF/bus_reg_dataout[2032] , 
        \DataPath/RF/bus_reg_dataout[2031] , 
        \DataPath/RF/bus_reg_dataout[2030] , 
        \DataPath/RF/bus_reg_dataout[2029] , 
        \DataPath/RF/bus_reg_dataout[2028] , 
        \DataPath/RF/bus_reg_dataout[2027] , 
        \DataPath/RF/bus_reg_dataout[2026] , 
        \DataPath/RF/bus_reg_dataout[2025] , 
        \DataPath/RF/bus_reg_dataout[2024] , 
        \DataPath/RF/bus_reg_dataout[2023] , 
        \DataPath/RF/bus_reg_dataout[2022] , 
        \DataPath/RF/bus_reg_dataout[2021] , 
        \DataPath/RF/bus_reg_dataout[2020] , 
        \DataPath/RF/bus_reg_dataout[2019] , 
        \DataPath/RF/bus_reg_dataout[2018] , 
        \DataPath/RF/bus_reg_dataout[2017] , 
        \DataPath/RF/bus_reg_dataout[2016] , 
        \DataPath/RF/bus_reg_dataout[2015] , 
        \DataPath/RF/bus_reg_dataout[2014] , 
        \DataPath/RF/bus_reg_dataout[2013] , 
        \DataPath/RF/bus_reg_dataout[2012] , 
        \DataPath/RF/bus_reg_dataout[2011] , 
        \DataPath/RF/bus_reg_dataout[2010] , 
        \DataPath/RF/bus_reg_dataout[2009] , 
        \DataPath/RF/bus_reg_dataout[2008] , 
        \DataPath/RF/bus_reg_dataout[2007] , 
        \DataPath/RF/bus_reg_dataout[2006] , 
        \DataPath/RF/bus_reg_dataout[2005] , 
        \DataPath/RF/bus_reg_dataout[2004] , 
        \DataPath/RF/bus_reg_dataout[2003] , 
        \DataPath/RF/bus_reg_dataout[2002] , 
        \DataPath/RF/bus_reg_dataout[2001] , 
        \DataPath/RF/bus_reg_dataout[2000] , 
        \DataPath/RF/bus_reg_dataout[1999] , 
        \DataPath/RF/bus_reg_dataout[1998] , 
        \DataPath/RF/bus_reg_dataout[1997] , 
        \DataPath/RF/bus_reg_dataout[1996] , 
        \DataPath/RF/bus_reg_dataout[1995] , 
        \DataPath/RF/bus_reg_dataout[1994] , 
        \DataPath/RF/bus_reg_dataout[1993] , 
        \DataPath/RF/bus_reg_dataout[1992] , 
        \DataPath/RF/bus_reg_dataout[1991] , 
        \DataPath/RF/bus_reg_dataout[1990] , 
        \DataPath/RF/bus_reg_dataout[1989] , 
        \DataPath/RF/bus_reg_dataout[1988] , 
        \DataPath/RF/bus_reg_dataout[1987] , 
        \DataPath/RF/bus_reg_dataout[1986] , 
        \DataPath/RF/bus_reg_dataout[1985] , 
        \DataPath/RF/bus_reg_dataout[1984] , 
        \DataPath/RF/bus_reg_dataout[1983] , 
        \DataPath/RF/bus_reg_dataout[1982] , 
        \DataPath/RF/bus_reg_dataout[1981] , 
        \DataPath/RF/bus_reg_dataout[1980] , 
        \DataPath/RF/bus_reg_dataout[1979] , 
        \DataPath/RF/bus_reg_dataout[1978] , 
        \DataPath/RF/bus_reg_dataout[1977] , 
        \DataPath/RF/bus_reg_dataout[1976] , 
        \DataPath/RF/bus_reg_dataout[1975] , 
        \DataPath/RF/bus_reg_dataout[1974] , 
        \DataPath/RF/bus_reg_dataout[1973] , 
        \DataPath/RF/bus_reg_dataout[1972] , 
        \DataPath/RF/bus_reg_dataout[1971] , 
        \DataPath/RF/bus_reg_dataout[1970] , 
        \DataPath/RF/bus_reg_dataout[1969] , 
        \DataPath/RF/bus_reg_dataout[1968] , 
        \DataPath/RF/bus_reg_dataout[1967] , 
        \DataPath/RF/bus_reg_dataout[1966] , 
        \DataPath/RF/bus_reg_dataout[1965] , 
        \DataPath/RF/bus_reg_dataout[1964] , 
        \DataPath/RF/bus_reg_dataout[1963] , 
        \DataPath/RF/bus_reg_dataout[1962] , 
        \DataPath/RF/bus_reg_dataout[1961] , 
        \DataPath/RF/bus_reg_dataout[1960] , 
        \DataPath/RF/bus_reg_dataout[1959] , 
        \DataPath/RF/bus_reg_dataout[1958] , 
        \DataPath/RF/bus_reg_dataout[1957] , 
        \DataPath/RF/bus_reg_dataout[1956] , 
        \DataPath/RF/bus_reg_dataout[1955] , 
        \DataPath/RF/bus_reg_dataout[1954] , 
        \DataPath/RF/bus_reg_dataout[1953] , 
        \DataPath/RF/bus_reg_dataout[1952] , 
        \DataPath/RF/bus_reg_dataout[1951] , 
        \DataPath/RF/bus_reg_dataout[1950] , 
        \DataPath/RF/bus_reg_dataout[1949] , 
        \DataPath/RF/bus_reg_dataout[1948] , 
        \DataPath/RF/bus_reg_dataout[1947] , 
        \DataPath/RF/bus_reg_dataout[1946] , 
        \DataPath/RF/bus_reg_dataout[1945] , 
        \DataPath/RF/bus_reg_dataout[1944] , 
        \DataPath/RF/bus_reg_dataout[1943] , 
        \DataPath/RF/bus_reg_dataout[1942] , 
        \DataPath/RF/bus_reg_dataout[1941] , 
        \DataPath/RF/bus_reg_dataout[1940] , 
        \DataPath/RF/bus_reg_dataout[1939] , 
        \DataPath/RF/bus_reg_dataout[1938] , 
        \DataPath/RF/bus_reg_dataout[1937] , 
        \DataPath/RF/bus_reg_dataout[1936] , 
        \DataPath/RF/bus_reg_dataout[1935] , 
        \DataPath/RF/bus_reg_dataout[1934] , 
        \DataPath/RF/bus_reg_dataout[1933] , 
        \DataPath/RF/bus_reg_dataout[1932] , 
        \DataPath/RF/bus_reg_dataout[1931] , 
        \DataPath/RF/bus_reg_dataout[1930] , 
        \DataPath/RF/bus_reg_dataout[1929] , 
        \DataPath/RF/bus_reg_dataout[1928] , 
        \DataPath/RF/bus_reg_dataout[1927] , 
        \DataPath/RF/bus_reg_dataout[1926] , 
        \DataPath/RF/bus_reg_dataout[1925] , 
        \DataPath/RF/bus_reg_dataout[1924] , 
        \DataPath/RF/bus_reg_dataout[1923] , 
        \DataPath/RF/bus_reg_dataout[1922] , 
        \DataPath/RF/bus_reg_dataout[1921] , 
        \DataPath/RF/bus_reg_dataout[1920] , 
        \DataPath/RF/bus_reg_dataout[1919] , 
        \DataPath/RF/bus_reg_dataout[1918] , 
        \DataPath/RF/bus_reg_dataout[1917] , 
        \DataPath/RF/bus_reg_dataout[1916] , 
        \DataPath/RF/bus_reg_dataout[1915] , 
        \DataPath/RF/bus_reg_dataout[1914] , 
        \DataPath/RF/bus_reg_dataout[1913] , 
        \DataPath/RF/bus_reg_dataout[1912] , 
        \DataPath/RF/bus_reg_dataout[1911] , 
        \DataPath/RF/bus_reg_dataout[1910] , 
        \DataPath/RF/bus_reg_dataout[1909] , 
        \DataPath/RF/bus_reg_dataout[1908] , 
        \DataPath/RF/bus_reg_dataout[1907] , 
        \DataPath/RF/bus_reg_dataout[1906] , 
        \DataPath/RF/bus_reg_dataout[1905] , 
        \DataPath/RF/bus_reg_dataout[1904] , 
        \DataPath/RF/bus_reg_dataout[1903] , 
        \DataPath/RF/bus_reg_dataout[1902] , 
        \DataPath/RF/bus_reg_dataout[1901] , 
        \DataPath/RF/bus_reg_dataout[1900] , 
        \DataPath/RF/bus_reg_dataout[1899] , 
        \DataPath/RF/bus_reg_dataout[1898] , 
        \DataPath/RF/bus_reg_dataout[1897] , 
        \DataPath/RF/bus_reg_dataout[1896] , 
        \DataPath/RF/bus_reg_dataout[1895] , 
        \DataPath/RF/bus_reg_dataout[1894] , 
        \DataPath/RF/bus_reg_dataout[1893] , 
        \DataPath/RF/bus_reg_dataout[1892] , 
        \DataPath/RF/bus_reg_dataout[1891] , 
        \DataPath/RF/bus_reg_dataout[1890] , 
        \DataPath/RF/bus_reg_dataout[1889] , 
        \DataPath/RF/bus_reg_dataout[1888] , 
        \DataPath/RF/bus_reg_dataout[1887] , 
        \DataPath/RF/bus_reg_dataout[1886] , 
        \DataPath/RF/bus_reg_dataout[1885] , 
        \DataPath/RF/bus_reg_dataout[1884] , 
        \DataPath/RF/bus_reg_dataout[1883] , 
        \DataPath/RF/bus_reg_dataout[1882] , 
        \DataPath/RF/bus_reg_dataout[1881] , 
        \DataPath/RF/bus_reg_dataout[1880] , 
        \DataPath/RF/bus_reg_dataout[1879] , 
        \DataPath/RF/bus_reg_dataout[1878] , 
        \DataPath/RF/bus_reg_dataout[1877] , 
        \DataPath/RF/bus_reg_dataout[1876] , 
        \DataPath/RF/bus_reg_dataout[1875] , 
        \DataPath/RF/bus_reg_dataout[1874] , 
        \DataPath/RF/bus_reg_dataout[1873] , 
        \DataPath/RF/bus_reg_dataout[1872] , 
        \DataPath/RF/bus_reg_dataout[1871] , 
        \DataPath/RF/bus_reg_dataout[1870] , 
        \DataPath/RF/bus_reg_dataout[1869] , 
        \DataPath/RF/bus_reg_dataout[1868] , 
        \DataPath/RF/bus_reg_dataout[1867] , 
        \DataPath/RF/bus_reg_dataout[1866] , 
        \DataPath/RF/bus_reg_dataout[1865] , 
        \DataPath/RF/bus_reg_dataout[1864] , 
        \DataPath/RF/bus_reg_dataout[1863] , 
        \DataPath/RF/bus_reg_dataout[1862] , 
        \DataPath/RF/bus_reg_dataout[1861] , 
        \DataPath/RF/bus_reg_dataout[1860] , 
        \DataPath/RF/bus_reg_dataout[1859] , 
        \DataPath/RF/bus_reg_dataout[1858] , 
        \DataPath/RF/bus_reg_dataout[1857] , 
        \DataPath/RF/bus_reg_dataout[1856] , 
        \DataPath/RF/bus_reg_dataout[1855] , 
        \DataPath/RF/bus_reg_dataout[1854] , 
        \DataPath/RF/bus_reg_dataout[1853] , 
        \DataPath/RF/bus_reg_dataout[1852] , 
        \DataPath/RF/bus_reg_dataout[1851] , 
        \DataPath/RF/bus_reg_dataout[1850] , 
        \DataPath/RF/bus_reg_dataout[1849] , 
        \DataPath/RF/bus_reg_dataout[1848] , 
        \DataPath/RF/bus_reg_dataout[1847] , 
        \DataPath/RF/bus_reg_dataout[1846] , 
        \DataPath/RF/bus_reg_dataout[1845] , 
        \DataPath/RF/bus_reg_dataout[1844] , 
        \DataPath/RF/bus_reg_dataout[1843] , 
        \DataPath/RF/bus_reg_dataout[1842] , 
        \DataPath/RF/bus_reg_dataout[1841] , 
        \DataPath/RF/bus_reg_dataout[1840] , 
        \DataPath/RF/bus_reg_dataout[1839] , 
        \DataPath/RF/bus_reg_dataout[1838] , 
        \DataPath/RF/bus_reg_dataout[1837] , 
        \DataPath/RF/bus_reg_dataout[1836] , 
        \DataPath/RF/bus_reg_dataout[1835] , 
        \DataPath/RF/bus_reg_dataout[1834] , 
        \DataPath/RF/bus_reg_dataout[1833] , 
        \DataPath/RF/bus_reg_dataout[1832] , 
        \DataPath/RF/bus_reg_dataout[1831] , 
        \DataPath/RF/bus_reg_dataout[1830] , 
        \DataPath/RF/bus_reg_dataout[1829] , 
        \DataPath/RF/bus_reg_dataout[1828] , 
        \DataPath/RF/bus_reg_dataout[1827] , 
        \DataPath/RF/bus_reg_dataout[1826] , 
        \DataPath/RF/bus_reg_dataout[1825] , 
        \DataPath/RF/bus_reg_dataout[1824] , 
        \DataPath/RF/bus_reg_dataout[1823] , 
        \DataPath/RF/bus_reg_dataout[1822] , 
        \DataPath/RF/bus_reg_dataout[1821] , 
        \DataPath/RF/bus_reg_dataout[1820] , 
        \DataPath/RF/bus_reg_dataout[1819] , 
        \DataPath/RF/bus_reg_dataout[1818] , 
        \DataPath/RF/bus_reg_dataout[1817] , 
        \DataPath/RF/bus_reg_dataout[1816] , 
        \DataPath/RF/bus_reg_dataout[1815] , 
        \DataPath/RF/bus_reg_dataout[1814] , 
        \DataPath/RF/bus_reg_dataout[1813] , 
        \DataPath/RF/bus_reg_dataout[1812] , 
        \DataPath/RF/bus_reg_dataout[1811] , 
        \DataPath/RF/bus_reg_dataout[1810] , 
        \DataPath/RF/bus_reg_dataout[1809] , 
        \DataPath/RF/bus_reg_dataout[1808] , 
        \DataPath/RF/bus_reg_dataout[1807] , 
        \DataPath/RF/bus_reg_dataout[1806] , 
        \DataPath/RF/bus_reg_dataout[1805] , 
        \DataPath/RF/bus_reg_dataout[1804] , 
        \DataPath/RF/bus_reg_dataout[1803] , 
        \DataPath/RF/bus_reg_dataout[1802] , 
        \DataPath/RF/bus_reg_dataout[1801] , 
        \DataPath/RF/bus_reg_dataout[1800] , 
        \DataPath/RF/bus_reg_dataout[1799] , 
        \DataPath/RF/bus_reg_dataout[1798] , 
        \DataPath/RF/bus_reg_dataout[1797] , 
        \DataPath/RF/bus_reg_dataout[1796] , 
        \DataPath/RF/bus_reg_dataout[1795] , 
        \DataPath/RF/bus_reg_dataout[1794] , 
        \DataPath/RF/bus_reg_dataout[1793] , 
        \DataPath/RF/bus_reg_dataout[1792] , 
        \DataPath/RF/bus_reg_dataout[1791] , 
        \DataPath/RF/bus_reg_dataout[1790] , 
        \DataPath/RF/bus_reg_dataout[1789] , 
        \DataPath/RF/bus_reg_dataout[1788] , 
        \DataPath/RF/bus_reg_dataout[1787] , 
        \DataPath/RF/bus_reg_dataout[1786] , 
        \DataPath/RF/bus_reg_dataout[1785] , 
        \DataPath/RF/bus_reg_dataout[1784] , 
        \DataPath/RF/bus_reg_dataout[1783] , 
        \DataPath/RF/bus_reg_dataout[1782] , 
        \DataPath/RF/bus_reg_dataout[1781] , 
        \DataPath/RF/bus_reg_dataout[1780] , 
        \DataPath/RF/bus_reg_dataout[1779] , 
        \DataPath/RF/bus_reg_dataout[1778] , 
        \DataPath/RF/bus_reg_dataout[1777] , 
        \DataPath/RF/bus_reg_dataout[1776] , 
        \DataPath/RF/bus_reg_dataout[1775] , 
        \DataPath/RF/bus_reg_dataout[1774] , 
        \DataPath/RF/bus_reg_dataout[1773] , 
        \DataPath/RF/bus_reg_dataout[1772] , 
        \DataPath/RF/bus_reg_dataout[1771] , 
        \DataPath/RF/bus_reg_dataout[1770] , 
        \DataPath/RF/bus_reg_dataout[1769] , 
        \DataPath/RF/bus_reg_dataout[1768] , 
        \DataPath/RF/bus_reg_dataout[1767] , 
        \DataPath/RF/bus_reg_dataout[1766] , 
        \DataPath/RF/bus_reg_dataout[1765] , 
        \DataPath/RF/bus_reg_dataout[1764] , 
        \DataPath/RF/bus_reg_dataout[1763] , 
        \DataPath/RF/bus_reg_dataout[1762] , 
        \DataPath/RF/bus_reg_dataout[1761] , 
        \DataPath/RF/bus_reg_dataout[1760] , 
        \DataPath/RF/bus_reg_dataout[1759] , 
        \DataPath/RF/bus_reg_dataout[1758] , 
        \DataPath/RF/bus_reg_dataout[1757] , 
        \DataPath/RF/bus_reg_dataout[1756] , 
        \DataPath/RF/bus_reg_dataout[1755] , 
        \DataPath/RF/bus_reg_dataout[1754] , 
        \DataPath/RF/bus_reg_dataout[1753] , 
        \DataPath/RF/bus_reg_dataout[1752] , 
        \DataPath/RF/bus_reg_dataout[1751] , 
        \DataPath/RF/bus_reg_dataout[1750] , 
        \DataPath/RF/bus_reg_dataout[1749] , 
        \DataPath/RF/bus_reg_dataout[1748] , 
        \DataPath/RF/bus_reg_dataout[1747] , 
        \DataPath/RF/bus_reg_dataout[1746] , 
        \DataPath/RF/bus_reg_dataout[1745] , 
        \DataPath/RF/bus_reg_dataout[1744] , 
        \DataPath/RF/bus_reg_dataout[1743] , 
        \DataPath/RF/bus_reg_dataout[1742] , 
        \DataPath/RF/bus_reg_dataout[1741] , 
        \DataPath/RF/bus_reg_dataout[1740] , 
        \DataPath/RF/bus_reg_dataout[1739] , 
        \DataPath/RF/bus_reg_dataout[1738] , 
        \DataPath/RF/bus_reg_dataout[1737] , 
        \DataPath/RF/bus_reg_dataout[1736] , 
        \DataPath/RF/bus_reg_dataout[1735] , 
        \DataPath/RF/bus_reg_dataout[1734] , 
        \DataPath/RF/bus_reg_dataout[1733] , 
        \DataPath/RF/bus_reg_dataout[1732] , 
        \DataPath/RF/bus_reg_dataout[1731] , 
        \DataPath/RF/bus_reg_dataout[1730] , 
        \DataPath/RF/bus_reg_dataout[1729] , 
        \DataPath/RF/bus_reg_dataout[1728] , 
        \DataPath/RF/bus_reg_dataout[1727] , 
        \DataPath/RF/bus_reg_dataout[1726] , 
        \DataPath/RF/bus_reg_dataout[1725] , 
        \DataPath/RF/bus_reg_dataout[1724] , 
        \DataPath/RF/bus_reg_dataout[1723] , 
        \DataPath/RF/bus_reg_dataout[1722] , 
        \DataPath/RF/bus_reg_dataout[1721] , 
        \DataPath/RF/bus_reg_dataout[1720] , 
        \DataPath/RF/bus_reg_dataout[1719] , 
        \DataPath/RF/bus_reg_dataout[1718] , 
        \DataPath/RF/bus_reg_dataout[1717] , 
        \DataPath/RF/bus_reg_dataout[1716] , 
        \DataPath/RF/bus_reg_dataout[1715] , 
        \DataPath/RF/bus_reg_dataout[1714] , 
        \DataPath/RF/bus_reg_dataout[1713] , 
        \DataPath/RF/bus_reg_dataout[1712] , 
        \DataPath/RF/bus_reg_dataout[1711] , 
        \DataPath/RF/bus_reg_dataout[1710] , 
        \DataPath/RF/bus_reg_dataout[1709] , 
        \DataPath/RF/bus_reg_dataout[1708] , 
        \DataPath/RF/bus_reg_dataout[1707] , 
        \DataPath/RF/bus_reg_dataout[1706] , 
        \DataPath/RF/bus_reg_dataout[1705] , 
        \DataPath/RF/bus_reg_dataout[1704] , 
        \DataPath/RF/bus_reg_dataout[1703] , 
        \DataPath/RF/bus_reg_dataout[1702] , 
        \DataPath/RF/bus_reg_dataout[1701] , 
        \DataPath/RF/bus_reg_dataout[1700] , 
        \DataPath/RF/bus_reg_dataout[1699] , 
        \DataPath/RF/bus_reg_dataout[1698] , 
        \DataPath/RF/bus_reg_dataout[1697] , 
        \DataPath/RF/bus_reg_dataout[1696] , 
        \DataPath/RF/bus_reg_dataout[1695] , 
        \DataPath/RF/bus_reg_dataout[1694] , 
        \DataPath/RF/bus_reg_dataout[1693] , 
        \DataPath/RF/bus_reg_dataout[1692] , 
        \DataPath/RF/bus_reg_dataout[1691] , 
        \DataPath/RF/bus_reg_dataout[1690] , 
        \DataPath/RF/bus_reg_dataout[1689] , 
        \DataPath/RF/bus_reg_dataout[1688] , 
        \DataPath/RF/bus_reg_dataout[1687] , 
        \DataPath/RF/bus_reg_dataout[1686] , 
        \DataPath/RF/bus_reg_dataout[1685] , 
        \DataPath/RF/bus_reg_dataout[1684] , 
        \DataPath/RF/bus_reg_dataout[1683] , 
        \DataPath/RF/bus_reg_dataout[1682] , 
        \DataPath/RF/bus_reg_dataout[1681] , 
        \DataPath/RF/bus_reg_dataout[1680] , 
        \DataPath/RF/bus_reg_dataout[1679] , 
        \DataPath/RF/bus_reg_dataout[1678] , 
        \DataPath/RF/bus_reg_dataout[1677] , 
        \DataPath/RF/bus_reg_dataout[1676] , 
        \DataPath/RF/bus_reg_dataout[1675] , 
        \DataPath/RF/bus_reg_dataout[1674] , 
        \DataPath/RF/bus_reg_dataout[1673] , 
        \DataPath/RF/bus_reg_dataout[1672] , 
        \DataPath/RF/bus_reg_dataout[1671] , 
        \DataPath/RF/bus_reg_dataout[1670] , 
        \DataPath/RF/bus_reg_dataout[1669] , 
        \DataPath/RF/bus_reg_dataout[1668] , 
        \DataPath/RF/bus_reg_dataout[1667] , 
        \DataPath/RF/bus_reg_dataout[1666] , 
        \DataPath/RF/bus_reg_dataout[1665] , 
        \DataPath/RF/bus_reg_dataout[1664] , 
        \DataPath/RF/bus_reg_dataout[1663] , 
        \DataPath/RF/bus_reg_dataout[1662] , 
        \DataPath/RF/bus_reg_dataout[1661] , 
        \DataPath/RF/bus_reg_dataout[1660] , 
        \DataPath/RF/bus_reg_dataout[1659] , 
        \DataPath/RF/bus_reg_dataout[1658] , 
        \DataPath/RF/bus_reg_dataout[1657] , 
        \DataPath/RF/bus_reg_dataout[1656] , 
        \DataPath/RF/bus_reg_dataout[1655] , 
        \DataPath/RF/bus_reg_dataout[1654] , 
        \DataPath/RF/bus_reg_dataout[1653] , 
        \DataPath/RF/bus_reg_dataout[1652] , 
        \DataPath/RF/bus_reg_dataout[1651] , 
        \DataPath/RF/bus_reg_dataout[1650] , 
        \DataPath/RF/bus_reg_dataout[1649] , 
        \DataPath/RF/bus_reg_dataout[1648] , 
        \DataPath/RF/bus_reg_dataout[1647] , 
        \DataPath/RF/bus_reg_dataout[1646] , 
        \DataPath/RF/bus_reg_dataout[1645] , 
        \DataPath/RF/bus_reg_dataout[1644] , 
        \DataPath/RF/bus_reg_dataout[1643] , 
        \DataPath/RF/bus_reg_dataout[1642] , 
        \DataPath/RF/bus_reg_dataout[1641] , 
        \DataPath/RF/bus_reg_dataout[1640] , 
        \DataPath/RF/bus_reg_dataout[1639] , 
        \DataPath/RF/bus_reg_dataout[1638] , 
        \DataPath/RF/bus_reg_dataout[1637] , 
        \DataPath/RF/bus_reg_dataout[1636] , 
        \DataPath/RF/bus_reg_dataout[1635] , 
        \DataPath/RF/bus_reg_dataout[1634] , 
        \DataPath/RF/bus_reg_dataout[1633] , 
        \DataPath/RF/bus_reg_dataout[1632] , 
        \DataPath/RF/bus_reg_dataout[1631] , 
        \DataPath/RF/bus_reg_dataout[1630] , 
        \DataPath/RF/bus_reg_dataout[1629] , 
        \DataPath/RF/bus_reg_dataout[1628] , 
        \DataPath/RF/bus_reg_dataout[1627] , 
        \DataPath/RF/bus_reg_dataout[1626] , 
        \DataPath/RF/bus_reg_dataout[1625] , 
        \DataPath/RF/bus_reg_dataout[1624] , 
        \DataPath/RF/bus_reg_dataout[1623] , 
        \DataPath/RF/bus_reg_dataout[1622] , 
        \DataPath/RF/bus_reg_dataout[1621] , 
        \DataPath/RF/bus_reg_dataout[1620] , 
        \DataPath/RF/bus_reg_dataout[1619] , 
        \DataPath/RF/bus_reg_dataout[1618] , 
        \DataPath/RF/bus_reg_dataout[1617] , 
        \DataPath/RF/bus_reg_dataout[1616] , 
        \DataPath/RF/bus_reg_dataout[1615] , 
        \DataPath/RF/bus_reg_dataout[1614] , 
        \DataPath/RF/bus_reg_dataout[1613] , 
        \DataPath/RF/bus_reg_dataout[1612] , 
        \DataPath/RF/bus_reg_dataout[1611] , 
        \DataPath/RF/bus_reg_dataout[1610] , 
        \DataPath/RF/bus_reg_dataout[1609] , 
        \DataPath/RF/bus_reg_dataout[1608] , 
        \DataPath/RF/bus_reg_dataout[1607] , 
        \DataPath/RF/bus_reg_dataout[1606] , 
        \DataPath/RF/bus_reg_dataout[1605] , 
        \DataPath/RF/bus_reg_dataout[1604] , 
        \DataPath/RF/bus_reg_dataout[1603] , 
        \DataPath/RF/bus_reg_dataout[1602] , 
        \DataPath/RF/bus_reg_dataout[1601] , 
        \DataPath/RF/bus_reg_dataout[1600] , 
        \DataPath/RF/bus_reg_dataout[1599] , 
        \DataPath/RF/bus_reg_dataout[1598] , 
        \DataPath/RF/bus_reg_dataout[1597] , 
        \DataPath/RF/bus_reg_dataout[1596] , 
        \DataPath/RF/bus_reg_dataout[1595] , 
        \DataPath/RF/bus_reg_dataout[1594] , 
        \DataPath/RF/bus_reg_dataout[1593] , 
        \DataPath/RF/bus_reg_dataout[1592] , 
        \DataPath/RF/bus_reg_dataout[1591] , 
        \DataPath/RF/bus_reg_dataout[1590] , 
        \DataPath/RF/bus_reg_dataout[1589] , 
        \DataPath/RF/bus_reg_dataout[1588] , 
        \DataPath/RF/bus_reg_dataout[1587] , 
        \DataPath/RF/bus_reg_dataout[1586] , 
        \DataPath/RF/bus_reg_dataout[1585] , 
        \DataPath/RF/bus_reg_dataout[1584] , 
        \DataPath/RF/bus_reg_dataout[1583] , 
        \DataPath/RF/bus_reg_dataout[1582] , 
        \DataPath/RF/bus_reg_dataout[1581] , 
        \DataPath/RF/bus_reg_dataout[1580] , 
        \DataPath/RF/bus_reg_dataout[1579] , 
        \DataPath/RF/bus_reg_dataout[1578] , 
        \DataPath/RF/bus_reg_dataout[1577] , 
        \DataPath/RF/bus_reg_dataout[1576] , 
        \DataPath/RF/bus_reg_dataout[1575] , 
        \DataPath/RF/bus_reg_dataout[1574] , 
        \DataPath/RF/bus_reg_dataout[1573] , 
        \DataPath/RF/bus_reg_dataout[1572] , 
        \DataPath/RF/bus_reg_dataout[1571] , 
        \DataPath/RF/bus_reg_dataout[1570] , 
        \DataPath/RF/bus_reg_dataout[1569] , 
        \DataPath/RF/bus_reg_dataout[1568] , 
        \DataPath/RF/bus_reg_dataout[1567] , 
        \DataPath/RF/bus_reg_dataout[1566] , 
        \DataPath/RF/bus_reg_dataout[1565] , 
        \DataPath/RF/bus_reg_dataout[1564] , 
        \DataPath/RF/bus_reg_dataout[1563] , 
        \DataPath/RF/bus_reg_dataout[1562] , 
        \DataPath/RF/bus_reg_dataout[1561] , 
        \DataPath/RF/bus_reg_dataout[1560] , 
        \DataPath/RF/bus_reg_dataout[1559] , 
        \DataPath/RF/bus_reg_dataout[1558] , 
        \DataPath/RF/bus_reg_dataout[1557] , 
        \DataPath/RF/bus_reg_dataout[1556] , 
        \DataPath/RF/bus_reg_dataout[1555] , 
        \DataPath/RF/bus_reg_dataout[1554] , 
        \DataPath/RF/bus_reg_dataout[1553] , 
        \DataPath/RF/bus_reg_dataout[1552] , 
        \DataPath/RF/bus_reg_dataout[1551] , 
        \DataPath/RF/bus_reg_dataout[1550] , 
        \DataPath/RF/bus_reg_dataout[1549] , 
        \DataPath/RF/bus_reg_dataout[1548] , 
        \DataPath/RF/bus_reg_dataout[1547] , 
        \DataPath/RF/bus_reg_dataout[1546] , 
        \DataPath/RF/bus_reg_dataout[1545] , 
        \DataPath/RF/bus_reg_dataout[1544] , 
        \DataPath/RF/bus_reg_dataout[1543] , 
        \DataPath/RF/bus_reg_dataout[1542] , 
        \DataPath/RF/bus_reg_dataout[1541] , 
        \DataPath/RF/bus_reg_dataout[1540] , 
        \DataPath/RF/bus_reg_dataout[1539] , 
        \DataPath/RF/bus_reg_dataout[1538] , 
        \DataPath/RF/bus_reg_dataout[1537] , 
        \DataPath/RF/bus_reg_dataout[1536] , 
        \DataPath/RF/bus_reg_dataout[1535] , 
        \DataPath/RF/bus_reg_dataout[1534] , 
        \DataPath/RF/bus_reg_dataout[1533] , 
        \DataPath/RF/bus_reg_dataout[1532] , 
        \DataPath/RF/bus_reg_dataout[1531] , 
        \DataPath/RF/bus_reg_dataout[1530] , 
        \DataPath/RF/bus_reg_dataout[1529] , 
        \DataPath/RF/bus_reg_dataout[1528] , 
        \DataPath/RF/bus_reg_dataout[1527] , 
        \DataPath/RF/bus_reg_dataout[1526] , 
        \DataPath/RF/bus_reg_dataout[1525] , 
        \DataPath/RF/bus_reg_dataout[1524] , 
        \DataPath/RF/bus_reg_dataout[1523] , 
        \DataPath/RF/bus_reg_dataout[1522] , 
        \DataPath/RF/bus_reg_dataout[1521] , 
        \DataPath/RF/bus_reg_dataout[1520] , 
        \DataPath/RF/bus_reg_dataout[1519] , 
        \DataPath/RF/bus_reg_dataout[1518] , 
        \DataPath/RF/bus_reg_dataout[1517] , 
        \DataPath/RF/bus_reg_dataout[1516] , 
        \DataPath/RF/bus_reg_dataout[1515] , 
        \DataPath/RF/bus_reg_dataout[1514] , 
        \DataPath/RF/bus_reg_dataout[1513] , 
        \DataPath/RF/bus_reg_dataout[1512] , 
        \DataPath/RF/bus_reg_dataout[1511] , 
        \DataPath/RF/bus_reg_dataout[1510] , 
        \DataPath/RF/bus_reg_dataout[1509] , 
        \DataPath/RF/bus_reg_dataout[1508] , 
        \DataPath/RF/bus_reg_dataout[1507] , 
        \DataPath/RF/bus_reg_dataout[1506] , 
        \DataPath/RF/bus_reg_dataout[1505] , 
        \DataPath/RF/bus_reg_dataout[1504] , 
        \DataPath/RF/bus_reg_dataout[1503] , 
        \DataPath/RF/bus_reg_dataout[1502] , 
        \DataPath/RF/bus_reg_dataout[1501] , 
        \DataPath/RF/bus_reg_dataout[1500] , 
        \DataPath/RF/bus_reg_dataout[1499] , 
        \DataPath/RF/bus_reg_dataout[1498] , 
        \DataPath/RF/bus_reg_dataout[1497] , 
        \DataPath/RF/bus_reg_dataout[1496] , 
        \DataPath/RF/bus_reg_dataout[1495] , 
        \DataPath/RF/bus_reg_dataout[1494] , 
        \DataPath/RF/bus_reg_dataout[1493] , 
        \DataPath/RF/bus_reg_dataout[1492] , 
        \DataPath/RF/bus_reg_dataout[1491] , 
        \DataPath/RF/bus_reg_dataout[1490] , 
        \DataPath/RF/bus_reg_dataout[1489] , 
        \DataPath/RF/bus_reg_dataout[1488] , 
        \DataPath/RF/bus_reg_dataout[1487] , 
        \DataPath/RF/bus_reg_dataout[1486] , 
        \DataPath/RF/bus_reg_dataout[1485] , 
        \DataPath/RF/bus_reg_dataout[1484] , 
        \DataPath/RF/bus_reg_dataout[1483] , 
        \DataPath/RF/bus_reg_dataout[1482] , 
        \DataPath/RF/bus_reg_dataout[1481] , 
        \DataPath/RF/bus_reg_dataout[1480] , 
        \DataPath/RF/bus_reg_dataout[1479] , 
        \DataPath/RF/bus_reg_dataout[1478] , 
        \DataPath/RF/bus_reg_dataout[1477] , 
        \DataPath/RF/bus_reg_dataout[1476] , 
        \DataPath/RF/bus_reg_dataout[1475] , 
        \DataPath/RF/bus_reg_dataout[1474] , 
        \DataPath/RF/bus_reg_dataout[1473] , 
        \DataPath/RF/bus_reg_dataout[1472] , 
        \DataPath/RF/bus_reg_dataout[1471] , 
        \DataPath/RF/bus_reg_dataout[1470] , 
        \DataPath/RF/bus_reg_dataout[1469] , 
        \DataPath/RF/bus_reg_dataout[1468] , 
        \DataPath/RF/bus_reg_dataout[1467] , 
        \DataPath/RF/bus_reg_dataout[1466] , 
        \DataPath/RF/bus_reg_dataout[1465] , 
        \DataPath/RF/bus_reg_dataout[1464] , 
        \DataPath/RF/bus_reg_dataout[1463] , 
        \DataPath/RF/bus_reg_dataout[1462] , 
        \DataPath/RF/bus_reg_dataout[1461] , 
        \DataPath/RF/bus_reg_dataout[1460] , 
        \DataPath/RF/bus_reg_dataout[1459] , 
        \DataPath/RF/bus_reg_dataout[1458] , 
        \DataPath/RF/bus_reg_dataout[1457] , 
        \DataPath/RF/bus_reg_dataout[1456] , 
        \DataPath/RF/bus_reg_dataout[1455] , 
        \DataPath/RF/bus_reg_dataout[1454] , 
        \DataPath/RF/bus_reg_dataout[1453] , 
        \DataPath/RF/bus_reg_dataout[1452] , 
        \DataPath/RF/bus_reg_dataout[1451] , 
        \DataPath/RF/bus_reg_dataout[1450] , 
        \DataPath/RF/bus_reg_dataout[1449] , 
        \DataPath/RF/bus_reg_dataout[1448] , 
        \DataPath/RF/bus_reg_dataout[1447] , 
        \DataPath/RF/bus_reg_dataout[1446] , 
        \DataPath/RF/bus_reg_dataout[1445] , 
        \DataPath/RF/bus_reg_dataout[1444] , 
        \DataPath/RF/bus_reg_dataout[1443] , 
        \DataPath/RF/bus_reg_dataout[1442] , 
        \DataPath/RF/bus_reg_dataout[1441] , 
        \DataPath/RF/bus_reg_dataout[1440] , 
        \DataPath/RF/bus_reg_dataout[1439] , 
        \DataPath/RF/bus_reg_dataout[1438] , 
        \DataPath/RF/bus_reg_dataout[1437] , 
        \DataPath/RF/bus_reg_dataout[1436] , 
        \DataPath/RF/bus_reg_dataout[1435] , 
        \DataPath/RF/bus_reg_dataout[1434] , 
        \DataPath/RF/bus_reg_dataout[1433] , 
        \DataPath/RF/bus_reg_dataout[1432] , 
        \DataPath/RF/bus_reg_dataout[1431] , 
        \DataPath/RF/bus_reg_dataout[1430] , 
        \DataPath/RF/bus_reg_dataout[1429] , 
        \DataPath/RF/bus_reg_dataout[1428] , 
        \DataPath/RF/bus_reg_dataout[1427] , 
        \DataPath/RF/bus_reg_dataout[1426] , 
        \DataPath/RF/bus_reg_dataout[1425] , 
        \DataPath/RF/bus_reg_dataout[1424] , 
        \DataPath/RF/bus_reg_dataout[1423] , 
        \DataPath/RF/bus_reg_dataout[1422] , 
        \DataPath/RF/bus_reg_dataout[1421] , 
        \DataPath/RF/bus_reg_dataout[1420] , 
        \DataPath/RF/bus_reg_dataout[1419] , 
        \DataPath/RF/bus_reg_dataout[1418] , 
        \DataPath/RF/bus_reg_dataout[1417] , 
        \DataPath/RF/bus_reg_dataout[1416] , 
        \DataPath/RF/bus_reg_dataout[1415] , 
        \DataPath/RF/bus_reg_dataout[1414] , 
        \DataPath/RF/bus_reg_dataout[1413] , 
        \DataPath/RF/bus_reg_dataout[1412] , 
        \DataPath/RF/bus_reg_dataout[1411] , 
        \DataPath/RF/bus_reg_dataout[1410] , 
        \DataPath/RF/bus_reg_dataout[1409] , 
        \DataPath/RF/bus_reg_dataout[1408] , 
        \DataPath/RF/bus_reg_dataout[1407] , 
        \DataPath/RF/bus_reg_dataout[1406] , 
        \DataPath/RF/bus_reg_dataout[1405] , 
        \DataPath/RF/bus_reg_dataout[1404] , 
        \DataPath/RF/bus_reg_dataout[1403] , 
        \DataPath/RF/bus_reg_dataout[1402] , 
        \DataPath/RF/bus_reg_dataout[1401] , 
        \DataPath/RF/bus_reg_dataout[1400] , 
        \DataPath/RF/bus_reg_dataout[1399] , 
        \DataPath/RF/bus_reg_dataout[1398] , 
        \DataPath/RF/bus_reg_dataout[1397] , 
        \DataPath/RF/bus_reg_dataout[1396] , 
        \DataPath/RF/bus_reg_dataout[1395] , 
        \DataPath/RF/bus_reg_dataout[1394] , 
        \DataPath/RF/bus_reg_dataout[1393] , 
        \DataPath/RF/bus_reg_dataout[1392] , 
        \DataPath/RF/bus_reg_dataout[1391] , 
        \DataPath/RF/bus_reg_dataout[1390] , 
        \DataPath/RF/bus_reg_dataout[1389] , 
        \DataPath/RF/bus_reg_dataout[1388] , 
        \DataPath/RF/bus_reg_dataout[1387] , 
        \DataPath/RF/bus_reg_dataout[1386] , 
        \DataPath/RF/bus_reg_dataout[1385] , 
        \DataPath/RF/bus_reg_dataout[1384] , 
        \DataPath/RF/bus_reg_dataout[1383] , 
        \DataPath/RF/bus_reg_dataout[1382] , 
        \DataPath/RF/bus_reg_dataout[1381] , 
        \DataPath/RF/bus_reg_dataout[1380] , 
        \DataPath/RF/bus_reg_dataout[1379] , 
        \DataPath/RF/bus_reg_dataout[1378] , 
        \DataPath/RF/bus_reg_dataout[1377] , 
        \DataPath/RF/bus_reg_dataout[1376] , 
        \DataPath/RF/bus_reg_dataout[1375] , 
        \DataPath/RF/bus_reg_dataout[1374] , 
        \DataPath/RF/bus_reg_dataout[1373] , 
        \DataPath/RF/bus_reg_dataout[1372] , 
        \DataPath/RF/bus_reg_dataout[1371] , 
        \DataPath/RF/bus_reg_dataout[1370] , 
        \DataPath/RF/bus_reg_dataout[1369] , 
        \DataPath/RF/bus_reg_dataout[1368] , 
        \DataPath/RF/bus_reg_dataout[1367] , 
        \DataPath/RF/bus_reg_dataout[1366] , 
        \DataPath/RF/bus_reg_dataout[1365] , 
        \DataPath/RF/bus_reg_dataout[1364] , 
        \DataPath/RF/bus_reg_dataout[1363] , 
        \DataPath/RF/bus_reg_dataout[1362] , 
        \DataPath/RF/bus_reg_dataout[1361] , 
        \DataPath/RF/bus_reg_dataout[1360] , 
        \DataPath/RF/bus_reg_dataout[1359] , 
        \DataPath/RF/bus_reg_dataout[1358] , 
        \DataPath/RF/bus_reg_dataout[1357] , 
        \DataPath/RF/bus_reg_dataout[1356] , 
        \DataPath/RF/bus_reg_dataout[1355] , 
        \DataPath/RF/bus_reg_dataout[1354] , 
        \DataPath/RF/bus_reg_dataout[1353] , 
        \DataPath/RF/bus_reg_dataout[1352] , 
        \DataPath/RF/bus_reg_dataout[1351] , 
        \DataPath/RF/bus_reg_dataout[1350] , 
        \DataPath/RF/bus_reg_dataout[1349] , 
        \DataPath/RF/bus_reg_dataout[1348] , 
        \DataPath/RF/bus_reg_dataout[1347] , 
        \DataPath/RF/bus_reg_dataout[1346] , 
        \DataPath/RF/bus_reg_dataout[1345] , 
        \DataPath/RF/bus_reg_dataout[1344] , 
        \DataPath/RF/bus_reg_dataout[1343] , 
        \DataPath/RF/bus_reg_dataout[1342] , 
        \DataPath/RF/bus_reg_dataout[1341] , 
        \DataPath/RF/bus_reg_dataout[1340] , 
        \DataPath/RF/bus_reg_dataout[1339] , 
        \DataPath/RF/bus_reg_dataout[1338] , 
        \DataPath/RF/bus_reg_dataout[1337] , 
        \DataPath/RF/bus_reg_dataout[1336] , 
        \DataPath/RF/bus_reg_dataout[1335] , 
        \DataPath/RF/bus_reg_dataout[1334] , 
        \DataPath/RF/bus_reg_dataout[1333] , 
        \DataPath/RF/bus_reg_dataout[1332] , 
        \DataPath/RF/bus_reg_dataout[1331] , 
        \DataPath/RF/bus_reg_dataout[1330] , 
        \DataPath/RF/bus_reg_dataout[1329] , 
        \DataPath/RF/bus_reg_dataout[1328] , 
        \DataPath/RF/bus_reg_dataout[1327] , 
        \DataPath/RF/bus_reg_dataout[1326] , 
        \DataPath/RF/bus_reg_dataout[1325] , 
        \DataPath/RF/bus_reg_dataout[1324] , 
        \DataPath/RF/bus_reg_dataout[1323] , 
        \DataPath/RF/bus_reg_dataout[1322] , 
        \DataPath/RF/bus_reg_dataout[1321] , 
        \DataPath/RF/bus_reg_dataout[1320] , 
        \DataPath/RF/bus_reg_dataout[1319] , 
        \DataPath/RF/bus_reg_dataout[1318] , 
        \DataPath/RF/bus_reg_dataout[1317] , 
        \DataPath/RF/bus_reg_dataout[1316] , 
        \DataPath/RF/bus_reg_dataout[1315] , 
        \DataPath/RF/bus_reg_dataout[1314] , 
        \DataPath/RF/bus_reg_dataout[1313] , 
        \DataPath/RF/bus_reg_dataout[1312] , 
        \DataPath/RF/bus_reg_dataout[1311] , 
        \DataPath/RF/bus_reg_dataout[1310] , 
        \DataPath/RF/bus_reg_dataout[1309] , 
        \DataPath/RF/bus_reg_dataout[1308] , 
        \DataPath/RF/bus_reg_dataout[1307] , 
        \DataPath/RF/bus_reg_dataout[1306] , 
        \DataPath/RF/bus_reg_dataout[1305] , 
        \DataPath/RF/bus_reg_dataout[1304] , 
        \DataPath/RF/bus_reg_dataout[1303] , 
        \DataPath/RF/bus_reg_dataout[1302] , 
        \DataPath/RF/bus_reg_dataout[1301] , 
        \DataPath/RF/bus_reg_dataout[1300] , 
        \DataPath/RF/bus_reg_dataout[1299] , 
        \DataPath/RF/bus_reg_dataout[1298] , 
        \DataPath/RF/bus_reg_dataout[1297] , 
        \DataPath/RF/bus_reg_dataout[1296] , 
        \DataPath/RF/bus_reg_dataout[1295] , 
        \DataPath/RF/bus_reg_dataout[1294] , 
        \DataPath/RF/bus_reg_dataout[1293] , 
        \DataPath/RF/bus_reg_dataout[1292] , 
        \DataPath/RF/bus_reg_dataout[1291] , 
        \DataPath/RF/bus_reg_dataout[1290] , 
        \DataPath/RF/bus_reg_dataout[1289] , 
        \DataPath/RF/bus_reg_dataout[1288] , 
        \DataPath/RF/bus_reg_dataout[1287] , 
        \DataPath/RF/bus_reg_dataout[1286] , 
        \DataPath/RF/bus_reg_dataout[1285] , 
        \DataPath/RF/bus_reg_dataout[1284] , 
        \DataPath/RF/bus_reg_dataout[1283] , 
        \DataPath/RF/bus_reg_dataout[1282] , 
        \DataPath/RF/bus_reg_dataout[1281] , 
        \DataPath/RF/bus_reg_dataout[1280] , 
        \DataPath/RF/bus_reg_dataout[1279] , 
        \DataPath/RF/bus_reg_dataout[1278] , 
        \DataPath/RF/bus_reg_dataout[1277] , 
        \DataPath/RF/bus_reg_dataout[1276] , 
        \DataPath/RF/bus_reg_dataout[1275] , 
        \DataPath/RF/bus_reg_dataout[1274] , 
        \DataPath/RF/bus_reg_dataout[1273] , 
        \DataPath/RF/bus_reg_dataout[1272] , 
        \DataPath/RF/bus_reg_dataout[1271] , 
        \DataPath/RF/bus_reg_dataout[1270] , 
        \DataPath/RF/bus_reg_dataout[1269] , 
        \DataPath/RF/bus_reg_dataout[1268] , 
        \DataPath/RF/bus_reg_dataout[1267] , 
        \DataPath/RF/bus_reg_dataout[1266] , 
        \DataPath/RF/bus_reg_dataout[1265] , 
        \DataPath/RF/bus_reg_dataout[1264] , 
        \DataPath/RF/bus_reg_dataout[1263] , 
        \DataPath/RF/bus_reg_dataout[1262] , 
        \DataPath/RF/bus_reg_dataout[1261] , 
        \DataPath/RF/bus_reg_dataout[1260] , 
        \DataPath/RF/bus_reg_dataout[1259] , 
        \DataPath/RF/bus_reg_dataout[1258] , 
        \DataPath/RF/bus_reg_dataout[1257] , 
        \DataPath/RF/bus_reg_dataout[1256] , 
        \DataPath/RF/bus_reg_dataout[1255] , 
        \DataPath/RF/bus_reg_dataout[1254] , 
        \DataPath/RF/bus_reg_dataout[1253] , 
        \DataPath/RF/bus_reg_dataout[1252] , 
        \DataPath/RF/bus_reg_dataout[1251] , 
        \DataPath/RF/bus_reg_dataout[1250] , 
        \DataPath/RF/bus_reg_dataout[1249] , 
        \DataPath/RF/bus_reg_dataout[1248] , 
        \DataPath/RF/bus_reg_dataout[1247] , 
        \DataPath/RF/bus_reg_dataout[1246] , 
        \DataPath/RF/bus_reg_dataout[1245] , 
        \DataPath/RF/bus_reg_dataout[1244] , 
        \DataPath/RF/bus_reg_dataout[1243] , 
        \DataPath/RF/bus_reg_dataout[1242] , 
        \DataPath/RF/bus_reg_dataout[1241] , 
        \DataPath/RF/bus_reg_dataout[1240] , 
        \DataPath/RF/bus_reg_dataout[1239] , 
        \DataPath/RF/bus_reg_dataout[1238] , 
        \DataPath/RF/bus_reg_dataout[1237] , 
        \DataPath/RF/bus_reg_dataout[1236] , 
        \DataPath/RF/bus_reg_dataout[1235] , 
        \DataPath/RF/bus_reg_dataout[1234] , 
        \DataPath/RF/bus_reg_dataout[1233] , 
        \DataPath/RF/bus_reg_dataout[1232] , 
        \DataPath/RF/bus_reg_dataout[1231] , 
        \DataPath/RF/bus_reg_dataout[1230] , 
        \DataPath/RF/bus_reg_dataout[1229] , 
        \DataPath/RF/bus_reg_dataout[1228] , 
        \DataPath/RF/bus_reg_dataout[1227] , 
        \DataPath/RF/bus_reg_dataout[1226] , 
        \DataPath/RF/bus_reg_dataout[1225] , 
        \DataPath/RF/bus_reg_dataout[1224] , 
        \DataPath/RF/bus_reg_dataout[1223] , 
        \DataPath/RF/bus_reg_dataout[1222] , 
        \DataPath/RF/bus_reg_dataout[1221] , 
        \DataPath/RF/bus_reg_dataout[1220] , 
        \DataPath/RF/bus_reg_dataout[1219] , 
        \DataPath/RF/bus_reg_dataout[1218] , 
        \DataPath/RF/bus_reg_dataout[1217] , 
        \DataPath/RF/bus_reg_dataout[1216] , 
        \DataPath/RF/bus_reg_dataout[1215] , 
        \DataPath/RF/bus_reg_dataout[1214] , 
        \DataPath/RF/bus_reg_dataout[1213] , 
        \DataPath/RF/bus_reg_dataout[1212] , 
        \DataPath/RF/bus_reg_dataout[1211] , 
        \DataPath/RF/bus_reg_dataout[1210] , 
        \DataPath/RF/bus_reg_dataout[1209] , 
        \DataPath/RF/bus_reg_dataout[1208] , 
        \DataPath/RF/bus_reg_dataout[1207] , 
        \DataPath/RF/bus_reg_dataout[1206] , 
        \DataPath/RF/bus_reg_dataout[1205] , 
        \DataPath/RF/bus_reg_dataout[1204] , 
        \DataPath/RF/bus_reg_dataout[1203] , 
        \DataPath/RF/bus_reg_dataout[1202] , 
        \DataPath/RF/bus_reg_dataout[1201] , 
        \DataPath/RF/bus_reg_dataout[1200] , 
        \DataPath/RF/bus_reg_dataout[1199] , 
        \DataPath/RF/bus_reg_dataout[1198] , 
        \DataPath/RF/bus_reg_dataout[1197] , 
        \DataPath/RF/bus_reg_dataout[1196] , 
        \DataPath/RF/bus_reg_dataout[1195] , 
        \DataPath/RF/bus_reg_dataout[1194] , 
        \DataPath/RF/bus_reg_dataout[1193] , 
        \DataPath/RF/bus_reg_dataout[1192] , 
        \DataPath/RF/bus_reg_dataout[1191] , 
        \DataPath/RF/bus_reg_dataout[1190] , 
        \DataPath/RF/bus_reg_dataout[1189] , 
        \DataPath/RF/bus_reg_dataout[1188] , 
        \DataPath/RF/bus_reg_dataout[1187] , 
        \DataPath/RF/bus_reg_dataout[1186] , 
        \DataPath/RF/bus_reg_dataout[1185] , 
        \DataPath/RF/bus_reg_dataout[1184] , 
        \DataPath/RF/bus_reg_dataout[1183] , 
        \DataPath/RF/bus_reg_dataout[1182] , 
        \DataPath/RF/bus_reg_dataout[1181] , 
        \DataPath/RF/bus_reg_dataout[1180] , 
        \DataPath/RF/bus_reg_dataout[1179] , 
        \DataPath/RF/bus_reg_dataout[1178] , 
        \DataPath/RF/bus_reg_dataout[1177] , 
        \DataPath/RF/bus_reg_dataout[1176] , 
        \DataPath/RF/bus_reg_dataout[1175] , 
        \DataPath/RF/bus_reg_dataout[1174] , 
        \DataPath/RF/bus_reg_dataout[1173] , 
        \DataPath/RF/bus_reg_dataout[1172] , 
        \DataPath/RF/bus_reg_dataout[1171] , 
        \DataPath/RF/bus_reg_dataout[1170] , 
        \DataPath/RF/bus_reg_dataout[1169] , 
        \DataPath/RF/bus_reg_dataout[1168] , 
        \DataPath/RF/bus_reg_dataout[1167] , 
        \DataPath/RF/bus_reg_dataout[1166] , 
        \DataPath/RF/bus_reg_dataout[1165] , 
        \DataPath/RF/bus_reg_dataout[1164] , 
        \DataPath/RF/bus_reg_dataout[1163] , 
        \DataPath/RF/bus_reg_dataout[1162] , 
        \DataPath/RF/bus_reg_dataout[1161] , 
        \DataPath/RF/bus_reg_dataout[1160] , 
        \DataPath/RF/bus_reg_dataout[1159] , 
        \DataPath/RF/bus_reg_dataout[1158] , 
        \DataPath/RF/bus_reg_dataout[1157] , 
        \DataPath/RF/bus_reg_dataout[1156] , 
        \DataPath/RF/bus_reg_dataout[1155] , 
        \DataPath/RF/bus_reg_dataout[1154] , 
        \DataPath/RF/bus_reg_dataout[1153] , 
        \DataPath/RF/bus_reg_dataout[1152] , 
        \DataPath/RF/bus_reg_dataout[1151] , 
        \DataPath/RF/bus_reg_dataout[1150] , 
        \DataPath/RF/bus_reg_dataout[1149] , 
        \DataPath/RF/bus_reg_dataout[1148] , 
        \DataPath/RF/bus_reg_dataout[1147] , 
        \DataPath/RF/bus_reg_dataout[1146] , 
        \DataPath/RF/bus_reg_dataout[1145] , 
        \DataPath/RF/bus_reg_dataout[1144] , 
        \DataPath/RF/bus_reg_dataout[1143] , 
        \DataPath/RF/bus_reg_dataout[1142] , 
        \DataPath/RF/bus_reg_dataout[1141] , 
        \DataPath/RF/bus_reg_dataout[1140] , 
        \DataPath/RF/bus_reg_dataout[1139] , 
        \DataPath/RF/bus_reg_dataout[1138] , 
        \DataPath/RF/bus_reg_dataout[1137] , 
        \DataPath/RF/bus_reg_dataout[1136] , 
        \DataPath/RF/bus_reg_dataout[1135] , 
        \DataPath/RF/bus_reg_dataout[1134] , 
        \DataPath/RF/bus_reg_dataout[1133] , 
        \DataPath/RF/bus_reg_dataout[1132] , 
        \DataPath/RF/bus_reg_dataout[1131] , 
        \DataPath/RF/bus_reg_dataout[1130] , 
        \DataPath/RF/bus_reg_dataout[1129] , 
        \DataPath/RF/bus_reg_dataout[1128] , 
        \DataPath/RF/bus_reg_dataout[1127] , 
        \DataPath/RF/bus_reg_dataout[1126] , 
        \DataPath/RF/bus_reg_dataout[1125] , 
        \DataPath/RF/bus_reg_dataout[1124] , 
        \DataPath/RF/bus_reg_dataout[1123] , 
        \DataPath/RF/bus_reg_dataout[1122] , 
        \DataPath/RF/bus_reg_dataout[1121] , 
        \DataPath/RF/bus_reg_dataout[1120] , 
        \DataPath/RF/bus_reg_dataout[1119] , 
        \DataPath/RF/bus_reg_dataout[1118] , 
        \DataPath/RF/bus_reg_dataout[1117] , 
        \DataPath/RF/bus_reg_dataout[1116] , 
        \DataPath/RF/bus_reg_dataout[1115] , 
        \DataPath/RF/bus_reg_dataout[1114] , 
        \DataPath/RF/bus_reg_dataout[1113] , 
        \DataPath/RF/bus_reg_dataout[1112] , 
        \DataPath/RF/bus_reg_dataout[1111] , 
        \DataPath/RF/bus_reg_dataout[1110] , 
        \DataPath/RF/bus_reg_dataout[1109] , 
        \DataPath/RF/bus_reg_dataout[1108] , 
        \DataPath/RF/bus_reg_dataout[1107] , 
        \DataPath/RF/bus_reg_dataout[1106] , 
        \DataPath/RF/bus_reg_dataout[1105] , 
        \DataPath/RF/bus_reg_dataout[1104] , 
        \DataPath/RF/bus_reg_dataout[1103] , 
        \DataPath/RF/bus_reg_dataout[1102] , 
        \DataPath/RF/bus_reg_dataout[1101] , 
        \DataPath/RF/bus_reg_dataout[1100] , 
        \DataPath/RF/bus_reg_dataout[1099] , 
        \DataPath/RF/bus_reg_dataout[1098] , 
        \DataPath/RF/bus_reg_dataout[1097] , 
        \DataPath/RF/bus_reg_dataout[1096] , 
        \DataPath/RF/bus_reg_dataout[1095] , 
        \DataPath/RF/bus_reg_dataout[1094] , 
        \DataPath/RF/bus_reg_dataout[1093] , 
        \DataPath/RF/bus_reg_dataout[1092] , 
        \DataPath/RF/bus_reg_dataout[1091] , 
        \DataPath/RF/bus_reg_dataout[1090] , 
        \DataPath/RF/bus_reg_dataout[1089] , 
        \DataPath/RF/bus_reg_dataout[1088] , 
        \DataPath/RF/bus_reg_dataout[1087] , 
        \DataPath/RF/bus_reg_dataout[1086] , 
        \DataPath/RF/bus_reg_dataout[1085] , 
        \DataPath/RF/bus_reg_dataout[1084] , 
        \DataPath/RF/bus_reg_dataout[1083] , 
        \DataPath/RF/bus_reg_dataout[1082] , 
        \DataPath/RF/bus_reg_dataout[1081] , 
        \DataPath/RF/bus_reg_dataout[1080] , 
        \DataPath/RF/bus_reg_dataout[1079] , 
        \DataPath/RF/bus_reg_dataout[1078] , 
        \DataPath/RF/bus_reg_dataout[1077] , 
        \DataPath/RF/bus_reg_dataout[1076] , 
        \DataPath/RF/bus_reg_dataout[1075] , 
        \DataPath/RF/bus_reg_dataout[1074] , 
        \DataPath/RF/bus_reg_dataout[1073] , 
        \DataPath/RF/bus_reg_dataout[1072] , 
        \DataPath/RF/bus_reg_dataout[1071] , 
        \DataPath/RF/bus_reg_dataout[1070] , 
        \DataPath/RF/bus_reg_dataout[1069] , 
        \DataPath/RF/bus_reg_dataout[1068] , 
        \DataPath/RF/bus_reg_dataout[1067] , 
        \DataPath/RF/bus_reg_dataout[1066] , 
        \DataPath/RF/bus_reg_dataout[1065] , 
        \DataPath/RF/bus_reg_dataout[1064] , 
        \DataPath/RF/bus_reg_dataout[1063] , 
        \DataPath/RF/bus_reg_dataout[1062] , 
        \DataPath/RF/bus_reg_dataout[1061] , 
        \DataPath/RF/bus_reg_dataout[1060] , 
        \DataPath/RF/bus_reg_dataout[1059] , 
        \DataPath/RF/bus_reg_dataout[1058] , 
        \DataPath/RF/bus_reg_dataout[1057] , 
        \DataPath/RF/bus_reg_dataout[1056] , 
        \DataPath/RF/bus_reg_dataout[1055] , 
        \DataPath/RF/bus_reg_dataout[1054] , 
        \DataPath/RF/bus_reg_dataout[1053] , 
        \DataPath/RF/bus_reg_dataout[1052] , 
        \DataPath/RF/bus_reg_dataout[1051] , 
        \DataPath/RF/bus_reg_dataout[1050] , 
        \DataPath/RF/bus_reg_dataout[1049] , 
        \DataPath/RF/bus_reg_dataout[1048] , 
        \DataPath/RF/bus_reg_dataout[1047] , 
        \DataPath/RF/bus_reg_dataout[1046] , 
        \DataPath/RF/bus_reg_dataout[1045] , 
        \DataPath/RF/bus_reg_dataout[1044] , 
        \DataPath/RF/bus_reg_dataout[1043] , 
        \DataPath/RF/bus_reg_dataout[1042] , 
        \DataPath/RF/bus_reg_dataout[1041] , 
        \DataPath/RF/bus_reg_dataout[1040] , 
        \DataPath/RF/bus_reg_dataout[1039] , 
        \DataPath/RF/bus_reg_dataout[1038] , 
        \DataPath/RF/bus_reg_dataout[1037] , 
        \DataPath/RF/bus_reg_dataout[1036] , 
        \DataPath/RF/bus_reg_dataout[1035] , 
        \DataPath/RF/bus_reg_dataout[1034] , 
        \DataPath/RF/bus_reg_dataout[1033] , 
        \DataPath/RF/bus_reg_dataout[1032] , 
        \DataPath/RF/bus_reg_dataout[1031] , 
        \DataPath/RF/bus_reg_dataout[1030] , 
        \DataPath/RF/bus_reg_dataout[1029] , 
        \DataPath/RF/bus_reg_dataout[1028] , 
        \DataPath/RF/bus_reg_dataout[1027] , 
        \DataPath/RF/bus_reg_dataout[1026] , 
        \DataPath/RF/bus_reg_dataout[1025] , 
        \DataPath/RF/bus_reg_dataout[1024] , 
        \DataPath/RF/bus_reg_dataout[1023] , 
        \DataPath/RF/bus_reg_dataout[1022] , 
        \DataPath/RF/bus_reg_dataout[1021] , 
        \DataPath/RF/bus_reg_dataout[1020] , 
        \DataPath/RF/bus_reg_dataout[1019] , 
        \DataPath/RF/bus_reg_dataout[1018] , 
        \DataPath/RF/bus_reg_dataout[1017] , 
        \DataPath/RF/bus_reg_dataout[1016] , 
        \DataPath/RF/bus_reg_dataout[1015] , 
        \DataPath/RF/bus_reg_dataout[1014] , 
        \DataPath/RF/bus_reg_dataout[1013] , 
        \DataPath/RF/bus_reg_dataout[1012] , 
        \DataPath/RF/bus_reg_dataout[1011] , 
        \DataPath/RF/bus_reg_dataout[1010] , 
        \DataPath/RF/bus_reg_dataout[1009] , 
        \DataPath/RF/bus_reg_dataout[1008] , 
        \DataPath/RF/bus_reg_dataout[1007] , 
        \DataPath/RF/bus_reg_dataout[1006] , 
        \DataPath/RF/bus_reg_dataout[1005] , 
        \DataPath/RF/bus_reg_dataout[1004] , 
        \DataPath/RF/bus_reg_dataout[1003] , 
        \DataPath/RF/bus_reg_dataout[1002] , 
        \DataPath/RF/bus_reg_dataout[1001] , 
        \DataPath/RF/bus_reg_dataout[1000] , 
        \DataPath/RF/bus_reg_dataout[999] , \DataPath/RF/bus_reg_dataout[998] , 
        \DataPath/RF/bus_reg_dataout[997] , \DataPath/RF/bus_reg_dataout[996] , 
        \DataPath/RF/bus_reg_dataout[995] , \DataPath/RF/bus_reg_dataout[994] , 
        \DataPath/RF/bus_reg_dataout[993] , \DataPath/RF/bus_reg_dataout[992] , 
        \DataPath/RF/bus_reg_dataout[991] , \DataPath/RF/bus_reg_dataout[990] , 
        \DataPath/RF/bus_reg_dataout[989] , \DataPath/RF/bus_reg_dataout[988] , 
        \DataPath/RF/bus_reg_dataout[987] , \DataPath/RF/bus_reg_dataout[986] , 
        \DataPath/RF/bus_reg_dataout[985] , \DataPath/RF/bus_reg_dataout[984] , 
        \DataPath/RF/bus_reg_dataout[983] , \DataPath/RF/bus_reg_dataout[982] , 
        \DataPath/RF/bus_reg_dataout[981] , \DataPath/RF/bus_reg_dataout[980] , 
        \DataPath/RF/bus_reg_dataout[979] , \DataPath/RF/bus_reg_dataout[978] , 
        \DataPath/RF/bus_reg_dataout[977] , \DataPath/RF/bus_reg_dataout[976] , 
        \DataPath/RF/bus_reg_dataout[975] , \DataPath/RF/bus_reg_dataout[974] , 
        \DataPath/RF/bus_reg_dataout[973] , \DataPath/RF/bus_reg_dataout[972] , 
        \DataPath/RF/bus_reg_dataout[971] , \DataPath/RF/bus_reg_dataout[970] , 
        \DataPath/RF/bus_reg_dataout[969] , \DataPath/RF/bus_reg_dataout[968] , 
        \DataPath/RF/bus_reg_dataout[967] , \DataPath/RF/bus_reg_dataout[966] , 
        \DataPath/RF/bus_reg_dataout[965] , \DataPath/RF/bus_reg_dataout[964] , 
        \DataPath/RF/bus_reg_dataout[963] , \DataPath/RF/bus_reg_dataout[962] , 
        \DataPath/RF/bus_reg_dataout[961] , \DataPath/RF/bus_reg_dataout[960] , 
        \DataPath/RF/bus_reg_dataout[959] , \DataPath/RF/bus_reg_dataout[958] , 
        \DataPath/RF/bus_reg_dataout[957] , \DataPath/RF/bus_reg_dataout[956] , 
        \DataPath/RF/bus_reg_dataout[955] , \DataPath/RF/bus_reg_dataout[954] , 
        \DataPath/RF/bus_reg_dataout[953] , \DataPath/RF/bus_reg_dataout[952] , 
        \DataPath/RF/bus_reg_dataout[951] , \DataPath/RF/bus_reg_dataout[950] , 
        \DataPath/RF/bus_reg_dataout[949] , \DataPath/RF/bus_reg_dataout[948] , 
        \DataPath/RF/bus_reg_dataout[947] , \DataPath/RF/bus_reg_dataout[946] , 
        \DataPath/RF/bus_reg_dataout[945] , \DataPath/RF/bus_reg_dataout[944] , 
        \DataPath/RF/bus_reg_dataout[943] , \DataPath/RF/bus_reg_dataout[942] , 
        \DataPath/RF/bus_reg_dataout[941] , \DataPath/RF/bus_reg_dataout[940] , 
        \DataPath/RF/bus_reg_dataout[939] , \DataPath/RF/bus_reg_dataout[938] , 
        \DataPath/RF/bus_reg_dataout[937] , \DataPath/RF/bus_reg_dataout[936] , 
        \DataPath/RF/bus_reg_dataout[935] , \DataPath/RF/bus_reg_dataout[934] , 
        \DataPath/RF/bus_reg_dataout[933] , \DataPath/RF/bus_reg_dataout[932] , 
        \DataPath/RF/bus_reg_dataout[931] , \DataPath/RF/bus_reg_dataout[930] , 
        \DataPath/RF/bus_reg_dataout[929] , \DataPath/RF/bus_reg_dataout[928] , 
        \DataPath/RF/bus_reg_dataout[927] , \DataPath/RF/bus_reg_dataout[926] , 
        \DataPath/RF/bus_reg_dataout[925] , \DataPath/RF/bus_reg_dataout[924] , 
        \DataPath/RF/bus_reg_dataout[923] , \DataPath/RF/bus_reg_dataout[922] , 
        \DataPath/RF/bus_reg_dataout[921] , \DataPath/RF/bus_reg_dataout[920] , 
        \DataPath/RF/bus_reg_dataout[919] , \DataPath/RF/bus_reg_dataout[918] , 
        \DataPath/RF/bus_reg_dataout[917] , \DataPath/RF/bus_reg_dataout[916] , 
        \DataPath/RF/bus_reg_dataout[915] , \DataPath/RF/bus_reg_dataout[914] , 
        \DataPath/RF/bus_reg_dataout[913] , \DataPath/RF/bus_reg_dataout[912] , 
        \DataPath/RF/bus_reg_dataout[911] , \DataPath/RF/bus_reg_dataout[910] , 
        \DataPath/RF/bus_reg_dataout[909] , \DataPath/RF/bus_reg_dataout[908] , 
        \DataPath/RF/bus_reg_dataout[907] , \DataPath/RF/bus_reg_dataout[906] , 
        \DataPath/RF/bus_reg_dataout[905] , \DataPath/RF/bus_reg_dataout[904] , 
        \DataPath/RF/bus_reg_dataout[903] , \DataPath/RF/bus_reg_dataout[902] , 
        \DataPath/RF/bus_reg_dataout[901] , \DataPath/RF/bus_reg_dataout[900] , 
        \DataPath/RF/bus_reg_dataout[899] , \DataPath/RF/bus_reg_dataout[898] , 
        \DataPath/RF/bus_reg_dataout[897] , \DataPath/RF/bus_reg_dataout[896] , 
        \DataPath/RF/bus_reg_dataout[895] , \DataPath/RF/bus_reg_dataout[894] , 
        \DataPath/RF/bus_reg_dataout[893] , \DataPath/RF/bus_reg_dataout[892] , 
        \DataPath/RF/bus_reg_dataout[891] , \DataPath/RF/bus_reg_dataout[890] , 
        \DataPath/RF/bus_reg_dataout[889] , \DataPath/RF/bus_reg_dataout[888] , 
        \DataPath/RF/bus_reg_dataout[887] , \DataPath/RF/bus_reg_dataout[886] , 
        \DataPath/RF/bus_reg_dataout[885] , \DataPath/RF/bus_reg_dataout[884] , 
        \DataPath/RF/bus_reg_dataout[883] , \DataPath/RF/bus_reg_dataout[882] , 
        \DataPath/RF/bus_reg_dataout[881] , \DataPath/RF/bus_reg_dataout[880] , 
        \DataPath/RF/bus_reg_dataout[879] , \DataPath/RF/bus_reg_dataout[878] , 
        \DataPath/RF/bus_reg_dataout[877] , \DataPath/RF/bus_reg_dataout[876] , 
        \DataPath/RF/bus_reg_dataout[875] , \DataPath/RF/bus_reg_dataout[874] , 
        \DataPath/RF/bus_reg_dataout[873] , \DataPath/RF/bus_reg_dataout[872] , 
        \DataPath/RF/bus_reg_dataout[871] , \DataPath/RF/bus_reg_dataout[870] , 
        \DataPath/RF/bus_reg_dataout[869] , \DataPath/RF/bus_reg_dataout[868] , 
        \DataPath/RF/bus_reg_dataout[867] , \DataPath/RF/bus_reg_dataout[866] , 
        \DataPath/RF/bus_reg_dataout[865] , \DataPath/RF/bus_reg_dataout[864] , 
        \DataPath/RF/bus_reg_dataout[863] , \DataPath/RF/bus_reg_dataout[862] , 
        \DataPath/RF/bus_reg_dataout[861] , \DataPath/RF/bus_reg_dataout[860] , 
        \DataPath/RF/bus_reg_dataout[859] , \DataPath/RF/bus_reg_dataout[858] , 
        \DataPath/RF/bus_reg_dataout[857] , \DataPath/RF/bus_reg_dataout[856] , 
        \DataPath/RF/bus_reg_dataout[855] , \DataPath/RF/bus_reg_dataout[854] , 
        \DataPath/RF/bus_reg_dataout[853] , \DataPath/RF/bus_reg_dataout[852] , 
        \DataPath/RF/bus_reg_dataout[851] , \DataPath/RF/bus_reg_dataout[850] , 
        \DataPath/RF/bus_reg_dataout[849] , \DataPath/RF/bus_reg_dataout[848] , 
        \DataPath/RF/bus_reg_dataout[847] , \DataPath/RF/bus_reg_dataout[846] , 
        \DataPath/RF/bus_reg_dataout[845] , \DataPath/RF/bus_reg_dataout[844] , 
        \DataPath/RF/bus_reg_dataout[843] , \DataPath/RF/bus_reg_dataout[842] , 
        \DataPath/RF/bus_reg_dataout[841] , \DataPath/RF/bus_reg_dataout[840] , 
        \DataPath/RF/bus_reg_dataout[839] , \DataPath/RF/bus_reg_dataout[838] , 
        \DataPath/RF/bus_reg_dataout[837] , \DataPath/RF/bus_reg_dataout[836] , 
        \DataPath/RF/bus_reg_dataout[835] , \DataPath/RF/bus_reg_dataout[834] , 
        \DataPath/RF/bus_reg_dataout[833] , \DataPath/RF/bus_reg_dataout[832] , 
        \DataPath/RF/bus_reg_dataout[831] , \DataPath/RF/bus_reg_dataout[830] , 
        \DataPath/RF/bus_reg_dataout[829] , \DataPath/RF/bus_reg_dataout[828] , 
        \DataPath/RF/bus_reg_dataout[827] , \DataPath/RF/bus_reg_dataout[826] , 
        \DataPath/RF/bus_reg_dataout[825] , \DataPath/RF/bus_reg_dataout[824] , 
        \DataPath/RF/bus_reg_dataout[823] , \DataPath/RF/bus_reg_dataout[822] , 
        \DataPath/RF/bus_reg_dataout[821] , \DataPath/RF/bus_reg_dataout[820] , 
        \DataPath/RF/bus_reg_dataout[819] , \DataPath/RF/bus_reg_dataout[818] , 
        \DataPath/RF/bus_reg_dataout[817] , \DataPath/RF/bus_reg_dataout[816] , 
        \DataPath/RF/bus_reg_dataout[815] , \DataPath/RF/bus_reg_dataout[814] , 
        \DataPath/RF/bus_reg_dataout[813] , \DataPath/RF/bus_reg_dataout[812] , 
        \DataPath/RF/bus_reg_dataout[811] , \DataPath/RF/bus_reg_dataout[810] , 
        \DataPath/RF/bus_reg_dataout[809] , \DataPath/RF/bus_reg_dataout[808] , 
        \DataPath/RF/bus_reg_dataout[807] , \DataPath/RF/bus_reg_dataout[806] , 
        \DataPath/RF/bus_reg_dataout[805] , \DataPath/RF/bus_reg_dataout[804] , 
        \DataPath/RF/bus_reg_dataout[803] , \DataPath/RF/bus_reg_dataout[802] , 
        \DataPath/RF/bus_reg_dataout[801] , \DataPath/RF/bus_reg_dataout[800] , 
        \DataPath/RF/bus_reg_dataout[799] , \DataPath/RF/bus_reg_dataout[798] , 
        \DataPath/RF/bus_reg_dataout[797] , \DataPath/RF/bus_reg_dataout[796] , 
        \DataPath/RF/bus_reg_dataout[795] , \DataPath/RF/bus_reg_dataout[794] , 
        \DataPath/RF/bus_reg_dataout[793] , \DataPath/RF/bus_reg_dataout[792] , 
        \DataPath/RF/bus_reg_dataout[791] , \DataPath/RF/bus_reg_dataout[790] , 
        \DataPath/RF/bus_reg_dataout[789] , \DataPath/RF/bus_reg_dataout[788] , 
        \DataPath/RF/bus_reg_dataout[787] , \DataPath/RF/bus_reg_dataout[786] , 
        \DataPath/RF/bus_reg_dataout[785] , \DataPath/RF/bus_reg_dataout[784] , 
        \DataPath/RF/bus_reg_dataout[783] , \DataPath/RF/bus_reg_dataout[782] , 
        \DataPath/RF/bus_reg_dataout[781] , \DataPath/RF/bus_reg_dataout[780] , 
        \DataPath/RF/bus_reg_dataout[779] , \DataPath/RF/bus_reg_dataout[778] , 
        \DataPath/RF/bus_reg_dataout[777] , \DataPath/RF/bus_reg_dataout[776] , 
        \DataPath/RF/bus_reg_dataout[775] , \DataPath/RF/bus_reg_dataout[774] , 
        \DataPath/RF/bus_reg_dataout[773] , \DataPath/RF/bus_reg_dataout[772] , 
        \DataPath/RF/bus_reg_dataout[771] , \DataPath/RF/bus_reg_dataout[770] , 
        \DataPath/RF/bus_reg_dataout[769] , \DataPath/RF/bus_reg_dataout[768] , 
        \DataPath/RF/bus_reg_dataout[767] , \DataPath/RF/bus_reg_dataout[766] , 
        \DataPath/RF/bus_reg_dataout[765] , \DataPath/RF/bus_reg_dataout[764] , 
        \DataPath/RF/bus_reg_dataout[763] , \DataPath/RF/bus_reg_dataout[762] , 
        \DataPath/RF/bus_reg_dataout[761] , \DataPath/RF/bus_reg_dataout[760] , 
        \DataPath/RF/bus_reg_dataout[759] , \DataPath/RF/bus_reg_dataout[758] , 
        \DataPath/RF/bus_reg_dataout[757] , \DataPath/RF/bus_reg_dataout[756] , 
        \DataPath/RF/bus_reg_dataout[755] , \DataPath/RF/bus_reg_dataout[754] , 
        \DataPath/RF/bus_reg_dataout[753] , \DataPath/RF/bus_reg_dataout[752] , 
        \DataPath/RF/bus_reg_dataout[751] , \DataPath/RF/bus_reg_dataout[750] , 
        \DataPath/RF/bus_reg_dataout[749] , \DataPath/RF/bus_reg_dataout[748] , 
        \DataPath/RF/bus_reg_dataout[747] , \DataPath/RF/bus_reg_dataout[746] , 
        \DataPath/RF/bus_reg_dataout[745] , \DataPath/RF/bus_reg_dataout[744] , 
        \DataPath/RF/bus_reg_dataout[743] , \DataPath/RF/bus_reg_dataout[742] , 
        \DataPath/RF/bus_reg_dataout[741] , \DataPath/RF/bus_reg_dataout[740] , 
        \DataPath/RF/bus_reg_dataout[739] , \DataPath/RF/bus_reg_dataout[738] , 
        \DataPath/RF/bus_reg_dataout[737] , \DataPath/RF/bus_reg_dataout[736] , 
        \DataPath/RF/bus_reg_dataout[735] , \DataPath/RF/bus_reg_dataout[734] , 
        \DataPath/RF/bus_reg_dataout[733] , \DataPath/RF/bus_reg_dataout[732] , 
        \DataPath/RF/bus_reg_dataout[731] , \DataPath/RF/bus_reg_dataout[730] , 
        \DataPath/RF/bus_reg_dataout[729] , \DataPath/RF/bus_reg_dataout[728] , 
        \DataPath/RF/bus_reg_dataout[727] , \DataPath/RF/bus_reg_dataout[726] , 
        \DataPath/RF/bus_reg_dataout[725] , \DataPath/RF/bus_reg_dataout[724] , 
        \DataPath/RF/bus_reg_dataout[723] , \DataPath/RF/bus_reg_dataout[722] , 
        \DataPath/RF/bus_reg_dataout[721] , \DataPath/RF/bus_reg_dataout[720] , 
        \DataPath/RF/bus_reg_dataout[719] , \DataPath/RF/bus_reg_dataout[718] , 
        \DataPath/RF/bus_reg_dataout[717] , \DataPath/RF/bus_reg_dataout[716] , 
        \DataPath/RF/bus_reg_dataout[715] , \DataPath/RF/bus_reg_dataout[714] , 
        \DataPath/RF/bus_reg_dataout[713] , \DataPath/RF/bus_reg_dataout[712] , 
        \DataPath/RF/bus_reg_dataout[711] , \DataPath/RF/bus_reg_dataout[710] , 
        \DataPath/RF/bus_reg_dataout[709] , \DataPath/RF/bus_reg_dataout[708] , 
        \DataPath/RF/bus_reg_dataout[707] , \DataPath/RF/bus_reg_dataout[706] , 
        \DataPath/RF/bus_reg_dataout[705] , \DataPath/RF/bus_reg_dataout[704] , 
        \DataPath/RF/bus_reg_dataout[703] , \DataPath/RF/bus_reg_dataout[702] , 
        \DataPath/RF/bus_reg_dataout[701] , \DataPath/RF/bus_reg_dataout[700] , 
        \DataPath/RF/bus_reg_dataout[699] , \DataPath/RF/bus_reg_dataout[698] , 
        \DataPath/RF/bus_reg_dataout[697] , \DataPath/RF/bus_reg_dataout[696] , 
        \DataPath/RF/bus_reg_dataout[695] , \DataPath/RF/bus_reg_dataout[694] , 
        \DataPath/RF/bus_reg_dataout[693] , \DataPath/RF/bus_reg_dataout[692] , 
        \DataPath/RF/bus_reg_dataout[691] , \DataPath/RF/bus_reg_dataout[690] , 
        \DataPath/RF/bus_reg_dataout[689] , \DataPath/RF/bus_reg_dataout[688] , 
        \DataPath/RF/bus_reg_dataout[687] , \DataPath/RF/bus_reg_dataout[686] , 
        \DataPath/RF/bus_reg_dataout[685] , \DataPath/RF/bus_reg_dataout[684] , 
        \DataPath/RF/bus_reg_dataout[683] , \DataPath/RF/bus_reg_dataout[682] , 
        \DataPath/RF/bus_reg_dataout[681] , \DataPath/RF/bus_reg_dataout[680] , 
        \DataPath/RF/bus_reg_dataout[679] , \DataPath/RF/bus_reg_dataout[678] , 
        \DataPath/RF/bus_reg_dataout[677] , \DataPath/RF/bus_reg_dataout[676] , 
        \DataPath/RF/bus_reg_dataout[675] , \DataPath/RF/bus_reg_dataout[674] , 
        \DataPath/RF/bus_reg_dataout[673] , \DataPath/RF/bus_reg_dataout[672] , 
        \DataPath/RF/bus_reg_dataout[671] , \DataPath/RF/bus_reg_dataout[670] , 
        \DataPath/RF/bus_reg_dataout[669] , \DataPath/RF/bus_reg_dataout[668] , 
        \DataPath/RF/bus_reg_dataout[667] , \DataPath/RF/bus_reg_dataout[666] , 
        \DataPath/RF/bus_reg_dataout[665] , \DataPath/RF/bus_reg_dataout[664] , 
        \DataPath/RF/bus_reg_dataout[663] , \DataPath/RF/bus_reg_dataout[662] , 
        \DataPath/RF/bus_reg_dataout[661] , \DataPath/RF/bus_reg_dataout[660] , 
        \DataPath/RF/bus_reg_dataout[659] , \DataPath/RF/bus_reg_dataout[658] , 
        \DataPath/RF/bus_reg_dataout[657] , \DataPath/RF/bus_reg_dataout[656] , 
        \DataPath/RF/bus_reg_dataout[655] , \DataPath/RF/bus_reg_dataout[654] , 
        \DataPath/RF/bus_reg_dataout[653] , \DataPath/RF/bus_reg_dataout[652] , 
        \DataPath/RF/bus_reg_dataout[651] , \DataPath/RF/bus_reg_dataout[650] , 
        \DataPath/RF/bus_reg_dataout[649] , \DataPath/RF/bus_reg_dataout[648] , 
        \DataPath/RF/bus_reg_dataout[647] , \DataPath/RF/bus_reg_dataout[646] , 
        \DataPath/RF/bus_reg_dataout[645] , \DataPath/RF/bus_reg_dataout[644] , 
        \DataPath/RF/bus_reg_dataout[643] , \DataPath/RF/bus_reg_dataout[642] , 
        \DataPath/RF/bus_reg_dataout[641] , \DataPath/RF/bus_reg_dataout[640] , 
        \DataPath/RF/bus_reg_dataout[639] , \DataPath/RF/bus_reg_dataout[638] , 
        \DataPath/RF/bus_reg_dataout[637] , \DataPath/RF/bus_reg_dataout[636] , 
        \DataPath/RF/bus_reg_dataout[635] , \DataPath/RF/bus_reg_dataout[634] , 
        \DataPath/RF/bus_reg_dataout[633] , \DataPath/RF/bus_reg_dataout[632] , 
        \DataPath/RF/bus_reg_dataout[631] , \DataPath/RF/bus_reg_dataout[630] , 
        \DataPath/RF/bus_reg_dataout[629] , \DataPath/RF/bus_reg_dataout[628] , 
        \DataPath/RF/bus_reg_dataout[627] , \DataPath/RF/bus_reg_dataout[626] , 
        \DataPath/RF/bus_reg_dataout[625] , \DataPath/RF/bus_reg_dataout[624] , 
        \DataPath/RF/bus_reg_dataout[623] , \DataPath/RF/bus_reg_dataout[622] , 
        \DataPath/RF/bus_reg_dataout[621] , \DataPath/RF/bus_reg_dataout[620] , 
        \DataPath/RF/bus_reg_dataout[619] , \DataPath/RF/bus_reg_dataout[618] , 
        \DataPath/RF/bus_reg_dataout[617] , \DataPath/RF/bus_reg_dataout[616] , 
        \DataPath/RF/bus_reg_dataout[615] , \DataPath/RF/bus_reg_dataout[614] , 
        \DataPath/RF/bus_reg_dataout[613] , \DataPath/RF/bus_reg_dataout[612] , 
        \DataPath/RF/bus_reg_dataout[611] , \DataPath/RF/bus_reg_dataout[610] , 
        \DataPath/RF/bus_reg_dataout[609] , \DataPath/RF/bus_reg_dataout[608] , 
        \DataPath/RF/bus_reg_dataout[607] , \DataPath/RF/bus_reg_dataout[606] , 
        \DataPath/RF/bus_reg_dataout[605] , \DataPath/RF/bus_reg_dataout[604] , 
        \DataPath/RF/bus_reg_dataout[603] , \DataPath/RF/bus_reg_dataout[602] , 
        \DataPath/RF/bus_reg_dataout[601] , \DataPath/RF/bus_reg_dataout[600] , 
        \DataPath/RF/bus_reg_dataout[599] , \DataPath/RF/bus_reg_dataout[598] , 
        \DataPath/RF/bus_reg_dataout[597] , \DataPath/RF/bus_reg_dataout[596] , 
        \DataPath/RF/bus_reg_dataout[595] , \DataPath/RF/bus_reg_dataout[594] , 
        \DataPath/RF/bus_reg_dataout[593] , \DataPath/RF/bus_reg_dataout[592] , 
        \DataPath/RF/bus_reg_dataout[591] , \DataPath/RF/bus_reg_dataout[590] , 
        \DataPath/RF/bus_reg_dataout[589] , \DataPath/RF/bus_reg_dataout[588] , 
        \DataPath/RF/bus_reg_dataout[587] , \DataPath/RF/bus_reg_dataout[586] , 
        \DataPath/RF/bus_reg_dataout[585] , \DataPath/RF/bus_reg_dataout[584] , 
        \DataPath/RF/bus_reg_dataout[583] , \DataPath/RF/bus_reg_dataout[582] , 
        \DataPath/RF/bus_reg_dataout[581] , \DataPath/RF/bus_reg_dataout[580] , 
        \DataPath/RF/bus_reg_dataout[579] , \DataPath/RF/bus_reg_dataout[578] , 
        \DataPath/RF/bus_reg_dataout[577] , \DataPath/RF/bus_reg_dataout[576] , 
        \DataPath/RF/bus_reg_dataout[575] , \DataPath/RF/bus_reg_dataout[574] , 
        \DataPath/RF/bus_reg_dataout[573] , \DataPath/RF/bus_reg_dataout[572] , 
        \DataPath/RF/bus_reg_dataout[571] , \DataPath/RF/bus_reg_dataout[570] , 
        \DataPath/RF/bus_reg_dataout[569] , \DataPath/RF/bus_reg_dataout[568] , 
        \DataPath/RF/bus_reg_dataout[567] , \DataPath/RF/bus_reg_dataout[566] , 
        \DataPath/RF/bus_reg_dataout[565] , \DataPath/RF/bus_reg_dataout[564] , 
        \DataPath/RF/bus_reg_dataout[563] , \DataPath/RF/bus_reg_dataout[562] , 
        \DataPath/RF/bus_reg_dataout[561] , \DataPath/RF/bus_reg_dataout[560] , 
        \DataPath/RF/bus_reg_dataout[559] , \DataPath/RF/bus_reg_dataout[558] , 
        \DataPath/RF/bus_reg_dataout[557] , \DataPath/RF/bus_reg_dataout[556] , 
        \DataPath/RF/bus_reg_dataout[555] , \DataPath/RF/bus_reg_dataout[554] , 
        \DataPath/RF/bus_reg_dataout[553] , \DataPath/RF/bus_reg_dataout[552] , 
        \DataPath/RF/bus_reg_dataout[551] , \DataPath/RF/bus_reg_dataout[550] , 
        \DataPath/RF/bus_reg_dataout[549] , \DataPath/RF/bus_reg_dataout[548] , 
        \DataPath/RF/bus_reg_dataout[547] , \DataPath/RF/bus_reg_dataout[546] , 
        \DataPath/RF/bus_reg_dataout[545] , \DataPath/RF/bus_reg_dataout[544] , 
        \DataPath/RF/bus_reg_dataout[543] , \DataPath/RF/bus_reg_dataout[542] , 
        \DataPath/RF/bus_reg_dataout[541] , \DataPath/RF/bus_reg_dataout[540] , 
        \DataPath/RF/bus_reg_dataout[539] , \DataPath/RF/bus_reg_dataout[538] , 
        \DataPath/RF/bus_reg_dataout[537] , \DataPath/RF/bus_reg_dataout[536] , 
        \DataPath/RF/bus_reg_dataout[535] , \DataPath/RF/bus_reg_dataout[534] , 
        \DataPath/RF/bus_reg_dataout[533] , \DataPath/RF/bus_reg_dataout[532] , 
        \DataPath/RF/bus_reg_dataout[531] , \DataPath/RF/bus_reg_dataout[530] , 
        \DataPath/RF/bus_reg_dataout[529] , \DataPath/RF/bus_reg_dataout[528] , 
        \DataPath/RF/bus_reg_dataout[527] , \DataPath/RF/bus_reg_dataout[526] , 
        \DataPath/RF/bus_reg_dataout[525] , \DataPath/RF/bus_reg_dataout[524] , 
        \DataPath/RF/bus_reg_dataout[523] , \DataPath/RF/bus_reg_dataout[522] , 
        \DataPath/RF/bus_reg_dataout[521] , \DataPath/RF/bus_reg_dataout[520] , 
        \DataPath/RF/bus_reg_dataout[519] , \DataPath/RF/bus_reg_dataout[518] , 
        \DataPath/RF/bus_reg_dataout[517] , \DataPath/RF/bus_reg_dataout[516] , 
        \DataPath/RF/bus_reg_dataout[515] , \DataPath/RF/bus_reg_dataout[514] , 
        \DataPath/RF/bus_reg_dataout[513] , \DataPath/RF/bus_reg_dataout[512] , 
        \DataPath/RF/bus_reg_dataout[511] , \DataPath/RF/bus_reg_dataout[510] , 
        \DataPath/RF/bus_reg_dataout[509] , \DataPath/RF/bus_reg_dataout[508] , 
        \DataPath/RF/bus_reg_dataout[507] , \DataPath/RF/bus_reg_dataout[506] , 
        \DataPath/RF/bus_reg_dataout[505] , \DataPath/RF/bus_reg_dataout[504] , 
        \DataPath/RF/bus_reg_dataout[503] , \DataPath/RF/bus_reg_dataout[502] , 
        \DataPath/RF/bus_reg_dataout[501] , \DataPath/RF/bus_reg_dataout[500] , 
        \DataPath/RF/bus_reg_dataout[499] , \DataPath/RF/bus_reg_dataout[498] , 
        \DataPath/RF/bus_reg_dataout[497] , \DataPath/RF/bus_reg_dataout[496] , 
        \DataPath/RF/bus_reg_dataout[495] , \DataPath/RF/bus_reg_dataout[494] , 
        \DataPath/RF/bus_reg_dataout[493] , \DataPath/RF/bus_reg_dataout[492] , 
        \DataPath/RF/bus_reg_dataout[491] , \DataPath/RF/bus_reg_dataout[490] , 
        \DataPath/RF/bus_reg_dataout[489] , \DataPath/RF/bus_reg_dataout[488] , 
        \DataPath/RF/bus_reg_dataout[487] , \DataPath/RF/bus_reg_dataout[486] , 
        \DataPath/RF/bus_reg_dataout[485] , \DataPath/RF/bus_reg_dataout[484] , 
        \DataPath/RF/bus_reg_dataout[483] , \DataPath/RF/bus_reg_dataout[482] , 
        \DataPath/RF/bus_reg_dataout[481] , \DataPath/RF/bus_reg_dataout[480] , 
        \DataPath/RF/bus_reg_dataout[479] , \DataPath/RF/bus_reg_dataout[478] , 
        \DataPath/RF/bus_reg_dataout[477] , \DataPath/RF/bus_reg_dataout[476] , 
        \DataPath/RF/bus_reg_dataout[475] , \DataPath/RF/bus_reg_dataout[474] , 
        \DataPath/RF/bus_reg_dataout[473] , \DataPath/RF/bus_reg_dataout[472] , 
        \DataPath/RF/bus_reg_dataout[471] , \DataPath/RF/bus_reg_dataout[470] , 
        \DataPath/RF/bus_reg_dataout[469] , \DataPath/RF/bus_reg_dataout[468] , 
        \DataPath/RF/bus_reg_dataout[467] , \DataPath/RF/bus_reg_dataout[466] , 
        \DataPath/RF/bus_reg_dataout[465] , \DataPath/RF/bus_reg_dataout[464] , 
        \DataPath/RF/bus_reg_dataout[463] , \DataPath/RF/bus_reg_dataout[462] , 
        \DataPath/RF/bus_reg_dataout[461] , \DataPath/RF/bus_reg_dataout[460] , 
        \DataPath/RF/bus_reg_dataout[459] , \DataPath/RF/bus_reg_dataout[458] , 
        \DataPath/RF/bus_reg_dataout[457] , \DataPath/RF/bus_reg_dataout[456] , 
        \DataPath/RF/bus_reg_dataout[455] , \DataPath/RF/bus_reg_dataout[454] , 
        \DataPath/RF/bus_reg_dataout[453] , \DataPath/RF/bus_reg_dataout[452] , 
        \DataPath/RF/bus_reg_dataout[451] , \DataPath/RF/bus_reg_dataout[450] , 
        \DataPath/RF/bus_reg_dataout[449] , \DataPath/RF/bus_reg_dataout[448] , 
        \DataPath/RF/bus_reg_dataout[447] , \DataPath/RF/bus_reg_dataout[446] , 
        \DataPath/RF/bus_reg_dataout[445] , \DataPath/RF/bus_reg_dataout[444] , 
        \DataPath/RF/bus_reg_dataout[443] , \DataPath/RF/bus_reg_dataout[442] , 
        \DataPath/RF/bus_reg_dataout[441] , \DataPath/RF/bus_reg_dataout[440] , 
        \DataPath/RF/bus_reg_dataout[439] , \DataPath/RF/bus_reg_dataout[438] , 
        \DataPath/RF/bus_reg_dataout[437] , \DataPath/RF/bus_reg_dataout[436] , 
        \DataPath/RF/bus_reg_dataout[435] , \DataPath/RF/bus_reg_dataout[434] , 
        \DataPath/RF/bus_reg_dataout[433] , \DataPath/RF/bus_reg_dataout[432] , 
        \DataPath/RF/bus_reg_dataout[431] , \DataPath/RF/bus_reg_dataout[430] , 
        \DataPath/RF/bus_reg_dataout[429] , \DataPath/RF/bus_reg_dataout[428] , 
        \DataPath/RF/bus_reg_dataout[427] , \DataPath/RF/bus_reg_dataout[426] , 
        \DataPath/RF/bus_reg_dataout[425] , \DataPath/RF/bus_reg_dataout[424] , 
        \DataPath/RF/bus_reg_dataout[423] , \DataPath/RF/bus_reg_dataout[422] , 
        \DataPath/RF/bus_reg_dataout[421] , \DataPath/RF/bus_reg_dataout[420] , 
        \DataPath/RF/bus_reg_dataout[419] , \DataPath/RF/bus_reg_dataout[418] , 
        \DataPath/RF/bus_reg_dataout[417] , \DataPath/RF/bus_reg_dataout[416] , 
        \DataPath/RF/bus_reg_dataout[415] , \DataPath/RF/bus_reg_dataout[414] , 
        \DataPath/RF/bus_reg_dataout[413] , \DataPath/RF/bus_reg_dataout[412] , 
        \DataPath/RF/bus_reg_dataout[411] , \DataPath/RF/bus_reg_dataout[410] , 
        \DataPath/RF/bus_reg_dataout[409] , \DataPath/RF/bus_reg_dataout[408] , 
        \DataPath/RF/bus_reg_dataout[407] , \DataPath/RF/bus_reg_dataout[406] , 
        \DataPath/RF/bus_reg_dataout[405] , \DataPath/RF/bus_reg_dataout[404] , 
        \DataPath/RF/bus_reg_dataout[403] , \DataPath/RF/bus_reg_dataout[402] , 
        \DataPath/RF/bus_reg_dataout[401] , \DataPath/RF/bus_reg_dataout[400] , 
        \DataPath/RF/bus_reg_dataout[399] , \DataPath/RF/bus_reg_dataout[398] , 
        \DataPath/RF/bus_reg_dataout[397] , \DataPath/RF/bus_reg_dataout[396] , 
        \DataPath/RF/bus_reg_dataout[395] , \DataPath/RF/bus_reg_dataout[394] , 
        \DataPath/RF/bus_reg_dataout[393] , \DataPath/RF/bus_reg_dataout[392] , 
        \DataPath/RF/bus_reg_dataout[391] , \DataPath/RF/bus_reg_dataout[390] , 
        \DataPath/RF/bus_reg_dataout[389] , \DataPath/RF/bus_reg_dataout[388] , 
        \DataPath/RF/bus_reg_dataout[387] , \DataPath/RF/bus_reg_dataout[386] , 
        \DataPath/RF/bus_reg_dataout[385] , \DataPath/RF/bus_reg_dataout[384] , 
        \DataPath/RF/bus_reg_dataout[383] , \DataPath/RF/bus_reg_dataout[382] , 
        \DataPath/RF/bus_reg_dataout[381] , \DataPath/RF/bus_reg_dataout[380] , 
        \DataPath/RF/bus_reg_dataout[379] , \DataPath/RF/bus_reg_dataout[378] , 
        \DataPath/RF/bus_reg_dataout[377] , \DataPath/RF/bus_reg_dataout[376] , 
        \DataPath/RF/bus_reg_dataout[375] , \DataPath/RF/bus_reg_dataout[374] , 
        \DataPath/RF/bus_reg_dataout[373] , \DataPath/RF/bus_reg_dataout[372] , 
        \DataPath/RF/bus_reg_dataout[371] , \DataPath/RF/bus_reg_dataout[370] , 
        \DataPath/RF/bus_reg_dataout[369] , \DataPath/RF/bus_reg_dataout[368] , 
        \DataPath/RF/bus_reg_dataout[367] , \DataPath/RF/bus_reg_dataout[366] , 
        \DataPath/RF/bus_reg_dataout[365] , \DataPath/RF/bus_reg_dataout[364] , 
        \DataPath/RF/bus_reg_dataout[363] , \DataPath/RF/bus_reg_dataout[362] , 
        \DataPath/RF/bus_reg_dataout[361] , \DataPath/RF/bus_reg_dataout[360] , 
        \DataPath/RF/bus_reg_dataout[359] , \DataPath/RF/bus_reg_dataout[358] , 
        \DataPath/RF/bus_reg_dataout[357] , \DataPath/RF/bus_reg_dataout[356] , 
        \DataPath/RF/bus_reg_dataout[355] , \DataPath/RF/bus_reg_dataout[354] , 
        \DataPath/RF/bus_reg_dataout[353] , \DataPath/RF/bus_reg_dataout[352] , 
        \DataPath/RF/bus_reg_dataout[351] , \DataPath/RF/bus_reg_dataout[350] , 
        \DataPath/RF/bus_reg_dataout[349] , \DataPath/RF/bus_reg_dataout[348] , 
        \DataPath/RF/bus_reg_dataout[347] , \DataPath/RF/bus_reg_dataout[346] , 
        \DataPath/RF/bus_reg_dataout[345] , \DataPath/RF/bus_reg_dataout[344] , 
        \DataPath/RF/bus_reg_dataout[343] , \DataPath/RF/bus_reg_dataout[342] , 
        \DataPath/RF/bus_reg_dataout[341] , \DataPath/RF/bus_reg_dataout[340] , 
        \DataPath/RF/bus_reg_dataout[339] , \DataPath/RF/bus_reg_dataout[338] , 
        \DataPath/RF/bus_reg_dataout[337] , \DataPath/RF/bus_reg_dataout[336] , 
        \DataPath/RF/bus_reg_dataout[335] , \DataPath/RF/bus_reg_dataout[334] , 
        \DataPath/RF/bus_reg_dataout[333] , \DataPath/RF/bus_reg_dataout[332] , 
        \DataPath/RF/bus_reg_dataout[331] , \DataPath/RF/bus_reg_dataout[330] , 
        \DataPath/RF/bus_reg_dataout[329] , \DataPath/RF/bus_reg_dataout[328] , 
        \DataPath/RF/bus_reg_dataout[327] , \DataPath/RF/bus_reg_dataout[326] , 
        \DataPath/RF/bus_reg_dataout[325] , \DataPath/RF/bus_reg_dataout[324] , 
        \DataPath/RF/bus_reg_dataout[323] , \DataPath/RF/bus_reg_dataout[322] , 
        \DataPath/RF/bus_reg_dataout[321] , \DataPath/RF/bus_reg_dataout[320] , 
        \DataPath/RF/bus_reg_dataout[319] , \DataPath/RF/bus_reg_dataout[318] , 
        \DataPath/RF/bus_reg_dataout[317] , \DataPath/RF/bus_reg_dataout[316] , 
        \DataPath/RF/bus_reg_dataout[315] , \DataPath/RF/bus_reg_dataout[314] , 
        \DataPath/RF/bus_reg_dataout[313] , \DataPath/RF/bus_reg_dataout[312] , 
        \DataPath/RF/bus_reg_dataout[311] , \DataPath/RF/bus_reg_dataout[310] , 
        \DataPath/RF/bus_reg_dataout[309] , \DataPath/RF/bus_reg_dataout[308] , 
        \DataPath/RF/bus_reg_dataout[307] , \DataPath/RF/bus_reg_dataout[306] , 
        \DataPath/RF/bus_reg_dataout[305] , \DataPath/RF/bus_reg_dataout[304] , 
        \DataPath/RF/bus_reg_dataout[303] , \DataPath/RF/bus_reg_dataout[302] , 
        \DataPath/RF/bus_reg_dataout[301] , \DataPath/RF/bus_reg_dataout[300] , 
        \DataPath/RF/bus_reg_dataout[299] , \DataPath/RF/bus_reg_dataout[298] , 
        \DataPath/RF/bus_reg_dataout[297] , \DataPath/RF/bus_reg_dataout[296] , 
        \DataPath/RF/bus_reg_dataout[295] , \DataPath/RF/bus_reg_dataout[294] , 
        \DataPath/RF/bus_reg_dataout[293] , \DataPath/RF/bus_reg_dataout[292] , 
        \DataPath/RF/bus_reg_dataout[291] , \DataPath/RF/bus_reg_dataout[290] , 
        \DataPath/RF/bus_reg_dataout[289] , \DataPath/RF/bus_reg_dataout[288] , 
        \DataPath/RF/bus_reg_dataout[287] , \DataPath/RF/bus_reg_dataout[286] , 
        \DataPath/RF/bus_reg_dataout[285] , \DataPath/RF/bus_reg_dataout[284] , 
        \DataPath/RF/bus_reg_dataout[283] , \DataPath/RF/bus_reg_dataout[282] , 
        \DataPath/RF/bus_reg_dataout[281] , \DataPath/RF/bus_reg_dataout[280] , 
        \DataPath/RF/bus_reg_dataout[279] , \DataPath/RF/bus_reg_dataout[278] , 
        \DataPath/RF/bus_reg_dataout[277] , \DataPath/RF/bus_reg_dataout[276] , 
        \DataPath/RF/bus_reg_dataout[275] , \DataPath/RF/bus_reg_dataout[274] , 
        \DataPath/RF/bus_reg_dataout[273] , \DataPath/RF/bus_reg_dataout[272] , 
        \DataPath/RF/bus_reg_dataout[271] , \DataPath/RF/bus_reg_dataout[270] , 
        \DataPath/RF/bus_reg_dataout[269] , \DataPath/RF/bus_reg_dataout[268] , 
        \DataPath/RF/bus_reg_dataout[267] , \DataPath/RF/bus_reg_dataout[266] , 
        \DataPath/RF/bus_reg_dataout[265] , \DataPath/RF/bus_reg_dataout[264] , 
        \DataPath/RF/bus_reg_dataout[263] , \DataPath/RF/bus_reg_dataout[262] , 
        \DataPath/RF/bus_reg_dataout[261] , \DataPath/RF/bus_reg_dataout[260] , 
        \DataPath/RF/bus_reg_dataout[259] , \DataPath/RF/bus_reg_dataout[258] , 
        \DataPath/RF/bus_reg_dataout[257] , \DataPath/RF/bus_reg_dataout[256] , 
        \DataPath/RF/bus_reg_dataout[255] , \DataPath/RF/bus_reg_dataout[254] , 
        \DataPath/RF/bus_reg_dataout[253] , \DataPath/RF/bus_reg_dataout[252] , 
        \DataPath/RF/bus_reg_dataout[251] , \DataPath/RF/bus_reg_dataout[250] , 
        \DataPath/RF/bus_reg_dataout[249] , \DataPath/RF/bus_reg_dataout[248] , 
        \DataPath/RF/bus_reg_dataout[247] , \DataPath/RF/bus_reg_dataout[246] , 
        \DataPath/RF/bus_reg_dataout[245] , \DataPath/RF/bus_reg_dataout[244] , 
        \DataPath/RF/bus_reg_dataout[243] , \DataPath/RF/bus_reg_dataout[242] , 
        \DataPath/RF/bus_reg_dataout[241] , \DataPath/RF/bus_reg_dataout[240] , 
        \DataPath/RF/bus_reg_dataout[239] , \DataPath/RF/bus_reg_dataout[238] , 
        \DataPath/RF/bus_reg_dataout[237] , \DataPath/RF/bus_reg_dataout[236] , 
        \DataPath/RF/bus_reg_dataout[235] , \DataPath/RF/bus_reg_dataout[234] , 
        \DataPath/RF/bus_reg_dataout[233] , \DataPath/RF/bus_reg_dataout[232] , 
        \DataPath/RF/bus_reg_dataout[231] , \DataPath/RF/bus_reg_dataout[230] , 
        \DataPath/RF/bus_reg_dataout[229] , \DataPath/RF/bus_reg_dataout[228] , 
        \DataPath/RF/bus_reg_dataout[227] , \DataPath/RF/bus_reg_dataout[226] , 
        \DataPath/RF/bus_reg_dataout[225] , \DataPath/RF/bus_reg_dataout[224] , 
        \DataPath/RF/bus_reg_dataout[223] , \DataPath/RF/bus_reg_dataout[222] , 
        \DataPath/RF/bus_reg_dataout[221] , \DataPath/RF/bus_reg_dataout[220] , 
        \DataPath/RF/bus_reg_dataout[219] , \DataPath/RF/bus_reg_dataout[218] , 
        \DataPath/RF/bus_reg_dataout[217] , \DataPath/RF/bus_reg_dataout[216] , 
        \DataPath/RF/bus_reg_dataout[215] , \DataPath/RF/bus_reg_dataout[214] , 
        \DataPath/RF/bus_reg_dataout[213] , \DataPath/RF/bus_reg_dataout[212] , 
        \DataPath/RF/bus_reg_dataout[211] , \DataPath/RF/bus_reg_dataout[210] , 
        \DataPath/RF/bus_reg_dataout[209] , \DataPath/RF/bus_reg_dataout[208] , 
        \DataPath/RF/bus_reg_dataout[207] , \DataPath/RF/bus_reg_dataout[206] , 
        \DataPath/RF/bus_reg_dataout[205] , \DataPath/RF/bus_reg_dataout[204] , 
        \DataPath/RF/bus_reg_dataout[203] , \DataPath/RF/bus_reg_dataout[202] , 
        \DataPath/RF/bus_reg_dataout[201] , \DataPath/RF/bus_reg_dataout[200] , 
        \DataPath/RF/bus_reg_dataout[199] , \DataPath/RF/bus_reg_dataout[198] , 
        \DataPath/RF/bus_reg_dataout[197] , \DataPath/RF/bus_reg_dataout[196] , 
        \DataPath/RF/bus_reg_dataout[195] , \DataPath/RF/bus_reg_dataout[194] , 
        \DataPath/RF/bus_reg_dataout[193] , \DataPath/RF/bus_reg_dataout[192] , 
        \DataPath/RF/bus_reg_dataout[191] , \DataPath/RF/bus_reg_dataout[190] , 
        \DataPath/RF/bus_reg_dataout[189] , \DataPath/RF/bus_reg_dataout[188] , 
        \DataPath/RF/bus_reg_dataout[187] , \DataPath/RF/bus_reg_dataout[186] , 
        \DataPath/RF/bus_reg_dataout[185] , \DataPath/RF/bus_reg_dataout[184] , 
        \DataPath/RF/bus_reg_dataout[183] , \DataPath/RF/bus_reg_dataout[182] , 
        \DataPath/RF/bus_reg_dataout[181] , \DataPath/RF/bus_reg_dataout[180] , 
        \DataPath/RF/bus_reg_dataout[179] , \DataPath/RF/bus_reg_dataout[178] , 
        \DataPath/RF/bus_reg_dataout[177] , \DataPath/RF/bus_reg_dataout[176] , 
        \DataPath/RF/bus_reg_dataout[175] , \DataPath/RF/bus_reg_dataout[174] , 
        \DataPath/RF/bus_reg_dataout[173] , \DataPath/RF/bus_reg_dataout[172] , 
        \DataPath/RF/bus_reg_dataout[171] , \DataPath/RF/bus_reg_dataout[170] , 
        \DataPath/RF/bus_reg_dataout[169] , \DataPath/RF/bus_reg_dataout[168] , 
        \DataPath/RF/bus_reg_dataout[167] , \DataPath/RF/bus_reg_dataout[166] , 
        \DataPath/RF/bus_reg_dataout[165] , \DataPath/RF/bus_reg_dataout[164] , 
        \DataPath/RF/bus_reg_dataout[163] , \DataPath/RF/bus_reg_dataout[162] , 
        \DataPath/RF/bus_reg_dataout[161] , \DataPath/RF/bus_reg_dataout[160] , 
        \DataPath/RF/bus_reg_dataout[159] , \DataPath/RF/bus_reg_dataout[158] , 
        \DataPath/RF/bus_reg_dataout[157] , \DataPath/RF/bus_reg_dataout[156] , 
        \DataPath/RF/bus_reg_dataout[155] , \DataPath/RF/bus_reg_dataout[154] , 
        \DataPath/RF/bus_reg_dataout[153] , \DataPath/RF/bus_reg_dataout[152] , 
        \DataPath/RF/bus_reg_dataout[151] , \DataPath/RF/bus_reg_dataout[150] , 
        \DataPath/RF/bus_reg_dataout[149] , \DataPath/RF/bus_reg_dataout[148] , 
        \DataPath/RF/bus_reg_dataout[147] , \DataPath/RF/bus_reg_dataout[146] , 
        \DataPath/RF/bus_reg_dataout[145] , \DataPath/RF/bus_reg_dataout[144] , 
        \DataPath/RF/bus_reg_dataout[143] , \DataPath/RF/bus_reg_dataout[142] , 
        \DataPath/RF/bus_reg_dataout[141] , \DataPath/RF/bus_reg_dataout[140] , 
        \DataPath/RF/bus_reg_dataout[139] , \DataPath/RF/bus_reg_dataout[138] , 
        \DataPath/RF/bus_reg_dataout[137] , \DataPath/RF/bus_reg_dataout[136] , 
        \DataPath/RF/bus_reg_dataout[135] , \DataPath/RF/bus_reg_dataout[134] , 
        \DataPath/RF/bus_reg_dataout[133] , \DataPath/RF/bus_reg_dataout[132] , 
        \DataPath/RF/bus_reg_dataout[131] , \DataPath/RF/bus_reg_dataout[130] , 
        \DataPath/RF/bus_reg_dataout[129] , \DataPath/RF/bus_reg_dataout[128] , 
        \DataPath/RF/bus_reg_dataout[127] , \DataPath/RF/bus_reg_dataout[126] , 
        \DataPath/RF/bus_reg_dataout[125] , \DataPath/RF/bus_reg_dataout[124] , 
        \DataPath/RF/bus_reg_dataout[123] , \DataPath/RF/bus_reg_dataout[122] , 
        \DataPath/RF/bus_reg_dataout[121] , \DataPath/RF/bus_reg_dataout[120] , 
        \DataPath/RF/bus_reg_dataout[119] , \DataPath/RF/bus_reg_dataout[118] , 
        \DataPath/RF/bus_reg_dataout[117] , \DataPath/RF/bus_reg_dataout[116] , 
        \DataPath/RF/bus_reg_dataout[115] , \DataPath/RF/bus_reg_dataout[114] , 
        \DataPath/RF/bus_reg_dataout[113] , \DataPath/RF/bus_reg_dataout[112] , 
        \DataPath/RF/bus_reg_dataout[111] , \DataPath/RF/bus_reg_dataout[110] , 
        \DataPath/RF/bus_reg_dataout[109] , \DataPath/RF/bus_reg_dataout[108] , 
        \DataPath/RF/bus_reg_dataout[107] , \DataPath/RF/bus_reg_dataout[106] , 
        \DataPath/RF/bus_reg_dataout[105] , \DataPath/RF/bus_reg_dataout[104] , 
        \DataPath/RF/bus_reg_dataout[103] , \DataPath/RF/bus_reg_dataout[102] , 
        \DataPath/RF/bus_reg_dataout[101] , \DataPath/RF/bus_reg_dataout[100] , 
        \DataPath/RF/bus_reg_dataout[99] , \DataPath/RF/bus_reg_dataout[98] , 
        \DataPath/RF/bus_reg_dataout[97] , \DataPath/RF/bus_reg_dataout[96] , 
        \DataPath/RF/bus_reg_dataout[95] , \DataPath/RF/bus_reg_dataout[94] , 
        \DataPath/RF/bus_reg_dataout[93] , \DataPath/RF/bus_reg_dataout[92] , 
        \DataPath/RF/bus_reg_dataout[91] , \DataPath/RF/bus_reg_dataout[90] , 
        \DataPath/RF/bus_reg_dataout[89] , \DataPath/RF/bus_reg_dataout[88] , 
        \DataPath/RF/bus_reg_dataout[87] , \DataPath/RF/bus_reg_dataout[86] , 
        \DataPath/RF/bus_reg_dataout[85] , \DataPath/RF/bus_reg_dataout[84] , 
        \DataPath/RF/bus_reg_dataout[83] , \DataPath/RF/bus_reg_dataout[82] , 
        \DataPath/RF/bus_reg_dataout[81] , \DataPath/RF/bus_reg_dataout[80] , 
        \DataPath/RF/bus_reg_dataout[79] , \DataPath/RF/bus_reg_dataout[78] , 
        \DataPath/RF/bus_reg_dataout[77] , \DataPath/RF/bus_reg_dataout[76] , 
        \DataPath/RF/bus_reg_dataout[75] , \DataPath/RF/bus_reg_dataout[74] , 
        \DataPath/RF/bus_reg_dataout[73] , \DataPath/RF/bus_reg_dataout[72] , 
        \DataPath/RF/bus_reg_dataout[71] , \DataPath/RF/bus_reg_dataout[70] , 
        \DataPath/RF/bus_reg_dataout[69] , \DataPath/RF/bus_reg_dataout[68] , 
        \DataPath/RF/bus_reg_dataout[67] , \DataPath/RF/bus_reg_dataout[66] , 
        \DataPath/RF/bus_reg_dataout[65] , \DataPath/RF/bus_reg_dataout[64] , 
        \DataPath/RF/bus_reg_dataout[63] , \DataPath/RF/bus_reg_dataout[62] , 
        \DataPath/RF/bus_reg_dataout[61] , \DataPath/RF/bus_reg_dataout[60] , 
        \DataPath/RF/bus_reg_dataout[59] , \DataPath/RF/bus_reg_dataout[58] , 
        \DataPath/RF/bus_reg_dataout[57] , \DataPath/RF/bus_reg_dataout[56] , 
        \DataPath/RF/bus_reg_dataout[55] , \DataPath/RF/bus_reg_dataout[54] , 
        \DataPath/RF/bus_reg_dataout[53] , \DataPath/RF/bus_reg_dataout[52] , 
        \DataPath/RF/bus_reg_dataout[51] , \DataPath/RF/bus_reg_dataout[50] , 
        \DataPath/RF/bus_reg_dataout[49] , \DataPath/RF/bus_reg_dataout[48] , 
        \DataPath/RF/bus_reg_dataout[47] , \DataPath/RF/bus_reg_dataout[46] , 
        \DataPath/RF/bus_reg_dataout[45] , \DataPath/RF/bus_reg_dataout[44] , 
        \DataPath/RF/bus_reg_dataout[43] , \DataPath/RF/bus_reg_dataout[42] , 
        \DataPath/RF/bus_reg_dataout[41] , \DataPath/RF/bus_reg_dataout[40] , 
        \DataPath/RF/bus_reg_dataout[39] , \DataPath/RF/bus_reg_dataout[38] , 
        \DataPath/RF/bus_reg_dataout[37] , \DataPath/RF/bus_reg_dataout[36] , 
        \DataPath/RF/bus_reg_dataout[35] , \DataPath/RF/bus_reg_dataout[34] , 
        \DataPath/RF/bus_reg_dataout[33] , \DataPath/RF/bus_reg_dataout[32] , 
        \DataPath/RF/bus_reg_dataout[31] , \DataPath/RF/bus_reg_dataout[30] , 
        \DataPath/RF/bus_reg_dataout[29] , \DataPath/RF/bus_reg_dataout[28] , 
        \DataPath/RF/bus_reg_dataout[27] , \DataPath/RF/bus_reg_dataout[26] , 
        \DataPath/RF/bus_reg_dataout[25] , \DataPath/RF/bus_reg_dataout[24] , 
        \DataPath/RF/bus_reg_dataout[23] , \DataPath/RF/bus_reg_dataout[22] , 
        \DataPath/RF/bus_reg_dataout[21] , \DataPath/RF/bus_reg_dataout[20] , 
        \DataPath/RF/bus_reg_dataout[19] , \DataPath/RF/bus_reg_dataout[18] , 
        \DataPath/RF/bus_reg_dataout[17] , \DataPath/RF/bus_reg_dataout[16] , 
        \DataPath/RF/bus_reg_dataout[15] , \DataPath/RF/bus_reg_dataout[14] , 
        \DataPath/RF/bus_reg_dataout[13] , \DataPath/RF/bus_reg_dataout[12] , 
        \DataPath/RF/bus_reg_dataout[11] , \DataPath/RF/bus_reg_dataout[10] , 
        \DataPath/RF/bus_reg_dataout[9] , \DataPath/RF/bus_reg_dataout[8] , 
        \DataPath/RF/bus_reg_dataout[7] , \DataPath/RF/bus_reg_dataout[6] , 
        \DataPath/RF/bus_reg_dataout[5] , \DataPath/RF/bus_reg_dataout[4] , 
        \DataPath/RF/bus_reg_dataout[3] , \DataPath/RF/bus_reg_dataout[2] , 
        \DataPath/RF/bus_reg_dataout[1] , \DataPath/RF/bus_reg_dataout[0] }), 
        .win({n7648, \DataPath/RF/c_win[3] , \DataPath/RF/c_win[2] , n8275, 
        \DataPath/RF/c_win[0] }), .curr_proc_regs({
        \DataPath/RF/bus_selected_win_data[767] , 
        \DataPath/RF/bus_selected_win_data[766] , 
        \DataPath/RF/bus_selected_win_data[765] , 
        \DataPath/RF/bus_selected_win_data[764] , 
        \DataPath/RF/bus_selected_win_data[763] , 
        \DataPath/RF/bus_selected_win_data[762] , 
        \DataPath/RF/bus_selected_win_data[761] , 
        \DataPath/RF/bus_selected_win_data[760] , 
        \DataPath/RF/bus_selected_win_data[759] , 
        \DataPath/RF/bus_selected_win_data[758] , 
        \DataPath/RF/bus_selected_win_data[757] , 
        \DataPath/RF/bus_selected_win_data[756] , 
        \DataPath/RF/bus_selected_win_data[755] , 
        \DataPath/RF/bus_selected_win_data[754] , 
        \DataPath/RF/bus_selected_win_data[753] , 
        \DataPath/RF/bus_selected_win_data[752] , 
        \DataPath/RF/bus_selected_win_data[751] , 
        \DataPath/RF/bus_selected_win_data[750] , 
        \DataPath/RF/bus_selected_win_data[749] , 
        \DataPath/RF/bus_selected_win_data[748] , 
        \DataPath/RF/bus_selected_win_data[747] , 
        \DataPath/RF/bus_selected_win_data[746] , 
        \DataPath/RF/bus_selected_win_data[745] , 
        \DataPath/RF/bus_selected_win_data[744] , 
        \DataPath/RF/bus_selected_win_data[743] , 
        \DataPath/RF/bus_selected_win_data[742] , 
        \DataPath/RF/bus_selected_win_data[741] , 
        \DataPath/RF/bus_selected_win_data[740] , 
        \DataPath/RF/bus_selected_win_data[739] , 
        \DataPath/RF/bus_selected_win_data[738] , 
        \DataPath/RF/bus_selected_win_data[737] , 
        \DataPath/RF/bus_selected_win_data[736] , 
        \DataPath/RF/bus_selected_win_data[735] , 
        \DataPath/RF/bus_selected_win_data[734] , 
        \DataPath/RF/bus_selected_win_data[733] , 
        \DataPath/RF/bus_selected_win_data[732] , 
        \DataPath/RF/bus_selected_win_data[731] , 
        \DataPath/RF/bus_selected_win_data[730] , 
        \DataPath/RF/bus_selected_win_data[729] , 
        \DataPath/RF/bus_selected_win_data[728] , 
        \DataPath/RF/bus_selected_win_data[727] , 
        \DataPath/RF/bus_selected_win_data[726] , 
        \DataPath/RF/bus_selected_win_data[725] , 
        \DataPath/RF/bus_selected_win_data[724] , 
        \DataPath/RF/bus_selected_win_data[723] , 
        \DataPath/RF/bus_selected_win_data[722] , 
        \DataPath/RF/bus_selected_win_data[721] , 
        \DataPath/RF/bus_selected_win_data[720] , 
        \DataPath/RF/bus_selected_win_data[719] , 
        \DataPath/RF/bus_selected_win_data[718] , 
        \DataPath/RF/bus_selected_win_data[717] , 
        \DataPath/RF/bus_selected_win_data[716] , 
        \DataPath/RF/bus_selected_win_data[715] , 
        \DataPath/RF/bus_selected_win_data[714] , 
        \DataPath/RF/bus_selected_win_data[713] , 
        \DataPath/RF/bus_selected_win_data[712] , 
        \DataPath/RF/bus_selected_win_data[711] , 
        \DataPath/RF/bus_selected_win_data[710] , 
        \DataPath/RF/bus_selected_win_data[709] , 
        \DataPath/RF/bus_selected_win_data[708] , 
        \DataPath/RF/bus_selected_win_data[707] , 
        \DataPath/RF/bus_selected_win_data[706] , 
        \DataPath/RF/bus_selected_win_data[705] , 
        \DataPath/RF/bus_selected_win_data[704] , 
        \DataPath/RF/bus_selected_win_data[703] , 
        \DataPath/RF/bus_selected_win_data[702] , 
        \DataPath/RF/bus_selected_win_data[701] , 
        \DataPath/RF/bus_selected_win_data[700] , 
        \DataPath/RF/bus_selected_win_data[699] , 
        \DataPath/RF/bus_selected_win_data[698] , 
        \DataPath/RF/bus_selected_win_data[697] , 
        \DataPath/RF/bus_selected_win_data[696] , 
        \DataPath/RF/bus_selected_win_data[695] , 
        \DataPath/RF/bus_selected_win_data[694] , 
        \DataPath/RF/bus_selected_win_data[693] , 
        \DataPath/RF/bus_selected_win_data[692] , 
        \DataPath/RF/bus_selected_win_data[691] , 
        \DataPath/RF/bus_selected_win_data[690] , 
        \DataPath/RF/bus_selected_win_data[689] , 
        \DataPath/RF/bus_selected_win_data[688] , 
        \DataPath/RF/bus_selected_win_data[687] , 
        \DataPath/RF/bus_selected_win_data[686] , 
        \DataPath/RF/bus_selected_win_data[685] , 
        \DataPath/RF/bus_selected_win_data[684] , 
        \DataPath/RF/bus_selected_win_data[683] , 
        \DataPath/RF/bus_selected_win_data[682] , 
        \DataPath/RF/bus_selected_win_data[681] , 
        \DataPath/RF/bus_selected_win_data[680] , 
        \DataPath/RF/bus_selected_win_data[679] , 
        \DataPath/RF/bus_selected_win_data[678] , 
        \DataPath/RF/bus_selected_win_data[677] , 
        \DataPath/RF/bus_selected_win_data[676] , 
        \DataPath/RF/bus_selected_win_data[675] , 
        \DataPath/RF/bus_selected_win_data[674] , 
        \DataPath/RF/bus_selected_win_data[673] , 
        \DataPath/RF/bus_selected_win_data[672] , 
        \DataPath/RF/bus_selected_win_data[671] , 
        \DataPath/RF/bus_selected_win_data[670] , 
        \DataPath/RF/bus_selected_win_data[669] , 
        \DataPath/RF/bus_selected_win_data[668] , 
        \DataPath/RF/bus_selected_win_data[667] , 
        \DataPath/RF/bus_selected_win_data[666] , 
        \DataPath/RF/bus_selected_win_data[665] , 
        \DataPath/RF/bus_selected_win_data[664] , 
        \DataPath/RF/bus_selected_win_data[663] , 
        \DataPath/RF/bus_selected_win_data[662] , 
        \DataPath/RF/bus_selected_win_data[661] , 
        \DataPath/RF/bus_selected_win_data[660] , 
        \DataPath/RF/bus_selected_win_data[659] , 
        \DataPath/RF/bus_selected_win_data[658] , 
        \DataPath/RF/bus_selected_win_data[657] , 
        \DataPath/RF/bus_selected_win_data[656] , 
        \DataPath/RF/bus_selected_win_data[655] , 
        \DataPath/RF/bus_selected_win_data[654] , 
        \DataPath/RF/bus_selected_win_data[653] , 
        \DataPath/RF/bus_selected_win_data[652] , 
        \DataPath/RF/bus_selected_win_data[651] , 
        \DataPath/RF/bus_selected_win_data[650] , 
        \DataPath/RF/bus_selected_win_data[649] , 
        \DataPath/RF/bus_selected_win_data[648] , 
        \DataPath/RF/bus_selected_win_data[647] , 
        \DataPath/RF/bus_selected_win_data[646] , 
        \DataPath/RF/bus_selected_win_data[645] , 
        \DataPath/RF/bus_selected_win_data[644] , 
        \DataPath/RF/bus_selected_win_data[643] , 
        \DataPath/RF/bus_selected_win_data[642] , 
        \DataPath/RF/bus_selected_win_data[641] , 
        \DataPath/RF/bus_selected_win_data[640] , 
        \DataPath/RF/bus_selected_win_data[639] , 
        \DataPath/RF/bus_selected_win_data[638] , 
        \DataPath/RF/bus_selected_win_data[637] , 
        \DataPath/RF/bus_selected_win_data[636] , 
        \DataPath/RF/bus_selected_win_data[635] , 
        \DataPath/RF/bus_selected_win_data[634] , 
        \DataPath/RF/bus_selected_win_data[633] , 
        \DataPath/RF/bus_selected_win_data[632] , 
        \DataPath/RF/bus_selected_win_data[631] , 
        \DataPath/RF/bus_selected_win_data[630] , 
        \DataPath/RF/bus_selected_win_data[629] , 
        \DataPath/RF/bus_selected_win_data[628] , 
        \DataPath/RF/bus_selected_win_data[627] , 
        \DataPath/RF/bus_selected_win_data[626] , 
        \DataPath/RF/bus_selected_win_data[625] , 
        \DataPath/RF/bus_selected_win_data[624] , 
        \DataPath/RF/bus_selected_win_data[623] , 
        \DataPath/RF/bus_selected_win_data[622] , 
        \DataPath/RF/bus_selected_win_data[621] , 
        \DataPath/RF/bus_selected_win_data[620] , 
        \DataPath/RF/bus_selected_win_data[619] , 
        \DataPath/RF/bus_selected_win_data[618] , 
        \DataPath/RF/bus_selected_win_data[617] , 
        \DataPath/RF/bus_selected_win_data[616] , 
        \DataPath/RF/bus_selected_win_data[615] , 
        \DataPath/RF/bus_selected_win_data[614] , 
        \DataPath/RF/bus_selected_win_data[613] , 
        \DataPath/RF/bus_selected_win_data[612] , 
        \DataPath/RF/bus_selected_win_data[611] , 
        \DataPath/RF/bus_selected_win_data[610] , 
        \DataPath/RF/bus_selected_win_data[609] , 
        \DataPath/RF/bus_selected_win_data[608] , 
        \DataPath/RF/bus_selected_win_data[607] , 
        \DataPath/RF/bus_selected_win_data[606] , 
        \DataPath/RF/bus_selected_win_data[605] , 
        \DataPath/RF/bus_selected_win_data[604] , 
        \DataPath/RF/bus_selected_win_data[603] , 
        \DataPath/RF/bus_selected_win_data[602] , 
        \DataPath/RF/bus_selected_win_data[601] , 
        \DataPath/RF/bus_selected_win_data[600] , 
        \DataPath/RF/bus_selected_win_data[599] , 
        \DataPath/RF/bus_selected_win_data[598] , 
        \DataPath/RF/bus_selected_win_data[597] , 
        \DataPath/RF/bus_selected_win_data[596] , 
        \DataPath/RF/bus_selected_win_data[595] , 
        \DataPath/RF/bus_selected_win_data[594] , 
        \DataPath/RF/bus_selected_win_data[593] , 
        \DataPath/RF/bus_selected_win_data[592] , 
        \DataPath/RF/bus_selected_win_data[591] , 
        \DataPath/RF/bus_selected_win_data[590] , 
        \DataPath/RF/bus_selected_win_data[589] , 
        \DataPath/RF/bus_selected_win_data[588] , 
        \DataPath/RF/bus_selected_win_data[587] , 
        \DataPath/RF/bus_selected_win_data[586] , 
        \DataPath/RF/bus_selected_win_data[585] , 
        \DataPath/RF/bus_selected_win_data[584] , 
        \DataPath/RF/bus_selected_win_data[583] , 
        \DataPath/RF/bus_selected_win_data[582] , 
        \DataPath/RF/bus_selected_win_data[581] , 
        \DataPath/RF/bus_selected_win_data[580] , 
        \DataPath/RF/bus_selected_win_data[579] , 
        \DataPath/RF/bus_selected_win_data[578] , 
        \DataPath/RF/bus_selected_win_data[577] , 
        \DataPath/RF/bus_selected_win_data[576] , 
        \DataPath/RF/bus_selected_win_data[575] , 
        \DataPath/RF/bus_selected_win_data[574] , 
        \DataPath/RF/bus_selected_win_data[573] , 
        \DataPath/RF/bus_selected_win_data[572] , 
        \DataPath/RF/bus_selected_win_data[571] , 
        \DataPath/RF/bus_selected_win_data[570] , 
        \DataPath/RF/bus_selected_win_data[569] , 
        \DataPath/RF/bus_selected_win_data[568] , 
        \DataPath/RF/bus_selected_win_data[567] , 
        \DataPath/RF/bus_selected_win_data[566] , 
        \DataPath/RF/bus_selected_win_data[565] , 
        \DataPath/RF/bus_selected_win_data[564] , 
        \DataPath/RF/bus_selected_win_data[563] , 
        \DataPath/RF/bus_selected_win_data[562] , 
        \DataPath/RF/bus_selected_win_data[561] , 
        \DataPath/RF/bus_selected_win_data[560] , 
        \DataPath/RF/bus_selected_win_data[559] , 
        \DataPath/RF/bus_selected_win_data[558] , 
        \DataPath/RF/bus_selected_win_data[557] , 
        \DataPath/RF/bus_selected_win_data[556] , 
        \DataPath/RF/bus_selected_win_data[555] , 
        \DataPath/RF/bus_selected_win_data[554] , 
        \DataPath/RF/bus_selected_win_data[553] , 
        \DataPath/RF/bus_selected_win_data[552] , 
        \DataPath/RF/bus_selected_win_data[551] , 
        \DataPath/RF/bus_selected_win_data[550] , 
        \DataPath/RF/bus_selected_win_data[549] , 
        \DataPath/RF/bus_selected_win_data[548] , 
        \DataPath/RF/bus_selected_win_data[547] , 
        \DataPath/RF/bus_selected_win_data[546] , 
        \DataPath/RF/bus_selected_win_data[545] , 
        \DataPath/RF/bus_selected_win_data[544] , 
        \DataPath/RF/bus_selected_win_data[543] , 
        \DataPath/RF/bus_selected_win_data[542] , 
        \DataPath/RF/bus_selected_win_data[541] , 
        \DataPath/RF/bus_selected_win_data[540] , 
        \DataPath/RF/bus_selected_win_data[539] , 
        \DataPath/RF/bus_selected_win_data[538] , 
        \DataPath/RF/bus_selected_win_data[537] , 
        \DataPath/RF/bus_selected_win_data[536] , 
        \DataPath/RF/bus_selected_win_data[535] , 
        \DataPath/RF/bus_selected_win_data[534] , 
        \DataPath/RF/bus_selected_win_data[533] , 
        \DataPath/RF/bus_selected_win_data[532] , 
        \DataPath/RF/bus_selected_win_data[531] , 
        \DataPath/RF/bus_selected_win_data[530] , 
        \DataPath/RF/bus_selected_win_data[529] , 
        \DataPath/RF/bus_selected_win_data[528] , 
        \DataPath/RF/bus_selected_win_data[527] , 
        \DataPath/RF/bus_selected_win_data[526] , 
        \DataPath/RF/bus_selected_win_data[525] , 
        \DataPath/RF/bus_selected_win_data[524] , 
        \DataPath/RF/bus_selected_win_data[523] , 
        \DataPath/RF/bus_selected_win_data[522] , 
        \DataPath/RF/bus_selected_win_data[521] , 
        \DataPath/RF/bus_selected_win_data[520] , 
        \DataPath/RF/bus_selected_win_data[519] , 
        \DataPath/RF/bus_selected_win_data[518] , 
        \DataPath/RF/bus_selected_win_data[517] , 
        \DataPath/RF/bus_selected_win_data[516] , 
        \DataPath/RF/bus_selected_win_data[515] , 
        \DataPath/RF/bus_selected_win_data[514] , 
        \DataPath/RF/bus_selected_win_data[513] , 
        \DataPath/RF/bus_selected_win_data[512] , 
        \DataPath/RF/bus_selected_win_data[511] , 
        \DataPath/RF/bus_selected_win_data[510] , 
        \DataPath/RF/bus_selected_win_data[509] , 
        \DataPath/RF/bus_selected_win_data[508] , 
        \DataPath/RF/bus_selected_win_data[507] , 
        \DataPath/RF/bus_selected_win_data[506] , 
        \DataPath/RF/bus_selected_win_data[505] , 
        \DataPath/RF/bus_selected_win_data[504] , 
        \DataPath/RF/bus_selected_win_data[503] , 
        \DataPath/RF/bus_selected_win_data[502] , 
        \DataPath/RF/bus_selected_win_data[501] , 
        \DataPath/RF/bus_selected_win_data[500] , 
        \DataPath/RF/bus_selected_win_data[499] , 
        \DataPath/RF/bus_selected_win_data[498] , 
        \DataPath/RF/bus_selected_win_data[497] , 
        \DataPath/RF/bus_selected_win_data[496] , 
        \DataPath/RF/bus_selected_win_data[495] , 
        \DataPath/RF/bus_selected_win_data[494] , 
        \DataPath/RF/bus_selected_win_data[493] , 
        \DataPath/RF/bus_selected_win_data[492] , 
        \DataPath/RF/bus_selected_win_data[491] , 
        \DataPath/RF/bus_selected_win_data[490] , 
        \DataPath/RF/bus_selected_win_data[489] , 
        \DataPath/RF/bus_selected_win_data[488] , 
        \DataPath/RF/bus_selected_win_data[487] , 
        \DataPath/RF/bus_selected_win_data[486] , 
        \DataPath/RF/bus_selected_win_data[485] , 
        \DataPath/RF/bus_selected_win_data[484] , 
        \DataPath/RF/bus_selected_win_data[483] , 
        \DataPath/RF/bus_selected_win_data[482] , 
        \DataPath/RF/bus_selected_win_data[481] , 
        \DataPath/RF/bus_selected_win_data[480] , 
        \DataPath/RF/bus_selected_win_data[479] , 
        \DataPath/RF/bus_selected_win_data[478] , 
        \DataPath/RF/bus_selected_win_data[477] , 
        \DataPath/RF/bus_selected_win_data[476] , 
        \DataPath/RF/bus_selected_win_data[475] , 
        \DataPath/RF/bus_selected_win_data[474] , 
        \DataPath/RF/bus_selected_win_data[473] , 
        \DataPath/RF/bus_selected_win_data[472] , 
        \DataPath/RF/bus_selected_win_data[471] , 
        \DataPath/RF/bus_selected_win_data[470] , 
        \DataPath/RF/bus_selected_win_data[469] , 
        \DataPath/RF/bus_selected_win_data[468] , 
        \DataPath/RF/bus_selected_win_data[467] , 
        \DataPath/RF/bus_selected_win_data[466] , 
        \DataPath/RF/bus_selected_win_data[465] , 
        \DataPath/RF/bus_selected_win_data[464] , 
        \DataPath/RF/bus_selected_win_data[463] , 
        \DataPath/RF/bus_selected_win_data[462] , 
        \DataPath/RF/bus_selected_win_data[461] , 
        \DataPath/RF/bus_selected_win_data[460] , 
        \DataPath/RF/bus_selected_win_data[459] , 
        \DataPath/RF/bus_selected_win_data[458] , 
        \DataPath/RF/bus_selected_win_data[457] , 
        \DataPath/RF/bus_selected_win_data[456] , 
        \DataPath/RF/bus_selected_win_data[455] , 
        \DataPath/RF/bus_selected_win_data[454] , 
        \DataPath/RF/bus_selected_win_data[453] , 
        \DataPath/RF/bus_selected_win_data[452] , 
        \DataPath/RF/bus_selected_win_data[451] , 
        \DataPath/RF/bus_selected_win_data[450] , 
        \DataPath/RF/bus_selected_win_data[449] , 
        \DataPath/RF/bus_selected_win_data[448] , 
        \DataPath/RF/bus_selected_win_data[447] , 
        \DataPath/RF/bus_selected_win_data[446] , 
        \DataPath/RF/bus_selected_win_data[445] , 
        \DataPath/RF/bus_selected_win_data[444] , 
        \DataPath/RF/bus_selected_win_data[443] , 
        \DataPath/RF/bus_selected_win_data[442] , 
        \DataPath/RF/bus_selected_win_data[441] , 
        \DataPath/RF/bus_selected_win_data[440] , 
        \DataPath/RF/bus_selected_win_data[439] , 
        \DataPath/RF/bus_selected_win_data[438] , 
        \DataPath/RF/bus_selected_win_data[437] , 
        \DataPath/RF/bus_selected_win_data[436] , 
        \DataPath/RF/bus_selected_win_data[435] , 
        \DataPath/RF/bus_selected_win_data[434] , 
        \DataPath/RF/bus_selected_win_data[433] , 
        \DataPath/RF/bus_selected_win_data[432] , 
        \DataPath/RF/bus_selected_win_data[431] , 
        \DataPath/RF/bus_selected_win_data[430] , 
        \DataPath/RF/bus_selected_win_data[429] , 
        \DataPath/RF/bus_selected_win_data[428] , 
        \DataPath/RF/bus_selected_win_data[427] , 
        \DataPath/RF/bus_selected_win_data[426] , 
        \DataPath/RF/bus_selected_win_data[425] , 
        \DataPath/RF/bus_selected_win_data[424] , 
        \DataPath/RF/bus_selected_win_data[423] , 
        \DataPath/RF/bus_selected_win_data[422] , 
        \DataPath/RF/bus_selected_win_data[421] , 
        \DataPath/RF/bus_selected_win_data[420] , 
        \DataPath/RF/bus_selected_win_data[419] , 
        \DataPath/RF/bus_selected_win_data[418] , 
        \DataPath/RF/bus_selected_win_data[417] , 
        \DataPath/RF/bus_selected_win_data[416] , 
        \DataPath/RF/bus_selected_win_data[415] , 
        \DataPath/RF/bus_selected_win_data[414] , 
        \DataPath/RF/bus_selected_win_data[413] , 
        \DataPath/RF/bus_selected_win_data[412] , 
        \DataPath/RF/bus_selected_win_data[411] , 
        \DataPath/RF/bus_selected_win_data[410] , 
        \DataPath/RF/bus_selected_win_data[409] , 
        \DataPath/RF/bus_selected_win_data[408] , 
        \DataPath/RF/bus_selected_win_data[407] , 
        \DataPath/RF/bus_selected_win_data[406] , 
        \DataPath/RF/bus_selected_win_data[405] , 
        \DataPath/RF/bus_selected_win_data[404] , 
        \DataPath/RF/bus_selected_win_data[403] , 
        \DataPath/RF/bus_selected_win_data[402] , 
        \DataPath/RF/bus_selected_win_data[401] , 
        \DataPath/RF/bus_selected_win_data[400] , 
        \DataPath/RF/bus_selected_win_data[399] , 
        \DataPath/RF/bus_selected_win_data[398] , 
        \DataPath/RF/bus_selected_win_data[397] , 
        \DataPath/RF/bus_selected_win_data[396] , 
        \DataPath/RF/bus_selected_win_data[395] , 
        \DataPath/RF/bus_selected_win_data[394] , 
        \DataPath/RF/bus_selected_win_data[393] , 
        \DataPath/RF/bus_selected_win_data[392] , 
        \DataPath/RF/bus_selected_win_data[391] , 
        \DataPath/RF/bus_selected_win_data[390] , 
        \DataPath/RF/bus_selected_win_data[389] , 
        \DataPath/RF/bus_selected_win_data[388] , 
        \DataPath/RF/bus_selected_win_data[387] , 
        \DataPath/RF/bus_selected_win_data[386] , 
        \DataPath/RF/bus_selected_win_data[385] , 
        \DataPath/RF/bus_selected_win_data[384] , 
        \DataPath/RF/bus_selected_win_data[383] , 
        \DataPath/RF/bus_selected_win_data[382] , 
        \DataPath/RF/bus_selected_win_data[381] , 
        \DataPath/RF/bus_selected_win_data[380] , 
        \DataPath/RF/bus_selected_win_data[379] , 
        \DataPath/RF/bus_selected_win_data[378] , 
        \DataPath/RF/bus_selected_win_data[377] , 
        \DataPath/RF/bus_selected_win_data[376] , 
        \DataPath/RF/bus_selected_win_data[375] , 
        \DataPath/RF/bus_selected_win_data[374] , 
        \DataPath/RF/bus_selected_win_data[373] , 
        \DataPath/RF/bus_selected_win_data[372] , 
        \DataPath/RF/bus_selected_win_data[371] , 
        \DataPath/RF/bus_selected_win_data[370] , 
        \DataPath/RF/bus_selected_win_data[369] , 
        \DataPath/RF/bus_selected_win_data[368] , 
        \DataPath/RF/bus_selected_win_data[367] , 
        \DataPath/RF/bus_selected_win_data[366] , 
        \DataPath/RF/bus_selected_win_data[365] , 
        \DataPath/RF/bus_selected_win_data[364] , 
        \DataPath/RF/bus_selected_win_data[363] , 
        \DataPath/RF/bus_selected_win_data[362] , 
        \DataPath/RF/bus_selected_win_data[361] , 
        \DataPath/RF/bus_selected_win_data[360] , 
        \DataPath/RF/bus_selected_win_data[359] , 
        \DataPath/RF/bus_selected_win_data[358] , 
        \DataPath/RF/bus_selected_win_data[357] , 
        \DataPath/RF/bus_selected_win_data[356] , 
        \DataPath/RF/bus_selected_win_data[355] , 
        \DataPath/RF/bus_selected_win_data[354] , 
        \DataPath/RF/bus_selected_win_data[353] , 
        \DataPath/RF/bus_selected_win_data[352] , 
        \DataPath/RF/bus_selected_win_data[351] , 
        \DataPath/RF/bus_selected_win_data[350] , 
        \DataPath/RF/bus_selected_win_data[349] , 
        \DataPath/RF/bus_selected_win_data[348] , 
        \DataPath/RF/bus_selected_win_data[347] , 
        \DataPath/RF/bus_selected_win_data[346] , 
        \DataPath/RF/bus_selected_win_data[345] , 
        \DataPath/RF/bus_selected_win_data[344] , 
        \DataPath/RF/bus_selected_win_data[343] , 
        \DataPath/RF/bus_selected_win_data[342] , 
        \DataPath/RF/bus_selected_win_data[341] , 
        \DataPath/RF/bus_selected_win_data[340] , 
        \DataPath/RF/bus_selected_win_data[339] , 
        \DataPath/RF/bus_selected_win_data[338] , 
        \DataPath/RF/bus_selected_win_data[337] , 
        \DataPath/RF/bus_selected_win_data[336] , 
        \DataPath/RF/bus_selected_win_data[335] , 
        \DataPath/RF/bus_selected_win_data[334] , 
        \DataPath/RF/bus_selected_win_data[333] , 
        \DataPath/RF/bus_selected_win_data[332] , 
        \DataPath/RF/bus_selected_win_data[331] , 
        \DataPath/RF/bus_selected_win_data[330] , 
        \DataPath/RF/bus_selected_win_data[329] , 
        \DataPath/RF/bus_selected_win_data[328] , 
        \DataPath/RF/bus_selected_win_data[327] , 
        \DataPath/RF/bus_selected_win_data[326] , 
        \DataPath/RF/bus_selected_win_data[325] , 
        \DataPath/RF/bus_selected_win_data[324] , 
        \DataPath/RF/bus_selected_win_data[323] , 
        \DataPath/RF/bus_selected_win_data[322] , 
        \DataPath/RF/bus_selected_win_data[321] , 
        \DataPath/RF/bus_selected_win_data[320] , 
        \DataPath/RF/bus_selected_win_data[319] , 
        \DataPath/RF/bus_selected_win_data[318] , 
        \DataPath/RF/bus_selected_win_data[317] , 
        \DataPath/RF/bus_selected_win_data[316] , 
        \DataPath/RF/bus_selected_win_data[315] , 
        \DataPath/RF/bus_selected_win_data[314] , 
        \DataPath/RF/bus_selected_win_data[313] , 
        \DataPath/RF/bus_selected_win_data[312] , 
        \DataPath/RF/bus_selected_win_data[311] , 
        \DataPath/RF/bus_selected_win_data[310] , 
        \DataPath/RF/bus_selected_win_data[309] , 
        \DataPath/RF/bus_selected_win_data[308] , 
        \DataPath/RF/bus_selected_win_data[307] , 
        \DataPath/RF/bus_selected_win_data[306] , 
        \DataPath/RF/bus_selected_win_data[305] , 
        \DataPath/RF/bus_selected_win_data[304] , 
        \DataPath/RF/bus_selected_win_data[303] , 
        \DataPath/RF/bus_selected_win_data[302] , 
        \DataPath/RF/bus_selected_win_data[301] , 
        \DataPath/RF/bus_selected_win_data[300] , 
        \DataPath/RF/bus_selected_win_data[299] , 
        \DataPath/RF/bus_selected_win_data[298] , 
        \DataPath/RF/bus_selected_win_data[297] , 
        \DataPath/RF/bus_selected_win_data[296] , 
        \DataPath/RF/bus_selected_win_data[295] , 
        \DataPath/RF/bus_selected_win_data[294] , 
        \DataPath/RF/bus_selected_win_data[293] , 
        \DataPath/RF/bus_selected_win_data[292] , 
        \DataPath/RF/bus_selected_win_data[291] , 
        \DataPath/RF/bus_selected_win_data[290] , 
        \DataPath/RF/bus_selected_win_data[289] , 
        \DataPath/RF/bus_selected_win_data[288] , 
        \DataPath/RF/bus_selected_win_data[287] , 
        \DataPath/RF/bus_selected_win_data[286] , 
        \DataPath/RF/bus_selected_win_data[285] , 
        \DataPath/RF/bus_selected_win_data[284] , 
        \DataPath/RF/bus_selected_win_data[283] , 
        \DataPath/RF/bus_selected_win_data[282] , 
        \DataPath/RF/bus_selected_win_data[281] , 
        \DataPath/RF/bus_selected_win_data[280] , 
        \DataPath/RF/bus_selected_win_data[279] , 
        \DataPath/RF/bus_selected_win_data[278] , 
        \DataPath/RF/bus_selected_win_data[277] , 
        \DataPath/RF/bus_selected_win_data[276] , 
        \DataPath/RF/bus_selected_win_data[275] , 
        \DataPath/RF/bus_selected_win_data[274] , 
        \DataPath/RF/bus_selected_win_data[273] , 
        \DataPath/RF/bus_selected_win_data[272] , 
        \DataPath/RF/bus_selected_win_data[271] , 
        \DataPath/RF/bus_selected_win_data[270] , 
        \DataPath/RF/bus_selected_win_data[269] , 
        \DataPath/RF/bus_selected_win_data[268] , 
        \DataPath/RF/bus_selected_win_data[267] , 
        \DataPath/RF/bus_selected_win_data[266] , 
        \DataPath/RF/bus_selected_win_data[265] , 
        \DataPath/RF/bus_selected_win_data[264] , 
        \DataPath/RF/bus_selected_win_data[263] , 
        \DataPath/RF/bus_selected_win_data[262] , 
        \DataPath/RF/bus_selected_win_data[261] , 
        \DataPath/RF/bus_selected_win_data[260] , 
        \DataPath/RF/bus_selected_win_data[259] , 
        \DataPath/RF/bus_selected_win_data[258] , 
        \DataPath/RF/bus_selected_win_data[257] , 
        \DataPath/RF/bus_selected_win_data[256] , 
        \DataPath/RF/bus_selected_win_data[255] , 
        \DataPath/RF/bus_selected_win_data[254] , 
        \DataPath/RF/bus_selected_win_data[253] , 
        \DataPath/RF/bus_selected_win_data[252] , 
        \DataPath/RF/bus_selected_win_data[251] , 
        \DataPath/RF/bus_selected_win_data[250] , 
        \DataPath/RF/bus_selected_win_data[249] , 
        \DataPath/RF/bus_selected_win_data[248] , 
        \DataPath/RF/bus_selected_win_data[247] , 
        \DataPath/RF/bus_selected_win_data[246] , 
        \DataPath/RF/bus_selected_win_data[245] , 
        \DataPath/RF/bus_selected_win_data[244] , 
        \DataPath/RF/bus_selected_win_data[243] , 
        \DataPath/RF/bus_selected_win_data[242] , 
        \DataPath/RF/bus_selected_win_data[241] , 
        \DataPath/RF/bus_selected_win_data[240] , 
        \DataPath/RF/bus_selected_win_data[239] , 
        \DataPath/RF/bus_selected_win_data[238] , 
        \DataPath/RF/bus_selected_win_data[237] , 
        \DataPath/RF/bus_selected_win_data[236] , 
        \DataPath/RF/bus_selected_win_data[235] , 
        \DataPath/RF/bus_selected_win_data[234] , 
        \DataPath/RF/bus_selected_win_data[233] , 
        \DataPath/RF/bus_selected_win_data[232] , 
        \DataPath/RF/bus_selected_win_data[231] , 
        \DataPath/RF/bus_selected_win_data[230] , 
        \DataPath/RF/bus_selected_win_data[229] , 
        \DataPath/RF/bus_selected_win_data[228] , 
        \DataPath/RF/bus_selected_win_data[227] , 
        \DataPath/RF/bus_selected_win_data[226] , 
        \DataPath/RF/bus_selected_win_data[225] , 
        \DataPath/RF/bus_selected_win_data[224] , 
        \DataPath/RF/bus_selected_win_data[223] , 
        \DataPath/RF/bus_selected_win_data[222] , 
        \DataPath/RF/bus_selected_win_data[221] , 
        \DataPath/RF/bus_selected_win_data[220] , 
        \DataPath/RF/bus_selected_win_data[219] , 
        \DataPath/RF/bus_selected_win_data[218] , 
        \DataPath/RF/bus_selected_win_data[217] , 
        \DataPath/RF/bus_selected_win_data[216] , 
        \DataPath/RF/bus_selected_win_data[215] , 
        \DataPath/RF/bus_selected_win_data[214] , 
        \DataPath/RF/bus_selected_win_data[213] , 
        \DataPath/RF/bus_selected_win_data[212] , 
        \DataPath/RF/bus_selected_win_data[211] , 
        \DataPath/RF/bus_selected_win_data[210] , 
        \DataPath/RF/bus_selected_win_data[209] , 
        \DataPath/RF/bus_selected_win_data[208] , 
        \DataPath/RF/bus_selected_win_data[207] , 
        \DataPath/RF/bus_selected_win_data[206] , 
        \DataPath/RF/bus_selected_win_data[205] , 
        \DataPath/RF/bus_selected_win_data[204] , 
        \DataPath/RF/bus_selected_win_data[203] , 
        \DataPath/RF/bus_selected_win_data[202] , 
        \DataPath/RF/bus_selected_win_data[201] , 
        \DataPath/RF/bus_selected_win_data[200] , 
        \DataPath/RF/bus_selected_win_data[199] , 
        \DataPath/RF/bus_selected_win_data[198] , 
        \DataPath/RF/bus_selected_win_data[197] , 
        \DataPath/RF/bus_selected_win_data[196] , 
        \DataPath/RF/bus_selected_win_data[195] , 
        \DataPath/RF/bus_selected_win_data[194] , 
        \DataPath/RF/bus_selected_win_data[193] , 
        \DataPath/RF/bus_selected_win_data[192] , 
        \DataPath/RF/bus_selected_win_data[191] , 
        \DataPath/RF/bus_selected_win_data[190] , 
        \DataPath/RF/bus_selected_win_data[189] , 
        \DataPath/RF/bus_selected_win_data[188] , 
        \DataPath/RF/bus_selected_win_data[187] , 
        \DataPath/RF/bus_selected_win_data[186] , 
        \DataPath/RF/bus_selected_win_data[185] , 
        \DataPath/RF/bus_selected_win_data[184] , 
        \DataPath/RF/bus_selected_win_data[183] , 
        \DataPath/RF/bus_selected_win_data[182] , 
        \DataPath/RF/bus_selected_win_data[181] , 
        \DataPath/RF/bus_selected_win_data[180] , 
        \DataPath/RF/bus_selected_win_data[179] , 
        \DataPath/RF/bus_selected_win_data[178] , 
        \DataPath/RF/bus_selected_win_data[177] , 
        \DataPath/RF/bus_selected_win_data[176] , 
        \DataPath/RF/bus_selected_win_data[175] , 
        \DataPath/RF/bus_selected_win_data[174] , 
        \DataPath/RF/bus_selected_win_data[173] , 
        \DataPath/RF/bus_selected_win_data[172] , 
        \DataPath/RF/bus_selected_win_data[171] , 
        \DataPath/RF/bus_selected_win_data[170] , 
        \DataPath/RF/bus_selected_win_data[169] , 
        \DataPath/RF/bus_selected_win_data[168] , 
        \DataPath/RF/bus_selected_win_data[167] , 
        \DataPath/RF/bus_selected_win_data[166] , 
        \DataPath/RF/bus_selected_win_data[165] , 
        \DataPath/RF/bus_selected_win_data[164] , 
        \DataPath/RF/bus_selected_win_data[163] , 
        \DataPath/RF/bus_selected_win_data[162] , 
        \DataPath/RF/bus_selected_win_data[161] , 
        \DataPath/RF/bus_selected_win_data[160] , 
        \DataPath/RF/bus_selected_win_data[159] , 
        \DataPath/RF/bus_selected_win_data[158] , 
        \DataPath/RF/bus_selected_win_data[157] , 
        \DataPath/RF/bus_selected_win_data[156] , 
        \DataPath/RF/bus_selected_win_data[155] , 
        \DataPath/RF/bus_selected_win_data[154] , 
        \DataPath/RF/bus_selected_win_data[153] , 
        \DataPath/RF/bus_selected_win_data[152] , 
        \DataPath/RF/bus_selected_win_data[151] , 
        \DataPath/RF/bus_selected_win_data[150] , 
        \DataPath/RF/bus_selected_win_data[149] , 
        \DataPath/RF/bus_selected_win_data[148] , 
        \DataPath/RF/bus_selected_win_data[147] , 
        \DataPath/RF/bus_selected_win_data[146] , 
        \DataPath/RF/bus_selected_win_data[145] , 
        \DataPath/RF/bus_selected_win_data[144] , 
        \DataPath/RF/bus_selected_win_data[143] , 
        \DataPath/RF/bus_selected_win_data[142] , 
        \DataPath/RF/bus_selected_win_data[141] , 
        \DataPath/RF/bus_selected_win_data[140] , 
        \DataPath/RF/bus_selected_win_data[139] , 
        \DataPath/RF/bus_selected_win_data[138] , 
        \DataPath/RF/bus_selected_win_data[137] , 
        \DataPath/RF/bus_selected_win_data[136] , 
        \DataPath/RF/bus_selected_win_data[135] , 
        \DataPath/RF/bus_selected_win_data[134] , 
        \DataPath/RF/bus_selected_win_data[133] , 
        \DataPath/RF/bus_selected_win_data[132] , 
        \DataPath/RF/bus_selected_win_data[131] , 
        \DataPath/RF/bus_selected_win_data[130] , 
        \DataPath/RF/bus_selected_win_data[129] , 
        \DataPath/RF/bus_selected_win_data[128] , 
        \DataPath/RF/bus_selected_win_data[127] , 
        \DataPath/RF/bus_selected_win_data[126] , 
        \DataPath/RF/bus_selected_win_data[125] , 
        \DataPath/RF/bus_selected_win_data[124] , 
        \DataPath/RF/bus_selected_win_data[123] , 
        \DataPath/RF/bus_selected_win_data[122] , 
        \DataPath/RF/bus_selected_win_data[121] , 
        \DataPath/RF/bus_selected_win_data[120] , 
        \DataPath/RF/bus_selected_win_data[119] , 
        \DataPath/RF/bus_selected_win_data[118] , 
        \DataPath/RF/bus_selected_win_data[117] , 
        \DataPath/RF/bus_selected_win_data[116] , 
        \DataPath/RF/bus_selected_win_data[115] , 
        \DataPath/RF/bus_selected_win_data[114] , 
        \DataPath/RF/bus_selected_win_data[113] , 
        \DataPath/RF/bus_selected_win_data[112] , 
        \DataPath/RF/bus_selected_win_data[111] , 
        \DataPath/RF/bus_selected_win_data[110] , 
        \DataPath/RF/bus_selected_win_data[109] , 
        \DataPath/RF/bus_selected_win_data[108] , 
        \DataPath/RF/bus_selected_win_data[107] , 
        \DataPath/RF/bus_selected_win_data[106] , 
        \DataPath/RF/bus_selected_win_data[105] , 
        \DataPath/RF/bus_selected_win_data[104] , 
        \DataPath/RF/bus_selected_win_data[103] , 
        \DataPath/RF/bus_selected_win_data[102] , 
        \DataPath/RF/bus_selected_win_data[101] , 
        \DataPath/RF/bus_selected_win_data[100] , 
        \DataPath/RF/bus_selected_win_data[99] , 
        \DataPath/RF/bus_selected_win_data[98] , 
        \DataPath/RF/bus_selected_win_data[97] , 
        \DataPath/RF/bus_selected_win_data[96] , 
        \DataPath/RF/bus_selected_win_data[95] , 
        \DataPath/RF/bus_selected_win_data[94] , 
        \DataPath/RF/bus_selected_win_data[93] , 
        \DataPath/RF/bus_selected_win_data[92] , 
        \DataPath/RF/bus_selected_win_data[91] , 
        \DataPath/RF/bus_selected_win_data[90] , 
        \DataPath/RF/bus_selected_win_data[89] , 
        \DataPath/RF/bus_selected_win_data[88] , 
        \DataPath/RF/bus_selected_win_data[87] , 
        \DataPath/RF/bus_selected_win_data[86] , 
        \DataPath/RF/bus_selected_win_data[85] , 
        \DataPath/RF/bus_selected_win_data[84] , 
        \DataPath/RF/bus_selected_win_data[83] , 
        \DataPath/RF/bus_selected_win_data[82] , 
        \DataPath/RF/bus_selected_win_data[81] , 
        \DataPath/RF/bus_selected_win_data[80] , 
        \DataPath/RF/bus_selected_win_data[79] , 
        \DataPath/RF/bus_selected_win_data[78] , 
        \DataPath/RF/bus_selected_win_data[77] , 
        \DataPath/RF/bus_selected_win_data[76] , 
        \DataPath/RF/bus_selected_win_data[75] , 
        \DataPath/RF/bus_selected_win_data[74] , 
        \DataPath/RF/bus_selected_win_data[73] , 
        \DataPath/RF/bus_selected_win_data[72] , 
        \DataPath/RF/bus_selected_win_data[71] , 
        \DataPath/RF/bus_selected_win_data[70] , 
        \DataPath/RF/bus_selected_win_data[69] , 
        \DataPath/RF/bus_selected_win_data[68] , 
        \DataPath/RF/bus_selected_win_data[67] , 
        \DataPath/RF/bus_selected_win_data[66] , 
        \DataPath/RF/bus_selected_win_data[65] , 
        \DataPath/RF/bus_selected_win_data[64] , 
        \DataPath/RF/bus_selected_win_data[63] , 
        \DataPath/RF/bus_selected_win_data[62] , 
        \DataPath/RF/bus_selected_win_data[61] , 
        \DataPath/RF/bus_selected_win_data[60] , 
        \DataPath/RF/bus_selected_win_data[59] , 
        \DataPath/RF/bus_selected_win_data[58] , 
        \DataPath/RF/bus_selected_win_data[57] , 
        \DataPath/RF/bus_selected_win_data[56] , 
        \DataPath/RF/bus_selected_win_data[55] , 
        \DataPath/RF/bus_selected_win_data[54] , 
        \DataPath/RF/bus_selected_win_data[53] , 
        \DataPath/RF/bus_selected_win_data[52] , 
        \DataPath/RF/bus_selected_win_data[51] , 
        \DataPath/RF/bus_selected_win_data[50] , 
        \DataPath/RF/bus_selected_win_data[49] , 
        \DataPath/RF/bus_selected_win_data[48] , 
        \DataPath/RF/bus_selected_win_data[47] , 
        \DataPath/RF/bus_selected_win_data[46] , 
        \DataPath/RF/bus_selected_win_data[45] , 
        \DataPath/RF/bus_selected_win_data[44] , 
        \DataPath/RF/bus_selected_win_data[43] , 
        \DataPath/RF/bus_selected_win_data[42] , 
        \DataPath/RF/bus_selected_win_data[41] , 
        \DataPath/RF/bus_selected_win_data[40] , 
        \DataPath/RF/bus_selected_win_data[39] , 
        \DataPath/RF/bus_selected_win_data[38] , 
        \DataPath/RF/bus_selected_win_data[37] , 
        \DataPath/RF/bus_selected_win_data[36] , 
        \DataPath/RF/bus_selected_win_data[35] , 
        \DataPath/RF/bus_selected_win_data[34] , 
        \DataPath/RF/bus_selected_win_data[33] , 
        \DataPath/RF/bus_selected_win_data[32] , 
        \DataPath/RF/bus_selected_win_data[31] , 
        \DataPath/RF/bus_selected_win_data[30] , 
        \DataPath/RF/bus_selected_win_data[29] , 
        \DataPath/RF/bus_selected_win_data[28] , 
        \DataPath/RF/bus_selected_win_data[27] , 
        \DataPath/RF/bus_selected_win_data[26] , 
        \DataPath/RF/bus_selected_win_data[25] , 
        \DataPath/RF/bus_selected_win_data[24] , 
        \DataPath/RF/bus_selected_win_data[23] , 
        \DataPath/RF/bus_selected_win_data[22] , 
        \DataPath/RF/bus_selected_win_data[21] , 
        \DataPath/RF/bus_selected_win_data[20] , 
        \DataPath/RF/bus_selected_win_data[19] , 
        \DataPath/RF/bus_selected_win_data[18] , 
        \DataPath/RF/bus_selected_win_data[17] , 
        \DataPath/RF/bus_selected_win_data[16] , 
        \DataPath/RF/bus_selected_win_data[15] , 
        \DataPath/RF/bus_selected_win_data[14] , 
        \DataPath/RF/bus_selected_win_data[13] , 
        \DataPath/RF/bus_selected_win_data[12] , 
        \DataPath/RF/bus_selected_win_data[11] , 
        \DataPath/RF/bus_selected_win_data[10] , 
        \DataPath/RF/bus_selected_win_data[9] , 
        \DataPath/RF/bus_selected_win_data[8] , 
        \DataPath/RF/bus_selected_win_data[7] , 
        \DataPath/RF/bus_selected_win_data[6] , 
        \DataPath/RF/bus_selected_win_data[5] , 
        \DataPath/RF/bus_selected_win_data[4] , 
        \DataPath/RF/bus_selected_win_data[3] , 
        \DataPath/RF/bus_selected_win_data[2] , 
        \DataPath/RF/bus_selected_win_data[1] , 
        \DataPath/RF/bus_selected_win_data[0] }) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[0]  ( .D(n3230), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[0] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[1]  ( .D(n3229), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[1] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[2]  ( .D(n3228), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[2] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[3]  ( .D(n3227), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[3] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[4]  ( .D(n3226), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[4] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[5]  ( .D(n3225), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[5] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[6]  ( .D(n3224), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[6] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[7]  ( .D(n3223), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[7] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[8]  ( .D(n3222), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[8] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[9]  ( .D(n3221), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[9] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[10]  ( .D(n3220), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[10] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[11]  ( .D(n3219), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[11] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[12]  ( .D(n3218), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[12] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[13]  ( .D(n3217), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[13] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[14]  ( .D(n3216), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[14] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[15]  ( .D(n3215), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[15] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[16]  ( .D(n3214), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[16] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[17]  ( .D(n3213), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[17] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[18]  ( .D(n3212), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[18] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[19]  ( .D(n3211), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[19] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[20]  ( .D(n3210), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[20] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[21]  ( .D(n3209), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[21] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[22]  ( .D(n3208), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[22] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[23]  ( .D(n3207), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[23] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[24]  ( .D(n3206), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[24] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[25]  ( .D(n3205), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[25] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[26]  ( .D(n3204), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[26] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[27]  ( .D(n3203), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[27] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[28]  ( .D(n3202), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[28] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[29]  ( .D(n3201), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[29] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[30]  ( .D(n3200), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[30] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_data_reg[31]  ( .D(n3197), .CK(CLK), .QN(
        \DataPath/WRF_CUhw/curr_data[31] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[0]  ( .D(n7169), .CK(CLK), 
        .QN(n555) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[1]  ( .D(n7168), .CK(CLK), 
        .QN(n556) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[3]  ( .D(n7166), .CK(CLK), 
        .QN(n558) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[5]  ( .D(n7164), .CK(CLK), 
        .QN(n560) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[6]  ( .D(n7163), .CK(CLK), 
        .Q(\DECODEhw/i_tickcounter[6] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[7]  ( .D(n7162), .CK(CLK), 
        .QN(n562) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[8]  ( .D(n7161), .CK(CLK), 
        .Q(\DECODEhw/i_tickcounter[8] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[9]  ( .D(n7160), .CK(CLK), 
        .QN(n564) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[10]  ( .D(n7159), .CK(CLK), .Q(\DECODEhw/i_tickcounter[10] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[11]  ( .D(n7158), .CK(CLK), .QN(n566) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[12]  ( .D(n7157), .CK(CLK), .Q(\DECODEhw/i_tickcounter[12] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[13]  ( .D(n7156), .CK(CLK), .QN(n568) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[14]  ( .D(n7155), .CK(CLK), .Q(\DECODEhw/i_tickcounter[14] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[15]  ( .D(n7154), .CK(CLK), .QN(n570) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[16]  ( .D(n7153), .CK(CLK), .Q(\DECODEhw/i_tickcounter[16] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[17]  ( .D(n7152), .CK(CLK), .QN(n572) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[18]  ( .D(n7151), .CK(CLK), .Q(\DECODEhw/i_tickcounter[18] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[19]  ( .D(n7150), .CK(CLK), .QN(n574) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[20]  ( .D(n7149), .CK(CLK), .Q(\DECODEhw/i_tickcounter[20] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[21]  ( .D(n7148), .CK(CLK), .QN(n576) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[22]  ( .D(n7147), .CK(CLK), .Q(\DECODEhw/i_tickcounter[22] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[23]  ( .D(n7146), .CK(CLK), .QN(n578) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[24]  ( .D(n7145), .CK(CLK), .Q(\DECODEhw/i_tickcounter[24] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[25]  ( .D(n7144), .CK(CLK), .QN(n580) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[26]  ( .D(n7143), .CK(CLK), .Q(\DECODEhw/i_tickcounter[26] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[27]  ( .D(n7142), .CK(CLK), .QN(n582) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[28]  ( .D(n7141), .CK(CLK), .QN(n583) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[29]  ( .D(n3153), .CK(CLK), .QN(\DECODEhw/i_tickcounter[29] ) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[30]  ( .D(n7140), .CK(CLK), .QN(n584) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[31]  ( .D(n7170), .CK(CLK), .Q(\DECODEhw/i_tickcounter[31] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[0]  ( .D(n5783), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2048] ) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[31]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N35 ), .Q(i_RD2[31]) );
  DFF_X1 \DataPath/REG_B/Q_reg[31]  ( .D(n2743), .CK(CLK), .Q(n8189), .QN(
        \DataPath/i_PIPLIN_B[31] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[31]  ( .D(n2712), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[31] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[7]  ( .D(n2216), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[7] ) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[31]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N35 ), .Q(i_RD1[31]) );
  DFFR_X1 \IR_reg[25]  ( .D(n7127), .CK(CLK), .RN(n8460), .QN(n173) );
  DFFR_X1 \IR_reg[24]  ( .D(n7128), .CK(CLK), .RN(n8466), .QN(n174) );
  DFFR_X1 \IR_reg[23]  ( .D(n7129), .CK(CLK), .RN(n8459), .QN(n175) );
  DFFR_X1 \IR_reg[17]  ( .D(n7135), .CK(CLK), .RN(n8461), .QN(n181) );
  DFFR_X1 \IR_reg[16]  ( .D(n7136), .CK(CLK), .RN(n8465), .QN(n182) );
  DFFS_X1 \IR_reg[8]  ( .D(n2890), .CK(CLK), .SN(n8462), .Q(n8139), .QN(IR[8])
         );
  DFFS_X1 \IR_reg[10]  ( .D(n2889), .CK(CLK), .SN(n8461), .Q(n8137), .QN(
        IR[10]) );
  DFFS_X1 \IR_reg[13]  ( .D(n2886), .CK(CLK), .SN(n8460), .Q(n8136), .QN(
        IR[13]) );
  DFF_X1 \DataPath/WRB1/Q_reg[0]  ( .D(n2870), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB1[0] ) );
  DFF_X1 \DataPath/WRB2/Q_reg[0]  ( .D(n2779), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB2[0] ) );
  DFF_X1 \DataPath/WRB3/Q_reg[0]  ( .D(n359), .CK(CLK), .Q(i_ADD_WB[0]), .QN(
        n537) );
  DFF_X1 \CU_I/CW_EX_reg[MEM_EN]  ( .D(n367), .CK(CLK), .QN(n8199) );
  DFF_X1 \CU_I/aluOpcode1_reg[0]  ( .D(n7090), .CK(CLK), .Q(i_ALU_OP[0]), .QN(
        n8182) );
  DFF_X1 \CU_I/setcmp_1_reg[1]  ( .D(n7084), .CK(CLK), .Q(\i_SEL_LGET[1] ), 
        .QN(n8198) );
  DFF_X1 \CU_I/i_FILL_delay_reg  ( .D(\CU_I/N314 ), .CK(CLK), .Q(
        \CU_I/i_FILL_delay ) );
  DFF_X1 \CU_I/i_SPILL_delay_reg  ( .D(\CU_I/N315 ), .CK(CLK), .QN(n8167) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_state_reg[0]  ( .D(n7064), .CK(CLK), 
        .Q(\DataPath/RF/PUSH_ADDRGEN/curr_state[0] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[1]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N47 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[1] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[2]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N48 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[2] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[3]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N49 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[3] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[4]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N50 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[4] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[5]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N51 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[5] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[6]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N52 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[6] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[7]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N53 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[7] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[8]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N54 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[8] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[9]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N55 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[9] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[10]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N56 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[10] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[11]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N57 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[11] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[12]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N58 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[12] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[13]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N59 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[13] ) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[14]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N60 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[14] ), .QN(n8104) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_state_reg[1]  ( .D(n90), .CK(CLK), 
        .QN(n849) );
  DFF_X1 \DataPath/WRF_CUhw/curr_state_reg[1]  ( .D(\DataPath/WRF_CUhw/N145 ), 
        .CK(CLK), .QN(n471) );
  DFF_X1 \DataPath/WRF_CUhw/curr_state_reg[0]  ( .D(n99), .CK(CLK), .Q(n8129), 
        .QN(n470) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_state_reg[1]  ( .D(n7057), .CK(CLK), 
        .Q(\DataPath/RF/POP_ADDRGEN/curr_state[1] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[1]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N47 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[1] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[2]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N48 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[2] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[3]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N49 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[3] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[4]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N50 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[4] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[5]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N51 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[5] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[6]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N52 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[6] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[7]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N53 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[7] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[9]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N55 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[9] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[10]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N56 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[10] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[11]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N57 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[11] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[12]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N58 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[12] ) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[14]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N60 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[14] ) );
  DLL_X1 \CU_I/CW_ID_reg[RF_RD1_EN]  ( .D(\CU_I/CW[RF_RD1_EN] ), .GN(n2872), 
        .Q(i_RF1) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[0]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N4 ), .Q(i_RD1[0]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[1]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N5 ), .Q(i_RD1[1]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[2]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N6 ), .Q(i_RD1[2]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[3]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N7 ), .Q(i_RD1[3]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[4]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N8 ), .Q(i_RD1[4]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[5]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N9 ), .Q(i_RD1[5]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[6]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N10 ), .Q(i_RD1[6]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[7]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N11 ), .Q(i_RD1[7]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[8]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N12 ), .Q(i_RD1[8]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[9]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N13 ), .Q(i_RD1[9]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[10]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N14 ), .Q(i_RD1[10]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[11]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N15 ), .Q(i_RD1[11]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[12]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N16 ), .Q(i_RD1[12]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[13]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N17 ), .Q(i_RD1[13]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[14]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N18 ), .Q(i_RD1[14]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[15]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N19 ), .Q(i_RD1[15]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[16]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N20 ), .Q(i_RD1[16]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[17]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N21 ), .Q(i_RD1[17]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[18]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N22 ), .Q(i_RD1[18]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[19]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N23 ), .Q(i_RD1[19]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[20]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N24 ), .Q(i_RD1[20]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[21]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N25 ), .Q(i_RD1[21]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[22]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N26 ), .Q(i_RD1[22]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[23]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N27 ), .Q(i_RD1[23]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[24]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N28 ), .Q(i_RD1[24]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[25]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N29 ), .Q(i_RD1[25]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[26]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N30 ), .Q(i_RD1[26]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[27]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N31 ), .Q(i_RD1[27]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[28]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N32 ), .Q(i_RD1[28]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[29]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N33 ), .Q(i_RD1[29]) );
  DLH_X1 \DataPath/RF/RDPORT0_OUTLATCH/q_mem_reg[30]  ( .G(
        \DataPath/RF/RDPORT0_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT0_OUTLATCH/N34 ), .Q(i_RD1[30]) );
  DLL_X1 \CU_I/CW_ID_reg[RF_RD2_EN]  ( .D(\CU_I/CW[RF_RD2_EN] ), .GN(n2872), 
        .Q(i_RF2) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[0]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N4 ), .Q(i_RD2[0]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[1]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N5 ), .Q(i_RD2[1]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[2]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N6 ), .Q(i_RD2[2]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[3]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N7 ), .Q(i_RD2[3]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[4]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N8 ), .Q(i_RD2[4]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[5]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N9 ), .Q(i_RD2[5]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[6]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N10 ), .Q(i_RD2[6]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[7]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N11 ), .Q(i_RD2[7]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[8]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N12 ), .Q(i_RD2[8]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[9]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N13 ), .Q(i_RD2[9]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[10]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N14 ), .Q(i_RD2[10]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[11]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N15 ), .Q(i_RD2[11]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[12]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N16 ), .Q(i_RD2[12]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[13]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N17 ), .Q(i_RD2[13]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[14]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N18 ), .Q(i_RD2[14]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[15]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N19 ), .Q(i_RD2[15]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[16]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N20 ), .Q(i_RD2[16]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[17]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N21 ), .Q(i_RD2[17]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[18]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N22 ), .Q(i_RD2[18]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[19]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N23 ), .Q(i_RD2[19]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[20]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N24 ), .Q(i_RD2[20]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[21]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N25 ), .Q(i_RD2[21]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[22]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N26 ), .Q(i_RD2[22]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[23]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N27 ), .Q(i_RD2[23]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[24]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N28 ), .Q(i_RD2[24]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[25]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N29 ), .Q(i_RD2[25]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[26]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N30 ), .Q(i_RD2[26]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[27]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N31 ), .Q(i_RD2[27]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[28]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N32 ), .Q(i_RD2[28]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[29]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N33 ), .Q(i_RD2[29]) );
  DLH_X1 \DataPath/RF/RDPORT1_OUTLATCH/q_mem_reg[30]  ( .G(
        \DataPath/RF/RDPORT1_OUTLATCH/N3 ), .D(
        \DataPath/RF/RDPORT1_OUTLATCH/N34 ), .Q(i_RD2[30]) );
  DLL_X1 \CU_I/CW_ID_reg[SEL_CMPB]  ( .D(\CU_I/CW[SEL_CMPB] ), .GN(n2872), .Q(
        i_SEL_CMPB) );
  DLL_X1 \CU_I/CW_ID_reg[UNSIGNED_ID]  ( .D(\CU_I/CW[UNSIGNED_ID] ), .GN(n2872), .Q(\CU_I/CW_ID[UNSIGNED_ID] ) );
  DFF_X1 \CU_I/unsigned_1_reg  ( .D(n7079), .CK(CLK), .QN(n218) );
  DFF_X1 \CU_I/unsigned_2_reg  ( .D(n7078), .CK(CLK), .QN(n217) );
  DLL_X1 \CU_I/CW_ID_reg[NPC_SEL]  ( .D(\CU_I/CW[NPC_SEL] ), .GN(n2872), .Q(
        i_NPC_SEL) );
  DFFR_X1 \PC_reg[0]  ( .D(n7056), .CK(CLK), .RN(n8467), .Q(IRAM_ADDRESS[0])
         );
  DFFR_X1 \PC_reg[6]  ( .D(n7050), .CK(CLK), .RN(n8464), .Q(IRAM_ADDRESS[6])
         );
  DFFR_X1 \PC_reg[10]  ( .D(n7046), .CK(CLK), .RN(n8463), .Q(IRAM_ADDRESS[10])
         );
  DFFR_X1 \PC_reg[16]  ( .D(n7040), .CK(CLK), .RN(n8457), .Q(IRAM_ADDRESS[16])
         );
  DFFR_X1 \PC_reg[18]  ( .D(n7038), .CK(CLK), .RN(n8469), .Q(IRAM_ADDRESS[18])
         );
  DFFR_X1 \PC_reg[21]  ( .D(n7035), .CK(CLK), .RN(n8468), .Q(IRAM_ADDRESS[21])
         );
  DFFR_X1 \PC_reg[22]  ( .D(n7034), .CK(CLK), .RN(n8469), .Q(IRAM_ADDRESS[22])
         );
  DFFR_X1 \PC_reg[23]  ( .D(n7033), .CK(CLK), .RN(n8464), .Q(IRAM_ADDRESS[23])
         );
  DFFR_X1 \PC_reg[24]  ( .D(n7032), .CK(CLK), .RN(n8460), .Q(IRAM_ADDRESS[24])
         );
  DFFR_X1 \PC_reg[25]  ( .D(n7031), .CK(CLK), .RN(n8465), .Q(IRAM_ADDRESS[25])
         );
  DFFR_X1 \PC_reg[29]  ( .D(n7027), .CK(CLK), .RN(n8463), .Q(IRAM_ADDRESS[29])
         );
  DLL_X1 \CU_I/CW_ID_reg[HAZARD_TABLE_WR1]  ( .D(n10296), .GN(n2872), .Q(n466)
         );
  DLL_X1 \CU_I/CW_ID_reg[MUXA_SEL]  ( .D(n10291), .GN(n2872), .Q(
        \CU_I/CW_ID[MUXA_SEL] ) );
  DFF_X1 \CU_I/CW_EX_reg[MUXA_SEL]  ( .D(n7080), .CK(CLK), .Q(n8444), .QN(n465) );
  DLL_X1 \CU_I/CW_ID_reg[MUXB_SEL]  ( .D(\CU_I/CW[MUXB_SEL] ), .GN(n2872), .Q(
        \CU_I/CW_ID[MUXB_SEL] ) );
  DFF_X1 \CU_I/CW_EX_reg[MUXB_SEL]  ( .D(n7081), .CK(CLK), .Q(i_S2), .QN(n8087) );
  DLL_X1 \CU_I/CW_ID_reg[DRAM_WE]  ( .D(\CU_I/CW[DRAM_WE] ), .GN(n2872), .Q(
        \CU_I/CW_ID[DRAM_WE] ) );
  DFF_X1 \CU_I/CW_EX_reg[DRAM_WE]  ( .D(n366), .CK(CLK), .QN(n8203) );
  DFF_X1 \CU_I/CW_MEM_reg[DRAM_WE]  ( .D(n7121), .CK(CLK), .QN(
        DRAM_READNOTWRITE) );
  DLL_X1 \CU_I/CW_ID_reg[DRAM_RE]  ( .D(\CU_I/CW[WB_MUX_SEL] ), .GN(n2872), 
        .Q(\CU_I/CW_ID[DRAM_RE] ) );
  DFF_X1 \CU_I/CW_EX_reg[DRAM_RE]  ( .D(n370), .CK(CLK), .QN(n8200) );
  DLL_X1 \CU_I/CW_ID_reg[DATA_SIZE][1]  ( .D(\CU_I/CW[DATA_SIZE][1] ), .GN(
        n2872), .Q(\CU_I/CW_ID[DATA_SIZE][1] ) );
  DFF_X1 \CU_I/CW_EX_reg[DATA_SIZE][1]  ( .D(n369), .CK(CLK), .QN(n8201) );
  DFF_X1 \CU_I/CW_MEM_reg[DATA_SIZE][1]  ( .D(n7092), .CK(CLK), .Q(
        DATA_SIZE[1]), .QN(n381) );
  DLL_X1 \CU_I/CW_ID_reg[DATA_SIZE][0]  ( .D(\CU_I/CW[DATA_SIZE][0] ), .GN(
        n2872), .Q(\CU_I/CW_ID[DATA_SIZE][0] ) );
  DFF_X1 \CU_I/CW_EX_reg[DATA_SIZE][0]  ( .D(n368), .CK(CLK), .QN(n8202) );
  DFF_X1 \CU_I/CW_MEM_reg[DATA_SIZE][0]  ( .D(n7093), .CK(CLK), .Q(
        DATA_SIZE[0]), .QN(n380) );
  DLL_X1 \CU_I/CW_ID_reg[WB_MUX_SEL]  ( .D(\CU_I/CW[WB_MUX_SEL] ), .GN(n2872), 
        .Q(\CU_I/CW_ID[WB_MUX_SEL] ) );
  DFF_X1 \CU_I/CW_EX_reg[WB_MUX_SEL]  ( .D(n2852), .CK(CLK), .QN(
        \CU_I/CW_EX[WB_MUX_SEL] ) );
  DFF_X1 \CU_I/CW_MEM_reg[WB_MUX_SEL]  ( .D(n2846), .CK(CLK), .QN(
        \CU_I/CW_MEM[WB_MUX_SEL] ) );
  DFF_X1 \CU_I/CW_WB_reg[WB_MUX_SEL]  ( .D(\CU_I/N302 ), .CK(CLK), .Q(i_S3) );
  DLL_X1 \CU_I/CW_ID_reg[WB_EN]  ( .D(\CU_I/CW_IF[WB_EN] ), .GN(n2872), .Q(
        \CU_I/CW_ID[WB_EN] ) );
  DFF_X1 \CU_I/CW_EX_reg[WB_EN]  ( .D(n2853), .CK(CLK), .QN(
        \CU_I/CW_EX[WB_EN] ) );
  DFF_X1 \CU_I/CW_MEM_reg[WB_EN]  ( .D(n2847), .CK(CLK), .QN(
        \CU_I/CW_MEM[WB_EN] ) );
  DFF_X1 \CU_I/CW_WB_reg[WB_EN]  ( .D(\CU_I/N301 ), .CK(CLK), .Q(i_WF), .QN(
        n8192) );
  DLL_X1 \CU_I/CW_ID_reg[EX_EN]  ( .D(n10274), .GN(n2872), .Q(
        \CU_I/CW_ID[EX_EN] ) );
  DFF_X1 \CU_I/CW_EX_reg[EX_EN]  ( .D(n2780), .CK(CLK), .Q(n8191), .QN(
        \CU_I/CW_EX[EX_EN] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[20]  ( .D(n7014), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[20] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[15]  ( .D(n7015), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[15] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[13]  ( .D(n7017), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[13] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[12]  ( .D(n7018), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[12] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[10]  ( .D(n7019), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[10] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[8]  ( .D(n7020), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[8] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[6]  ( .D(n7021), .CK(CLK), .QN(n497) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[4]  ( .D(n7022), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[4] ), .QN(n8211) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[3]  ( .D(n7023), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[3] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[0]  ( .D(n7024), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[0] ), .QN(n8221) );
  DFF_X1 \DataPath/REG_B/Q_reg[14]  ( .D(n7071), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_B[14] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[14]  ( .D(n2729), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[14] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[13]  ( .D(n7072), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_B[13] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[13]  ( .D(n2730), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[13] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[8]  ( .D(n7073), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_B[8] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[8]  ( .D(n2735), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[8] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[6]  ( .D(n7070), .CK(CLK), .Q(
        \DataPath/i_REG_ME_DATA_DATAMEM[6] ), .QN(n8223) );
  DFF_X1 \DataPath/REG_ME/Q_reg[4]  ( .D(n2738), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[4] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[3]  ( .D(n7076), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_B[3] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[3]  ( .D(n2739), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[3] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[0]  ( .D(n7077), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_B[0] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[0]  ( .D(n2742), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[0] ) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[2]  ( .D(n7117), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[2] ) );
  DFF_X1 \DataPath/REG_CMP/Q_reg[1]  ( .D(n7120), .CK(CLK), .Q(n8106), .QN(
        n506) );
  DFF_X1 \DataPath/REG_A/Q_reg[20]  ( .D(n6723), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_A[20] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[14]  ( .D(n6724), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_A[14] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[13]  ( .D(n6725), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_A[13] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[8]  ( .D(n6726), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_A[8] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[3]  ( .D(n6727), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_A[3] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[1]  ( .D(n6728), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_A[1] ) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[9]  ( .D(n7111), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[9] ), .QN(n8220) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[7]  ( .D(n7112), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[7] ), .QN(n8219) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[6]  ( .D(n7113), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[6] ), .QN(n8218) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[5]  ( .D(n7114), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[5] ), .QN(n8217) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[4]  ( .D(n7115), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[4] ), .QN(n8216) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[3]  ( .D(n7116), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[3] ), .QN(n8215) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[1]  ( .D(n7118), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[1] ), .QN(n8214) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[0]  ( .D(n7119), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN1[0] ), .QN(n8213) );
  DFF_X1 \DataPath/REG_A/Q_reg[0]  ( .D(n3256), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[0] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[2]  ( .D(n3255), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[2] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[4]  ( .D(n3254), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[4] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[5]  ( .D(n3253), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[5] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[6]  ( .D(n3252), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[6] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[7]  ( .D(n3251), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[7] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[9]  ( .D(n3250), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[9] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[10]  ( .D(n3249), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[10] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[11]  ( .D(n3248), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[11] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[12]  ( .D(n3247), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[12] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[15]  ( .D(n3246), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[15] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[16]  ( .D(n3245), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[16] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[17]  ( .D(n3244), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[17] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[18]  ( .D(n3243), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[18] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[19]  ( .D(n3242), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[19] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[21]  ( .D(n3241), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[21] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[22]  ( .D(n3240), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[22] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[23]  ( .D(n3239), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[23] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[24]  ( .D(n3238), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[24] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[25]  ( .D(n3237), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[25] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[26]  ( .D(n3236), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[26] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[27]  ( .D(n3235), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[27] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[28]  ( .D(n3234), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[28] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[29]  ( .D(n3233), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[29] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[30]  ( .D(n3232), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[30] ) );
  DFF_X1 \DataPath/REG_A/Q_reg[31]  ( .D(n3231), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_A[31] ) );
  DFF_X1 \DataPath/WRB1/Q_reg[1]  ( .D(n2869), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB1[1] ) );
  DFF_X1 \DataPath/WRB2/Q_reg[1]  ( .D(n2778), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB2[1] ) );
  DFF_X1 \DataPath/WRB3/Q_reg[1]  ( .D(n360), .CK(CLK), .Q(i_ADD_WB[1]), .QN(
        n8170) );
  DFF_X1 \DataPath/WRB1/Q_reg[2]  ( .D(n2868), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB1[2] ) );
  DFF_X1 \DataPath/WRB2/Q_reg[2]  ( .D(n2777), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB2[2] ) );
  DFF_X1 \DataPath/WRB3/Q_reg[2]  ( .D(n361), .CK(CLK), .Q(i_ADD_WB[2]), .QN(
        n539) );
  DFF_X1 \DataPath/WRB1/Q_reg[3]  ( .D(n2867), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB1[3] ) );
  DFF_X1 \DataPath/WRB2/Q_reg[3]  ( .D(n2776), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB2[3] ) );
  DFF_X1 \DataPath/WRB3/Q_reg[3]  ( .D(n362), .CK(CLK), .Q(i_ADD_WB[3]) );
  DFF_X1 \DataPath/WRB1/Q_reg[4]  ( .D(n2866), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB1[4] ) );
  DFF_X1 \DataPath/WRB2/Q_reg[4]  ( .D(n2775), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_WRB2[4] ) );
  DFF_X1 \DataPath/WRB3/Q_reg[4]  ( .D(n363), .CK(CLK), .Q(i_ADD_WB[4]), .QN(
        n8102) );
  DFF_X1 \DataPath/REG_CMP/Q_reg[0]  ( .D(n102), .CK(CLK), .Q(
        \DataPath/i_LGET[0] ), .QN(n8197) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[8]  ( .D(n2861), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN1[8] ) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[10]  ( .D(n2859), .CK(CLK), .Q(n8162), .QN(
        \DataPath/i_PIPLIN_IN1[10] ) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[13]  ( .D(n2856), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN1[13] ) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[14]  ( .D(n2855), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN1[14] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[1]  ( .D(n2767), .CK(CLK), .Q(n7711), .QN(
        \DataPath/i_PIPLIN_B[1] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[1]  ( .D(n2741), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[1] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[2]  ( .D(n2766), .CK(CLK), .Q(n8141), .QN(
        \DataPath/i_PIPLIN_B[2] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[2]  ( .D(n2740), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[2] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[5]  ( .D(n2765), .CK(CLK), .Q(n8142), .QN(
        \DataPath/i_PIPLIN_B[5] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[5]  ( .D(n2737), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[5] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[7]  ( .D(n2764), .CK(CLK), .Q(n8143), .QN(
        \DataPath/i_PIPLIN_B[7] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[7]  ( .D(n2736), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[7] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[9]  ( .D(n2763), .CK(CLK), .Q(n8144), .QN(
        \DataPath/i_PIPLIN_B[9] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[9]  ( .D(n2734), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[9] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[10]  ( .D(n2762), .CK(CLK), .Q(n8146), .QN(
        \DataPath/i_PIPLIN_B[10] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[10]  ( .D(n2733), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[10] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[11]  ( .D(n2761), .CK(CLK), .Q(n8145), .QN(
        \DataPath/i_PIPLIN_B[11] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[11]  ( .D(n2732), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[11] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[12]  ( .D(n2760), .CK(CLK), .Q(n8147), .QN(
        \DataPath/i_PIPLIN_B[12] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[12]  ( .D(n2731), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[12] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[15]  ( .D(n2759), .CK(CLK), .Q(n8148), .QN(
        \DataPath/i_PIPLIN_B[15] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[15]  ( .D(n2728), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[15] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[16]  ( .D(n2758), .CK(CLK), .Q(n8150), .QN(
        \DataPath/i_PIPLIN_B[16] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[16]  ( .D(n2727), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[16] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[17]  ( .D(n2757), .CK(CLK), .Q(n8149), .QN(
        \DataPath/i_PIPLIN_B[17] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[17]  ( .D(n2726), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[17] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[18]  ( .D(n2756), .CK(CLK), .Q(n8152), .QN(
        \DataPath/i_PIPLIN_B[18] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[18]  ( .D(n2725), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[18] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[19]  ( .D(n2755), .CK(CLK), .Q(n8151), .QN(
        \DataPath/i_PIPLIN_B[19] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[19]  ( .D(n2724), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[19] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[20]  ( .D(n2754), .CK(CLK), .Q(n8153), .QN(
        \DataPath/i_PIPLIN_B[20] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[20]  ( .D(n2723), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[20] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[21]  ( .D(n2753), .CK(CLK), .Q(n8131), .QN(
        \DataPath/i_PIPLIN_B[21] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[21]  ( .D(n2722), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[21] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[22]  ( .D(n2752), .CK(CLK), .Q(n8155), .QN(
        \DataPath/i_PIPLIN_B[22] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[22]  ( .D(n2721), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[22] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[23]  ( .D(n2751), .CK(CLK), .Q(n8154), .QN(
        \DataPath/i_PIPLIN_B[23] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[23]  ( .D(n2720), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[23] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[24]  ( .D(n2750), .CK(CLK), .Q(n8157), .QN(
        \DataPath/i_PIPLIN_B[24] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[24]  ( .D(n2719), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[24] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[25]  ( .D(n2749), .CK(CLK), .Q(n8156), .QN(
        \DataPath/i_PIPLIN_B[25] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[25]  ( .D(n2718), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[25] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[26]  ( .D(n2748), .CK(CLK), .Q(n8186), .QN(
        \DataPath/i_PIPLIN_B[26] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[26]  ( .D(n2717), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[26] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[27]  ( .D(n2747), .CK(CLK), .Q(n8132), .QN(
        \DataPath/i_PIPLIN_B[27] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[27]  ( .D(n2716), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[27] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[28]  ( .D(n2746), .CK(CLK), .Q(n8188), .QN(
        \DataPath/i_PIPLIN_B[28] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[28]  ( .D(n2715), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[28] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[29]  ( .D(n2745), .CK(CLK), .Q(n8187), .QN(
        \DataPath/i_PIPLIN_B[29] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[29]  ( .D(n2714), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[29] ) );
  DFF_X1 \DataPath/REG_B/Q_reg[30]  ( .D(n2744), .CK(CLK), .Q(n8190), .QN(
        \DataPath/i_PIPLIN_B[30] ) );
  DFF_X1 \DataPath/REG_ME/Q_reg[30]  ( .D(n2713), .CK(CLK), .QN(
        \DataPath/i_REG_ME_DATA_DATAMEM[30] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[1]  ( .D(n2398), .CK(CLK), .Q(n7710), .QN(
        \DataPath/i_PIPLIN_IN2[1] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[2]  ( .D(n2396), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[2] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[5]  ( .D(n2392), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[5] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[7]  ( .D(n2389), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[7] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[9]  ( .D(n2386), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[9] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[11]  ( .D(n2383), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[11] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[16]  ( .D(n2377), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[16] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[17]  ( .D(n2375), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[17] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[18]  ( .D(n2373), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[18] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[19]  ( .D(n2371), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[19] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[21]  ( .D(n2366), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[21] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[22]  ( .D(n2364), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[22] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[23]  ( .D(n2362), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[23] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[24]  ( .D(n2360), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[24] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[25]  ( .D(n2358), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[25] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[26]  ( .D(n2356), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[26] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[27]  ( .D(n2354), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[27] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[28]  ( .D(n2352), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[28] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[29]  ( .D(n2350), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[29] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[30]  ( .D(n2348), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[30] ) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[31]  ( .D(n2346), .CK(CLK), .QN(
        \DataPath/i_PIPLIN_IN2[31] ) );
  DFF_X1 \CU_I/setcmp_1_reg[0]  ( .D(n7085), .CK(CLK), .QN(n222) );
  DFF_X1 \CU_I/setcmp_1_reg[2]  ( .D(n7083), .CK(CLK), .QN(n223) );
  DFF_X1 \CU_I/aluOpcode1_reg[4]  ( .D(n7086), .CK(CLK), .Q(i_ALU_OP[4]), .QN(
        n8085) );
  DFF_X1 \CU_I/aluOpcode1_reg[3]  ( .D(n7087), .CK(CLK), .Q(i_ALU_OP[3]), .QN(
        n8095) );
  DFF_X1 \CU_I/aluOpcode1_reg[1]  ( .D(n7089), .CK(CLK), .Q(i_ALU_OP[1]), .QN(
        n8174) );
  DFF_X1 \CU_I/sel_alu_setcmp_1_reg  ( .D(n7082), .CK(CLK), .Q(
        i_SEL_ALU_SETCMP), .QN(n8105) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[7]  ( .D(n2011), .CK(CLK), .QN(
        DRAM_ADDRESS[7]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[7]  ( .D(n1156), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[7] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[3]  ( .D(n2133), .CK(CLK), .QN(
        DRAM_ADDRESS[3]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[3]  ( .D(n1160), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[3] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[2]  ( .D(n2165), .CK(CLK), .QN(
        DRAM_ADDRESS[2]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[2]  ( .D(n1161), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[2] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[17]  ( .D(n6999), .CK(CLK), .Q(
        DRAM_ADDRESS[17]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[17]  ( .D(n1146), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[17] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[13]  ( .D(n7003), .CK(CLK), .Q(
        DRAM_ADDRESS[13]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[13]  ( .D(n1150), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[13] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[9]  ( .D(n7007), .CK(CLK), .Q(
        DRAM_ADDRESS[9]), .QN(n8206) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[9]  ( .D(n1154), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[9] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[5]  ( .D(n7010), .CK(CLK), .Q(
        DRAM_ADDRESS[5]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[5]  ( .D(n1158), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[5] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[1]  ( .D(n7012), .CK(CLK), .Q(n8168), 
        .QN(n508) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[1]  ( .D(n1162), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[1] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[23]  ( .D(n2200), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[23] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[31]  ( .D(n2192), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[31] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[15]  ( .D(n2208), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[15] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[21]  ( .D(n6995), .CK(CLK), .Q(
        DRAM_ADDRESS[21]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[21]  ( .D(n1142), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[21] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[25]  ( .D(n6991), .CK(CLK), .Q(
        DRAM_ADDRESS[25]), .QN(n8222) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[25]  ( .D(n1138), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[25] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[29]  ( .D(n6987), .CK(CLK), .Q(
        DRAM_ADDRESS[29]) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[29]  ( .D(n1134), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[29] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[4]  ( .D(n7011), .CK(CLK), .Q(
        DRAM_ADDRESS[4]), .QN(n509) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[4]  ( .D(n1159), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[4] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[6]  ( .D(n7009), .CK(CLK), .Q(
        DRAM_ADDRESS[6]), .QN(n510) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[6]  ( .D(n1157), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[6] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[8]  ( .D(n7008), .CK(CLK), .Q(
        DRAM_ADDRESS[8]), .QN(n511) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[8]  ( .D(n1155), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[8] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[10]  ( .D(n7006), .CK(CLK), .Q(
        DRAM_ADDRESS[10]), .QN(n512) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[10]  ( .D(n1153), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[10] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[11]  ( .D(n7005), .CK(CLK), .Q(
        DRAM_ADDRESS[11]), .QN(n513) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[11]  ( .D(n1152), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[11] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[12]  ( .D(n7004), .CK(CLK), .Q(
        DRAM_ADDRESS[12]), .QN(n514) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[12]  ( .D(n1151), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[12] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[14]  ( .D(n7002), .CK(CLK), .Q(
        DRAM_ADDRESS[14]), .QN(n515) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[14]  ( .D(n1149), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[14] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[15]  ( .D(n7001), .CK(CLK), .Q(
        DRAM_ADDRESS[15]), .QN(n516) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[15]  ( .D(n1148), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[15] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[15]  ( .D(n6777), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[47] ), .QN(n625) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[15]  ( .D(n6809), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[79] ), .QN(n657) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[15]  ( .D(n6841), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[111] ), .QN(n689) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[15]  ( .D(n6873), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[143] ), .QN(n721) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[15]  ( .D(n6905), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[175] ), .QN(n753) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[15]  ( .D(n6937), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[207] ), .QN(n785) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[15]  ( .D(n6969), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[239] ), .QN(n817) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[15]  ( .D(n3337), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[15] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[15]  ( .D(n3392), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[47] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[15]  ( .D(n3430), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[79] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[15]  ( .D(n3468), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[111] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[15]  ( .D(n3506), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[143] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[15]  ( .D(n3544), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[175] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[15]  ( .D(n3582), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[207] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[15]  ( .D(n3620), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[239] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[15]  ( .D(n3658), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[271] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[15]  ( .D(n3695), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[303] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[15]  ( .D(n3732), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[335] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[15]  ( .D(n3769), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[367] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[15]  ( .D(n3804), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[399] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[15]  ( .D(n3839), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[431] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[15]  ( .D(n3874), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[463] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[15]  ( .D(n3925), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[495] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[15]  ( .D(n3993), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[527] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[15]  ( .D(n4045), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[559] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[15]  ( .D(n4080), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[591] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[15]  ( .D(n4115), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[623] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[15]  ( .D(n4150), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[655] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[15]  ( .D(n4185), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[687] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[15]  ( .D(n4220), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[719] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[15]  ( .D(n4255), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[751] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[15]  ( .D(n4290), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[783] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[15]  ( .D(n4325), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[815] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[15]  ( .D(n4360), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[847] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[15]  ( .D(n4395), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[879] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[15]  ( .D(n4430), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[911] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[15]  ( .D(n4465), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[943] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[15]  ( .D(n4500), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[975] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[15]  ( .D(n4535), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1007] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[15]  ( .D(n4586), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1039] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[15]  ( .D(n4638), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1071] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[15]  ( .D(n4673), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1103] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[15]  ( .D(n4708), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1135] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[15]  ( .D(n4743), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1167] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[15]  ( .D(n4778), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1199] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[15]  ( .D(n4813), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1231] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[15]  ( .D(n4848), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1263] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[15]  ( .D(n4883), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1295] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[15]  ( .D(n4918), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1327] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[15]  ( .D(n4953), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1359] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[15]  ( .D(n4988), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1391] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[15]  ( .D(n5023), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1423] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[15]  ( .D(n5058), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1455] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[15]  ( .D(n5093), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1487] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[15]  ( .D(n5128), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1519] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[15]  ( .D(n5179), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1551] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[15]  ( .D(n5230), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1583] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[15]  ( .D(n5266), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1615] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[15]  ( .D(n5301), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1647] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[15]  ( .D(n5336), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1679] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[15]  ( .D(n5371), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1711] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[15]  ( .D(n5406), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1743] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[15]  ( .D(n5441), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1775] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[15]  ( .D(n5476), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1807] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[15]  ( .D(n5511), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1839] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[15]  ( .D(n5546), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1871] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[15]  ( .D(n5581), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1903] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[15]  ( .D(n5620), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1935] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[15]  ( .D(n5657), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1967] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[15]  ( .D(n5694), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1999] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[15]  ( .D(n5731), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2031] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[15]  ( .D(n898), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2383] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[15]  ( .D(n962), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2415] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[15]  ( .D(n1000), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2447] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[15]  ( .D(n1037), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2479] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[15]  ( .D(n1074), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2511] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[15]  ( .D(n1111), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2543] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[15]  ( .D(n5768), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2063] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[15]  ( .D(n5807), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2095] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[15]  ( .D(n5843), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2127] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[15]  ( .D(n5879), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2159] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[15]  ( .D(n5915), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2191] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[15]  ( .D(n5951), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2223] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[15]  ( .D(n5987), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2255] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[15]  ( .D(n6023), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2287] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[15]  ( .D(n6060), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2319] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[15]  ( .D(n6096), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2351] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[16]  ( .D(n7000), .CK(CLK), .Q(
        DRAM_ADDRESS[16]), .QN(n517) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[16]  ( .D(n1147), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[16] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[18]  ( .D(n6998), .CK(CLK), .Q(
        DRAM_ADDRESS[18]), .QN(n518) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[18]  ( .D(n1145), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[18] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[19]  ( .D(n6997), .CK(CLK), .Q(
        DRAM_ADDRESS[19]), .QN(n519) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[19]  ( .D(n1144), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[19] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[20]  ( .D(n6996), .CK(CLK), .Q(
        DRAM_ADDRESS[20]), .QN(n520) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[20]  ( .D(n1143), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[20] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[22]  ( .D(n6994), .CK(CLK), .Q(
        DRAM_ADDRESS[22]), .QN(n521) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[22]  ( .D(n1141), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[22] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[23]  ( .D(n6993), .CK(CLK), .Q(
        DRAM_ADDRESS[23]), .QN(n522) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[23]  ( .D(n1140), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[23] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[23]  ( .D(n3321), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[23] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[23]  ( .D(n3384), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[55] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[23]  ( .D(n3422), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[87] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[23]  ( .D(n3460), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[119] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[23]  ( .D(n3498), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[151] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[23]  ( .D(n3536), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[183] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[23]  ( .D(n3574), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[215] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[23]  ( .D(n3612), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[247] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[23]  ( .D(n3650), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[279] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[23]  ( .D(n3687), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[311] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[23]  ( .D(n3724), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[343] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[23]  ( .D(n3761), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[375] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[23]  ( .D(n3796), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[407] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[23]  ( .D(n3831), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[439] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[23]  ( .D(n3866), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[471] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[23]  ( .D(n3909), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[503] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[23]  ( .D(n3977), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[535] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[23]  ( .D(n4037), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[567] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[23]  ( .D(n4072), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[599] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[23]  ( .D(n4107), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[631] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[23]  ( .D(n4142), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[663] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[23]  ( .D(n4177), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[695] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[23]  ( .D(n4212), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[727] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[23]  ( .D(n4247), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[759] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[23]  ( .D(n4282), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[791] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[23]  ( .D(n4317), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[823] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[23]  ( .D(n4352), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[855] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[23]  ( .D(n4387), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[887] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[23]  ( .D(n4422), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[919] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[23]  ( .D(n4457), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[951] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[23]  ( .D(n4492), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[983] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[23]  ( .D(n4527), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1015] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[23]  ( .D(n4570), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1047] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[23]  ( .D(n4630), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1079] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[23]  ( .D(n4665), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1111] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[23]  ( .D(n4700), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1143] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[23]  ( .D(n4735), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1175] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[23]  ( .D(n4770), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1207] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[23]  ( .D(n4805), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1239] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[23]  ( .D(n4840), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1271] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[23]  ( .D(n4875), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1303] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[23]  ( .D(n4910), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1335] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[23]  ( .D(n4945), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1367] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[23]  ( .D(n4980), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1399] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[23]  ( .D(n5015), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1431] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[23]  ( .D(n5050), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1463] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[23]  ( .D(n5085), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1495] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[23]  ( .D(n5120), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1527] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[23]  ( .D(n5163), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1559] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[23]  ( .D(n5222), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1591] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[23]  ( .D(n5258), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1623] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[23]  ( .D(n5293), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1655] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[23]  ( .D(n5328), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1687] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[23]  ( .D(n5363), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1719] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[23]  ( .D(n5398), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1751] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[23]  ( .D(n5433), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1783] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[23]  ( .D(n5468), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1815] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[23]  ( .D(n5503), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1847] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[23]  ( .D(n5538), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1879] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[23]  ( .D(n5573), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1911] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[23]  ( .D(n5612), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1943] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[23]  ( .D(n5649), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1975] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[23]  ( .D(n5686), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2007] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[23]  ( .D(n5723), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2039] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[23]  ( .D(n948), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2423] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[23]  ( .D(n992), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2455] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[23]  ( .D(n1029), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2487] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[23]  ( .D(n1066), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2519] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[23]  ( .D(n1103), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2551] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[23]  ( .D(n5760), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2071] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[23]  ( .D(n5799), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2103] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[23]  ( .D(n5835), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2135] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[23]  ( .D(n5871), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2167] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[23]  ( .D(n5907), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2199] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[23]  ( .D(n5943), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2231] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[23]  ( .D(n5979), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2263] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[23]  ( .D(n6015), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2295] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[23]  ( .D(n6052), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2327] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[23]  ( .D(n6088), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2359] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[23]  ( .D(n6122), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2391] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[24]  ( .D(n6992), .CK(CLK), .Q(
        DRAM_ADDRESS[24]), .QN(n523) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[24]  ( .D(n1139), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[24] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[26]  ( .D(n6990), .CK(CLK), .Q(
        DRAM_ADDRESS[26]), .QN(n524) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[26]  ( .D(n1137), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[26] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[27]  ( .D(n6989), .CK(CLK), .Q(
        DRAM_ADDRESS[27]), .QN(n525) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[27]  ( .D(n1136), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[27] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[28]  ( .D(n6988), .CK(CLK), .Q(
        DRAM_ADDRESS[28]), .QN(n526) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[28]  ( .D(n1135), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[28] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[30]  ( .D(n6986), .CK(CLK), .Q(
        DRAM_ADDRESS[30]), .QN(n527) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[30]  ( .D(n1133), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[30] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[31]  ( .D(n6985), .CK(CLK), .Q(
        DRAM_ADDRESS[31]), .QN(n528) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[31]  ( .D(n1130), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[31] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[31]  ( .D(n6761), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[63] ), .QN(n641) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[31]  ( .D(n6793), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[95] ), .QN(n673) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[31]  ( .D(n6825), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[127] ), .QN(n705) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[31]  ( .D(n6857), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[159] ), .QN(n737) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[31]  ( .D(n6889), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[191] ), .QN(n769) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[31]  ( .D(n6921), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[223] ), .QN(n801) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[31]  ( .D(n6953), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[255] ), .QN(n833) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[31]  ( .D(n3147), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[31] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[31]  ( .D(n3374), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[63] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[31]  ( .D(n3412), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[95] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[31]  ( .D(n3450), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[127] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[31]  ( .D(n3488), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[159] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[31]  ( .D(n3526), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[191] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[31]  ( .D(n3564), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[223] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[31]  ( .D(n3602), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[255] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[31]  ( .D(n3640), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[287] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[31]  ( .D(n3677), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[319] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[31]  ( .D(n3714), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[351] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[31]  ( .D(n3751), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[383] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[31]  ( .D(n3786), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[415] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[31]  ( .D(n3821), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[447] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[31]  ( .D(n3856), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[479] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[31]  ( .D(n3891), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[511] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[31]  ( .D(n3959), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[543] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[31]  ( .D(n4027), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[575] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[31]  ( .D(n4062), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[607] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[31]  ( .D(n4097), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[639] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[31]  ( .D(n4132), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[671] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[31]  ( .D(n4167), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[703] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[31]  ( .D(n4202), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[735] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[31]  ( .D(n4237), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[767] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[31]  ( .D(n4272), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[799] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[31]  ( .D(n4307), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[831] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[31]  ( .D(n4342), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[863] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[31]  ( .D(n4377), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[895] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[31]  ( .D(n4412), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[927] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[31]  ( .D(n4447), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[959] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[31]  ( .D(n4482), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[991] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[31]  ( .D(n4517), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1023] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[31]  ( .D(n4552), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1055] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[31]  ( .D(n4620), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1087] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[31]  ( .D(n4655), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1119] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[31]  ( .D(n4690), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1151] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[31]  ( .D(n4725), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1183] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[31]  ( .D(n4760), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1215] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[31]  ( .D(n4795), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1247] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[31]  ( .D(n4830), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1279] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[31]  ( .D(n4865), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1311] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[31]  ( .D(n4900), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1343] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[31]  ( .D(n4935), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1375] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[31]  ( .D(n4970), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1407] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[31]  ( .D(n5005), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1439] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[31]  ( .D(n5040), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1471] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[31]  ( .D(n5075), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1503] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[31]  ( .D(n5110), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1535] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[31]  ( .D(n5145), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1567] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[31]  ( .D(n5212), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1599] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[31]  ( .D(n5248), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1631] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[31]  ( .D(n5283), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1663] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[31]  ( .D(n5318), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1695] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[31]  ( .D(n5353), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1727] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[31]  ( .D(n5388), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1759] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[31]  ( .D(n5423), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1791] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[31]  ( .D(n5458), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1823] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[31]  ( .D(n5493), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1855] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[31]  ( .D(n5528), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1887] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[31]  ( .D(n5563), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1919] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[31]  ( .D(n5602), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1951] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[31]  ( .D(n5639), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1983] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[31]  ( .D(n5676), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2015] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[31]  ( .D(n5713), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2047] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[31]  ( .D(n930), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2431] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[31]  ( .D(n982), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2463] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[31]  ( .D(n1019), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2495] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[31]  ( .D(n1056), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2527] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[31]  ( .D(n1093), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2559] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[31]  ( .D(n5750), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2079] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[31]  ( .D(n5789), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2111] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[31]  ( .D(n5825), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2143] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[31]  ( .D(n5861), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2175] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[31]  ( .D(n5897), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2207] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[31]  ( .D(n5933), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2239] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[31]  ( .D(n5969), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2271] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[31]  ( .D(n6005), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2303] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[31]  ( .D(n6042), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2335] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[31]  ( .D(n6078), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2367] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[31]  ( .D(n6114), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2399] ) );
  DFF_X1 \DataPath/REG_ALU_OUT/Q_reg[0]  ( .D(n7013), .CK(CLK), .Q(n8208), 
        .QN(n507) );
  DFF_X1 \DataPath/REG_MEM_ALUOUT/Q_reg[0]  ( .D(n1163), .CK(CLK), .QN(
        \DataPath/i_REG_MEM_ALUOUT[0] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[17]  ( .D(n2206), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[17] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[17]  ( .D(n6775), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[49] ), .QN(n627) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[17]  ( .D(n6807), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[81] ), .QN(n659) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[17]  ( .D(n6839), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[113] ), .QN(n691) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[17]  ( .D(n6871), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[145] ), .QN(n723) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[17]  ( .D(n6903), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[177] ), .QN(n755) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[17]  ( .D(n6935), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[209] ), .QN(n787) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[17]  ( .D(n6967), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[241] ), .QN(n819) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[17]  ( .D(n3333), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[17] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[17]  ( .D(n3390), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[49] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[17]  ( .D(n3428), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[81] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[17]  ( .D(n3466), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[113] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[17]  ( .D(n3504), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[145] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[17]  ( .D(n3542), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[177] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[17]  ( .D(n3580), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[209] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[17]  ( .D(n3618), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[241] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[17]  ( .D(n3656), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[273] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[17]  ( .D(n3693), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[305] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[17]  ( .D(n3730), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[337] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[17]  ( .D(n3767), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[369] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[17]  ( .D(n3802), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[401] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[17]  ( .D(n3837), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[433] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[17]  ( .D(n3872), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[465] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[17]  ( .D(n3921), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[497] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[17]  ( .D(n3989), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[529] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[17]  ( .D(n4043), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[561] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[17]  ( .D(n4078), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[593] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[17]  ( .D(n4113), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[625] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[17]  ( .D(n4148), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[657] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[17]  ( .D(n4183), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[689] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[17]  ( .D(n4218), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[721] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[17]  ( .D(n4253), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[753] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[17]  ( .D(n4288), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[785] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[17]  ( .D(n4323), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[817] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[17]  ( .D(n4358), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[849] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[17]  ( .D(n4393), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[881] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[17]  ( .D(n4428), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[913] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[17]  ( .D(n4463), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[945] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[17]  ( .D(n4498), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[977] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[17]  ( .D(n4533), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1009] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[17]  ( .D(n4582), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1041] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[17]  ( .D(n4636), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1073] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[17]  ( .D(n4671), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1105] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[17]  ( .D(n4706), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1137] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[17]  ( .D(n4741), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1169] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[17]  ( .D(n4776), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1201] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[17]  ( .D(n4811), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1233] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[17]  ( .D(n4846), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1265] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[17]  ( .D(n4881), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1297] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[17]  ( .D(n4916), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1329] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[17]  ( .D(n4951), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1361] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[17]  ( .D(n4986), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1393] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[17]  ( .D(n5021), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1425] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[17]  ( .D(n5056), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1457] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[17]  ( .D(n5091), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1489] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[17]  ( .D(n5126), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1521] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[17]  ( .D(n5175), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1553] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[17]  ( .D(n5228), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1585] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[17]  ( .D(n5264), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1617] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[17]  ( .D(n5299), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1649] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[17]  ( .D(n5334), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1681] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[17]  ( .D(n5369), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1713] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[17]  ( .D(n5404), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1745] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[17]  ( .D(n5439), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1777] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[17]  ( .D(n5474), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1809] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[17]  ( .D(n5509), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1841] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[17]  ( .D(n5544), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1873] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[17]  ( .D(n5579), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1905] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[17]  ( .D(n5618), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1937] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[17]  ( .D(n5655), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1969] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[17]  ( .D(n5692), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2001] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[17]  ( .D(n5729), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2033] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[17]  ( .D(n892), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2385] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[17]  ( .D(n960), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2417] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[17]  ( .D(n998), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2449] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[17]  ( .D(n1035), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2481] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[17]  ( .D(n1072), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2513] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[17]  ( .D(n1109), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2545] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[17]  ( .D(n5766), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2065] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[17]  ( .D(n5805), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2097] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[17]  ( .D(n5841), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2129] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[17]  ( .D(n5877), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2161] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[17]  ( .D(n5913), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2193] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[17]  ( .D(n5949), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2225] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[17]  ( .D(n5985), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2257] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[17]  ( .D(n6021), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2289] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[17]  ( .D(n6058), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2321] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[17]  ( .D(n6094), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2353] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[25]  ( .D(n2198), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[25] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[25]  ( .D(n3317), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[25] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[25]  ( .D(n3382), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[57] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[25]  ( .D(n3420), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[89] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[25]  ( .D(n3458), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[121] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[25]  ( .D(n3496), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[153] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[25]  ( .D(n3534), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[185] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[25]  ( .D(n3572), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[217] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[25]  ( .D(n3610), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[249] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[25]  ( .D(n3648), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[281] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[25]  ( .D(n3685), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[313] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[25]  ( .D(n3722), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[345] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[25]  ( .D(n3759), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[377] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[25]  ( .D(n3794), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[409] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[25]  ( .D(n3829), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[441] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[25]  ( .D(n3864), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[473] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[25]  ( .D(n3905), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[505] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[25]  ( .D(n3973), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[537] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[25]  ( .D(n4035), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[569] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[25]  ( .D(n4070), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[601] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[25]  ( .D(n4105), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[633] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[25]  ( .D(n4140), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[665] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[25]  ( .D(n4175), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[697] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[25]  ( .D(n4210), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[729] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[25]  ( .D(n4245), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[761] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[25]  ( .D(n4280), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[793] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[25]  ( .D(n4315), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[825] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[25]  ( .D(n4350), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[857] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[25]  ( .D(n4385), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[889] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[25]  ( .D(n4420), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[921] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[25]  ( .D(n4455), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[953] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[25]  ( .D(n4490), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[985] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[25]  ( .D(n4525), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1017] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[25]  ( .D(n4566), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1049] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[25]  ( .D(n4628), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1081] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[25]  ( .D(n4663), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1113] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[25]  ( .D(n4698), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1145] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[25]  ( .D(n4733), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1177] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[25]  ( .D(n4768), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1209] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[25]  ( .D(n4803), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1241] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[25]  ( .D(n4838), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1273] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[25]  ( .D(n4873), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1305] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[25]  ( .D(n4908), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1337] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[25]  ( .D(n4943), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1369] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[25]  ( .D(n4978), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1401] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[25]  ( .D(n5013), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1433] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[25]  ( .D(n5048), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1465] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[25]  ( .D(n5083), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1497] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[25]  ( .D(n5118), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1529] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[25]  ( .D(n5159), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1561] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[25]  ( .D(n5220), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1593] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[25]  ( .D(n5256), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1625] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[25]  ( .D(n5291), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1657] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[25]  ( .D(n5326), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1689] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[25]  ( .D(n5361), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1721] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[25]  ( .D(n5396), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1753] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[25]  ( .D(n5431), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1785] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[25]  ( .D(n5466), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1817] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[25]  ( .D(n5501), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1849] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[25]  ( .D(n5536), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1881] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[25]  ( .D(n5571), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1913] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[25]  ( .D(n5610), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1945] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[25]  ( .D(n5647), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1977] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[25]  ( .D(n5684), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2009] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[25]  ( .D(n5721), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2041] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[25]  ( .D(n944), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2425] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[25]  ( .D(n990), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2457] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[25]  ( .D(n1027), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2489] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[25]  ( .D(n1064), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2521] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[25]  ( .D(n1101), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2553] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[25]  ( .D(n5758), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2073] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[25]  ( .D(n5797), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2105] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[25]  ( .D(n5833), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2137] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[25]  ( .D(n5869), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2169] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[25]  ( .D(n5905), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2201] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[25]  ( .D(n5941), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2233] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[25]  ( .D(n5977), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2265] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[25]  ( .D(n6013), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2297] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[25]  ( .D(n6050), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2329] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[25]  ( .D(n6086), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2361] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[25]  ( .D(n6120), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2393] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[9]  ( .D(n2214), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[9] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[9]  ( .D(n3349), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[9] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[9]  ( .D(n3398), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[41] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[9]  ( .D(n3436), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[73] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[9]  ( .D(n3474), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[105] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[9]  ( .D(n3512), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[137] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[9]  ( .D(n3550), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[169] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[9]  ( .D(n3588), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[201] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[9]  ( .D(n3626), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[233] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[9]  ( .D(n3664), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[265] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[9]  ( .D(n3701), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[297] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[9]  ( .D(n3738), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[329] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[9]  ( .D(n3775), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[361] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[9]  ( .D(n3810), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[393] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[9]  ( .D(n3845), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[425] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[9]  ( .D(n3880), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[457] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[9]  ( .D(n3937), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[489] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[9]  ( .D(n4005), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[521] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[9]  ( .D(n4051), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[553] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[9]  ( .D(n4086), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[585] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[9]  ( .D(n4121), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[617] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[9]  ( .D(n4156), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[649] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[9]  ( .D(n4191), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[681] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[9]  ( .D(n4226), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[713] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[9]  ( .D(n4261), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[745] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[9]  ( .D(n4296), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[777] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[9]  ( .D(n4331), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[809] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[9]  ( .D(n4366), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[841] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[9]  ( .D(n4401), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[873] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[9]  ( .D(n4436), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[905] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[9]  ( .D(n4471), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[937] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[9]  ( .D(n4506), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[969] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[9]  ( .D(n4541), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1001] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[9]  ( .D(n4598), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1033] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[9]  ( .D(n4644), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1065] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[9]  ( .D(n4679), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1097] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[9]  ( .D(n4714), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1129] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[9]  ( .D(n4749), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1161] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[9]  ( .D(n4784), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1193] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[9]  ( .D(n4819), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1225] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[9]  ( .D(n4854), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1257] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[9]  ( .D(n4889), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1289] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[9]  ( .D(n4924), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1321] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[9]  ( .D(n4959), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1353] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[9]  ( .D(n4994), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1385] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[9]  ( .D(n5029), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1417] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[9]  ( .D(n5064), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1449] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[9]  ( .D(n5099), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1481] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[9]  ( .D(n5134), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1513] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[9]  ( .D(n5191), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1545] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[9]  ( .D(n5236), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1577] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[9]  ( .D(n5272), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1609] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[9]  ( .D(n5307), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1641] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[9]  ( .D(n5342), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1673] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[9]  ( .D(n5377), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1705] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[9]  ( .D(n5412), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1737] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[9]  ( .D(n5447), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1769] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[9]  ( .D(n5482), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1801] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[9]  ( .D(n5517), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1833] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[9]  ( .D(n5552), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1865] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[9]  ( .D(n5587), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1897] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[9]  ( .D(n5626), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1929] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[9]  ( .D(n5663), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1961] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[9]  ( .D(n5700), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1993] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[9]  ( .D(n5737), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2025] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[9]  ( .D(n910), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2377] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[9]  ( .D(n968), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2409] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[9]  ( .D(n1006), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2441] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[9]  ( .D(n1043), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2473] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[9]  ( .D(n1080), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2505] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[9]  ( .D(n1117), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2537] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[9]  ( .D(n5774), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2057] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[9]  ( .D(n5813), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2089] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[9]  ( .D(n5849), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2121] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[9]  ( .D(n5885), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2153] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[9]  ( .D(n5921), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2185] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[9]  ( .D(n5957), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2217] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[9]  ( .D(n5993), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2249] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[9]  ( .D(n6029), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2281] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[9]  ( .D(n6066), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2313] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[9]  ( .D(n6102), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2345] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[1]  ( .D(n2222), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[1] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[1]  ( .D(n3365), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[1]  ( .D(n3406), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[33] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[1]  ( .D(n3444), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[65] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[1]  ( .D(n3482), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[97] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[1]  ( .D(n3520), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[129] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[1]  ( .D(n3558), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[161] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[1]  ( .D(n3596), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[193] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[1]  ( .D(n3634), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[225] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[1]  ( .D(n3672), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[257] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[1]  ( .D(n3709), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[289] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[1]  ( .D(n3746), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[321] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[1]  ( .D(n3783), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[353] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[1]  ( .D(n3818), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[385] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[1]  ( .D(n3853), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[417] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[1]  ( .D(n3888), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[449] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[1]  ( .D(n3953), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[481] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[1]  ( .D(n4021), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[513] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[1]  ( .D(n4059), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[545] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[1]  ( .D(n4094), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[577] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[1]  ( .D(n4129), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[609] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[1]  ( .D(n4164), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[641] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[1]  ( .D(n4199), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[673] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[1]  ( .D(n4234), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[705] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[1]  ( .D(n4269), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[737] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[1]  ( .D(n4304), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[769] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[1]  ( .D(n4339), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[801] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[1]  ( .D(n4374), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[833] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[1]  ( .D(n4409), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[865] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[1]  ( .D(n4444), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[897] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[1]  ( .D(n4479), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[929] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[1]  ( .D(n4514), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[961] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[1]  ( .D(n4549), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[993] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[1]  ( .D(n4614), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1025] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[1]  ( .D(n4652), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1057] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[1]  ( .D(n4687), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1089] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[1]  ( .D(n4722), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1121] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[1]  ( .D(n4757), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1153] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[1]  ( .D(n4792), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1185] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[1]  ( .D(n4827), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1217] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[1]  ( .D(n4862), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1249] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[1]  ( .D(n4897), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1281] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[1]  ( .D(n4932), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1313] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[1]  ( .D(n4967), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1345] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[1]  ( .D(n5002), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1377] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[1]  ( .D(n5037), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1409] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[1]  ( .D(n5072), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1441] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[1]  ( .D(n5107), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1473] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[1]  ( .D(n5142), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1505] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[1]  ( .D(n5207), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1537] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[1]  ( .D(n5244), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1569] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[1]  ( .D(n5280), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1601] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[1]  ( .D(n5315), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1633] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[1]  ( .D(n5350), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1665] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[1]  ( .D(n5385), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1697] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[1]  ( .D(n5420), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1729] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[1]  ( .D(n5455), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1761] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[1]  ( .D(n5490), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1793] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[1]  ( .D(n5525), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1825] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[1]  ( .D(n5560), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1857] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[1]  ( .D(n5595), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1889] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[1]  ( .D(n5634), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1921] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[1]  ( .D(n5671), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1953] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[1]  ( .D(n5708), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1985] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[1]  ( .D(n5745), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2017] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[1]  ( .D(n926), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2369] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[1]  ( .D(n976), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2401] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[1]  ( .D(n1014), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2433] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[1]  ( .D(n1051), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2465] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[1]  ( .D(n1088), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2497] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[1]  ( .D(n1125), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2529] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[1]  ( .D(n5782), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2049] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[1]  ( .D(n5821), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2081] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[1]  ( .D(n5857), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2113] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[1]  ( .D(n5893), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2145] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[1]  ( .D(n5929), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2177] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[1]  ( .D(n5965), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2209] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[1]  ( .D(n6001), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2241] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[1]  ( .D(n6037), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2273] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[1]  ( .D(n6074), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2305] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[1]  ( .D(n6110), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2337] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[14]  ( .D(n2209), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[14] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[14]  ( .D(n6778), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[46] ), .QN(n624) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[14]  ( .D(n6810), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[78] ), .QN(n656) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[14]  ( .D(n6842), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[110] ), .QN(n688) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[14]  ( .D(n6874), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[142] ), .QN(n720) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[14]  ( .D(n6906), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[174] ), .QN(n752) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[14]  ( .D(n6938), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[206] ), .QN(n784) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[14]  ( .D(n6970), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[238] ), .QN(n816) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[14]  ( .D(n3339), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[14] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[14]  ( .D(n3393), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[46] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[14]  ( .D(n3431), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[78] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[14]  ( .D(n3469), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[110] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[14]  ( .D(n3507), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[142] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[14]  ( .D(n3545), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[174] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[14]  ( .D(n3583), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[206] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[14]  ( .D(n3621), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[238] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[14]  ( .D(n3659), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[270] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[14]  ( .D(n3696), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[302] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[14]  ( .D(n3733), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[334] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[14]  ( .D(n3770), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[366] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[14]  ( .D(n3805), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[398] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[14]  ( .D(n3840), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[430] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[14]  ( .D(n3875), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[462] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[14]  ( .D(n3927), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[494] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[14]  ( .D(n3995), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[526] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[14]  ( .D(n4046), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[558] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[14]  ( .D(n4081), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[590] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[14]  ( .D(n4116), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[622] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[14]  ( .D(n4151), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[654] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[14]  ( .D(n4186), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[686] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[14]  ( .D(n4221), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[718] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[14]  ( .D(n4256), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[750] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[14]  ( .D(n4291), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[782] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[14]  ( .D(n4326), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[814] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[14]  ( .D(n4361), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[846] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[14]  ( .D(n4396), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[878] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[14]  ( .D(n4431), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[910] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[14]  ( .D(n4466), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[942] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[14]  ( .D(n4501), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[974] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[14]  ( .D(n4536), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1006] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[14]  ( .D(n4588), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1038] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[14]  ( .D(n4639), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1070] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[14]  ( .D(n4674), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1102] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[14]  ( .D(n4709), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1134] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[14]  ( .D(n4744), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1166] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[14]  ( .D(n4779), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1198] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[14]  ( .D(n4814), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1230] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[14]  ( .D(n4849), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1262] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[14]  ( .D(n4884), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1294] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[14]  ( .D(n4919), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1326] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[14]  ( .D(n4954), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1358] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[14]  ( .D(n4989), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1390] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[14]  ( .D(n5024), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1422] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[14]  ( .D(n5059), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1454] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[14]  ( .D(n5094), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1486] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[14]  ( .D(n5129), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1518] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[14]  ( .D(n5181), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1550] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[14]  ( .D(n5231), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1582] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[14]  ( .D(n5267), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1614] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[14]  ( .D(n5302), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1646] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[14]  ( .D(n5337), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1678] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[14]  ( .D(n5372), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1710] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[14]  ( .D(n5407), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1742] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[14]  ( .D(n5442), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1774] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[14]  ( .D(n5477), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1806] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[14]  ( .D(n5512), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1838] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[14]  ( .D(n5547), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1870] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[14]  ( .D(n5582), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1902] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[14]  ( .D(n5621), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1934] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[14]  ( .D(n5658), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1966] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[14]  ( .D(n5695), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1998] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[14]  ( .D(n5732), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2030] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[14]  ( .D(n900), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2382] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[14]  ( .D(n963), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2414] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[14]  ( .D(n1001), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2446] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[14]  ( .D(n1038), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2478] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[14]  ( .D(n1075), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2510] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[14]  ( .D(n1112), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2542] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[14]  ( .D(n5769), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2062] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[14]  ( .D(n5808), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2094] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[14]  ( .D(n5844), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2126] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[14]  ( .D(n5880), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2158] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[14]  ( .D(n5916), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2190] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[14]  ( .D(n5952), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2222] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[14]  ( .D(n5988), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2254] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[14]  ( .D(n6024), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2286] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[14]  ( .D(n6061), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2318] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[14]  ( .D(n6097), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2350] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[22]  ( .D(n2201), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[22] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[22]  ( .D(n3323), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[22] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[22]  ( .D(n3385), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[54] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[22]  ( .D(n3423), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[86] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[22]  ( .D(n3461), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[118] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[22]  ( .D(n3499), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[150] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[22]  ( .D(n3537), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[182] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[22]  ( .D(n3575), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[214] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[22]  ( .D(n3613), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[246] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[22]  ( .D(n3651), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[278] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[22]  ( .D(n3688), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[310] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[22]  ( .D(n3725), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[342] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[22]  ( .D(n3762), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[374] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[22]  ( .D(n3797), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[406] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[22]  ( .D(n3832), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[438] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[22]  ( .D(n3867), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[470] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[22]  ( .D(n3911), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[502] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[22]  ( .D(n3979), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[534] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[22]  ( .D(n4038), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[566] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[22]  ( .D(n4073), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[598] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[22]  ( .D(n4108), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[630] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[22]  ( .D(n4143), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[662] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[22]  ( .D(n4178), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[694] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[22]  ( .D(n4213), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[726] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[22]  ( .D(n4248), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[758] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[22]  ( .D(n4283), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[790] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[22]  ( .D(n4318), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[822] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[22]  ( .D(n4353), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[854] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[22]  ( .D(n4388), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[886] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[22]  ( .D(n4423), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[918] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[22]  ( .D(n4458), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[950] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[22]  ( .D(n4493), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[982] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[22]  ( .D(n4528), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1014] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[22]  ( .D(n4572), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1046] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[22]  ( .D(n4631), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1078] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[22]  ( .D(n4666), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1110] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[22]  ( .D(n4701), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1142] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[22]  ( .D(n4736), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1174] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[22]  ( .D(n4771), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1206] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[22]  ( .D(n4806), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1238] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[22]  ( .D(n4841), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1270] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[22]  ( .D(n4876), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1302] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[22]  ( .D(n4911), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1334] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[22]  ( .D(n4946), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1366] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[22]  ( .D(n4981), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1398] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[22]  ( .D(n5016), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1430] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[22]  ( .D(n5051), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1462] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[22]  ( .D(n5086), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1494] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[22]  ( .D(n5121), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1526] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[22]  ( .D(n5165), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1558] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[22]  ( .D(n5223), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1590] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[22]  ( .D(n5259), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1622] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[22]  ( .D(n5294), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1654] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[22]  ( .D(n5329), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1686] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[22]  ( .D(n5364), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1718] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[22]  ( .D(n5399), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1750] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[22]  ( .D(n5434), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1782] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[22]  ( .D(n5469), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1814] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[22]  ( .D(n5504), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1846] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[22]  ( .D(n5539), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1878] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[22]  ( .D(n5574), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1910] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[22]  ( .D(n5613), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1942] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[22]  ( .D(n5650), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1974] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[22]  ( .D(n5687), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2006] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[22]  ( .D(n5724), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2038] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[22]  ( .D(n950), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2422] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[22]  ( .D(n993), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2454] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[22]  ( .D(n1030), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2486] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[22]  ( .D(n1067), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2518] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[22]  ( .D(n1104), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2550] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[22]  ( .D(n5761), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2070] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[22]  ( .D(n5800), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2102] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[22]  ( .D(n5836), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2134] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[22]  ( .D(n5872), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2166] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[22]  ( .D(n5908), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2198] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[22]  ( .D(n5944), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2230] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[22]  ( .D(n5980), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2262] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[22]  ( .D(n6016), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2294] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[22]  ( .D(n6053), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2326] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[22]  ( .D(n6089), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2358] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[22]  ( .D(n6123), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2390] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[30]  ( .D(n2193), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[30] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[30]  ( .D(n6762), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[62] ), .QN(n640) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[30]  ( .D(n6794), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[94] ), .QN(n672) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[30]  ( .D(n6826), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[126] ), .QN(n704) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[30]  ( .D(n6858), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[158] ), .QN(n736) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[30]  ( .D(n6890), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[190] ), .QN(n768) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[30]  ( .D(n6922), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[222] ), .QN(n800) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[30]  ( .D(n6954), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[254] ), .QN(n832) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[30]  ( .D(n3307), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[30] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[30]  ( .D(n3377), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[62] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[30]  ( .D(n3415), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[94] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[30]  ( .D(n3453), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[126] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[30]  ( .D(n3491), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[158] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[30]  ( .D(n3529), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[190] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[30]  ( .D(n3567), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[222] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[30]  ( .D(n3605), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[254] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[30]  ( .D(n3643), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[286] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[30]  ( .D(n3680), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[318] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[30]  ( .D(n3717), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[350] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[30]  ( .D(n3754), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[382] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[30]  ( .D(n3789), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[414] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[30]  ( .D(n3824), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[446] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[30]  ( .D(n3859), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[478] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[30]  ( .D(n3895), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[510] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[30]  ( .D(n3963), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[542] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[30]  ( .D(n4030), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[574] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[30]  ( .D(n4065), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[606] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[30]  ( .D(n4100), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[638] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[30]  ( .D(n4135), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[670] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[30]  ( .D(n4170), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[702] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[30]  ( .D(n4205), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[734] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[30]  ( .D(n4240), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[766] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[30]  ( .D(n4275), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[798] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[30]  ( .D(n4310), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[830] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[30]  ( .D(n4345), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[862] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[30]  ( .D(n4380), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[894] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[30]  ( .D(n4415), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[926] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[30]  ( .D(n4450), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[958] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[30]  ( .D(n4485), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[990] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[30]  ( .D(n4520), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1022] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[30]  ( .D(n4556), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1054] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[30]  ( .D(n4623), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1086] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[30]  ( .D(n4658), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1118] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[30]  ( .D(n4693), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1150] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[30]  ( .D(n4728), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1182] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[30]  ( .D(n4763), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1214] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[30]  ( .D(n4798), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1246] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[30]  ( .D(n4833), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1278] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[30]  ( .D(n4868), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1310] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[30]  ( .D(n4903), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1342] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[30]  ( .D(n4938), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1374] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[30]  ( .D(n4973), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1406] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[30]  ( .D(n5008), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1438] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[30]  ( .D(n5043), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1470] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[30]  ( .D(n5078), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1502] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[30]  ( .D(n5113), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1534] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[30]  ( .D(n5149), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1566] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[30]  ( .D(n5215), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1598] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[30]  ( .D(n5251), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1630] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[30]  ( .D(n5286), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1662] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[30]  ( .D(n5321), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1694] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[30]  ( .D(n5356), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1726] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[30]  ( .D(n5391), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1758] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[30]  ( .D(n5426), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1790] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[30]  ( .D(n5461), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1822] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[30]  ( .D(n5496), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1854] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[30]  ( .D(n5531), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1886] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[30]  ( .D(n5566), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1918] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[30]  ( .D(n5605), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1950] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[30]  ( .D(n5642), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1982] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[30]  ( .D(n5679), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2014] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[30]  ( .D(n5716), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2046] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[30]  ( .D(n934), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2430] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[30]  ( .D(n985), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2462] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[30]  ( .D(n1022), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2494] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[30]  ( .D(n1059), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2526] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[30]  ( .D(n1096), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2558] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[30]  ( .D(n5753), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2078] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[30]  ( .D(n5792), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2110] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[30]  ( .D(n5828), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2142] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[30]  ( .D(n5864), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2174] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[30]  ( .D(n5900), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2206] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[30]  ( .D(n5936), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2238] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[30]  ( .D(n5972), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2270] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[30]  ( .D(n6008), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2302] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[30]  ( .D(n6045), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2334] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[30]  ( .D(n6081), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2366] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[30]  ( .D(n6115), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2398] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[6]  ( .D(n2217), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[6] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[6]  ( .D(n3355), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[6] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[6]  ( .D(n3401), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[38] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[6]  ( .D(n3439), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[70] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[6]  ( .D(n3477), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[102] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[6]  ( .D(n3515), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[134] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[6]  ( .D(n3553), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[166] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[6]  ( .D(n3591), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[198] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[6]  ( .D(n3629), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[230] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[6]  ( .D(n3667), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[262] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[6]  ( .D(n3704), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[294] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[6]  ( .D(n3741), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[326] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[6]  ( .D(n3778), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[358] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[6]  ( .D(n3813), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[390] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[6]  ( .D(n3848), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[422] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[6]  ( .D(n3883), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[454] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[6]  ( .D(n3943), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[486] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[6]  ( .D(n4011), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[518] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[6]  ( .D(n4054), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[550] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[6]  ( .D(n4089), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[582] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[6]  ( .D(n4124), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[614] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[6]  ( .D(n4159), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[646] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[6]  ( .D(n4194), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[678] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[6]  ( .D(n4229), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[710] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[6]  ( .D(n4264), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[742] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[6]  ( .D(n4299), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[774] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[6]  ( .D(n4334), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[806] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[6]  ( .D(n4369), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[838] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[6]  ( .D(n4404), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[870] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[6]  ( .D(n4439), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[902] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[6]  ( .D(n4474), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[934] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[6]  ( .D(n4509), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[966] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[6]  ( .D(n4544), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[998] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[6]  ( .D(n4604), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1030] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[6]  ( .D(n4647), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1062] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[6]  ( .D(n4682), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1094] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[6]  ( .D(n4717), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1126] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[6]  ( .D(n4752), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1158] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[6]  ( .D(n4787), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1190] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[6]  ( .D(n4822), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1222] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[6]  ( .D(n4857), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1254] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[6]  ( .D(n4892), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1286] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[6]  ( .D(n4927), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1318] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[6]  ( .D(n4962), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1350] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[6]  ( .D(n4997), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1382] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[6]  ( .D(n5032), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1414] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[6]  ( .D(n5067), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1446] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[6]  ( .D(n5102), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1478] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[6]  ( .D(n5137), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1510] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[6]  ( .D(n5197), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1542] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[6]  ( .D(n5239), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1574] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[6]  ( .D(n5275), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1606] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[6]  ( .D(n5310), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1638] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[6]  ( .D(n5345), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1670] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[6]  ( .D(n5380), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1702] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[6]  ( .D(n5415), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1734] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[6]  ( .D(n5450), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1766] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[6]  ( .D(n5485), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1798] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[6]  ( .D(n5520), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1830] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[6]  ( .D(n5555), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1862] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[6]  ( .D(n5590), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1894] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[6]  ( .D(n5629), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1926] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[6]  ( .D(n5666), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1958] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[6]  ( .D(n5703), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1990] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[6]  ( .D(n5740), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2022] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[6]  ( .D(n916), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2374] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[6]  ( .D(n971), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2406] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[6]  ( .D(n1009), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2438] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[6]  ( .D(n1046), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2470] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[6]  ( .D(n1083), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2502] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[6]  ( .D(n1120), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2534] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[6]  ( .D(n5777), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2054] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[6]  ( .D(n5816), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2086] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[6]  ( .D(n5852), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2118] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[6]  ( .D(n5888), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2150] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[6]  ( .D(n5924), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2182] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[6]  ( .D(n5960), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2214] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[6]  ( .D(n5996), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2246] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[6]  ( .D(n6032), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2278] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[6]  ( .D(n6069), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2310] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[6]  ( .D(n6105), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2342] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[13]  ( .D(n2210), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[13] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[13]  ( .D(n6779), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[45] ), .QN(n623) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[13]  ( .D(n6811), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[77] ), .QN(n655) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[13]  ( .D(n6843), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[109] ), .QN(n687) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[13]  ( .D(n6875), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[141] ), .QN(n719) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[13]  ( .D(n6907), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[173] ), .QN(n751) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[13]  ( .D(n6939), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[205] ), .QN(n783) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[13]  ( .D(n6971), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[237] ), .QN(n815) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[13]  ( .D(n3341), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[13] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[13]  ( .D(n3394), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[45] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[13]  ( .D(n3432), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[77] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[13]  ( .D(n3470), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[109] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[13]  ( .D(n3508), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[141] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[13]  ( .D(n3546), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[173] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[13]  ( .D(n3584), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[205] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[13]  ( .D(n3622), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[237] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[13]  ( .D(n3660), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[269] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[13]  ( .D(n3697), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[301] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[13]  ( .D(n3734), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[333] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[13]  ( .D(n3771), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[365] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[13]  ( .D(n3806), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[397] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[13]  ( .D(n3841), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[429] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[13]  ( .D(n3876), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[461] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[13]  ( .D(n3929), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[493] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[13]  ( .D(n3997), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[525] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[13]  ( .D(n4047), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[557] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[13]  ( .D(n4082), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[589] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[13]  ( .D(n4117), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[621] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[13]  ( .D(n4152), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[653] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[13]  ( .D(n4187), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[685] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[13]  ( .D(n4222), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[717] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[13]  ( .D(n4257), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[749] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[13]  ( .D(n4292), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[781] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[13]  ( .D(n4327), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[813] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[13]  ( .D(n4362), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[845] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[13]  ( .D(n4397), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[877] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[13]  ( .D(n4432), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[909] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[13]  ( .D(n4467), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[941] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[13]  ( .D(n4502), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[973] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[13]  ( .D(n4537), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1005] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[13]  ( .D(n4590), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1037] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[13]  ( .D(n4640), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1069] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[13]  ( .D(n4675), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1101] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[13]  ( .D(n4710), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1133] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[13]  ( .D(n4745), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1165] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[13]  ( .D(n4780), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1197] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[13]  ( .D(n4815), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1229] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[13]  ( .D(n4850), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1261] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[13]  ( .D(n4885), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1293] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[13]  ( .D(n4920), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1325] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[13]  ( .D(n4955), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1357] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[13]  ( .D(n4990), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1389] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[13]  ( .D(n5025), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1421] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[13]  ( .D(n5060), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1453] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[13]  ( .D(n5095), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1485] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[13]  ( .D(n5130), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1517] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[13]  ( .D(n5183), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1549] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[13]  ( .D(n5232), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1581] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[13]  ( .D(n5268), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1613] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[13]  ( .D(n5303), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1645] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[13]  ( .D(n5338), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1677] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[13]  ( .D(n5373), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1709] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[13]  ( .D(n5408), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1741] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[13]  ( .D(n5443), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1773] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[13]  ( .D(n5478), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1805] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[13]  ( .D(n5513), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1837] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[13]  ( .D(n5548), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1869] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[13]  ( .D(n5583), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1901] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[13]  ( .D(n5622), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1933] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[13]  ( .D(n5659), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1965] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[13]  ( .D(n5696), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1997] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[13]  ( .D(n5733), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2029] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[13]  ( .D(n902), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2381] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[13]  ( .D(n964), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2413] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[13]  ( .D(n1002), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2445] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[13]  ( .D(n1039), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2477] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[13]  ( .D(n1076), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2509] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[13]  ( .D(n1113), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2541] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[13]  ( .D(n5770), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2061] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[13]  ( .D(n5809), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2093] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[13]  ( .D(n5845), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2125] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[13]  ( .D(n5881), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2157] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[13]  ( .D(n5917), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2189] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[13]  ( .D(n5953), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2221] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[13]  ( .D(n5989), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2253] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[13]  ( .D(n6025), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2285] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[13]  ( .D(n6062), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2317] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[13]  ( .D(n6098), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2349] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[21]  ( .D(n2202), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[21] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[21]  ( .D(n6771), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[53] ), .QN(n631) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[21]  ( .D(n6803), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[85] ), .QN(n663) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[21]  ( .D(n6835), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[117] ), .QN(n695) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[21]  ( .D(n6867), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[149] ), .QN(n727) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[21]  ( .D(n6899), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[181] ), .QN(n759) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[21]  ( .D(n6931), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[213] ), .QN(n791) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[21]  ( .D(n6963), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[245] ), .QN(n823) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[21]  ( .D(n3325), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[21] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[21]  ( .D(n3386), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[53] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[21]  ( .D(n3424), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[85] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[21]  ( .D(n3462), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[117] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[21]  ( .D(n3500), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[149] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[21]  ( .D(n3538), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[181] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[21]  ( .D(n3576), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[213] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[21]  ( .D(n3614), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[245] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[21]  ( .D(n3652), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[277] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[21]  ( .D(n3689), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[309] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[21]  ( .D(n3726), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[341] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[21]  ( .D(n3763), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[373] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[21]  ( .D(n3798), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[405] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[21]  ( .D(n3833), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[437] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[21]  ( .D(n3868), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[469] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[21]  ( .D(n3913), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[501] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[21]  ( .D(n3981), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[533] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[21]  ( .D(n4039), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[565] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[21]  ( .D(n4074), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[597] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[21]  ( .D(n4109), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[629] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[21]  ( .D(n4144), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[661] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[21]  ( .D(n4179), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[693] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[21]  ( .D(n4214), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[725] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[21]  ( .D(n4249), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[757] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[21]  ( .D(n4284), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[789] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[21]  ( .D(n4319), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[821] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[21]  ( .D(n4354), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[853] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[21]  ( .D(n4389), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[885] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[21]  ( .D(n4424), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[917] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[21]  ( .D(n4459), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[949] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[21]  ( .D(n4494), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[981] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[21]  ( .D(n4529), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1013] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[21]  ( .D(n4574), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1045] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[21]  ( .D(n4632), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1077] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[21]  ( .D(n4667), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1109] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[21]  ( .D(n4702), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1141] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[21]  ( .D(n4737), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1173] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[21]  ( .D(n4772), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1205] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[21]  ( .D(n4807), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1237] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[21]  ( .D(n4842), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1269] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[21]  ( .D(n4877), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1301] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[21]  ( .D(n4912), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1333] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[21]  ( .D(n4947), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1365] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[21]  ( .D(n4982), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1397] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[21]  ( .D(n5017), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1429] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[21]  ( .D(n5052), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1461] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[21]  ( .D(n5087), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1493] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[21]  ( .D(n5122), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1525] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[21]  ( .D(n5167), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1557] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[21]  ( .D(n5224), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1589] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[21]  ( .D(n5260), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1621] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[21]  ( .D(n5295), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1653] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[21]  ( .D(n5330), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1685] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[21]  ( .D(n5365), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1717] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[21]  ( .D(n5400), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1749] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[21]  ( .D(n5435), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1781] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[21]  ( .D(n5470), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1813] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[21]  ( .D(n5505), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1845] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[21]  ( .D(n5540), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1877] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[21]  ( .D(n5575), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1909] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[21]  ( .D(n5614), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1941] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[21]  ( .D(n5651), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1973] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[21]  ( .D(n5688), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2005] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[21]  ( .D(n5725), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2037] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[21]  ( .D(n952), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2421] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[21]  ( .D(n994), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2453] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[21]  ( .D(n1031), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2485] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[21]  ( .D(n1068), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2517] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[21]  ( .D(n1105), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2549] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[21]  ( .D(n5762), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2069] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[21]  ( .D(n5801), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2101] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[21]  ( .D(n5837), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2133] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[21]  ( .D(n5873), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2165] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[21]  ( .D(n5909), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2197] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[21]  ( .D(n5945), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2229] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[21]  ( .D(n5981), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2261] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[21]  ( .D(n6017), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2293] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[21]  ( .D(n6054), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2325] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[21]  ( .D(n6090), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2357] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[21]  ( .D(n6124), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2389] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[29]  ( .D(n2194), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[29] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[29]  ( .D(n6763), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[61] ), .QN(n639) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[29]  ( .D(n6795), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[93] ), .QN(n671) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[29]  ( .D(n6827), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[125] ), .QN(n703) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[29]  ( .D(n6859), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[157] ), .QN(n735) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[29]  ( .D(n6891), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[189] ), .QN(n767) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[29]  ( .D(n6923), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[221] ), .QN(n799) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[29]  ( .D(n6955), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[253] ), .QN(n831) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[29]  ( .D(n3309), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[29] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[29]  ( .D(n3378), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[61] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[29]  ( .D(n3416), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[93] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[29]  ( .D(n3454), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[125] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[29]  ( .D(n3492), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[157] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[29]  ( .D(n3530), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[189] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[29]  ( .D(n3568), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[221] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[29]  ( .D(n3606), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[253] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[29]  ( .D(n3644), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[285] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[29]  ( .D(n3681), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[317] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[29]  ( .D(n3718), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[349] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[29]  ( .D(n3755), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[381] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[29]  ( .D(n3790), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[413] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[29]  ( .D(n3825), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[445] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[29]  ( .D(n3860), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[477] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[29]  ( .D(n3897), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[509] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[29]  ( .D(n3965), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[541] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[29]  ( .D(n4031), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[573] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[29]  ( .D(n4066), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[605] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[29]  ( .D(n4101), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[637] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[29]  ( .D(n4136), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[669] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[29]  ( .D(n4171), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[701] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[29]  ( .D(n4206), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[733] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[29]  ( .D(n4241), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[765] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[29]  ( .D(n4276), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[797] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[29]  ( .D(n4311), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[829] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[29]  ( .D(n4346), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[861] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[29]  ( .D(n4381), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[893] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[29]  ( .D(n4416), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[925] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[29]  ( .D(n4451), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[957] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[29]  ( .D(n4486), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[989] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[29]  ( .D(n4521), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1021] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[29]  ( .D(n4558), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1053] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[29]  ( .D(n4624), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1085] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[29]  ( .D(n4659), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1117] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[29]  ( .D(n4694), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1149] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[29]  ( .D(n4729), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1181] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[29]  ( .D(n4764), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1213] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[29]  ( .D(n4799), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1245] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[29]  ( .D(n4834), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1277] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[29]  ( .D(n4869), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1309] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[29]  ( .D(n4904), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1341] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[29]  ( .D(n4939), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1373] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[29]  ( .D(n4974), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1405] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[29]  ( .D(n5009), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1437] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[29]  ( .D(n5044), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1469] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[29]  ( .D(n5079), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1501] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[29]  ( .D(n5114), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1533] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[29]  ( .D(n5151), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1565] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[29]  ( .D(n5216), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1597] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[29]  ( .D(n5252), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1629] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[29]  ( .D(n5287), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1661] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[29]  ( .D(n5322), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1693] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[29]  ( .D(n5357), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1725] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[29]  ( .D(n5392), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1757] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[29]  ( .D(n5427), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1789] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[29]  ( .D(n5462), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1821] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[29]  ( .D(n5497), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1853] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[29]  ( .D(n5532), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1885] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[29]  ( .D(n5567), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1917] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[29]  ( .D(n5606), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1949] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[29]  ( .D(n5643), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1981] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[29]  ( .D(n5680), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2013] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[29]  ( .D(n5717), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2045] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[29]  ( .D(n936), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2429] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[29]  ( .D(n986), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2461] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[29]  ( .D(n1023), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2493] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[29]  ( .D(n1060), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2525] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[29]  ( .D(n1097), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2557] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[29]  ( .D(n5754), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2077] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[29]  ( .D(n5793), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2109] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[29]  ( .D(n5829), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2141] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[29]  ( .D(n5865), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2173] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[29]  ( .D(n5901), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2205] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[29]  ( .D(n5937), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2237] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[29]  ( .D(n5973), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2269] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[29]  ( .D(n6009), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2301] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[29]  ( .D(n6046), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2333] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[29]  ( .D(n6082), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2365] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[29]  ( .D(n6116), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2397] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[5]  ( .D(n2218), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[5] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[5]  ( .D(n3357), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[5] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[5]  ( .D(n3402), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[37] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[5]  ( .D(n3440), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[69] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[5]  ( .D(n3478), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[101] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[5]  ( .D(n3516), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[133] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[5]  ( .D(n3554), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[165] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[5]  ( .D(n3592), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[197] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[5]  ( .D(n3630), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[229] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[5]  ( .D(n3668), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[261] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[5]  ( .D(n3705), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[293] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[5]  ( .D(n3742), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[325] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[5]  ( .D(n3779), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[357] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[5]  ( .D(n3814), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[389] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[5]  ( .D(n3849), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[421] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[5]  ( .D(n3884), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[453] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[5]  ( .D(n3945), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[485] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[5]  ( .D(n4013), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[517] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[5]  ( .D(n4055), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[549] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[5]  ( .D(n4090), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[581] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[5]  ( .D(n4125), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[613] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[5]  ( .D(n4160), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[645] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[5]  ( .D(n4195), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[677] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[5]  ( .D(n4230), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[709] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[5]  ( .D(n4265), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[741] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[5]  ( .D(n4300), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[773] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[5]  ( .D(n4335), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[805] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[5]  ( .D(n4370), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[837] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[5]  ( .D(n4405), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[869] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[5]  ( .D(n4440), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[901] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[5]  ( .D(n4475), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[933] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[5]  ( .D(n4510), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[965] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[5]  ( .D(n4545), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[997] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[5]  ( .D(n4606), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1029] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[5]  ( .D(n4648), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1061] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[5]  ( .D(n4683), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1093] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[5]  ( .D(n4718), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1125] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[5]  ( .D(n4753), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1157] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[5]  ( .D(n4788), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1189] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[5]  ( .D(n4823), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1221] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[5]  ( .D(n4858), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1253] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[5]  ( .D(n4893), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1285] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[5]  ( .D(n4928), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1317] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[5]  ( .D(n4963), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1349] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[5]  ( .D(n4998), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1381] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[5]  ( .D(n5033), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1413] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[5]  ( .D(n5068), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1445] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[5]  ( .D(n5103), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1477] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[5]  ( .D(n5138), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1509] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[5]  ( .D(n5199), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1541] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[5]  ( .D(n5240), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1573] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[5]  ( .D(n5276), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1605] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[5]  ( .D(n5311), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1637] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[5]  ( .D(n5346), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1669] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[5]  ( .D(n5381), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1701] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[5]  ( .D(n5416), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1733] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[5]  ( .D(n5451), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1765] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[5]  ( .D(n5486), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1797] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[5]  ( .D(n5521), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1829] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[5]  ( .D(n5556), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1861] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[5]  ( .D(n5591), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1893] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[5]  ( .D(n5630), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1925] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[5]  ( .D(n5667), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1957] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[5]  ( .D(n5704), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1989] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[5]  ( .D(n5741), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2021] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[5]  ( .D(n918), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2373] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[5]  ( .D(n972), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2405] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[5]  ( .D(n1010), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2437] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[5]  ( .D(n1047), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2469] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[5]  ( .D(n1084), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2501] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[5]  ( .D(n1121), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2533] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[5]  ( .D(n5778), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2053] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[5]  ( .D(n5817), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2085] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[5]  ( .D(n5853), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2117] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[5]  ( .D(n5889), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2149] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[5]  ( .D(n5925), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2181] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[5]  ( .D(n5961), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2213] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[5]  ( .D(n5997), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2245] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[5]  ( .D(n6033), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2277] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[5]  ( .D(n6070), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2309] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[5]  ( .D(n6106), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2341] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[12]  ( .D(n2211), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[12] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[12]  ( .D(n6780), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[44] ), .QN(n622) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[12]  ( .D(n6812), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[76] ), .QN(n654) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[12]  ( .D(n6844), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[108] ), .QN(n686) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[12]  ( .D(n6876), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[140] ), .QN(n718) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[12]  ( .D(n6908), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[172] ), .QN(n750) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[12]  ( .D(n6940), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[204] ), .QN(n782) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[12]  ( .D(n6972), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[236] ), .QN(n814) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[12]  ( .D(n3343), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[12] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[12]  ( .D(n3395), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[44] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[12]  ( .D(n3433), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[76] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[12]  ( .D(n3471), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[108] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[12]  ( .D(n3509), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[140] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[12]  ( .D(n3547), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[172] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[12]  ( .D(n3585), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[204] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[12]  ( .D(n3623), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[236] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[12]  ( .D(n3661), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[268] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[12]  ( .D(n3698), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[300] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[12]  ( .D(n3735), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[332] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[12]  ( .D(n3772), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[364] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[12]  ( .D(n3807), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[396] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[12]  ( .D(n3842), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[428] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[12]  ( .D(n3877), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[460] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[12]  ( .D(n3931), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[492] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[12]  ( .D(n3999), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[524] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[12]  ( .D(n4048), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[556] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[12]  ( .D(n4083), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[588] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[12]  ( .D(n4118), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[620] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[12]  ( .D(n4153), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[652] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[12]  ( .D(n4188), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[684] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[12]  ( .D(n4223), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[716] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[12]  ( .D(n4258), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[748] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[12]  ( .D(n4293), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[780] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[12]  ( .D(n4328), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[812] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[12]  ( .D(n4363), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[844] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[12]  ( .D(n4398), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[876] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[12]  ( .D(n4433), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[908] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[12]  ( .D(n4468), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[940] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[12]  ( .D(n4503), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[972] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[12]  ( .D(n4538), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1004] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[12]  ( .D(n4592), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1036] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[12]  ( .D(n4641), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1068] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[12]  ( .D(n4676), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1100] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[12]  ( .D(n4711), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1132] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[12]  ( .D(n4746), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1164] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[12]  ( .D(n4781), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1196] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[12]  ( .D(n4816), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1228] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[12]  ( .D(n4851), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1260] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[12]  ( .D(n4886), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1292] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[12]  ( .D(n4921), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1324] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[12]  ( .D(n4956), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1356] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[12]  ( .D(n4991), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1388] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[12]  ( .D(n5026), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1420] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[12]  ( .D(n5061), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1452] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[12]  ( .D(n5096), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1484] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[12]  ( .D(n5131), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1516] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[12]  ( .D(n5185), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1548] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[12]  ( .D(n5233), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1580] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[12]  ( .D(n5269), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1612] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[12]  ( .D(n5304), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1644] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[12]  ( .D(n5339), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1676] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[12]  ( .D(n5374), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1708] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[12]  ( .D(n5409), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1740] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[12]  ( .D(n5444), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1772] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[12]  ( .D(n5479), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1804] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[12]  ( .D(n5514), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1836] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[12]  ( .D(n5549), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1868] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[12]  ( .D(n5584), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1900] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[12]  ( .D(n5623), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1932] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[12]  ( .D(n5660), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1964] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[12]  ( .D(n5697), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1996] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[12]  ( .D(n5734), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2028] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[12]  ( .D(n904), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2380] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[12]  ( .D(n965), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2412] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[12]  ( .D(n1003), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2444] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[12]  ( .D(n1040), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2476] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[12]  ( .D(n1077), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2508] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[12]  ( .D(n1114), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2540] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[12]  ( .D(n5771), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2060] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[12]  ( .D(n5810), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2092] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[12]  ( .D(n5846), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2124] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[12]  ( .D(n5882), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2156] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[12]  ( .D(n5918), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2188] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[12]  ( .D(n5954), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2220] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[12]  ( .D(n5990), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2252] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[12]  ( .D(n6026), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2284] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[12]  ( .D(n6063), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2316] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[12]  ( .D(n6099), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2348] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[20]  ( .D(n2203), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[20] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[20]  ( .D(n6772), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[52] ), .QN(n630) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[20]  ( .D(n6804), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[84] ), .QN(n662) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[20]  ( .D(n6836), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[116] ), .QN(n694) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[20]  ( .D(n6868), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[148] ), .QN(n726) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[20]  ( .D(n6900), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[180] ), .QN(n758) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[20]  ( .D(n6932), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[212] ), .QN(n790) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[20]  ( .D(n6964), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[244] ), .QN(n822) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[20]  ( .D(n3327), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[20] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[20]  ( .D(n3387), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[52] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[20]  ( .D(n3425), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[84] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[20]  ( .D(n3463), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[116] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[20]  ( .D(n3501), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[148] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[20]  ( .D(n3539), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[180] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[20]  ( .D(n3577), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[212] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[20]  ( .D(n3615), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[244] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[20]  ( .D(n3653), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[276] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[20]  ( .D(n3690), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[308] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[20]  ( .D(n3727), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[340] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[20]  ( .D(n3764), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[372] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[20]  ( .D(n3799), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[404] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[20]  ( .D(n3834), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[436] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[20]  ( .D(n3869), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[468] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[20]  ( .D(n3915), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[500] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[20]  ( .D(n3983), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[532] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[20]  ( .D(n4040), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[564] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[20]  ( .D(n4075), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[596] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[20]  ( .D(n4110), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[628] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[20]  ( .D(n4145), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[660] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[20]  ( .D(n4180), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[692] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[20]  ( .D(n4215), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[724] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[20]  ( .D(n4250), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[756] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[20]  ( .D(n4285), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[788] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[20]  ( .D(n4320), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[820] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[20]  ( .D(n4355), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[852] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[20]  ( .D(n4390), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[884] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[20]  ( .D(n4425), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[916] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[20]  ( .D(n4460), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[948] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[20]  ( .D(n4495), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[980] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[20]  ( .D(n4530), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1012] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[20]  ( .D(n4576), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1044] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[20]  ( .D(n4633), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1076] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[20]  ( .D(n4668), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1108] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[20]  ( .D(n4703), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1140] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[20]  ( .D(n4738), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1172] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[20]  ( .D(n4773), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1204] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[20]  ( .D(n4808), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1236] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[20]  ( .D(n4843), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1268] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[20]  ( .D(n4878), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1300] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[20]  ( .D(n4913), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1332] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[20]  ( .D(n4948), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1364] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[20]  ( .D(n4983), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1396] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[20]  ( .D(n5018), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1428] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[20]  ( .D(n5053), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1460] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[20]  ( .D(n5088), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1492] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[20]  ( .D(n5123), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1524] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[20]  ( .D(n5169), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1556] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[20]  ( .D(n5225), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1588] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[20]  ( .D(n5261), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1620] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[20]  ( .D(n5296), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1652] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[20]  ( .D(n5331), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1684] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[20]  ( .D(n5366), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1716] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[20]  ( .D(n5401), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1748] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[20]  ( .D(n5436), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1780] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[20]  ( .D(n5471), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1812] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[20]  ( .D(n5506), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1844] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[20]  ( .D(n5541), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1876] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[20]  ( .D(n5576), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1908] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[20]  ( .D(n5615), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1940] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[20]  ( .D(n5652), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1972] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[20]  ( .D(n5689), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2004] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[20]  ( .D(n5726), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2036] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[20]  ( .D(n954), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2420] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[20]  ( .D(n995), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2452] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[20]  ( .D(n1032), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2484] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[20]  ( .D(n1069), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2516] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[20]  ( .D(n1106), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2548] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[20]  ( .D(n5763), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2068] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[20]  ( .D(n5802), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2100] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[20]  ( .D(n5838), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2132] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[20]  ( .D(n5874), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2164] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[20]  ( .D(n5910), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2196] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[20]  ( .D(n5946), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2228] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[20]  ( .D(n5982), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2260] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[20]  ( .D(n6018), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2292] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[20]  ( .D(n6055), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2324] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[20]  ( .D(n6091), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2356] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[20]  ( .D(n6125), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2388] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[28]  ( .D(n2195), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[28] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[28]  ( .D(n6764), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[60] ), .QN(n638) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[28]  ( .D(n6796), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[92] ), .QN(n670) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[28]  ( .D(n6828), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[124] ), .QN(n702) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[28]  ( .D(n6860), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[156] ), .QN(n734) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[28]  ( .D(n6892), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[188] ), .QN(n766) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[28]  ( .D(n6924), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[220] ), .QN(n798) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[28]  ( .D(n6956), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[252] ), .QN(n830) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[28]  ( .D(n3311), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[28] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[28]  ( .D(n3379), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[60] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[28]  ( .D(n3417), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[92] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[28]  ( .D(n3455), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[124] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[28]  ( .D(n3493), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[156] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[28]  ( .D(n3531), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[188] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[28]  ( .D(n3569), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[220] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[28]  ( .D(n3607), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[252] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[28]  ( .D(n3645), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[284] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[28]  ( .D(n3682), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[316] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[28]  ( .D(n3719), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[348] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[28]  ( .D(n3756), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[380] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[28]  ( .D(n3791), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[412] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[28]  ( .D(n3826), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[444] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[28]  ( .D(n3861), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[476] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[28]  ( .D(n3899), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[508] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[28]  ( .D(n3967), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[540] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[28]  ( .D(n4032), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[572] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[28]  ( .D(n4067), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[604] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[28]  ( .D(n4102), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[636] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[28]  ( .D(n4137), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[668] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[28]  ( .D(n4172), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[700] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[28]  ( .D(n4207), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[732] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[28]  ( .D(n4242), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[764] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[28]  ( .D(n4277), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[796] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[28]  ( .D(n4312), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[828] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[28]  ( .D(n4347), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[860] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[28]  ( .D(n4382), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[892] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[28]  ( .D(n4417), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[924] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[28]  ( .D(n4452), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[956] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[28]  ( .D(n4487), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[988] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[28]  ( .D(n4522), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1020] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[28]  ( .D(n4560), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1052] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[28]  ( .D(n4625), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1084] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[28]  ( .D(n4660), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1116] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[28]  ( .D(n4695), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1148] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[28]  ( .D(n4730), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1180] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[28]  ( .D(n4765), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1212] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[28]  ( .D(n4800), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1244] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[28]  ( .D(n4835), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1276] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[28]  ( .D(n4870), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1308] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[28]  ( .D(n4905), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1340] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[28]  ( .D(n4940), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1372] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[28]  ( .D(n4975), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1404] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[28]  ( .D(n5010), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1436] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[28]  ( .D(n5045), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1468] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[28]  ( .D(n5080), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1500] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[28]  ( .D(n5115), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1532] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[28]  ( .D(n5153), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1564] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[28]  ( .D(n5217), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1596] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[28]  ( .D(n5253), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1628] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[28]  ( .D(n5288), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1660] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[28]  ( .D(n5323), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1692] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[28]  ( .D(n5358), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1724] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[28]  ( .D(n5393), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1756] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[28]  ( .D(n5428), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1788] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[28]  ( .D(n5463), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1820] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[28]  ( .D(n5498), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1852] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[28]  ( .D(n5533), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1884] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[28]  ( .D(n5568), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1916] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[28]  ( .D(n5607), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1948] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[28]  ( .D(n5644), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1980] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[28]  ( .D(n5681), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2012] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[28]  ( .D(n5718), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2044] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[28]  ( .D(n938), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2428] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[28]  ( .D(n987), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2460] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[28]  ( .D(n1024), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2492] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[28]  ( .D(n1061), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2524] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[28]  ( .D(n1098), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2556] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[28]  ( .D(n5755), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2076] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[28]  ( .D(n5794), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2108] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[28]  ( .D(n5830), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2140] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[28]  ( .D(n5866), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2172] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[28]  ( .D(n5902), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2204] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[28]  ( .D(n5938), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2236] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[28]  ( .D(n5974), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2268] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[28]  ( .D(n6010), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2300] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[28]  ( .D(n6047), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2332] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[28]  ( .D(n6083), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2364] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[28]  ( .D(n6117), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2396] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[4]  ( .D(n2219), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[4] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[4]  ( .D(n3359), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[4] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[4]  ( .D(n3403), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[36] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[4]  ( .D(n3441), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[68] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[4]  ( .D(n3479), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[100] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[4]  ( .D(n3517), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[132] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[4]  ( .D(n3555), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[164] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[4]  ( .D(n3593), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[196] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[4]  ( .D(n3631), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[228] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[4]  ( .D(n3669), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[260] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[4]  ( .D(n3706), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[292] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[4]  ( .D(n3743), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[324] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[4]  ( .D(n3780), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[356] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[4]  ( .D(n3815), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[388] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[4]  ( .D(n3850), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[420] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[4]  ( .D(n3885), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[452] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[4]  ( .D(n3947), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[484] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[4]  ( .D(n4015), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[516] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[4]  ( .D(n4056), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[548] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[4]  ( .D(n4091), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[580] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[4]  ( .D(n4126), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[612] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[4]  ( .D(n4161), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[644] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[4]  ( .D(n4196), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[676] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[4]  ( .D(n4231), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[708] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[4]  ( .D(n4266), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[740] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[4]  ( .D(n4301), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[772] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[4]  ( .D(n4336), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[804] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[4]  ( .D(n4371), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[836] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[4]  ( .D(n4406), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[868] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[4]  ( .D(n4441), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[900] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[4]  ( .D(n4476), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[932] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[4]  ( .D(n4511), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[964] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[4]  ( .D(n4546), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[996] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[4]  ( .D(n4608), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1028] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[4]  ( .D(n4649), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1060] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[4]  ( .D(n4684), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1092] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[4]  ( .D(n4719), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1124] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[4]  ( .D(n4754), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1156] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[4]  ( .D(n4789), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1188] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[4]  ( .D(n4824), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1220] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[4]  ( .D(n4859), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1252] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[4]  ( .D(n4894), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1284] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[4]  ( .D(n4929), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1316] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[4]  ( .D(n4964), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1348] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[4]  ( .D(n4999), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1380] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[4]  ( .D(n5034), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1412] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[4]  ( .D(n5069), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1444] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[4]  ( .D(n5104), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1476] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[4]  ( .D(n5139), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1508] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[4]  ( .D(n5201), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1540] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[4]  ( .D(n5241), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1572] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[4]  ( .D(n5277), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1604] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[4]  ( .D(n5312), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1636] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[4]  ( .D(n5347), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1668] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[4]  ( .D(n5382), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1700] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[4]  ( .D(n5417), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1732] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[4]  ( .D(n5452), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1764] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[4]  ( .D(n5487), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1796] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[4]  ( .D(n5522), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1828] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[4]  ( .D(n5557), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1860] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[4]  ( .D(n5592), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1892] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[4]  ( .D(n5631), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1924] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[4]  ( .D(n5668), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1956] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[4]  ( .D(n5705), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1988] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[4]  ( .D(n5742), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2020] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[4]  ( .D(n920), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2372] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[4]  ( .D(n973), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2404] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[4]  ( .D(n1011), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2436] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[4]  ( .D(n1048), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2468] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[4]  ( .D(n1085), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2500] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[4]  ( .D(n1122), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2532] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[4]  ( .D(n5779), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2052] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[4]  ( .D(n5818), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2084] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[4]  ( .D(n5854), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2116] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[4]  ( .D(n5890), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2148] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[4]  ( .D(n5926), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2180] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[4]  ( .D(n5962), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2212] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[4]  ( .D(n5998), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2244] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[4]  ( .D(n6034), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2276] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[4]  ( .D(n6071), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2308] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[4]  ( .D(n6107), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2340] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[11]  ( .D(n2212), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[11] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[11]  ( .D(n6781), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[43] ), .QN(n621) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[11]  ( .D(n6813), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[75] ), .QN(n653) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[11]  ( .D(n6845), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[107] ), .QN(n685) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[11]  ( .D(n6877), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[139] ), .QN(n717) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[11]  ( .D(n6909), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[171] ), .QN(n749) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[11]  ( .D(n6941), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[203] ), .QN(n781) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[11]  ( .D(n6973), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[235] ), .QN(n813) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[11]  ( .D(n3345), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[11] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[11]  ( .D(n3396), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[43] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[11]  ( .D(n3434), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[75] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[11]  ( .D(n3472), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[107] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[11]  ( .D(n3510), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[139] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[11]  ( .D(n3548), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[171] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[11]  ( .D(n3586), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[203] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[11]  ( .D(n3624), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[235] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[11]  ( .D(n3662), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[267] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[11]  ( .D(n3699), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[299] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[11]  ( .D(n3736), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[331] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[11]  ( .D(n3773), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[363] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[11]  ( .D(n3808), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[395] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[11]  ( .D(n3843), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[427] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[11]  ( .D(n3878), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[459] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[11]  ( .D(n3933), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[491] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[11]  ( .D(n4001), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[523] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[11]  ( .D(n4049), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[555] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[11]  ( .D(n4084), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[587] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[11]  ( .D(n4119), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[619] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[11]  ( .D(n4154), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[651] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[11]  ( .D(n4189), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[683] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[11]  ( .D(n4224), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[715] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[11]  ( .D(n4259), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[747] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[11]  ( .D(n4294), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[779] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[11]  ( .D(n4329), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[811] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[11]  ( .D(n4364), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[843] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[11]  ( .D(n4399), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[875] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[11]  ( .D(n4434), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[907] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[11]  ( .D(n4469), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[939] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[11]  ( .D(n4504), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[971] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[11]  ( .D(n4539), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1003] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[11]  ( .D(n4594), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1035] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[11]  ( .D(n4642), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1067] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[11]  ( .D(n4677), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1099] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[11]  ( .D(n4712), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1131] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[11]  ( .D(n4747), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1163] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[11]  ( .D(n4782), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1195] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[11]  ( .D(n4817), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1227] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[11]  ( .D(n4852), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1259] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[11]  ( .D(n4887), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1291] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[11]  ( .D(n4922), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1323] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[11]  ( .D(n4957), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1355] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[11]  ( .D(n4992), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1387] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[11]  ( .D(n5027), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1419] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[11]  ( .D(n5062), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1451] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[11]  ( .D(n5097), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1483] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[11]  ( .D(n5132), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1515] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[11]  ( .D(n5187), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1547] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[11]  ( .D(n5234), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1579] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[11]  ( .D(n5270), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1611] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[11]  ( .D(n5305), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1643] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[11]  ( .D(n5340), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1675] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[11]  ( .D(n5375), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1707] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[11]  ( .D(n5410), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1739] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[11]  ( .D(n5445), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1771] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[11]  ( .D(n5480), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1803] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[11]  ( .D(n5515), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1835] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[11]  ( .D(n5550), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1867] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[11]  ( .D(n5585), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1899] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[11]  ( .D(n5624), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1931] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[11]  ( .D(n5661), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1963] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[11]  ( .D(n5698), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1995] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[11]  ( .D(n5735), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2027] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[11]  ( .D(n906), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2379] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[11]  ( .D(n966), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2411] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[11]  ( .D(n1004), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2443] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[11]  ( .D(n1041), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2475] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[11]  ( .D(n1078), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2507] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[11]  ( .D(n1115), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2539] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[11]  ( .D(n5772), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2059] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[11]  ( .D(n5811), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2091] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[11]  ( .D(n5847), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2123] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[11]  ( .D(n5883), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2155] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[11]  ( .D(n5919), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2187] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[11]  ( .D(n5955), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2219] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[11]  ( .D(n5991), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2251] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[11]  ( .D(n6027), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2283] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[11]  ( .D(n6064), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2315] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[11]  ( .D(n6100), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2347] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[19]  ( .D(n2204), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[19] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[19]  ( .D(n6773), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[51] ), .QN(n629) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[19]  ( .D(n6805), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[83] ), .QN(n661) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[19]  ( .D(n6837), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[115] ), .QN(n693) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[19]  ( .D(n6869), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[147] ), .QN(n725) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[19]  ( .D(n6901), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[179] ), .QN(n757) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[19]  ( .D(n6933), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[211] ), .QN(n789) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[19]  ( .D(n6965), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[243] ), .QN(n821) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[19]  ( .D(n3329), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[19] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[19]  ( .D(n3388), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[51] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[19]  ( .D(n3426), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[83] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[19]  ( .D(n3464), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[115] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[19]  ( .D(n3502), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[147] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[19]  ( .D(n3540), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[179] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[19]  ( .D(n3578), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[211] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[19]  ( .D(n3616), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[243] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[19]  ( .D(n3654), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[275] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[19]  ( .D(n3691), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[307] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[19]  ( .D(n3728), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[339] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[19]  ( .D(n3765), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[371] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[19]  ( .D(n3800), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[403] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[19]  ( .D(n3835), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[435] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[19]  ( .D(n3870), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[467] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[19]  ( .D(n3917), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[499] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[19]  ( .D(n3985), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[531] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[19]  ( .D(n4041), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[563] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[19]  ( .D(n4076), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[595] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[19]  ( .D(n4111), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[627] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[19]  ( .D(n4146), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[659] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[19]  ( .D(n4181), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[691] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[19]  ( .D(n4216), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[723] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[19]  ( .D(n4251), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[755] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[19]  ( .D(n4286), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[787] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[19]  ( .D(n4321), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[819] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[19]  ( .D(n4356), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[851] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[19]  ( .D(n4391), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[883] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[19]  ( .D(n4426), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[915] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[19]  ( .D(n4461), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[947] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[19]  ( .D(n4496), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[979] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[19]  ( .D(n4531), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1011] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[19]  ( .D(n4578), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1043] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[19]  ( .D(n4634), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1075] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[19]  ( .D(n4669), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1107] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[19]  ( .D(n4704), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1139] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[19]  ( .D(n4739), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1171] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[19]  ( .D(n4774), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1203] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[19]  ( .D(n4809), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1235] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[19]  ( .D(n4844), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1267] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[19]  ( .D(n4879), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1299] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[19]  ( .D(n4914), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1331] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[19]  ( .D(n4949), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1363] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[19]  ( .D(n4984), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1395] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[19]  ( .D(n5019), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1427] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[19]  ( .D(n5054), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1459] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[19]  ( .D(n5089), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1491] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[19]  ( .D(n5124), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1523] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[19]  ( .D(n5171), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1555] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[19]  ( .D(n5226), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1587] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[19]  ( .D(n5262), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1619] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[19]  ( .D(n5297), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1651] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[19]  ( .D(n5332), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1683] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[19]  ( .D(n5367), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1715] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[19]  ( .D(n5402), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1747] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[19]  ( .D(n5437), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1779] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[19]  ( .D(n5472), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1811] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[19]  ( .D(n5507), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1843] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[19]  ( .D(n5542), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1875] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[19]  ( .D(n5577), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1907] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[19]  ( .D(n5616), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1939] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[19]  ( .D(n5653), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1971] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[19]  ( .D(n5690), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2003] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[19]  ( .D(n5727), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2035] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[19]  ( .D(n956), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2419] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[19]  ( .D(n996), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2451] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[19]  ( .D(n1033), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2483] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[19]  ( .D(n1070), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2515] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[19]  ( .D(n1107), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2547] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[19]  ( .D(n5764), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2067] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[19]  ( .D(n5803), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2099] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[19]  ( .D(n5839), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2131] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[19]  ( .D(n5875), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2163] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[19]  ( .D(n5911), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2195] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[19]  ( .D(n5947), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2227] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[19]  ( .D(n5983), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2259] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[19]  ( .D(n6019), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2291] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[19]  ( .D(n6056), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2323] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[19]  ( .D(n6092), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2355] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[19]  ( .D(n6126), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2387] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[27]  ( .D(n2196), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[27] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[27]  ( .D(n3313), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[27] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[27]  ( .D(n3380), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[59] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[27]  ( .D(n3418), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[91] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[27]  ( .D(n3456), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[123] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[27]  ( .D(n3494), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[155] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[27]  ( .D(n3532), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[187] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[27]  ( .D(n3570), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[219] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[27]  ( .D(n3608), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[251] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[27]  ( .D(n3646), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[283] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[27]  ( .D(n3683), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[315] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[27]  ( .D(n3720), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[347] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[27]  ( .D(n3757), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[379] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[27]  ( .D(n3792), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[411] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[27]  ( .D(n3827), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[443] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[27]  ( .D(n3862), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[475] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[27]  ( .D(n3901), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[507] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[27]  ( .D(n3969), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[539] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[27]  ( .D(n4033), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[571] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[27]  ( .D(n4068), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[603] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[27]  ( .D(n4103), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[635] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[27]  ( .D(n4138), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[667] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[27]  ( .D(n4173), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[699] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[27]  ( .D(n4208), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[731] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[27]  ( .D(n4243), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[763] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[27]  ( .D(n4278), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[795] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[27]  ( .D(n4313), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[827] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[27]  ( .D(n4348), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[859] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[27]  ( .D(n4383), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[891] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[27]  ( .D(n4418), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[923] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[27]  ( .D(n4453), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[955] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[27]  ( .D(n4488), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[987] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[27]  ( .D(n4523), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1019] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[27]  ( .D(n4562), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1051] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[27]  ( .D(n4626), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1083] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[27]  ( .D(n4661), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1115] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[27]  ( .D(n4696), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1147] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[27]  ( .D(n4731), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1179] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[27]  ( .D(n4766), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1211] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[27]  ( .D(n4801), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1243] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[27]  ( .D(n4836), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1275] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[27]  ( .D(n4871), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1307] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[27]  ( .D(n4906), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1339] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[27]  ( .D(n4941), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1371] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[27]  ( .D(n4976), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1403] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[27]  ( .D(n5011), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1435] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[27]  ( .D(n5046), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1467] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[27]  ( .D(n5081), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1499] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[27]  ( .D(n5116), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1531] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[27]  ( .D(n5155), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1563] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[27]  ( .D(n5218), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1595] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[27]  ( .D(n5254), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1627] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[27]  ( .D(n5289), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1659] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[27]  ( .D(n5324), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1691] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[27]  ( .D(n5359), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1723] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[27]  ( .D(n5394), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1755] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[27]  ( .D(n5429), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1787] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[27]  ( .D(n5464), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1819] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[27]  ( .D(n5499), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1851] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[27]  ( .D(n5534), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1883] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[27]  ( .D(n5569), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1915] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[27]  ( .D(n5608), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1947] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[27]  ( .D(n5645), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1979] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[27]  ( .D(n5682), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2011] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[27]  ( .D(n5719), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2043] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[27]  ( .D(n940), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2427] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[27]  ( .D(n988), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2459] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[27]  ( .D(n1025), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2491] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[27]  ( .D(n1062), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2523] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[27]  ( .D(n1099), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2555] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[27]  ( .D(n5756), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2075] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[27]  ( .D(n5795), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2107] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[27]  ( .D(n5831), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2139] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[27]  ( .D(n5867), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2171] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[27]  ( .D(n5903), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2203] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[27]  ( .D(n5939), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2235] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[27]  ( .D(n5975), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2267] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[27]  ( .D(n6011), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2299] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[27]  ( .D(n6048), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2331] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[27]  ( .D(n6084), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2363] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[27]  ( .D(n6118), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2395] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[3]  ( .D(n2220), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[3] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[3]  ( .D(n3361), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[3] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[3]  ( .D(n3404), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[35] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[3]  ( .D(n3442), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[67] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[3]  ( .D(n3480), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[99] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[3]  ( .D(n3518), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[131] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[3]  ( .D(n3556), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[163] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[3]  ( .D(n3594), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[195] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[3]  ( .D(n3632), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[227] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[3]  ( .D(n3670), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[259] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[3]  ( .D(n3707), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[291] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[3]  ( .D(n3744), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[323] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[3]  ( .D(n3781), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[355] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[3]  ( .D(n3816), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[387] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[3]  ( .D(n3851), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[419] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[3]  ( .D(n3886), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[451] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[3]  ( .D(n3949), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[483] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[3]  ( .D(n4017), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[515] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[3]  ( .D(n4057), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[547] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[3]  ( .D(n4092), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[579] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[3]  ( .D(n4127), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[611] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[3]  ( .D(n4162), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[643] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[3]  ( .D(n4197), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[675] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[3]  ( .D(n4232), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[707] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[3]  ( .D(n4267), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[739] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[3]  ( .D(n4302), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[771] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[3]  ( .D(n4337), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[803] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[3]  ( .D(n4372), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[835] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[3]  ( .D(n4407), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[867] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[3]  ( .D(n4442), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[899] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[3]  ( .D(n4477), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[931] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[3]  ( .D(n4512), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[963] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[3]  ( .D(n4547), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[995] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[3]  ( .D(n4610), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1027] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[3]  ( .D(n4650), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1059] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[3]  ( .D(n4685), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1091] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[3]  ( .D(n4720), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1123] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[3]  ( .D(n4755), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1155] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[3]  ( .D(n4790), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1187] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[3]  ( .D(n4825), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1219] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[3]  ( .D(n4860), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1251] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[3]  ( .D(n4895), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1283] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[3]  ( .D(n4930), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1315] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[3]  ( .D(n4965), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1347] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[3]  ( .D(n5000), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1379] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[3]  ( .D(n5035), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1411] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[3]  ( .D(n5070), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1443] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[3]  ( .D(n5105), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1475] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[3]  ( .D(n5140), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1507] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[3]  ( .D(n5203), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1539] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[3]  ( .D(n5242), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1571] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[3]  ( .D(n5278), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1603] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[3]  ( .D(n5313), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1635] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[3]  ( .D(n5348), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1667] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[3]  ( .D(n5383), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1699] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[3]  ( .D(n5418), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1731] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[3]  ( .D(n5453), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1763] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[3]  ( .D(n5488), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1795] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[3]  ( .D(n5523), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1827] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[3]  ( .D(n5558), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1859] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[3]  ( .D(n5593), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1891] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[3]  ( .D(n5632), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1923] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[3]  ( .D(n5669), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1955] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[3]  ( .D(n5706), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1987] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[3]  ( .D(n5743), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2019] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[3]  ( .D(n922), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2371] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[3]  ( .D(n974), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2403] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[3]  ( .D(n1012), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2435] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[3]  ( .D(n1049), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2467] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[3]  ( .D(n1086), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2499] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[3]  ( .D(n1123), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2531] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[3]  ( .D(n5780), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2051] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[3]  ( .D(n5819), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2083] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[3]  ( .D(n5855), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2115] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[3]  ( .D(n5891), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2147] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[3]  ( .D(n5927), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2179] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[3]  ( .D(n5963), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2211] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[3]  ( .D(n5999), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2243] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[3]  ( .D(n6035), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2275] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[3]  ( .D(n6072), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2307] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[3]  ( .D(n6108), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2339] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[10]  ( .D(n2213), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[10] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[10]  ( .D(n6814), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[74] ), .QN(n652) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[10]  ( .D(n6846), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[106] ), .QN(n684) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[10]  ( .D(n6942), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[202] ), .QN(n780) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[10]  ( .D(n6974), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[234] ), .QN(n812) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[10]  ( .D(n3347), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[10] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[10]  ( .D(n3397), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[42] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[10]  ( .D(n3435), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[74] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[10]  ( .D(n3473), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[106] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[10]  ( .D(n3511), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[138] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[10]  ( .D(n3549), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[170] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[10]  ( .D(n3587), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[202] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[10]  ( .D(n3625), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[234] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[10]  ( .D(n3663), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[266] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[10]  ( .D(n3700), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[298] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[10]  ( .D(n3737), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[330] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[10]  ( .D(n3774), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[362] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[10]  ( .D(n3809), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[394] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[10]  ( .D(n3844), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[426] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[10]  ( .D(n3879), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[458] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[10]  ( .D(n3935), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[490] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[10]  ( .D(n4003), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[522] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[10]  ( .D(n4050), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[554] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[10]  ( .D(n4085), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[586] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[10]  ( .D(n4120), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[618] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[10]  ( .D(n4155), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[650] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[10]  ( .D(n4190), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[682] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[10]  ( .D(n4225), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[714] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[10]  ( .D(n4260), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[746] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[10]  ( .D(n4295), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[778] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[10]  ( .D(n4330), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[810] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[10]  ( .D(n4365), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[842] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[10]  ( .D(n4400), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[874] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[10]  ( .D(n4435), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[906] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[10]  ( .D(n4470), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[938] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[10]  ( .D(n4505), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[970] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[10]  ( .D(n4540), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1002] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[10]  ( .D(n4596), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1034] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[10]  ( .D(n4643), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1066] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[10]  ( .D(n4678), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1098] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[10]  ( .D(n4713), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1130] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[10]  ( .D(n4748), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1162] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[10]  ( .D(n4783), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1194] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[10]  ( .D(n4818), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1226] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[10]  ( .D(n4853), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1258] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[10]  ( .D(n4888), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1290] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[10]  ( .D(n4923), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1322] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[10]  ( .D(n4958), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1354] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[10]  ( .D(n4993), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1386] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[10]  ( .D(n5028), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1418] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[10]  ( .D(n5063), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1450] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[10]  ( .D(n5098), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1482] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[10]  ( .D(n5133), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1514] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[10]  ( .D(n5189), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1546] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[10]  ( .D(n5235), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1578] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[10]  ( .D(n5271), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1610] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[10]  ( .D(n5306), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1642] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[10]  ( .D(n5341), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1674] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[10]  ( .D(n5376), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1706] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[10]  ( .D(n5411), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1738] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[10]  ( .D(n5446), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1770] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[10]  ( .D(n5481), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1802] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[10]  ( .D(n5516), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1834] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[10]  ( .D(n5551), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1866] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[10]  ( .D(n5586), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1898] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[10]  ( .D(n5625), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1930] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[10]  ( .D(n5662), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1962] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[10]  ( .D(n5699), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1994] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[10]  ( .D(n5736), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2026] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[10]  ( .D(n908), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2378] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[10]  ( .D(n967), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2410] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[10]  ( .D(n1005), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2442] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[10]  ( .D(n1042), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2474] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[10]  ( .D(n1079), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2506] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[10]  ( .D(n1116), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2538] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[10]  ( .D(n5773), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2058] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[10]  ( .D(n5812), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2090] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[10]  ( .D(n5848), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2122] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[10]  ( .D(n5884), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2154] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[10]  ( .D(n5920), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2186] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[10]  ( .D(n5956), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2218] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[10]  ( .D(n5992), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2250] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[10]  ( .D(n6028), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2282] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[10]  ( .D(n6065), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2314] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[10]  ( .D(n6101), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2346] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[18]  ( .D(n2205), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[18] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[18]  ( .D(n6774), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[50] ), .QN(n628) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[18]  ( .D(n6806), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[82] ), .QN(n660) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[18]  ( .D(n6838), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[114] ), .QN(n692) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[18]  ( .D(n6870), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[146] ), .QN(n724) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[18]  ( .D(n6902), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[178] ), .QN(n756) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[18]  ( .D(n6934), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[210] ), .QN(n788) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[18]  ( .D(n6966), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[242] ), .QN(n820) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[18]  ( .D(n3331), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[18] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[18]  ( .D(n3389), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[50] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[18]  ( .D(n3427), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[82] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[18]  ( .D(n3465), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[114] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[18]  ( .D(n3503), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[146] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[18]  ( .D(n3541), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[178] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[18]  ( .D(n3579), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[210] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[18]  ( .D(n3617), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[242] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[18]  ( .D(n3655), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[274] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[18]  ( .D(n3692), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[306] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[18]  ( .D(n3729), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[338] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[18]  ( .D(n3766), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[370] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[18]  ( .D(n3801), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[402] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[18]  ( .D(n3836), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[434] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[18]  ( .D(n3871), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[466] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[18]  ( .D(n3919), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[498] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[18]  ( .D(n3987), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[530] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[18]  ( .D(n4042), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[562] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[18]  ( .D(n4077), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[594] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[18]  ( .D(n4112), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[626] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[18]  ( .D(n4147), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[658] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[18]  ( .D(n4182), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[690] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[18]  ( .D(n4217), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[722] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[18]  ( .D(n4252), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[754] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[18]  ( .D(n4287), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[786] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[18]  ( .D(n4322), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[818] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[18]  ( .D(n4357), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[850] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[18]  ( .D(n4392), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[882] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[18]  ( .D(n4427), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[914] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[18]  ( .D(n4462), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[946] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[18]  ( .D(n4497), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[978] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[18]  ( .D(n4532), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1010] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[18]  ( .D(n4580), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1042] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[18]  ( .D(n4635), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1074] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[18]  ( .D(n4670), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1106] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[18]  ( .D(n4705), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1138] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[18]  ( .D(n4740), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1170] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[18]  ( .D(n4775), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1202] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[18]  ( .D(n4810), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1234] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[18]  ( .D(n4845), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1266] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[18]  ( .D(n4880), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1298] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[18]  ( .D(n4915), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1330] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[18]  ( .D(n4950), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1362] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[18]  ( .D(n4985), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1394] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[18]  ( .D(n5020), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1426] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[18]  ( .D(n5055), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1458] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[18]  ( .D(n5090), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1490] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[18]  ( .D(n5125), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1522] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[18]  ( .D(n5173), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1554] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[18]  ( .D(n5227), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1586] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[18]  ( .D(n5263), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1618] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[18]  ( .D(n5298), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1650] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[18]  ( .D(n5333), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1682] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[18]  ( .D(n5368), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1714] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[18]  ( .D(n5403), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1746] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[18]  ( .D(n5438), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1778] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[18]  ( .D(n5473), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1810] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[18]  ( .D(n5508), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1842] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[18]  ( .D(n5543), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1874] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[18]  ( .D(n5578), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1906] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[18]  ( .D(n5617), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1938] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[18]  ( .D(n5654), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1970] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[18]  ( .D(n5691), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2002] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[18]  ( .D(n5728), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2034] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[18]  ( .D(n958), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2418] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[18]  ( .D(n997), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2450] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[18]  ( .D(n1034), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2482] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[18]  ( .D(n1071), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2514] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[18]  ( .D(n1108), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2546] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[18]  ( .D(n5765), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2066] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[18]  ( .D(n5804), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2098] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[18]  ( .D(n5840), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2130] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[18]  ( .D(n5876), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2162] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[18]  ( .D(n5912), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2194] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[18]  ( .D(n5948), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2226] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[18]  ( .D(n5984), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2258] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[18]  ( .D(n6020), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2290] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[18]  ( .D(n6057), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2322] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[18]  ( .D(n6093), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2354] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[18]  ( .D(n6127), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2386] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[26]  ( .D(n2197), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[26] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[26]  ( .D(n6766), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[58] ), .QN(n636) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[26]  ( .D(n6798), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[90] ), .QN(n668) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[26]  ( .D(n6830), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[122] ), .QN(n700) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[26]  ( .D(n6862), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[154] ), .QN(n732) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[26]  ( .D(n6894), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[186] ), .QN(n764) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[26]  ( .D(n6926), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[218] ), .QN(n796) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[26]  ( .D(n6958), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[250] ), .QN(n828) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[26]  ( .D(n3315), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[26] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[26]  ( .D(n3381), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[58] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[26]  ( .D(n3419), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[90] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[26]  ( .D(n3457), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[122] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[26]  ( .D(n3495), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[154] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[26]  ( .D(n3533), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[186] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[26]  ( .D(n3571), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[218] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[26]  ( .D(n3609), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[250] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[26]  ( .D(n3647), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[282] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[26]  ( .D(n3684), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[314] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[26]  ( .D(n3721), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[346] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[26]  ( .D(n3758), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[378] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[26]  ( .D(n3793), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[410] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[26]  ( .D(n3828), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[442] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[26]  ( .D(n3863), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[474] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[26]  ( .D(n3903), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[506] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[26]  ( .D(n3971), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[538] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[26]  ( .D(n4034), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[570] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[26]  ( .D(n4069), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[602] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[26]  ( .D(n4104), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[634] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[26]  ( .D(n4139), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[666] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[26]  ( .D(n4174), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[698] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[26]  ( .D(n4209), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[730] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[26]  ( .D(n4244), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[762] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[26]  ( .D(n4279), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[794] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[26]  ( .D(n4314), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[826] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[26]  ( .D(n4349), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[858] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[26]  ( .D(n4384), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[890] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[26]  ( .D(n4419), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[922] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[26]  ( .D(n4454), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[954] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[26]  ( .D(n4489), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[986] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[26]  ( .D(n4524), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1018] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[26]  ( .D(n4564), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1050] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[26]  ( .D(n4627), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1082] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[26]  ( .D(n4662), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1114] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[26]  ( .D(n4697), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1146] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[26]  ( .D(n4732), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1178] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[26]  ( .D(n4767), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1210] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[26]  ( .D(n4802), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1242] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[26]  ( .D(n4837), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1274] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[26]  ( .D(n4872), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1306] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[26]  ( .D(n4907), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1338] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[26]  ( .D(n4942), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1370] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[26]  ( .D(n4977), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1402] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[26]  ( .D(n5012), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1434] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[26]  ( .D(n5047), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1466] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[26]  ( .D(n5082), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1498] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[26]  ( .D(n5117), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1530] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[26]  ( .D(n5157), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1562] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[26]  ( .D(n5219), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1594] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[26]  ( .D(n5255), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1626] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[26]  ( .D(n5290), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1658] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[26]  ( .D(n5325), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1690] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[26]  ( .D(n5360), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1722] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[26]  ( .D(n5395), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1754] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[26]  ( .D(n5430), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1786] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[26]  ( .D(n5465), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1818] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[26]  ( .D(n5500), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1850] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[26]  ( .D(n5535), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1882] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[26]  ( .D(n5570), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1914] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[26]  ( .D(n5609), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1946] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[26]  ( .D(n5646), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1978] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[26]  ( .D(n5683), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2010] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[26]  ( .D(n5720), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2042] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[26]  ( .D(n942), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2426] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[26]  ( .D(n989), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2458] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[26]  ( .D(n1026), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2490] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[26]  ( .D(n1063), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2522] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[26]  ( .D(n1100), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2554] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[26]  ( .D(n5757), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2074] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[26]  ( .D(n5796), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2106] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[26]  ( .D(n5832), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2138] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[26]  ( .D(n5868), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2170] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[26]  ( .D(n5904), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2202] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[26]  ( .D(n5940), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2234] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[26]  ( .D(n5976), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2266] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[26]  ( .D(n6012), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2298] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[26]  ( .D(n6049), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2330] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[26]  ( .D(n6085), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2362] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[26]  ( .D(n6119), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2394] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[2]  ( .D(n2221), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[2] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[2]  ( .D(n3363), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[2]  ( .D(n3405), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[34] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[2]  ( .D(n3443), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[66] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[2]  ( .D(n3481), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[98] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[2]  ( .D(n3519), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[130] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[2]  ( .D(n3557), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[162] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[2]  ( .D(n3595), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[194] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[2]  ( .D(n3633), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[226] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[2]  ( .D(n3671), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[258] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[2]  ( .D(n3708), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[290] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[2]  ( .D(n3745), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[322] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[2]  ( .D(n3782), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[354] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[2]  ( .D(n3817), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[386] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[2]  ( .D(n3852), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[418] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[2]  ( .D(n3887), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[450] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[2]  ( .D(n3951), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[482] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[2]  ( .D(n4019), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[514] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[2]  ( .D(n4058), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[546] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[2]  ( .D(n4093), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[578] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[2]  ( .D(n4128), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[610] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[2]  ( .D(n4163), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[642] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[2]  ( .D(n4198), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[674] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[2]  ( .D(n4233), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[706] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[2]  ( .D(n4268), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[738] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[2]  ( .D(n4303), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[770] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[2]  ( .D(n4338), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[802] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[2]  ( .D(n4373), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[834] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[2]  ( .D(n4408), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[866] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[2]  ( .D(n4443), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[898] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[2]  ( .D(n4478), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[930] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[2]  ( .D(n4513), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[962] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[2]  ( .D(n4548), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[994] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[2]  ( .D(n4612), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1026] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[2]  ( .D(n4651), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1058] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[2]  ( .D(n4686), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1090] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[2]  ( .D(n4721), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1122] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[2]  ( .D(n4756), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1154] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[2]  ( .D(n4791), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1186] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[2]  ( .D(n4826), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1218] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[2]  ( .D(n4861), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1250] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[2]  ( .D(n4896), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1282] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[2]  ( .D(n4931), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1314] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[2]  ( .D(n4966), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1346] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[2]  ( .D(n5001), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1378] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[2]  ( .D(n5036), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1410] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[2]  ( .D(n5071), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1442] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[2]  ( .D(n5106), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1474] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[2]  ( .D(n5141), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1506] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[2]  ( .D(n5205), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1538] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[2]  ( .D(n5243), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1570] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[2]  ( .D(n5279), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1602] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[2]  ( .D(n5314), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1634] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[2]  ( .D(n5349), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1666] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[2]  ( .D(n5384), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1698] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[2]  ( .D(n5419), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1730] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[2]  ( .D(n5454), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1762] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[2]  ( .D(n5489), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1794] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[2]  ( .D(n5524), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1826] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[2]  ( .D(n5559), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1858] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[2]  ( .D(n5594), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1890] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[2]  ( .D(n5633), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1922] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[2]  ( .D(n5670), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1954] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[2]  ( .D(n5707), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1986] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[2]  ( .D(n5744), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2018] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[2]  ( .D(n924), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2370] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[2]  ( .D(n975), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2402] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[2]  ( .D(n1013), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2434] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[2]  ( .D(n1050), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2466] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[2]  ( .D(n1087), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2498] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[2]  ( .D(n1124), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2530] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[2]  ( .D(n5781), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2050] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[2]  ( .D(n5820), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2082] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[2]  ( .D(n5856), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2114] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[2]  ( .D(n5892), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2146] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[2]  ( .D(n5928), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2178] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[2]  ( .D(n5964), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2210] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[2]  ( .D(n6000), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2242] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[2]  ( .D(n6036), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2274] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[2]  ( .D(n6073), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2306] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[2]  ( .D(n6109), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2338] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[16]  ( .D(n2207), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[16] ) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[16]  ( .D(n6776), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[48] ), .QN(n626) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[16]  ( .D(n6808), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[80] ), .QN(n658) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[16]  ( .D(n6840), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[112] ), .QN(n690) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[16]  ( .D(n6872), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[144] ), .QN(n722) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[16]  ( .D(n6904), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[176] ), .QN(n754) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[16]  ( .D(n6936), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[208] ), .QN(n786) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[16]  ( .D(n6968), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[240] ), .QN(n818) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[16]  ( .D(n3335), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[16] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[16]  ( .D(n3391), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[48] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[16]  ( .D(n3429), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[80] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[16]  ( .D(n3467), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[112] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[16]  ( .D(n3505), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[144] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[16]  ( .D(n3543), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[176] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[16]  ( .D(n3581), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[208] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[16]  ( .D(n3619), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[240] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[16]  ( .D(n3657), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[272] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[16]  ( .D(n3694), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[304] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[16]  ( .D(n3731), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[336] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[16]  ( .D(n3768), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[368] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[16]  ( .D(n3803), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[400] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[16]  ( .D(n3838), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[432] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[16]  ( .D(n3873), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[464] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[16]  ( .D(n3923), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[496] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[16]  ( .D(n3991), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[528] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[16]  ( .D(n4044), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[560] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[16]  ( .D(n4079), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[592] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[16]  ( .D(n4114), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[624] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[16]  ( .D(n4149), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[656] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[16]  ( .D(n4184), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[688] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[16]  ( .D(n4219), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[720] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[16]  ( .D(n4254), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[752] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[16]  ( .D(n4289), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[784] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[16]  ( .D(n4324), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[816] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[16]  ( .D(n4359), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[848] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[16]  ( .D(n4394), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[880] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[16]  ( .D(n4429), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[912] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[16]  ( .D(n4464), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[944] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[16]  ( .D(n4499), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[976] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[16]  ( .D(n4534), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1008] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[16]  ( .D(n4584), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1040] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[16]  ( .D(n4637), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1072] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[16]  ( .D(n4672), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1104] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[16]  ( .D(n4707), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1136] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[16]  ( .D(n4742), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1168] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[16]  ( .D(n4777), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1200] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[16]  ( .D(n4812), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1232] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[16]  ( .D(n4847), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1264] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[16]  ( .D(n4882), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1296] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[16]  ( .D(n4917), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1328] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[16]  ( .D(n4952), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1360] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[16]  ( .D(n4987), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1392] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[16]  ( .D(n5022), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1424] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[16]  ( .D(n5057), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1456] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[16]  ( .D(n5092), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1488] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[16]  ( .D(n5127), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1520] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[16]  ( .D(n5177), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1552] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[16]  ( .D(n5229), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1584] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[16]  ( .D(n5265), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1616] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[16]  ( .D(n5300), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1648] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[16]  ( .D(n5335), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1680] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[16]  ( .D(n5370), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1712] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[16]  ( .D(n5405), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1744] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[16]  ( .D(n5440), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1776] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[16]  ( .D(n5475), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1808] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[16]  ( .D(n5510), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1840] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[16]  ( .D(n5545), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1872] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[16]  ( .D(n5580), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1904] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[16]  ( .D(n5619), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1936] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[16]  ( .D(n5656), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1968] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[16]  ( .D(n5693), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2000] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[16]  ( .D(n5730), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2032] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[16]  ( .D(n896), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2384] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[16]  ( .D(n961), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2416] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[16]  ( .D(n999), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2448] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[16]  ( .D(n1036), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2480] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[16]  ( .D(n1073), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2512] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[16]  ( .D(n1110), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2544] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[16]  ( .D(n5767), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2064] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[16]  ( .D(n5806), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2096] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[16]  ( .D(n5842), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2128] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[16]  ( .D(n5878), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2160] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[16]  ( .D(n5914), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2192] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[16]  ( .D(n5950), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2224] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[16]  ( .D(n5986), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2256] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[16]  ( .D(n6022), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2288] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[16]  ( .D(n6059), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2320] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[16]  ( .D(n6095), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2352] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[24]  ( .D(n2199), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[24] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[24]  ( .D(n3319), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[24] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[24]  ( .D(n3383), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[56] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[24]  ( .D(n3421), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[88] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[24]  ( .D(n3459), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[120] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[24]  ( .D(n3497), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[152] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[24]  ( .D(n3535), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[184] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[24]  ( .D(n3573), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[216] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[24]  ( .D(n3611), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[248] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[24]  ( .D(n3649), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[280] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[24]  ( .D(n3686), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[312] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[24]  ( .D(n3723), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[344] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[24]  ( .D(n3760), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[376] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[24]  ( .D(n3795), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[408] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[24]  ( .D(n3830), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[440] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[24]  ( .D(n3865), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[472] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[24]  ( .D(n3907), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[504] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[24]  ( .D(n3975), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[536] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[24]  ( .D(n4036), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[568] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[24]  ( .D(n4071), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[600] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[24]  ( .D(n4106), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[632] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[24]  ( .D(n4141), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[664] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[24]  ( .D(n4176), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[696] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[24]  ( .D(n4211), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[728] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[24]  ( .D(n4246), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[760] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[24]  ( .D(n4281), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[792] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[24]  ( .D(n4316), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[824] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[24]  ( .D(n4351), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[856] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[24]  ( .D(n4386), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[888] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[24]  ( .D(n4421), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[920] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[24]  ( .D(n4456), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[952] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[24]  ( .D(n4491), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[984] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[24]  ( .D(n4526), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1016] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[24]  ( .D(n4568), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1048] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[24]  ( .D(n4629), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1080] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[24]  ( .D(n4664), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1112] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[24]  ( .D(n4699), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1144] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[24]  ( .D(n4734), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1176] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[24]  ( .D(n4769), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1208] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[24]  ( .D(n4804), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1240] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[24]  ( .D(n4839), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1272] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[24]  ( .D(n4874), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1304] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[24]  ( .D(n4909), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1336] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[24]  ( .D(n4944), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1368] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[24]  ( .D(n4979), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1400] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[24]  ( .D(n5014), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1432] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[24]  ( .D(n5049), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1464] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[24]  ( .D(n5084), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1496] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[24]  ( .D(n5119), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1528] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[24]  ( .D(n5161), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1560] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[24]  ( .D(n5221), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1592] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[24]  ( .D(n5257), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1624] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[24]  ( .D(n5292), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1656] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[24]  ( .D(n5327), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1688] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[24]  ( .D(n5362), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1720] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[24]  ( .D(n5397), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1752] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[24]  ( .D(n5432), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1784] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[24]  ( .D(n5467), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1816] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[24]  ( .D(n5502), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1848] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[24]  ( .D(n5537), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1880] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[24]  ( .D(n5572), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1912] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[24]  ( .D(n5611), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1944] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[24]  ( .D(n5648), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1976] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[24]  ( .D(n5685), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2008] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[24]  ( .D(n5722), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2040] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[24]  ( .D(n946), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2424] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[24]  ( .D(n991), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2456] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[24]  ( .D(n1028), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2488] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[24]  ( .D(n1065), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2520] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[24]  ( .D(n1102), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2552] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[24]  ( .D(n5759), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2072] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[24]  ( .D(n5798), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2104] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[24]  ( .D(n5834), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2136] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[24]  ( .D(n5870), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2168] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[24]  ( .D(n5906), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2200] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[24]  ( .D(n5942), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2232] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[24]  ( .D(n5978), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2264] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[24]  ( .D(n6014), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2296] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[24]  ( .D(n6051), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2328] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[24]  ( .D(n6087), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2360] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[24]  ( .D(n6121), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2392] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[8]  ( .D(n2215), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[8] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[8]  ( .D(n3351), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[8] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[8]  ( .D(n3399), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[40] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[8]  ( .D(n3437), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[72] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[8]  ( .D(n3475), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[104] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[8]  ( .D(n3513), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[136] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[8]  ( .D(n3551), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[168] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[8]  ( .D(n3589), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[200] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[8]  ( .D(n3627), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[232] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[8]  ( .D(n3665), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[264] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[8]  ( .D(n3702), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[296] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[8]  ( .D(n3739), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[328] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[8]  ( .D(n3776), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[360] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[8]  ( .D(n3811), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[392] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[8]  ( .D(n3846), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[424] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[8]  ( .D(n3881), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[456] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[8]  ( .D(n3939), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[488] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[8]  ( .D(n4007), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[520] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[8]  ( .D(n4052), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[552] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[8]  ( .D(n4087), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[584] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[8]  ( .D(n4122), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[616] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[8]  ( .D(n4157), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[648] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[8]  ( .D(n4192), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[680] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[8]  ( .D(n4227), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[712] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[8]  ( .D(n4262), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[744] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[8]  ( .D(n4297), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[776] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[8]  ( .D(n4332), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[808] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[8]  ( .D(n4367), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[840] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[8]  ( .D(n4402), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[872] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[8]  ( .D(n4437), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[904] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[8]  ( .D(n4472), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[936] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[8]  ( .D(n4507), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[968] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[8]  ( .D(n4542), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1000] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[8]  ( .D(n4600), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1032] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[8]  ( .D(n4645), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1064] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[8]  ( .D(n4680), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1096] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[8]  ( .D(n4715), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1128] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[8]  ( .D(n4750), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1160] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[8]  ( .D(n4785), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1192] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[8]  ( .D(n4820), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1224] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[8]  ( .D(n4855), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1256] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[8]  ( .D(n4890), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1288] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[8]  ( .D(n4925), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1320] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[8]  ( .D(n4960), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1352] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[8]  ( .D(n4995), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1384] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[8]  ( .D(n5030), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1416] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[8]  ( .D(n5065), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1448] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[8]  ( .D(n5100), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1480] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[8]  ( .D(n5135), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1512] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[8]  ( .D(n5193), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1544] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[8]  ( .D(n5237), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1576] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[8]  ( .D(n5273), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1608] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[8]  ( .D(n5308), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1640] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[8]  ( .D(n5343), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1672] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[8]  ( .D(n5378), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1704] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[8]  ( .D(n5413), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1736] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[8]  ( .D(n5448), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1768] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[8]  ( .D(n5483), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1800] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[8]  ( .D(n5518), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1832] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[8]  ( .D(n5553), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1864] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[8]  ( .D(n5588), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1896] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[8]  ( .D(n5627), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1928] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[8]  ( .D(n5664), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1960] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[8]  ( .D(n5701), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1992] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[8]  ( .D(n5738), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2024] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[8]  ( .D(n912), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2376] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[8]  ( .D(n969), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2408] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[8]  ( .D(n1007), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2440] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[8]  ( .D(n1044), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2472] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[8]  ( .D(n1081), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2504] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[8]  ( .D(n1118), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2536] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[8]  ( .D(n5775), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2056] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[8]  ( .D(n5814), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2088] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[8]  ( .D(n5850), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2120] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[8]  ( .D(n5886), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2152] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[8]  ( .D(n5922), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2184] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[8]  ( .D(n5958), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2216] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[8]  ( .D(n5994), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2248] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[8]  ( .D(n6030), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2280] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[8]  ( .D(n6067), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2312] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[8]  ( .D(n6103), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2344] ) );
  DFF_X1 \DataPath/REG_MEM_LDSTR_OUT/Q_reg[0]  ( .D(n2223), .CK(CLK), .QN(
        \DataPath/i_REG_LDSTR_OUT[0] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[0]  ( .D(n3367), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[0] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[0]  ( .D(n3407), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[32] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[0]  ( .D(n3445), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[64] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[0]  ( .D(n3483), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[96] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[0]  ( .D(n3521), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[128] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[0]  ( .D(n3559), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[160] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[0]  ( .D(n3597), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[192] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[0]  ( .D(n3635), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[224] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[0]  ( .D(n3673), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[256] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[0]  ( .D(n3710), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[288] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[0]  ( .D(n3747), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[320] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[0]  ( .D(n3784), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[352] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[0]  ( .D(n3819), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[384] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[0]  ( .D(n3854), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[416] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[0]  ( .D(n3889), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[448] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[0]  ( .D(n3955), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[480] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[0]  ( .D(n4023), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[512] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[0]  ( .D(n4060), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[544] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[0]  ( .D(n4095), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[576] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[0]  ( .D(n4130), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[608] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[0]  ( .D(n4165), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[640] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[0]  ( .D(n4200), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[672] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[0]  ( .D(n4235), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[704] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[0]  ( .D(n4270), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[736] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[0]  ( .D(n4305), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[768] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[0]  ( .D(n4340), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[800] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[0]  ( .D(n4375), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[832] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[0]  ( .D(n4410), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[864] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[0]  ( .D(n4445), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[896] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[0]  ( .D(n4480), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[928] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[0]  ( .D(n4515), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[960] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[0]  ( .D(n4550), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[992] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[0]  ( .D(n4616), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1024] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[0]  ( .D(n4653), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1056] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[0]  ( .D(n4688), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1088] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[0]  ( .D(n4723), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1120] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[0]  ( .D(n4758), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1152] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[0]  ( .D(n4793), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1184] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[0]  ( .D(n4828), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1216] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[0]  ( .D(n4863), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1248] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[0]  ( .D(n4898), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1280] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[0]  ( .D(n4933), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1312] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[0]  ( .D(n4968), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1344] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[0]  ( .D(n5003), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1376] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[0]  ( .D(n5038), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1408] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[0]  ( .D(n5073), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1440] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[0]  ( .D(n5108), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1472] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[0]  ( .D(n5143), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1504] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[0]  ( .D(n5209), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1536] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[0]  ( .D(n5245), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1568] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[0]  ( .D(n5281), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1600] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[0]  ( .D(n5316), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1632] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[0]  ( .D(n5351), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1664] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[0]  ( .D(n5386), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1696] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[0]  ( .D(n5421), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1728] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[0]  ( .D(n5456), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1760] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[0]  ( .D(n5491), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1792] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[0]  ( .D(n5526), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1824] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[0]  ( .D(n5561), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1856] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[0]  ( .D(n5596), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1888] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[0]  ( .D(n5635), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1920] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[0]  ( .D(n5672), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1952] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[0]  ( .D(n5709), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1984] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[0]  ( .D(n5746), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2016] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[0]  ( .D(n928), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2368] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[0]  ( .D(n977), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2400] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[0]  ( .D(n1015), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2432] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[0]  ( .D(n1052), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2464] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[0]  ( .D(n1089), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2496] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[0]  ( .D(n1126), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2528] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[0]  ( .D(n5822), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2080] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[0]  ( .D(n5858), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2112] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[0]  ( .D(n5894), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2144] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[0]  ( .D(n5930), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2176] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[0]  ( .D(n5966), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2208] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[0]  ( .D(n6002), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2240] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[0]  ( .D(n6038), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2272] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[0]  ( .D(n6075), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2304] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[0]  ( .D(n6111), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2336] ) );
  DFF_X1 \DataPath/RF/BLOCKi_8/Q_reg[7]  ( .D(n3353), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[7] ) );
  DFF_X1 \DataPath/RF/BLOCKi_9/Q_reg[7]  ( .D(n3400), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[39] ) );
  DFF_X1 \DataPath/RF/BLOCKi_10/Q_reg[7]  ( .D(n3438), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[71] ) );
  DFF_X1 \DataPath/RF/BLOCKi_11/Q_reg[7]  ( .D(n3476), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[103] ) );
  DFF_X1 \DataPath/RF/BLOCKi_12/Q_reg[7]  ( .D(n3514), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[135] ) );
  DFF_X1 \DataPath/RF/BLOCKi_13/Q_reg[7]  ( .D(n3552), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[167] ) );
  DFF_X1 \DataPath/RF/BLOCKi_14/Q_reg[7]  ( .D(n3590), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[199] ) );
  DFF_X1 \DataPath/RF/BLOCKi_15/Q_reg[7]  ( .D(n3628), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[231] ) );
  DFF_X1 \DataPath/RF/BLOCKi_16/Q_reg[7]  ( .D(n3666), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[263] ) );
  DFF_X1 \DataPath/RF/BLOCKi_17/Q_reg[7]  ( .D(n3703), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[295] ) );
  DFF_X1 \DataPath/RF/BLOCKi_18/Q_reg[7]  ( .D(n3740), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[327] ) );
  DFF_X1 \DataPath/RF/BLOCKi_19/Q_reg[7]  ( .D(n3777), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[359] ) );
  DFF_X1 \DataPath/RF/BLOCKi_20/Q_reg[7]  ( .D(n3812), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[391] ) );
  DFF_X1 \DataPath/RF/BLOCKi_21/Q_reg[7]  ( .D(n3847), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[423] ) );
  DFF_X1 \DataPath/RF/BLOCKi_22/Q_reg[7]  ( .D(n3882), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[455] ) );
  DFF_X1 \DataPath/RF/BLOCKi_23/Q_reg[7]  ( .D(n3941), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[487] ) );
  DFF_X1 \DataPath/RF/BLOCKi_24/Q_reg[7]  ( .D(n4009), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[519] ) );
  DFF_X1 \DataPath/RF/BLOCKi_25/Q_reg[7]  ( .D(n4053), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[551] ) );
  DFF_X1 \DataPath/RF/BLOCKi_26/Q_reg[7]  ( .D(n4088), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[583] ) );
  DFF_X1 \DataPath/RF/BLOCKi_27/Q_reg[7]  ( .D(n4123), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[615] ) );
  DFF_X1 \DataPath/RF/BLOCKi_28/Q_reg[7]  ( .D(n4158), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[647] ) );
  DFF_X1 \DataPath/RF/BLOCKi_29/Q_reg[7]  ( .D(n4193), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[679] ) );
  DFF_X1 \DataPath/RF/BLOCKi_30/Q_reg[7]  ( .D(n4228), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[711] ) );
  DFF_X1 \DataPath/RF/BLOCKi_31/Q_reg[7]  ( .D(n4263), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[743] ) );
  DFF_X1 \DataPath/RF/BLOCKi_32/Q_reg[7]  ( .D(n4298), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[775] ) );
  DFF_X1 \DataPath/RF/BLOCKi_33/Q_reg[7]  ( .D(n4333), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[807] ) );
  DFF_X1 \DataPath/RF/BLOCKi_34/Q_reg[7]  ( .D(n4368), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[839] ) );
  DFF_X1 \DataPath/RF/BLOCKi_35/Q_reg[7]  ( .D(n4403), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[871] ) );
  DFF_X1 \DataPath/RF/BLOCKi_36/Q_reg[7]  ( .D(n4438), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[903] ) );
  DFF_X1 \DataPath/RF/BLOCKi_37/Q_reg[7]  ( .D(n4473), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[935] ) );
  DFF_X1 \DataPath/RF/BLOCKi_38/Q_reg[7]  ( .D(n4508), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[967] ) );
  DFF_X1 \DataPath/RF/BLOCKi_39/Q_reg[7]  ( .D(n4543), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[999] ) );
  DFF_X1 \DataPath/RF/BLOCKi_40/Q_reg[7]  ( .D(n4602), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1031] ) );
  DFF_X1 \DataPath/RF/BLOCKi_41/Q_reg[7]  ( .D(n4646), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1063] ) );
  DFF_X1 \DataPath/RF/BLOCKi_42/Q_reg[7]  ( .D(n4681), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1095] ) );
  DFF_X1 \DataPath/RF/BLOCKi_43/Q_reg[7]  ( .D(n4716), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1127] ) );
  DFF_X1 \DataPath/RF/BLOCKi_44/Q_reg[7]  ( .D(n4751), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1159] ) );
  DFF_X1 \DataPath/RF/BLOCKi_45/Q_reg[7]  ( .D(n4786), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1191] ) );
  DFF_X1 \DataPath/RF/BLOCKi_46/Q_reg[7]  ( .D(n4821), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1223] ) );
  DFF_X1 \DataPath/RF/BLOCKi_47/Q_reg[7]  ( .D(n4856), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1255] ) );
  DFF_X1 \DataPath/RF/BLOCKi_48/Q_reg[7]  ( .D(n4891), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1287] ) );
  DFF_X1 \DataPath/RF/BLOCKi_49/Q_reg[7]  ( .D(n4926), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1319] ) );
  DFF_X1 \DataPath/RF/BLOCKi_50/Q_reg[7]  ( .D(n4961), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1351] ) );
  DFF_X1 \DataPath/RF/BLOCKi_51/Q_reg[7]  ( .D(n4996), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1383] ) );
  DFF_X1 \DataPath/RF/BLOCKi_52/Q_reg[7]  ( .D(n5031), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1415] ) );
  DFF_X1 \DataPath/RF/BLOCKi_53/Q_reg[7]  ( .D(n5066), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1447] ) );
  DFF_X1 \DataPath/RF/BLOCKi_54/Q_reg[7]  ( .D(n5101), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1479] ) );
  DFF_X1 \DataPath/RF/BLOCKi_55/Q_reg[7]  ( .D(n5136), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1511] ) );
  DFF_X1 \DataPath/RF/BLOCKi_56/Q_reg[7]  ( .D(n5195), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1543] ) );
  DFF_X1 \DataPath/RF/BLOCKi_57/Q_reg[7]  ( .D(n5238), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1575] ) );
  DFF_X1 \DataPath/RF/BLOCKi_58/Q_reg[7]  ( .D(n5274), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1607] ) );
  DFF_X1 \DataPath/RF/BLOCKi_59/Q_reg[7]  ( .D(n5309), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1639] ) );
  DFF_X1 \DataPath/RF/BLOCKi_60/Q_reg[7]  ( .D(n5344), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1671] ) );
  DFF_X1 \DataPath/RF/BLOCKi_61/Q_reg[7]  ( .D(n5379), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1703] ) );
  DFF_X1 \DataPath/RF/BLOCKi_62/Q_reg[7]  ( .D(n5414), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1735] ) );
  DFF_X1 \DataPath/RF/BLOCKi_63/Q_reg[7]  ( .D(n5449), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1767] ) );
  DFF_X1 \DataPath/RF/BLOCKi_64/Q_reg[7]  ( .D(n5484), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1799] ) );
  DFF_X1 \DataPath/RF/BLOCKi_65/Q_reg[7]  ( .D(n5519), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1831] ) );
  DFF_X1 \DataPath/RF/BLOCKi_66/Q_reg[7]  ( .D(n5554), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1863] ) );
  DFF_X1 \DataPath/RF/BLOCKi_67/Q_reg[7]  ( .D(n5589), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1895] ) );
  DFF_X1 \DataPath/RF/BLOCKi_68/Q_reg[7]  ( .D(n5628), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1927] ) );
  DFF_X1 \DataPath/RF/BLOCKi_69/Q_reg[7]  ( .D(n5665), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1959] ) );
  DFF_X1 \DataPath/RF/BLOCKi_70/Q_reg[7]  ( .D(n5702), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[1991] ) );
  DFF_X1 \DataPath/RF/BLOCKi_71/Q_reg[7]  ( .D(n5739), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2023] ) );
  DFF_X1 \DataPath/RF/BLOCKi_82/Q_reg[7]  ( .D(n914), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2375] ) );
  DFF_X1 \DataPath/RF/BLOCKi_83/Q_reg[7]  ( .D(n970), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2407] ) );
  DFF_X1 \DataPath/RF/BLOCKi_84/Q_reg[7]  ( .D(n1008), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2439] ) );
  DFF_X1 \DataPath/RF/BLOCKi_85/Q_reg[7]  ( .D(n1045), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2471] ) );
  DFF_X1 \DataPath/RF/BLOCKi_86/Q_reg[7]  ( .D(n1082), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2503] ) );
  DFF_X1 \DataPath/RF/BLOCKi_87/Q_reg[7]  ( .D(n1119), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2535] ) );
  DFF_X1 \DataPath/RF/BLOCKi_72/Q_reg[7]  ( .D(n5776), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2055] ) );
  DFF_X1 \DataPath/RF/BLOCKi_73/Q_reg[7]  ( .D(n5815), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2087] ) );
  DFF_X1 \DataPath/RF/BLOCKi_74/Q_reg[7]  ( .D(n5851), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2119] ) );
  DFF_X1 \DataPath/RF/BLOCKi_75/Q_reg[7]  ( .D(n5887), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2151] ) );
  DFF_X1 \DataPath/RF/BLOCKi_76/Q_reg[7]  ( .D(n5923), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2183] ) );
  DFF_X1 \DataPath/RF/BLOCKi_77/Q_reg[7]  ( .D(n5959), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2215] ) );
  DFF_X1 \DataPath/RF/BLOCKi_78/Q_reg[7]  ( .D(n5995), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2247] ) );
  DFF_X1 \DataPath/RF/BLOCKi_79/Q_reg[7]  ( .D(n6031), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2279] ) );
  DFF_X1 \DataPath/RF/BLOCKi_80/Q_reg[7]  ( .D(n6068), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2311] ) );
  DFF_X1 \DataPath/RF/BLOCKi_81/Q_reg[7]  ( .D(n6104), .CK(CLK), .QN(
        \DataPath/RF/bus_reg_dataout[2343] ) );
  DFFS_X1 \IR_reg[28]  ( .D(n7124), .CK(CLK), .SN(n8460), .Q(n8130), .QN(n167)
         );
  DFF_X1 \DataPath/RF/CWP/Q_reg[1]  ( .D(n7068), .CK(CLK), .Q(
        \DataPath/RF/c_win[1] ), .QN(n8274) );
  DFFS_X1 \IR_reg[30]  ( .D(n7122), .CK(CLK), .SN(n8460), .Q(n8279), .QN(n165)
         );
  DFF_X1 \CU_I/CW_MEM_reg[DRAM_RE]  ( .D(n7091), .CK(CLK), .Q(i_DATAMEM_RM), 
        .QN(n8277) );
  DFF_X1 \DataPath/RF/CWP/Q_reg[0]  ( .D(n7069), .CK(CLK), .Q(
        \DataPath/RF/c_win[0] ), .QN(n8273) );
  DFF_X1 \DataPath/RF/CWP/Q_reg[2]  ( .D(n7067), .CK(CLK), .Q(
        \DataPath/RF/c_win[2] ), .QN(n589) );
  DLL_X1 \CU_I/CW_ID_reg[MEM_EN]  ( .D(n10274), .GN(n2872), .Q(
        \CU_I/CW_ID[MEM_EN] ) );
  DLL_X1 \CU_I/CW_ID_reg[ID_EN]  ( .D(n10274), .GN(n2872), .Q(
        \CU_I/CW_ID[ID_EN] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[30]  ( .D(n8258), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[30] ) );
  DFFS_X1 \PC_reg[30]  ( .D(n8256), .CK(CLK), .SN(n8457), .Q(n10263), .QN(
        IRAM_ADDRESS[30]) );
  NOR2_X1 \intadd_1/U33  ( .A1(\intadd_1/B[1] ), .A2(\intadd_1/A[1] ), .ZN(
        \intadd_1/n25 ) );
  AOI21_X1 \intadd_1/U22  ( .B1(\intadd_1/n20 ), .B2(\intadd_1/n28 ), .A(
        \intadd_1/n21 ), .ZN(\intadd_1/n19 ) );
  NOR2_X1 \intadd_1/U10  ( .A1(\intadd_1/B[4] ), .A2(\intadd_1/A[4] ), .ZN(
        \intadd_1/n11 ) );
  NAND2_X1 \intadd_1/U11  ( .A1(\intadd_1/B[4] ), .A2(\intadd_1/A[4] ), .ZN(
        \intadd_1/n12 ) );
  OAI21_X1 \intadd_1/U7  ( .B1(\intadd_1/n17 ), .B2(\intadd_1/n11 ), .A(
        \intadd_1/n12 ), .ZN(\intadd_1/n10 ) );
  NOR2_X1 \intadd_0/U30  ( .A1(\intadd_0/B[2] ), .A2(n8127), .ZN(
        \intadd_0/n25 ) );
  NOR2_X1 \intadd_0/U24  ( .A1(\intadd_0/B[3] ), .A2(n8126), .ZN(
        \intadd_0/n22 ) );
  NAND2_X1 \intadd_0/U36  ( .A1(n8122), .A2(n8091), .ZN(\intadd_0/n30 ) );
  NOR2_X1 \intadd_0/U16  ( .A1(n8124), .A2(\intadd_0/n30 ), .ZN(\intadd_0/n16 ) );
  NAND2_X1 \intadd_0/U51  ( .A1(\intadd_0/B[0] ), .A2(\intadd_0/A[0] ), .ZN(
        \intadd_0/n40 ) );
  NAND2_X1 \intadd_0/U43  ( .A1(\intadd_0/B[1] ), .A2(n8128), .ZN(
        \intadd_0/n35 ) );
  AOI21_X1 \intadd_0/U37  ( .B1(n8091), .B2(\intadd_0/n38 ), .A(\intadd_0/n33 ), .ZN(\intadd_0/n31 ) );
  NAND2_X1 \intadd_0/U31  ( .A1(\intadd_0/B[2] ), .A2(n8127), .ZN(
        \intadd_0/n26 ) );
  NAND2_X1 \intadd_0/U25  ( .A1(\intadd_0/B[3] ), .A2(n8126), .ZN(
        \intadd_0/n23 ) );
  OAI21_X1 \intadd_0/U21  ( .B1(\intadd_0/n22 ), .B2(\intadd_0/n26 ), .A(
        \intadd_0/n23 ), .ZN(\intadd_0/n21 ) );
  OAI21_X1 \intadd_0/U17  ( .B1(n8124), .B2(\intadd_0/n31 ), .A(\intadd_0/n19 ), .ZN(\intadd_0/n17 ) );
  NAND2_X1 \intadd_0/U13  ( .A1(\intadd_0/B[4] ), .A2(n8125), .ZN(
        \intadd_0/n14 ) );
  NAND2_X1 \intadd_2/U26  ( .A1(n8123), .A2(n8092), .ZN(\intadd_2/n22 ) );
  NOR2_X1 \intadd_2/U20  ( .A1(\intadd_2/B[2] ), .A2(IRAM_ADDRESS[23]), .ZN(
        \intadd_2/n17 ) );
  NOR2_X1 \intadd_2/U16  ( .A1(\intadd_2/n22 ), .A2(\intadd_2/n17 ), .ZN(
        \intadd_2/n15 ) );
  NAND2_X1 \intadd_2/U41  ( .A1(\intadd_2/B[0] ), .A2(IRAM_ADDRESS[21]), .ZN(
        \intadd_2/n32 ) );
  NAND2_X1 \intadd_2/U33  ( .A1(\intadd_2/B[1] ), .A2(IRAM_ADDRESS[22]), .ZN(
        \intadd_2/n27 ) );
  AOI21_X1 \intadd_2/U27  ( .B1(n8092), .B2(\intadd_2/n30 ), .A(\intadd_2/n25 ), .ZN(\intadd_2/n23 ) );
  NAND2_X1 \intadd_2/U21  ( .A1(\intadd_2/B[2] ), .A2(IRAM_ADDRESS[23]), .ZN(
        \intadd_2/n18 ) );
  OAI21_X1 \intadd_2/U17  ( .B1(\intadd_2/n23 ), .B2(\intadd_2/n17 ), .A(
        \intadd_2/n18 ), .ZN(\intadd_2/n16 ) );
  NAND2_X1 \intadd_2/U13  ( .A1(\intadd_2/B[3] ), .A2(IRAM_ADDRESS[24]), .ZN(
        \intadd_2/n13 ) );
  AOI21_X1 \intadd_2/U7  ( .B1(\intadd_2/n16 ), .B2(n8120), .A(\intadd_2/n11 ), 
        .ZN(\intadd_2/n9 ) );
  NAND2_X1 \intadd_2/U10  ( .A1(n8120), .A2(\intadd_2/n13 ), .ZN(\intadd_2/n1 ) );
  XOR2_X1 \intadd_2/U2  ( .A(\intadd_2/n14 ), .B(\intadd_2/n1 ), .Z(
        \intadd_2/SUM[3] ) );
  NAND2_X1 \intadd_2/U30  ( .A1(n8092), .A2(\intadd_2/n27 ), .ZN(\intadd_2/n3 ) );
  XOR2_X1 \intadd_2/U22  ( .A(\intadd_2/n28 ), .B(\intadd_2/n3 ), .Z(
        \intadd_2/SUM[1] ) );
  NAND2_X1 \intadd_2/U38  ( .A1(n8123), .A2(\intadd_2/n32 ), .ZN(\intadd_2/n4 ) );
  OAI21_X1 \intadd_0/U27  ( .B1(\intadd_0/n27 ), .B2(\intadd_0/n25 ), .A(
        \intadd_0/n26 ), .ZN(\intadd_0/n24 ) );
  NAND2_X1 \intadd_0/U22  ( .A1(\intadd_0/n44 ), .A2(\intadd_0/n23 ), .ZN(
        \intadd_0/n2 ) );
  XNOR2_X1 \intadd_0/U14  ( .A(\intadd_0/n24 ), .B(\intadd_0/n2 ), .ZN(
        \intadd_0/SUM[3] ) );
  NAND2_X1 \intadd_0/U28  ( .A1(\intadd_0/n45 ), .A2(\intadd_0/n26 ), .ZN(
        \intadd_0/n3 ) );
  XOR2_X1 \intadd_0/U26  ( .A(\intadd_0/n27 ), .B(\intadd_0/n3 ), .Z(
        \intadd_0/SUM[2] ) );
  NAND2_X1 \intadd_0/U40  ( .A1(n8091), .A2(\intadd_0/n35 ), .ZN(\intadd_0/n4 ) );
  XOR2_X1 \intadd_0/U32  ( .A(\intadd_0/n36 ), .B(\intadd_0/n4 ), .Z(
        \intadd_0/SUM[1] ) );
  NAND2_X1 \intadd_0/U10  ( .A1(n8093), .A2(\intadd_0/n14 ), .ZN(\intadd_0/n1 ) );
  XOR2_X1 \intadd_0/U2  ( .A(\intadd_0/n15 ), .B(\intadd_0/n1 ), .Z(
        \intadd_0/SUM[4] ) );
  NAND2_X1 \intadd_1/U31  ( .A1(\intadd_1/n35 ), .A2(\intadd_1/n26 ), .ZN(
        \intadd_1/n4 ) );
  XOR2_X1 \intadd_1/U29  ( .A(\intadd_1/n27 ), .B(\intadd_1/n4 ), .Z(
        \intadd_1/SUM[1] ) );
  XNOR2_X1 \intadd_1/U35  ( .A(\intadd_1/n5 ), .B(\intadd_1/CI ), .ZN(
        \intadd_1/SUM[0] ) );
  NAND2_X1 \intadd_0/U48  ( .A1(n8122), .A2(\intadd_0/n40 ), .ZN(\intadd_0/n5 ) );
  OAI21_X1 \intadd_1/U30  ( .B1(\intadd_1/n27 ), .B2(n7939), .A(\intadd_1/n26 ), .ZN(\intadd_1/n24 ) );
  NAND2_X1 \intadd_1/U25  ( .A1(\intadd_1/n34 ), .A2(\intadd_1/n23 ), .ZN(
        \intadd_1/n3 ) );
  XNOR2_X1 \intadd_1/U20  ( .A(\intadd_1/n24 ), .B(\intadd_1/n3 ), .ZN(
        \intadd_1/SUM[2] ) );
  AOI21_X1 \intadd_1/U13  ( .B1(\intadd_1/n18 ), .B2(\intadd_1/n33 ), .A(
        \intadd_1/n15 ), .ZN(\intadd_1/n13 ) );
  NAND2_X1 \intadd_1/U8  ( .A1(\intadd_1/n32 ), .A2(\intadd_1/n12 ), .ZN(
        \intadd_1/n1 ) );
  XOR2_X1 \intadd_1/U2  ( .A(\intadd_1/n13 ), .B(\intadd_1/n1 ), .Z(
        \intadd_1/SUM[4] ) );
  NAND2_X1 \intadd_1/U16  ( .A1(\intadd_1/n33 ), .A2(n7719), .ZN(\intadd_1/n2 ) );
  XNOR2_X1 \intadd_1/U12  ( .A(\intadd_1/n18 ), .B(\intadd_1/n2 ), .ZN(
        \intadd_1/SUM[3] ) );
  FA_X1 \DP_OP_1091J1_126_6973/U31  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[2] ), .CI(\DP_OP_1091J1_126_6973/n37 ), 
        .CO(\DP_OP_1091J1_126_6973/n30 ), .S(\C620/DATA2_2 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U30  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[3] ), .CI(\DP_OP_1091J1_126_6973/n30 ), 
        .CO(\DP_OP_1091J1_126_6973/n29 ), .S(\C620/DATA2_3 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U27  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[6] ), .CI(\DP_OP_1091J1_126_6973/n27 ), 
        .CO(\DP_OP_1091J1_126_6973/n26 ), .S(\C620/DATA2_6 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U26  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[7] ), .CI(\DP_OP_1091J1_126_6973/n26 ), 
        .CO(\DP_OP_1091J1_126_6973/n25 ), .S(\C620/DATA2_7 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U25  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[8] ), .CI(\DP_OP_1091J1_126_6973/n25 ), 
        .CO(\DP_OP_1091J1_126_6973/n24 ), .S(\C620/DATA2_8 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U24  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[9] ), .CI(\DP_OP_1091J1_126_6973/n24 ), 
        .CO(\DP_OP_1091J1_126_6973/n23 ), .S(\C620/DATA2_9 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U23  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[10] ), .CI(\DP_OP_1091J1_126_6973/n23 ), 
        .CO(\DP_OP_1091J1_126_6973/n22 ), .S(\C620/DATA2_10 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U10  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[23] ), .CI(\DP_OP_1091J1_126_6973/n10 ), 
        .CO(\DP_OP_1091J1_126_6973/n9 ), .S(\C620/DATA2_23 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U9  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[24] ), .CI(\DP_OP_1091J1_126_6973/n9 ), 
        .CO(\DP_OP_1091J1_126_6973/n8 ), .S(\C620/DATA2_24 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U8  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[25] ), .CI(\DP_OP_1091J1_126_6973/n8 ), 
        .CO(\DP_OP_1091J1_126_6973/n7 ), .S(\C620/DATA2_25 ) );
  FA_X1 \DP_OP_1091J1_126_6973/U7  ( .A(n7776), .B(
        \DataPath/WRF_CUhw/curr_addr[26] ), .CI(\DP_OP_1091J1_126_6973/n7 ), 
        .CO(\DP_OP_1091J1_126_6973/n6 ), .S(\C620/DATA2_26 ) );
  XOR2_X1 \DP_OP_751_130_6421/U167  ( .A(\DP_OP_751_130_6421/n20 ), .B(
        \DP_OP_751_130_6421/n140 ), .Z(\DataPath/ALUhw/i_Q_EXTENDED[38] ) );
  NAND2_X1 \DP_OP_751_130_6421/U169  ( .A1(\DP_OP_751_130_6421/n183 ), .A2(
        \DP_OP_751_130_6421/n139 ), .ZN(\DP_OP_751_130_6421/n20 ) );
  NAND2_X1 \DP_OP_751_130_6421/U155  ( .A1(\DP_OP_751_130_6421/n181 ), .A2(
        \DP_OP_751_130_6421/n131 ), .ZN(\DP_OP_751_130_6421/n18 ) );
  NAND2_X1 \DP_OP_751_130_6421/U149  ( .A1(n8065), .A2(
        \DP_OP_751_130_6421/n128 ), .ZN(\DP_OP_751_130_6421/n17 ) );
  XOR2_X1 \DP_OP_751_130_6421/U181  ( .A(\DP_OP_751_130_6421/n22 ), .B(
        \DP_OP_751_130_6421/n148 ), .Z(\DataPath/ALUhw/i_Q_EXTENDED[36] ) );
  NAND2_X1 \DP_OP_751_130_6421/U183  ( .A1(\DP_OP_751_130_6421/n185 ), .A2(
        \DP_OP_751_130_6421/n147 ), .ZN(\DP_OP_751_130_6421/n22 ) );
  XNOR2_X1 \DP_OP_751_130_6421/U136  ( .A(\DP_OP_751_130_6421/n16 ), .B(
        \DP_OP_751_130_6421/n123 ), .ZN(\DataPath/ALUhw/i_Q_EXTENDED[42] ) );
  NAND2_X1 \DP_OP_751_130_6421/U140  ( .A1(n8071), .A2(
        \DP_OP_751_130_6421/n122 ), .ZN(\DP_OP_751_130_6421/n16 ) );
  NAND2_X1 \DP_OP_751_130_6421/U118  ( .A1(\DP_OP_751_130_6421/n176 ), .A2(
        \DP_OP_751_130_6421/n109 ), .ZN(\DP_OP_751_130_6421/n13 ) );
  XOR2_X1 \DP_OP_751_130_6421/U95  ( .A(\DP_OP_751_130_6421/n10 ), .B(
        \DP_OP_751_130_6421/n98 ), .Z(\DataPath/ALUhw/i_Q_EXTENDED[48] ) );
  NAND2_X1 \DP_OP_751_130_6421/U97  ( .A1(\DP_OP_751_130_6421/n173 ), .A2(
        \DP_OP_751_130_6421/n97 ), .ZN(\DP_OP_751_130_6421/n10 ) );
  XNOR2_X1 \DP_OP_751_130_6421/U87  ( .A(\DP_OP_751_130_6421/n9 ), .B(
        \DP_OP_751_130_6421/n95 ), .ZN(\DataPath/ALUhw/i_Q_EXTENDED[49] ) );
  NAND2_X1 \DP_OP_751_130_6421/U91  ( .A1(n8069), .A2(\DP_OP_751_130_6421/n94 ), .ZN(\DP_OP_751_130_6421/n9 ) );
  XOR2_X1 \DP_OP_751_130_6421/U81  ( .A(\DP_OP_751_130_6421/n8 ), .B(n7643), 
        .Z(\DataPath/ALUhw/i_Q_EXTENDED[50] ) );
  NAND2_X1 \DP_OP_751_130_6421/U83  ( .A1(\DP_OP_751_130_6421/n171 ), .A2(
        \DP_OP_751_130_6421/n89 ), .ZN(\DP_OP_751_130_6421/n8 ) );
  NAND2_X1 \DP_OP_751_130_6421/U77  ( .A1(n8068), .A2(\DP_OP_751_130_6421/n86 ), .ZN(\DP_OP_751_130_6421/n7 ) );
  NAND2_X1 \DP_OP_751_130_6421/U69  ( .A1(\DP_OP_751_130_6421/n169 ), .A2(
        \DP_OP_751_130_6421/n81 ), .ZN(\DP_OP_751_130_6421/n6 ) );
  NAND2_X1 \DP_OP_751_130_6421/U63  ( .A1(n8064), .A2(\DP_OP_751_130_6421/n78 ), .ZN(\DP_OP_751_130_6421/n5 ) );
  XNOR2_X1 \DP_OP_751_130_6421/U48  ( .A(\DP_OP_751_130_6421/n4 ), .B(n7629), 
        .ZN(\DataPath/ALUhw/i_Q_EXTENDED[56] ) );
  NAND2_X1 \DP_OP_751_130_6421/U52  ( .A1(n8070), .A2(\DP_OP_751_130_6421/n71 ), .ZN(\DP_OP_751_130_6421/n4 ) );
  NAND2_X1 \DP_OP_751_130_6421/U55  ( .A1(\DP_OP_751_130_6421/n562 ), .A2(
        \DP_OP_751_130_6421/n660 ), .ZN(\DP_OP_751_130_6421/n71 ) );
  NAND2_X1 \DP_OP_751_130_6421/U72  ( .A1(\DP_OP_751_130_6421/n766 ), .A2(
        \DP_OP_751_130_6421/n864 ), .ZN(\DP_OP_751_130_6421/n81 ) );
  NAND2_X1 \DP_OP_751_130_6421/U80  ( .A1(\DP_OP_751_130_6421/n866 ), .A2(
        \DP_OP_751_130_6421/n867 ), .ZN(\DP_OP_751_130_6421/n86 ) );
  NAND2_X1 \DP_OP_751_130_6421/U86  ( .A1(\DP_OP_751_130_6421/n868 ), .A2(
        \DP_OP_751_130_6421/n966 ), .ZN(\DP_OP_751_130_6421/n89 ) );
  NOR2_X1 \DP_OP_751_130_6421/U85  ( .A1(\DP_OP_751_130_6421/n868 ), .A2(
        \DP_OP_751_130_6421/n966 ), .ZN(\DP_OP_751_130_6421/n88 ) );
  XOR2_X1 \DP_OP_751_130_6421/U703  ( .A(\DataPath/ALUhw/MULT/mux_out[9][18] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n902 ) );
  NAND2_X1 \DP_OP_751_130_6421/U94  ( .A1(\DP_OP_751_130_6421/n968 ), .A2(
        \DP_OP_751_130_6421/n969 ), .ZN(\DP_OP_751_130_6421/n94 ) );
  XOR2_X1 \DP_OP_751_130_6421/U772  ( .A(\DataPath/ALUhw/MULT/mux_out[8][17] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n1003 ) );
  NAND2_X1 \DP_OP_751_130_6421/U100  ( .A1(\DP_OP_751_130_6421/n970 ), .A2(
        \DP_OP_751_130_6421/n1068 ), .ZN(\DP_OP_751_130_6421/n97 ) );
  NOR2_X1 \DP_OP_751_130_6421/U99  ( .A1(\DP_OP_751_130_6421/n970 ), .A2(
        \DP_OP_751_130_6421/n1068 ), .ZN(\DP_OP_751_130_6421/n96 ) );
  XOR2_X1 \DP_OP_751_130_6421/U841  ( .A(\DataPath/ALUhw/MULT/mux_out[7][16] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1104 ) );
  XOR2_X1 \DP_OP_751_130_6421/U773  ( .A(\DataPath/ALUhw/MULT/mux_out[8][16] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n1004 ) );
  NAND2_X1 \DP_OP_751_130_6421/U107  ( .A1(\DP_OP_751_130_6421/n1070 ), .A2(
        \DP_OP_751_130_6421/n1071 ), .ZN(\DP_OP_751_130_6421/n101 ) );
  NAND2_X1 \DP_OP_751_130_6421/U115  ( .A1(\DP_OP_751_130_6421/n1072 ), .A2(
        \DP_OP_751_130_6421/n1170 ), .ZN(\DP_OP_751_130_6421/n106 ) );
  NAND2_X1 \DP_OP_751_130_6421/U121  ( .A1(\DP_OP_751_130_6421/n1172 ), .A2(
        \DP_OP_751_130_6421/n1173 ), .ZN(\DP_OP_751_130_6421/n109 ) );
  NAND2_X1 \DP_OP_751_130_6421/U129  ( .A1(\DP_OP_751_130_6421/n1174 ), .A2(
        \DP_OP_751_130_6421/n1272 ), .ZN(\DP_OP_751_130_6421/n114 ) );
  NAND2_X1 \DP_OP_751_130_6421/U135  ( .A1(\DP_OP_751_130_6421/n1274 ), .A2(
        \DP_OP_751_130_6421/n1275 ), .ZN(\DP_OP_751_130_6421/n117 ) );
  AOI21_X1 \DP_OP_751_130_6421/U137  ( .B1(n8071), .B2(
        \DP_OP_751_130_6421/n123 ), .A(\DP_OP_751_130_6421/n120 ), .ZN(
        \DP_OP_751_130_6421/n118 ) );
  NAND2_X1 \DP_OP_751_130_6421/U143  ( .A1(\DP_OP_751_130_6421/n1276 ), .A2(
        \DP_OP_751_130_6421/n1374 ), .ZN(\DP_OP_751_130_6421/n122 ) );
  NAND2_X1 \DP_OP_751_130_6421/U152  ( .A1(\DP_OP_751_130_6421/n1376 ), .A2(
        \DP_OP_751_130_6421/n1377 ), .ZN(\DP_OP_751_130_6421/n128 ) );
  NAND2_X1 \DP_OP_751_130_6421/U158  ( .A1(\DP_OP_751_130_6421/n1378 ), .A2(
        \DP_OP_751_130_6421/n1476 ), .ZN(\DP_OP_751_130_6421/n131 ) );
  AOI21_X1 \DP_OP_751_130_6421/U160  ( .B1(n8072), .B2(
        \DP_OP_751_130_6421/n137 ), .A(\DP_OP_751_130_6421/n134 ), .ZN(
        \DP_OP_751_130_6421/n132 ) );
  NAND2_X1 \DP_OP_751_130_6421/U166  ( .A1(\DP_OP_751_130_6421/n1478 ), .A2(
        \DP_OP_751_130_6421/n1479 ), .ZN(\DP_OP_751_130_6421/n136 ) );
  OAI21_X1 \DP_OP_751_130_6421/U168  ( .B1(\DP_OP_751_130_6421/n138 ), .B2(
        \DP_OP_751_130_6421/n140 ), .A(\DP_OP_751_130_6421/n139 ), .ZN(
        \DP_OP_751_130_6421/n137 ) );
  NAND2_X1 \DP_OP_751_130_6421/U172  ( .A1(\DP_OP_751_130_6421/n1480 ), .A2(
        \DP_OP_751_130_6421/n1578 ), .ZN(\DP_OP_751_130_6421/n139 ) );
  AOI21_X1 \DP_OP_751_130_6421/U174  ( .B1(\DP_OP_751_130_6421/n145 ), .B2(
        n8073), .A(\DP_OP_751_130_6421/n142 ), .ZN(\DP_OP_751_130_6421/n140 )
         );
  NAND2_X1 \DP_OP_751_130_6421/U180  ( .A1(\DP_OP_751_130_6421/n1580 ), .A2(
        \DP_OP_751_130_6421/n1581 ), .ZN(\DP_OP_751_130_6421/n144 ) );
  OAI21_X1 \DP_OP_751_130_6421/U182  ( .B1(\DP_OP_751_130_6421/n146 ), .B2(
        \DP_OP_751_130_6421/n148 ), .A(\DP_OP_751_130_6421/n147 ), .ZN(
        \DP_OP_751_130_6421/n145 ) );
  NAND2_X1 \DP_OP_751_130_6421/U186  ( .A1(\DP_OP_751_130_6421/n1582 ), .A2(
        \DP_OP_751_130_6421/n1680 ), .ZN(\DP_OP_751_130_6421/n147 ) );
  AOI21_X1 \DP_OP_751_130_6421/U188  ( .B1(\DP_OP_751_130_6421/n151 ), .B2(
        \DP_OP_751_130_6421/n153 ), .A(\DP_OP_751_130_6421/n150 ), .ZN(
        \DP_OP_751_130_6421/n148 ) );
  NAND2_X1 \DP_OP_751_130_6421/U194  ( .A1(\DP_OP_751_130_6421/n1682 ), .A2(
        \DP_OP_751_130_6421/n1683 ), .ZN(\DP_OP_751_130_6421/n152 ) );
  OAI21_X1 \DP_OP_751_130_6421/U196  ( .B1(\DP_OP_751_130_6421/n154 ), .B2(
        \DP_OP_751_130_6421/n158 ), .A(\DP_OP_751_130_6421/n155 ), .ZN(
        \DP_OP_751_130_6421/n153 ) );
  NAND2_X1 \DP_OP_751_130_6421/U200  ( .A1(\DP_OP_751_130_6421/n1684 ), .A2(
        \DP_OP_751_130_6421/n1685 ), .ZN(\DP_OP_751_130_6421/n155 ) );
  NAND2_X1 \DP_OP_751_130_6421/U204  ( .A1(\DP_OP_751_130_6421/n159 ), .A2(
        \DP_OP_751_130_6421/n161 ), .ZN(\DP_OP_751_130_6421/n158 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1299  ( .A(n7766), .B(
        \DataPath/ALUhw/MULT/mux_out[0][0] ), .S(n8060), .Z(
        \DP_OP_751_130_6421/n1753 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1265  ( .A(\DataPath/ALUhw/MULT/mux_out[1][2] ), 
        .B(n7690), .Z(\DP_OP_751_130_6421/n1685 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1264  ( .A(\DataPath/ALUhw/MULT/mux_out[1][3] ), 
        .B(n7690), .Z(\DP_OP_751_130_6421/n1683 ) );
  NOR2_X1 \DP_OP_751_130_6421/U185  ( .A1(\DP_OP_751_130_6421/n1582 ), .A2(
        \DP_OP_751_130_6421/n1680 ), .ZN(\DP_OP_751_130_6421/n146 ) );
  NOR2_X1 \DP_OP_751_130_6421/U171  ( .A1(\DP_OP_751_130_6421/n1480 ), .A2(
        \DP_OP_751_130_6421/n1578 ), .ZN(\DP_OP_751_130_6421/n138 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1192  ( .A(\DataPath/ALUhw/MULT/mux_out[2][5] ), 
        .B(n8057), .Z(\DP_OP_751_130_6421/n1615 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1123  ( .A(\DataPath/ALUhw/MULT/mux_out[3][6] ), 
        .B(\DP_OP_751_130_6421/n1515 ), .Z(\DP_OP_751_130_6421/n1514 ) );
  NOR2_X1 \DP_OP_751_130_6421/U157  ( .A1(\DP_OP_751_130_6421/n1378 ), .A2(
        \DP_OP_751_130_6421/n1476 ), .ZN(\DP_OP_751_130_6421/n130 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1122  ( .A(\DataPath/ALUhw/MULT/mux_out[3][7] ), 
        .B(n8056), .Z(\DP_OP_751_130_6421/n1513 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1191  ( .A(\DataPath/ALUhw/MULT/mux_out[2][6] ), 
        .B(n8057), .Z(\DP_OP_751_130_6421/n1614 ) );
  NOR2_X1 \DP_OP_751_130_6421/U134  ( .A1(\DP_OP_751_130_6421/n1274 ), .A2(
        \DP_OP_751_130_6421/n1275 ), .ZN(\DP_OP_751_130_6421/n116 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1052  ( .A(\DataPath/ALUhw/MULT/mux_out[4][9] ), 
        .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1411 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1121  ( .A(\DataPath/ALUhw/MULT/mux_out[3][8] ), 
        .B(n8056), .Z(\DP_OP_751_130_6421/n1512 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1190  ( .A(\DataPath/ALUhw/MULT/mux_out[2][7] ), 
        .B(n8057), .Z(\DP_OP_751_130_6421/n1613 ) );
  XOR2_X1 \DP_OP_751_130_6421/U983  ( .A(\DataPath/ALUhw/MULT/mux_out[5][10] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1310 ) );
  NOR2_X1 \DP_OP_751_130_6421/U120  ( .A1(\DP_OP_751_130_6421/n1172 ), .A2(
        \DP_OP_751_130_6421/n1173 ), .ZN(\DP_OP_751_130_6421/n108 ) );
  XOR2_X1 \DP_OP_751_130_6421/U982  ( .A(\DataPath/ALUhw/MULT/mux_out[5][11] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1309 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1051  ( .A(\DataPath/ALUhw/MULT/mux_out[4][10] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1410 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1120  ( .A(\DataPath/ALUhw/MULT/mux_out[3][9] ), 
        .B(n8056), .Z(\DP_OP_751_130_6421/n1511 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1189  ( .A(\DataPath/ALUhw/MULT/mux_out[2][8] ), 
        .B(n8057), .Z(\DP_OP_751_130_6421/n1612 ) );
  XOR2_X1 \DP_OP_751_130_6421/U913  ( .A(\DataPath/ALUhw/MULT/mux_out[6][12] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1208 ) );
  NOR2_X1 \DP_OP_751_130_6421/U106  ( .A1(\DP_OP_751_130_6421/n1070 ), .A2(
        \DP_OP_751_130_6421/n1071 ), .ZN(\DP_OP_751_130_6421/n100 ) );
  XOR2_X1 \DP_OP_751_130_6421/U912  ( .A(\DataPath/ALUhw/MULT/mux_out[6][13] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1207 ) );
  XOR2_X1 \DP_OP_751_130_6421/U981  ( .A(\DataPath/ALUhw/MULT/mux_out[5][12] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1308 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1050  ( .A(\DataPath/ALUhw/MULT/mux_out[4][11] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1409 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1119  ( .A(\DataPath/ALUhw/MULT/mux_out[3][10] ), .B(\DP_OP_751_130_6421/n1515 ), .Z(\DP_OP_751_130_6421/n1510 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1188  ( .A(\DataPath/ALUhw/MULT/mux_out[2][9] ), 
        .B(n8057), .Z(\DP_OP_751_130_6421/n1611 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1291  ( .A(\DP_OP_751_130_6421/n1779 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][8] ), .S(n8060), .Z(
        \DP_OP_751_130_6421/n1744 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1259  ( .A(\DataPath/ALUhw/MULT/mux_out[1][8] ), 
        .B(n7690), .Z(\DP_OP_751_130_6421/n1714 ) );
  XOR2_X1 \DP_OP_751_130_6421/U843  ( .A(\DataPath/ALUhw/MULT/mux_out[7][14] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1106 ) );
  XOR2_X1 \DP_OP_751_130_6421/U910  ( .A(\DataPath/ALUhw/MULT/mux_out[6][15] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1205 ) );
  XOR2_X1 \DP_OP_751_130_6421/U842  ( .A(\DataPath/ALUhw/MULT/mux_out[7][15] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1105 ) );
  XOR2_X1 \DP_OP_751_130_6421/U979  ( .A(\DataPath/ALUhw/MULT/mux_out[5][14] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1306 ) );
  XOR2_X1 \DP_OP_751_130_6421/U911  ( .A(\DataPath/ALUhw/MULT/mux_out[6][14] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1206 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1048  ( .A(\DataPath/ALUhw/MULT/mux_out[4][13] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1407 ) );
  XOR2_X1 \DP_OP_751_130_6421/U980  ( .A(\DataPath/ALUhw/MULT/mux_out[5][13] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1307 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1117  ( .A(\DataPath/ALUhw/MULT/mux_out[3][12] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1508 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1049  ( .A(\DataPath/ALUhw/MULT/mux_out[4][12] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1408 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1186  ( .A(\DataPath/ALUhw/MULT/mux_out[2][11] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1609 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1118  ( .A(\DataPath/ALUhw/MULT/mux_out[3][11] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1509 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1289  ( .A(\DP_OP_751_130_6421/n1777 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][10] ), .S(n7974), .Z(
        \DP_OP_751_130_6421/n1742 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1257  ( .A(\DataPath/ALUhw/MULT/mux_out[1][10] ), .B(n8059), .Z(\DP_OP_751_130_6421/n1712 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1187  ( .A(\DataPath/ALUhw/MULT/mux_out[2][10] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1610 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1290  ( .A(\DP_OP_751_130_6421/n1778 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][9] ), .S(n8060), .Z(
        \DP_OP_751_130_6421/n1743 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1258  ( .A(\DataPath/ALUhw/MULT/mux_out[1][9] ), 
        .B(n7690), .Z(\DP_OP_751_130_6421/n1713 ) );
  NOR2_X1 \DP_OP_751_130_6421/U71  ( .A1(\DP_OP_751_130_6421/n766 ), .A2(
        \DP_OP_751_130_6421/n864 ), .ZN(\DP_OP_751_130_6421/n80 ) );
  XOR2_X1 \DP_OP_751_130_6421/U702  ( .A(\DataPath/ALUhw/MULT/mux_out[9][19] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n901 ) );
  XOR2_X1 \DP_OP_751_130_6421/U771  ( .A(\DataPath/ALUhw/MULT/mux_out[8][18] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n1002 ) );
  XOR2_X1 \DP_OP_751_130_6421/U840  ( .A(\DataPath/ALUhw/MULT/mux_out[7][17] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1103 ) );
  XOR2_X1 \DP_OP_751_130_6421/U909  ( .A(\DataPath/ALUhw/MULT/mux_out[6][16] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1204 ) );
  XOR2_X1 \DP_OP_751_130_6421/U978  ( .A(\DataPath/ALUhw/MULT/mux_out[5][15] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1305 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1047  ( .A(\DataPath/ALUhw/MULT/mux_out[4][14] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1406 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1116  ( .A(\DataPath/ALUhw/MULT/mux_out[3][13] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1507 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1185  ( .A(\DataPath/ALUhw/MULT/mux_out[2][12] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1608 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1288  ( .A(\DP_OP_751_130_6421/n1776 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][11] ), .S(n8060), .Z(
        \DP_OP_751_130_6421/n1741 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1256  ( .A(\DataPath/ALUhw/MULT/mux_out[1][11] ), .B(n7690), .Z(\DP_OP_751_130_6421/n1711 ) );
  XOR2_X1 \DP_OP_751_130_6421/U633  ( .A(\DataPath/ALUhw/MULT/mux_out[10][20] ), .B(n8062), .Z(\DP_OP_751_130_6421/n800 ) );
  XOR2_X1 \DP_OP_751_130_6421/U632  ( .A(\DataPath/ALUhw/MULT/mux_out[10][21] ), .B(n8062), .Z(\DP_OP_751_130_6421/n799 ) );
  XOR2_X1 \DP_OP_751_130_6421/U701  ( .A(\DataPath/ALUhw/MULT/mux_out[9][20] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n900 ) );
  XOR2_X1 \DP_OP_751_130_6421/U770  ( .A(\DataPath/ALUhw/MULT/mux_out[8][19] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n1001 ) );
  XOR2_X1 \DP_OP_751_130_6421/U839  ( .A(\DataPath/ALUhw/MULT/mux_out[7][18] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1102 ) );
  XOR2_X1 \DP_OP_751_130_6421/U908  ( .A(\DataPath/ALUhw/MULT/mux_out[6][17] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1203 ) );
  XOR2_X1 \DP_OP_751_130_6421/U977  ( .A(\DataPath/ALUhw/MULT/mux_out[5][16] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1304 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1046  ( .A(\DataPath/ALUhw/MULT/mux_out[4][15] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1405 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1115  ( .A(\DataPath/ALUhw/MULT/mux_out[3][14] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1506 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1184  ( .A(\DataPath/ALUhw/MULT/mux_out[2][13] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1607 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1287  ( .A(\DP_OP_751_130_6421/n1775 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][12] ), .S(n7974), .Z(
        \DP_OP_751_130_6421/n1740 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1255  ( .A(\DataPath/ALUhw/MULT/mux_out[1][12] ), .B(n8059), .Z(\DP_OP_751_130_6421/n1710 ) );
  XOR2_X1 \DP_OP_751_130_6421/U563  ( .A(\DataPath/ALUhw/MULT/mux_out[11][22] ), .B(n7782), .Z(\DP_OP_751_130_6421/n698 ) );
  XOR2_X1 \DP_OP_751_130_6421/U562  ( .A(\DataPath/ALUhw/MULT/mux_out[11][23] ), .B(n7782), .Z(\DP_OP_751_130_6421/n697 ) );
  XOR2_X1 \DP_OP_751_130_6421/U631  ( .A(\DataPath/ALUhw/MULT/mux_out[10][22] ), .B(n8062), .Z(\DP_OP_751_130_6421/n798 ) );
  XOR2_X1 \DP_OP_751_130_6421/U700  ( .A(\DataPath/ALUhw/MULT/mux_out[9][21] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n899 ) );
  XOR2_X1 \DP_OP_751_130_6421/U769  ( .A(\DataPath/ALUhw/MULT/mux_out[8][20] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n1000 ) );
  XOR2_X1 \DP_OP_751_130_6421/U838  ( .A(\DataPath/ALUhw/MULT/mux_out[7][19] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1101 ) );
  XOR2_X1 \DP_OP_751_130_6421/U907  ( .A(\DataPath/ALUhw/MULT/mux_out[6][18] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1202 ) );
  XOR2_X1 \DP_OP_751_130_6421/U976  ( .A(\DataPath/ALUhw/MULT/mux_out[5][17] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1303 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1045  ( .A(\DataPath/ALUhw/MULT/mux_out[4][16] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1404 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1114  ( .A(\DataPath/ALUhw/MULT/mux_out[3][15] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1505 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1183  ( .A(\DataPath/ALUhw/MULT/mux_out[2][14] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1606 ) );
  XOR2_X1 \DP_OP_751_130_6421/U493  ( .A(\DataPath/ALUhw/MULT/mux_out[12][24] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n596 ) );
  XOR2_X1 \DP_OP_751_130_6421/U492  ( .A(\DataPath/ALUhw/MULT/mux_out[12][25] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n595 ) );
  XOR2_X1 \DP_OP_751_130_6421/U561  ( .A(\DataPath/ALUhw/MULT/mux_out[11][24] ), .B(n7782), .Z(\DP_OP_751_130_6421/n696 ) );
  XOR2_X1 \DP_OP_751_130_6421/U630  ( .A(\DataPath/ALUhw/MULT/mux_out[10][23] ), .B(n8062), .Z(\DP_OP_751_130_6421/n797 ) );
  XOR2_X1 \DP_OP_751_130_6421/U699  ( .A(\DataPath/ALUhw/MULT/mux_out[9][22] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n898 ) );
  XOR2_X1 \DP_OP_751_130_6421/U768  ( .A(\DataPath/ALUhw/MULT/mux_out[8][21] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n999 ) );
  XOR2_X1 \DP_OP_751_130_6421/U837  ( .A(\DataPath/ALUhw/MULT/mux_out[7][20] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1100 ) );
  XOR2_X1 \DP_OP_751_130_6421/U906  ( .A(\DataPath/ALUhw/MULT/mux_out[6][19] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1201 ) );
  XOR2_X1 \DP_OP_751_130_6421/U975  ( .A(\DataPath/ALUhw/MULT/mux_out[5][18] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1302 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1044  ( .A(\DataPath/ALUhw/MULT/mux_out[4][17] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1403 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1113  ( .A(\DataPath/ALUhw/MULT/mux_out[3][16] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1504 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1182  ( .A(\DataPath/ALUhw/MULT/mux_out[2][15] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1605 ) );
  XOR2_X1 \DP_OP_751_130_6421/U423  ( .A(\DataPath/ALUhw/MULT/mux_out[13][26] ), .B(\DP_OP_751_130_6421/n495 ), .Z(\DP_OP_751_130_6421/n494 ) );
  XOR2_X1 \DP_OP_751_130_6421/U422  ( .A(\DataPath/ALUhw/MULT/mux_out[13][27] ), .B(\DP_OP_751_130_6421/n495 ), .Z(\DP_OP_751_130_6421/n493 ) );
  XOR2_X1 \DP_OP_751_130_6421/U491  ( .A(\DataPath/ALUhw/MULT/mux_out[12][26] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n594 ) );
  XOR2_X1 \DP_OP_751_130_6421/U560  ( .A(\DataPath/ALUhw/MULT/mux_out[11][25] ), .B(n7782), .Z(\DP_OP_751_130_6421/n695 ) );
  XOR2_X1 \DP_OP_751_130_6421/U629  ( .A(\DataPath/ALUhw/MULT/mux_out[10][24] ), .B(n8062), .Z(\DP_OP_751_130_6421/n796 ) );
  XOR2_X1 \DP_OP_751_130_6421/U698  ( .A(\DataPath/ALUhw/MULT/mux_out[9][23] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n897 ) );
  XOR2_X1 \DP_OP_751_130_6421/U767  ( .A(\DataPath/ALUhw/MULT/mux_out[8][22] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n998 ) );
  XOR2_X1 \DP_OP_751_130_6421/U836  ( .A(\DataPath/ALUhw/MULT/mux_out[7][21] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1099 ) );
  XOR2_X1 \DP_OP_751_130_6421/U905  ( .A(\DataPath/ALUhw/MULT/mux_out[6][20] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1200 ) );
  XOR2_X1 \DP_OP_751_130_6421/U974  ( .A(\DataPath/ALUhw/MULT/mux_out[5][19] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1301 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1043  ( .A(\DataPath/ALUhw/MULT/mux_out[4][18] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1402 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1112  ( .A(\DataPath/ALUhw/MULT/mux_out[3][17] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1503 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1181  ( .A(\DataPath/ALUhw/MULT/mux_out[2][16] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1604 ) );
  XOR2_X1 \DP_OP_751_130_6421/U353  ( .A(\DataPath/ALUhw/MULT/mux_out[14][28] ), .B(\DP_OP_751_130_6421/n393 ), .Z(\DP_OP_751_130_6421/n392 ) );
  XOR2_X1 \DP_OP_751_130_6421/U352  ( .A(\DataPath/ALUhw/MULT/mux_out[14][29] ), .B(\DP_OP_751_130_6421/n393 ), .Z(\DP_OP_751_130_6421/n391 ) );
  XOR2_X1 \DP_OP_751_130_6421/U421  ( .A(\DataPath/ALUhw/MULT/mux_out[13][28] ), .B(\DP_OP_751_130_6421/n495 ), .Z(\DP_OP_751_130_6421/n492 ) );
  XOR2_X1 \DP_OP_751_130_6421/U490  ( .A(\DataPath/ALUhw/MULT/mux_out[12][27] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n593 ) );
  XOR2_X1 \DP_OP_751_130_6421/U559  ( .A(\DataPath/ALUhw/MULT/mux_out[11][26] ), .B(n7782), .Z(\DP_OP_751_130_6421/n694 ) );
  XOR2_X1 \DP_OP_751_130_6421/U628  ( .A(\DataPath/ALUhw/MULT/mux_out[10][25] ), .B(n8062), .Z(\DP_OP_751_130_6421/n795 ) );
  XOR2_X1 \DP_OP_751_130_6421/U697  ( .A(\DataPath/ALUhw/MULT/mux_out[9][24] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n896 ) );
  XOR2_X1 \DP_OP_751_130_6421/U766  ( .A(\DataPath/ALUhw/MULT/mux_out[8][23] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n997 ) );
  XOR2_X1 \DP_OP_751_130_6421/U835  ( .A(\DataPath/ALUhw/MULT/mux_out[7][22] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1098 ) );
  XOR2_X1 \DP_OP_751_130_6421/U904  ( .A(\DataPath/ALUhw/MULT/mux_out[6][21] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1199 ) );
  XOR2_X1 \DP_OP_751_130_6421/U973  ( .A(\DataPath/ALUhw/MULT/mux_out[5][20] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1300 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1042  ( .A(\DataPath/ALUhw/MULT/mux_out[4][19] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1401 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1111  ( .A(\DataPath/ALUhw/MULT/mux_out[3][18] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1502 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1180  ( .A(\DataPath/ALUhw/MULT/mux_out[2][17] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1603 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1283  ( .A(\DP_OP_751_130_6421/n1771 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][16] ), .S(n7974), .Z(
        \DP_OP_751_130_6421/n1736 ) );
  XOR2_X1 \DP_OP_751_130_6421/U283  ( .A(\DataPath/ALUhw/MULT/mux_out[15][30] ), .B(\DP_OP_751_130_6421/n291 ), .Z(\DP_OP_751_130_6421/n290 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1268  ( .A(\DP_OP_751_130_6421/n1756 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][31] ), .S(n7880), .Z(
        \DP_OP_751_130_6421/n1721 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1236  ( .A(\DataPath/ALUhw/MULT/mux_out[1][31] ), .B(n7690), .Z(\DP_OP_751_130_6421/n1691 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1098  ( .A(\DataPath/ALUhw/MULT/mux_out[3][31] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1489 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1030  ( .A(\DataPath/ALUhw/MULT/mux_out[4][31] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1389 ) );
  XOR2_X1 \DP_OP_751_130_6421/U962  ( .A(\DataPath/ALUhw/MULT/mux_out[5][31] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1289 ) );
  XOR2_X1 \DP_OP_751_130_6421/U894  ( .A(\DataPath/ALUhw/MULT/mux_out[6][31] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1189 ) );
  XOR2_X1 \DP_OP_751_130_6421/U826  ( .A(\DataPath/ALUhw/MULT/mux_out[7][31] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1089 ) );
  XOR2_X1 \DP_OP_751_130_6421/U758  ( .A(\DataPath/ALUhw/MULT/mux_out[8][31] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n989 ) );
  XOR2_X1 \DP_OP_751_130_6421/U690  ( .A(\DataPath/ALUhw/MULT/mux_out[9][31] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n889 ) );
  XOR2_X1 \DP_OP_751_130_6421/U622  ( .A(\DataPath/ALUhw/MULT/mux_out[10][31] ), .B(n8062), .Z(\DP_OP_751_130_6421/n789 ) );
  XOR2_X1 \DP_OP_751_130_6421/U554  ( .A(\DataPath/ALUhw/MULT/mux_out[11][31] ), .B(n7782), .Z(\DP_OP_751_130_6421/n689 ) );
  XOR2_X1 \DP_OP_751_130_6421/U486  ( .A(\DataPath/ALUhw/MULT/mux_out[12][31] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n589 ) );
  XOR2_X1 \DP_OP_751_130_6421/U418  ( .A(\DataPath/ALUhw/MULT/mux_out[13][31] ), .B(\DP_OP_751_130_6421/n495 ), .Z(\DP_OP_751_130_6421/n489 ) );
  XOR2_X1 \DP_OP_751_130_6421/U350  ( .A(\DataPath/ALUhw/MULT/mux_out[14][31] ), .B(\DP_OP_751_130_6421/n393 ), .Z(\DP_OP_751_130_6421/n389 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1237  ( .A(\DataPath/ALUhw/MULT/mux_out[1][30] ), .B(n7690), .Z(\DP_OP_751_130_6421/n1692 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1167  ( .A(\DataPath/ALUhw/MULT/mux_out[2][30] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1590 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1099  ( .A(\DataPath/ALUhw/MULT/mux_out[3][30] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1490 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1031  ( .A(\DataPath/ALUhw/MULT/mux_out[4][30] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1390 ) );
  XOR2_X1 \DP_OP_751_130_6421/U963  ( .A(\DataPath/ALUhw/MULT/mux_out[5][30] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1290 ) );
  XOR2_X1 \DP_OP_751_130_6421/U895  ( .A(\DataPath/ALUhw/MULT/mux_out[6][30] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1190 ) );
  XOR2_X1 \DP_OP_751_130_6421/U827  ( .A(\DataPath/ALUhw/MULT/mux_out[7][30] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1090 ) );
  XOR2_X1 \DP_OP_751_130_6421/U759  ( .A(\DataPath/ALUhw/MULT/mux_out[8][30] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n990 ) );
  XOR2_X1 \DP_OP_751_130_6421/U691  ( .A(\DataPath/ALUhw/MULT/mux_out[9][30] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n890 ) );
  XOR2_X1 \DP_OP_751_130_6421/U623  ( .A(\DataPath/ALUhw/MULT/mux_out[10][30] ), .B(n8062), .Z(\DP_OP_751_130_6421/n790 ) );
  XOR2_X1 \DP_OP_751_130_6421/U555  ( .A(\DataPath/ALUhw/MULT/mux_out[11][30] ), .B(n7782), .Z(\DP_OP_751_130_6421/n690 ) );
  XOR2_X1 \DP_OP_751_130_6421/U487  ( .A(\DataPath/ALUhw/MULT/mux_out[12][30] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n590 ) );
  XOR2_X1 \DP_OP_751_130_6421/U419  ( .A(\DataPath/ALUhw/MULT/mux_out[13][30] ), .B(\DP_OP_751_130_6421/n495 ), .Z(\DP_OP_751_130_6421/n490 ) );
  XOR2_X1 \DP_OP_751_130_6421/U351  ( .A(\DataPath/ALUhw/MULT/mux_out[14][30] ), .B(\DP_OP_751_130_6421/n393 ), .Z(\DP_OP_751_130_6421/n390 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1168  ( .A(\DataPath/ALUhw/MULT/mux_out[2][29] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1591 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1100  ( .A(\DataPath/ALUhw/MULT/mux_out[3][29] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1491 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1032  ( .A(\DataPath/ALUhw/MULT/mux_out[4][29] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1391 ) );
  XOR2_X1 \DP_OP_751_130_6421/U964  ( .A(\DataPath/ALUhw/MULT/mux_out[5][29] ), 
        .B(\DP_OP_751_130_6421/n1311 ), .Z(\DP_OP_751_130_6421/n1291 ) );
  XOR2_X1 \DP_OP_751_130_6421/U896  ( .A(\DataPath/ALUhw/MULT/mux_out[6][29] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1191 ) );
  XOR2_X1 \DP_OP_751_130_6421/U828  ( .A(\DataPath/ALUhw/MULT/mux_out[7][29] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1091 ) );
  XOR2_X1 \DP_OP_751_130_6421/U760  ( .A(\DataPath/ALUhw/MULT/mux_out[8][29] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n991 ) );
  XOR2_X1 \DP_OP_751_130_6421/U692  ( .A(\DataPath/ALUhw/MULT/mux_out[9][29] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n891 ) );
  XOR2_X1 \DP_OP_751_130_6421/U624  ( .A(\DataPath/ALUhw/MULT/mux_out[10][29] ), .B(n8062), .Z(\DP_OP_751_130_6421/n791 ) );
  XOR2_X1 \DP_OP_751_130_6421/U556  ( .A(\DataPath/ALUhw/MULT/mux_out[11][29] ), .B(n7782), .Z(\DP_OP_751_130_6421/n691 ) );
  XOR2_X1 \DP_OP_751_130_6421/U488  ( .A(\DataPath/ALUhw/MULT/mux_out[12][29] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n591 ) );
  XOR2_X1 \DP_OP_751_130_6421/U420  ( .A(\DataPath/ALUhw/MULT/mux_out[13][29] ), .B(\DP_OP_751_130_6421/n495 ), .Z(\DP_OP_751_130_6421/n491 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1101  ( .A(\DataPath/ALUhw/MULT/mux_out[3][28] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1492 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1033  ( .A(\DataPath/ALUhw/MULT/mux_out[4][28] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1392 ) );
  XOR2_X1 \DP_OP_751_130_6421/U965  ( .A(\DataPath/ALUhw/MULT/mux_out[5][28] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1292 ) );
  XOR2_X1 \DP_OP_751_130_6421/U897  ( .A(\DataPath/ALUhw/MULT/mux_out[6][28] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1192 ) );
  XOR2_X1 \DP_OP_751_130_6421/U829  ( .A(\DataPath/ALUhw/MULT/mux_out[7][28] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1092 ) );
  XOR2_X1 \DP_OP_751_130_6421/U761  ( .A(\DataPath/ALUhw/MULT/mux_out[8][28] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n992 ) );
  XOR2_X1 \DP_OP_751_130_6421/U693  ( .A(\DataPath/ALUhw/MULT/mux_out[9][28] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n892 ) );
  XOR2_X1 \DP_OP_751_130_6421/U625  ( .A(\DataPath/ALUhw/MULT/mux_out[10][28] ), .B(n8062), .Z(\DP_OP_751_130_6421/n792 ) );
  XOR2_X1 \DP_OP_751_130_6421/U557  ( .A(\DataPath/ALUhw/MULT/mux_out[11][28] ), .B(n7782), .Z(\DP_OP_751_130_6421/n692 ) );
  XOR2_X1 \DP_OP_751_130_6421/U489  ( .A(\DataPath/ALUhw/MULT/mux_out[12][28] ), .B(\DP_OP_751_130_6421/n597 ), .Z(\DP_OP_751_130_6421/n592 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1102  ( .A(\DataPath/ALUhw/MULT/mux_out[3][27] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1493 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1034  ( .A(\DataPath/ALUhw/MULT/mux_out[4][27] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1393 ) );
  XOR2_X1 \DP_OP_751_130_6421/U966  ( .A(\DataPath/ALUhw/MULT/mux_out[5][27] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1293 ) );
  XOR2_X1 \DP_OP_751_130_6421/U898  ( .A(\DataPath/ALUhw/MULT/mux_out[6][27] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1193 ) );
  XOR2_X1 \DP_OP_751_130_6421/U830  ( .A(\DataPath/ALUhw/MULT/mux_out[7][27] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1093 ) );
  XOR2_X1 \DP_OP_751_130_6421/U762  ( .A(\DataPath/ALUhw/MULT/mux_out[8][27] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n993 ) );
  XOR2_X1 \DP_OP_751_130_6421/U694  ( .A(\DataPath/ALUhw/MULT/mux_out[9][27] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n893 ) );
  XOR2_X1 \DP_OP_751_130_6421/U626  ( .A(\DataPath/ALUhw/MULT/mux_out[10][27] ), .B(n8062), .Z(\DP_OP_751_130_6421/n793 ) );
  XOR2_X1 \DP_OP_751_130_6421/U558  ( .A(\DataPath/ALUhw/MULT/mux_out[11][27] ), .B(n7782), .Z(\DP_OP_751_130_6421/n693 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1273  ( .A(\DP_OP_751_130_6421/n1761 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][26] ), .S(n7880), .Z(
        \DP_OP_751_130_6421/n1726 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1171  ( .A(\DataPath/ALUhw/MULT/mux_out[2][26] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1594 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1103  ( .A(\DataPath/ALUhw/MULT/mux_out[3][26] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1494 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1035  ( .A(\DataPath/ALUhw/MULT/mux_out[4][26] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1394 ) );
  XOR2_X1 \DP_OP_751_130_6421/U967  ( .A(\DataPath/ALUhw/MULT/mux_out[5][26] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1294 ) );
  XOR2_X1 \DP_OP_751_130_6421/U899  ( .A(\DataPath/ALUhw/MULT/mux_out[6][26] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1194 ) );
  XOR2_X1 \DP_OP_751_130_6421/U831  ( .A(\DataPath/ALUhw/MULT/mux_out[7][26] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1094 ) );
  XOR2_X1 \DP_OP_751_130_6421/U763  ( .A(\DataPath/ALUhw/MULT/mux_out[8][26] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n994 ) );
  XOR2_X1 \DP_OP_751_130_6421/U695  ( .A(\DataPath/ALUhw/MULT/mux_out[9][26] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n894 ) );
  XOR2_X1 \DP_OP_751_130_6421/U627  ( .A(\DataPath/ALUhw/MULT/mux_out[10][26] ), .B(n8062), .Z(\DP_OP_751_130_6421/n794 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1274  ( .A(\DP_OP_751_130_6421/n1762 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][25] ), .S(n7880), .Z(
        \DP_OP_751_130_6421/n1727 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1172  ( .A(\DataPath/ALUhw/MULT/mux_out[2][25] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1595 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1104  ( .A(\DataPath/ALUhw/MULT/mux_out[3][25] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1495 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1036  ( .A(\DataPath/ALUhw/MULT/mux_out[4][25] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1395 ) );
  XOR2_X1 \DP_OP_751_130_6421/U968  ( .A(\DataPath/ALUhw/MULT/mux_out[5][25] ), 
        .B(\DP_OP_751_130_6421/n1311 ), .Z(\DP_OP_751_130_6421/n1295 ) );
  XOR2_X1 \DP_OP_751_130_6421/U900  ( .A(\DataPath/ALUhw/MULT/mux_out[6][25] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1195 ) );
  XOR2_X1 \DP_OP_751_130_6421/U832  ( .A(\DataPath/ALUhw/MULT/mux_out[7][25] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1095 ) );
  XOR2_X1 \DP_OP_751_130_6421/U764  ( .A(\DataPath/ALUhw/MULT/mux_out[8][25] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n995 ) );
  XOR2_X1 \DP_OP_751_130_6421/U696  ( .A(\DataPath/ALUhw/MULT/mux_out[9][25] ), 
        .B(n8061), .Z(\DP_OP_751_130_6421/n895 ) );
  MUX2_X1 \DP_OP_751_130_6421/U1275  ( .A(\DP_OP_751_130_6421/n1763 ), .B(
        \DataPath/ALUhw/MULT/mux_out[0][24] ), .S(n7880), .Z(
        \DP_OP_751_130_6421/n1728 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1173  ( .A(\DataPath/ALUhw/MULT/mux_out[2][24] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1596 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1105  ( .A(\DataPath/ALUhw/MULT/mux_out[3][24] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1496 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1037  ( .A(\DataPath/ALUhw/MULT/mux_out[4][24] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1396 ) );
  XOR2_X1 \DP_OP_751_130_6421/U969  ( .A(\DataPath/ALUhw/MULT/mux_out[5][24] ), 
        .B(\DP_OP_751_130_6421/n1311 ), .Z(\DP_OP_751_130_6421/n1296 ) );
  XOR2_X1 \DP_OP_751_130_6421/U901  ( .A(\DataPath/ALUhw/MULT/mux_out[6][24] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1196 ) );
  XOR2_X1 \DP_OP_751_130_6421/U833  ( .A(\DataPath/ALUhw/MULT/mux_out[7][24] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1096 ) );
  XOR2_X1 \DP_OP_751_130_6421/U765  ( .A(\DataPath/ALUhw/MULT/mux_out[8][24] ), 
        .B(\DP_OP_751_130_6421/n1005 ), .Z(\DP_OP_751_130_6421/n996 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1174  ( .A(\DataPath/ALUhw/MULT/mux_out[2][23] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1597 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1106  ( .A(\DataPath/ALUhw/MULT/mux_out[3][23] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1497 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1038  ( .A(\DataPath/ALUhw/MULT/mux_out[4][23] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1397 ) );
  XOR2_X1 \DP_OP_751_130_6421/U970  ( .A(\DataPath/ALUhw/MULT/mux_out[5][23] ), 
        .B(\DP_OP_751_130_6421/n1311 ), .Z(\DP_OP_751_130_6421/n1297 ) );
  XOR2_X1 \DP_OP_751_130_6421/U902  ( .A(\DataPath/ALUhw/MULT/mux_out[6][23] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1197 ) );
  XOR2_X1 \DP_OP_751_130_6421/U834  ( .A(\DataPath/ALUhw/MULT/mux_out[7][23] ), 
        .B(\DP_OP_751_130_6421/n1107 ), .Z(\DP_OP_751_130_6421/n1097 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1175  ( .A(\DataPath/ALUhw/MULT/mux_out[2][22] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1598 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1107  ( .A(\DataPath/ALUhw/MULT/mux_out[3][22] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1498 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1039  ( .A(\DataPath/ALUhw/MULT/mux_out[4][22] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1398 ) );
  XOR2_X1 \DP_OP_751_130_6421/U971  ( .A(\DataPath/ALUhw/MULT/mux_out[5][22] ), 
        .B(\DP_OP_751_130_6421/n1311 ), .Z(\DP_OP_751_130_6421/n1298 ) );
  XOR2_X1 \DP_OP_751_130_6421/U903  ( .A(\DataPath/ALUhw/MULT/mux_out[6][22] ), 
        .B(\DP_OP_751_130_6421/n1209 ), .Z(\DP_OP_751_130_6421/n1198 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1246  ( .A(\DataPath/ALUhw/MULT/mux_out[1][21] ), .B(n7690), .Z(\DP_OP_751_130_6421/n1701 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1176  ( .A(\DataPath/ALUhw/MULT/mux_out[2][21] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1599 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1108  ( .A(\DataPath/ALUhw/MULT/mux_out[3][21] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1499 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1040  ( .A(\DataPath/ALUhw/MULT/mux_out[4][21] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1399 ) );
  XOR2_X1 \DP_OP_751_130_6421/U972  ( .A(\DataPath/ALUhw/MULT/mux_out[5][21] ), 
        .B(n8055), .Z(\DP_OP_751_130_6421/n1299 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1247  ( .A(\DataPath/ALUhw/MULT/mux_out[1][20] ), .B(n7690), .Z(\DP_OP_751_130_6421/n1702 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1177  ( .A(\DataPath/ALUhw/MULT/mux_out[2][20] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1600 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1109  ( .A(\DataPath/ALUhw/MULT/mux_out[3][20] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1500 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1041  ( .A(\DataPath/ALUhw/MULT/mux_out[4][20] ), .B(\DP_OP_751_130_6421/n1413 ), .Z(\DP_OP_751_130_6421/n1400 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1178  ( .A(\DataPath/ALUhw/MULT/mux_out[2][19] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1601 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1110  ( .A(\DataPath/ALUhw/MULT/mux_out[3][19] ), .B(n8056), .Z(\DP_OP_751_130_6421/n1501 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1249  ( .A(\DataPath/ALUhw/MULT/mux_out[1][18] ), .B(n7690), .Z(\DP_OP_751_130_6421/n1704 ) );
  XOR2_X1 \DP_OP_751_130_6421/U1179  ( .A(\DataPath/ALUhw/MULT/mux_out[2][18] ), .B(n8057), .Z(\DP_OP_751_130_6421/n1602 ) );
  HA_X1 \DP_OP_751_130_6421/U1225  ( .A(\DP_OP_751_130_6421/n1714 ), .B(
        \DP_OP_751_130_6421/n1744 ), .CO(\DP_OP_751_130_6421/n1671 ), .S(
        \DP_OP_751_130_6421/n1672 ) );
  HA_X1 \DP_OP_751_130_6421/U1224  ( .A(\DP_OP_751_130_6421/n1713 ), .B(
        \DP_OP_751_130_6421/n1743 ), .CO(\DP_OP_751_130_6421/n1669 ), .S(
        \DP_OP_751_130_6421/n1670 ) );
  HA_X1 \DP_OP_751_130_6421/U1223  ( .A(\DP_OP_751_130_6421/n1712 ), .B(
        \DP_OP_751_130_6421/n1742 ), .CO(\DP_OP_751_130_6421/n1667 ), .S(
        \DP_OP_751_130_6421/n1668 ) );
  HA_X1 \DP_OP_751_130_6421/U1222  ( .A(\DP_OP_751_130_6421/n1711 ), .B(
        \DP_OP_751_130_6421/n1741 ), .CO(\DP_OP_751_130_6421/n1665 ), .S(
        \DP_OP_751_130_6421/n1666 ) );
  HA_X1 \DP_OP_751_130_6421/U1221  ( .A(\DP_OP_751_130_6421/n1710 ), .B(
        \DP_OP_751_130_6421/n1740 ), .CO(\DP_OP_751_130_6421/n1663 ), .S(
        \DP_OP_751_130_6421/n1664 ) );
  HA_X1 \DP_OP_751_130_6421/U1217  ( .A(\DP_OP_751_130_6421/n1706 ), .B(
        \DP_OP_751_130_6421/n1736 ), .CO(\DP_OP_751_130_6421/n1655 ), .S(
        \DP_OP_751_130_6421/n1656 ) );
  HA_X1 \DP_OP_751_130_6421/U1216  ( .A(\DP_OP_751_130_6421/n1705 ), .B(
        \DP_OP_751_130_6421/n1735 ), .CO(\DP_OP_751_130_6421/n1653 ), .S(
        \DP_OP_751_130_6421/n1654 ) );
  HA_X1 \DP_OP_751_130_6421/U1215  ( .A(\DP_OP_751_130_6421/n1704 ), .B(
        \DP_OP_751_130_6421/n1734 ), .CO(\DP_OP_751_130_6421/n1651 ), .S(
        \DP_OP_751_130_6421/n1652 ) );
  HA_X1 \DP_OP_751_130_6421/U1214  ( .A(\DP_OP_751_130_6421/n1703 ), .B(
        \DP_OP_751_130_6421/n1733 ), .CO(\DP_OP_751_130_6421/n1649 ), .S(
        \DP_OP_751_130_6421/n1650 ) );
  HA_X1 \DP_OP_751_130_6421/U1213  ( .A(\DP_OP_751_130_6421/n1702 ), .B(
        \DP_OP_751_130_6421/n1732 ), .CO(\DP_OP_751_130_6421/n1647 ), .S(
        \DP_OP_751_130_6421/n1648 ) );
  HA_X1 \DP_OP_751_130_6421/U1212  ( .A(\DP_OP_751_130_6421/n1701 ), .B(
        \DP_OP_751_130_6421/n1731 ), .CO(\DP_OP_751_130_6421/n1645 ), .S(
        \DP_OP_751_130_6421/n1646 ) );
  HA_X1 \DP_OP_751_130_6421/U1210  ( .A(\DP_OP_751_130_6421/n1699 ), .B(
        \DP_OP_751_130_6421/n1729 ), .CO(\DP_OP_751_130_6421/n1641 ), .S(
        \DP_OP_751_130_6421/n1642 ) );
  HA_X1 \DP_OP_751_130_6421/U1209  ( .A(\DP_OP_751_130_6421/n1698 ), .B(
        \DP_OP_751_130_6421/n1728 ), .CO(\DP_OP_751_130_6421/n1639 ), .S(
        \DP_OP_751_130_6421/n1640 ) );
  HA_X1 \DP_OP_751_130_6421/U1202  ( .A(\DP_OP_751_130_6421/n1691 ), .B(
        \DP_OP_751_130_6421/n1721 ), .S(\DP_OP_751_130_6421/n1626 ) );
  FA_X1 \DP_OP_751_130_6421/U1158  ( .A(\DP_OP_751_130_6421/n1679 ), .B(
        \DP_OP_751_130_6421/n1615 ), .CI(\DP_OP_751_130_6421/n1678 ), .CO(
        \DP_OP_751_130_6421/n1579 ), .S(\DP_OP_751_130_6421/n1580 ) );
  FA_X1 \DP_OP_751_130_6421/U1157  ( .A(\DP_OP_751_130_6421/n1677 ), .B(
        \DP_OP_751_130_6421/n1614 ), .CI(\DP_OP_751_130_6421/n1676 ), .CO(
        \DP_OP_751_130_6421/n1577 ), .S(\DP_OP_751_130_6421/n1578 ) );
  FA_X1 \DP_OP_751_130_6421/U1156  ( .A(\DP_OP_751_130_6421/n1675 ), .B(
        \DP_OP_751_130_6421/n1613 ), .CI(\DP_OP_751_130_6421/n1674 ), .CO(
        \DP_OP_751_130_6421/n1575 ), .S(\DP_OP_751_130_6421/n1576 ) );
  FA_X1 \DP_OP_751_130_6421/U1155  ( .A(\DP_OP_751_130_6421/n1673 ), .B(
        \DP_OP_751_130_6421/n1612 ), .CI(\DP_OP_751_130_6421/n1672 ), .CO(
        \DP_OP_751_130_6421/n1573 ), .S(\DP_OP_751_130_6421/n1574 ) );
  FA_X1 \DP_OP_751_130_6421/U1154  ( .A(\DP_OP_751_130_6421/n1671 ), .B(
        \DP_OP_751_130_6421/n1611 ), .CI(\DP_OP_751_130_6421/n1670 ), .CO(
        \DP_OP_751_130_6421/n1571 ), .S(\DP_OP_751_130_6421/n1572 ) );
  FA_X1 \DP_OP_751_130_6421/U1153  ( .A(\DP_OP_751_130_6421/n1669 ), .B(
        \DP_OP_751_130_6421/n1610 ), .CI(\DP_OP_751_130_6421/n1668 ), .CO(
        \DP_OP_751_130_6421/n1569 ), .S(\DP_OP_751_130_6421/n1570 ) );
  FA_X1 \DP_OP_751_130_6421/U1152  ( .A(\DP_OP_751_130_6421/n1667 ), .B(
        \DP_OP_751_130_6421/n1609 ), .CI(\DP_OP_751_130_6421/n1666 ), .CO(
        \DP_OP_751_130_6421/n1567 ), .S(\DP_OP_751_130_6421/n1568 ) );
  FA_X1 \DP_OP_751_130_6421/U1151  ( .A(\DP_OP_751_130_6421/n1665 ), .B(
        \DP_OP_751_130_6421/n1608 ), .CI(\DP_OP_751_130_6421/n1664 ), .CO(
        \DP_OP_751_130_6421/n1565 ), .S(\DP_OP_751_130_6421/n1566 ) );
  FA_X1 \DP_OP_751_130_6421/U1150  ( .A(\DP_OP_751_130_6421/n1663 ), .B(
        \DP_OP_751_130_6421/n1607 ), .CI(\DP_OP_751_130_6421/n1662 ), .CO(
        \DP_OP_751_130_6421/n1563 ), .S(\DP_OP_751_130_6421/n1564 ) );
  FA_X1 \DP_OP_751_130_6421/U1149  ( .A(\DP_OP_751_130_6421/n1661 ), .B(
        \DP_OP_751_130_6421/n1606 ), .CI(\DP_OP_751_130_6421/n1660 ), .CO(
        \DP_OP_751_130_6421/n1561 ), .S(\DP_OP_751_130_6421/n1562 ) );
  FA_X1 \DP_OP_751_130_6421/U1148  ( .A(\DP_OP_751_130_6421/n1659 ), .B(
        \DP_OP_751_130_6421/n1605 ), .CI(\DP_OP_751_130_6421/n1658 ), .CO(
        \DP_OP_751_130_6421/n1559 ), .S(\DP_OP_751_130_6421/n1560 ) );
  FA_X1 \DP_OP_751_130_6421/U1147  ( .A(\DP_OP_751_130_6421/n1657 ), .B(
        \DP_OP_751_130_6421/n1604 ), .CI(\DP_OP_751_130_6421/n1656 ), .CO(
        \DP_OP_751_130_6421/n1557 ), .S(\DP_OP_751_130_6421/n1558 ) );
  FA_X1 \DP_OP_751_130_6421/U1146  ( .A(\DP_OP_751_130_6421/n1655 ), .B(
        \DP_OP_751_130_6421/n1603 ), .CI(\DP_OP_751_130_6421/n1654 ), .CO(
        \DP_OP_751_130_6421/n1555 ), .S(\DP_OP_751_130_6421/n1556 ) );
  FA_X1 \DP_OP_751_130_6421/U1145  ( .A(\DP_OP_751_130_6421/n1653 ), .B(
        \DP_OP_751_130_6421/n1602 ), .CI(\DP_OP_751_130_6421/n1652 ), .CO(
        \DP_OP_751_130_6421/n1553 ), .S(\DP_OP_751_130_6421/n1554 ) );
  FA_X1 \DP_OP_751_130_6421/U1144  ( .A(\DP_OP_751_130_6421/n1651 ), .B(
        \DP_OP_751_130_6421/n1601 ), .CI(\DP_OP_751_130_6421/n1650 ), .CO(
        \DP_OP_751_130_6421/n1551 ), .S(\DP_OP_751_130_6421/n1552 ) );
  FA_X1 \DP_OP_751_130_6421/U1143  ( .A(\DP_OP_751_130_6421/n1649 ), .B(
        \DP_OP_751_130_6421/n1600 ), .CI(\DP_OP_751_130_6421/n1648 ), .CO(
        \DP_OP_751_130_6421/n1549 ), .S(\DP_OP_751_130_6421/n1550 ) );
  FA_X1 \DP_OP_751_130_6421/U1142  ( .A(\DP_OP_751_130_6421/n1599 ), .B(
        \DP_OP_751_130_6421/n1647 ), .CI(\DP_OP_751_130_6421/n1646 ), .CO(
        \DP_OP_751_130_6421/n1547 ), .S(\DP_OP_751_130_6421/n1548 ) );
  FA_X1 \DP_OP_751_130_6421/U1141  ( .A(\DP_OP_751_130_6421/n1645 ), .B(
        \DP_OP_751_130_6421/n1598 ), .CI(\DP_OP_751_130_6421/n1644 ), .CO(
        \DP_OP_751_130_6421/n1545 ), .S(\DP_OP_751_130_6421/n1546 ) );
  FA_X1 \DP_OP_751_130_6421/U1140  ( .A(\DP_OP_751_130_6421/n1643 ), .B(
        \DP_OP_751_130_6421/n1597 ), .CI(\DP_OP_751_130_6421/n1642 ), .CO(
        \DP_OP_751_130_6421/n1543 ), .S(\DP_OP_751_130_6421/n1544 ) );
  FA_X1 \DP_OP_751_130_6421/U1139  ( .A(\DP_OP_751_130_6421/n1641 ), .B(
        \DP_OP_751_130_6421/n1596 ), .CI(\DP_OP_751_130_6421/n1640 ), .CO(
        \DP_OP_751_130_6421/n1541 ), .S(\DP_OP_751_130_6421/n1542 ) );
  FA_X1 \DP_OP_751_130_6421/U1138  ( .A(\DP_OP_751_130_6421/n1639 ), .B(
        \DP_OP_751_130_6421/n1595 ), .CI(\DP_OP_751_130_6421/n1638 ), .CO(
        \DP_OP_751_130_6421/n1539 ), .S(\DP_OP_751_130_6421/n1540 ) );
  FA_X1 \DP_OP_751_130_6421/U1137  ( .A(\DP_OP_751_130_6421/n1637 ), .B(
        \DP_OP_751_130_6421/n1594 ), .CI(\DP_OP_751_130_6421/n1636 ), .CO(
        \DP_OP_751_130_6421/n1537 ), .S(\DP_OP_751_130_6421/n1538 ) );
  FA_X1 \DP_OP_751_130_6421/U1136  ( .A(\DP_OP_751_130_6421/n1635 ), .B(
        \DP_OP_751_130_6421/n1593 ), .CI(\DP_OP_751_130_6421/n1634 ), .CO(
        \DP_OP_751_130_6421/n1535 ), .S(\DP_OP_751_130_6421/n1536 ) );
  FA_X1 \DP_OP_751_130_6421/U1135  ( .A(\DP_OP_751_130_6421/n1632 ), .B(
        \DP_OP_751_130_6421/n1592 ), .CI(\DP_OP_751_130_6421/n1633 ), .CO(
        \DP_OP_751_130_6421/n1533 ), .S(\DP_OP_751_130_6421/n1534 ) );
  FA_X1 \DP_OP_751_130_6421/U1134  ( .A(\DP_OP_751_130_6421/n1591 ), .B(
        \DP_OP_751_130_6421/n1631 ), .CI(\DP_OP_751_130_6421/n1630 ), .CO(
        \DP_OP_751_130_6421/n1531 ), .S(\DP_OP_751_130_6421/n1532 ) );
  FA_X1 \DP_OP_751_130_6421/U1133  ( .A(\DP_OP_751_130_6421/n1629 ), .B(
        \DP_OP_751_130_6421/n1590 ), .CI(\DP_OP_751_130_6421/n1628 ), .CO(
        \DP_OP_751_130_6421/n1529 ), .S(\DP_OP_751_130_6421/n1530 ) );
  FA_X1 \DP_OP_751_130_6421/U1089  ( .A(\DP_OP_751_130_6421/n1514 ), .B(n8056), 
        .CI(\DP_OP_751_130_6421/n1579 ), .CO(\DP_OP_751_130_6421/n1479 ), .S(
        \DP_OP_751_130_6421/n1480 ) );
  FA_X1 \DP_OP_751_130_6421/U1088  ( .A(\DP_OP_751_130_6421/n1577 ), .B(
        \DP_OP_751_130_6421/n1513 ), .CI(\DP_OP_751_130_6421/n1576 ), .CO(
        \DP_OP_751_130_6421/n1477 ), .S(\DP_OP_751_130_6421/n1478 ) );
  FA_X1 \DP_OP_751_130_6421/U1087  ( .A(\DP_OP_751_130_6421/n1575 ), .B(
        \DP_OP_751_130_6421/n1512 ), .CI(\DP_OP_751_130_6421/n1574 ), .CO(
        \DP_OP_751_130_6421/n1475 ), .S(\DP_OP_751_130_6421/n1476 ) );
  FA_X1 \DP_OP_751_130_6421/U1086  ( .A(\DP_OP_751_130_6421/n1573 ), .B(
        \DP_OP_751_130_6421/n1511 ), .CI(\DP_OP_751_130_6421/n1572 ), .CO(
        \DP_OP_751_130_6421/n1473 ), .S(\DP_OP_751_130_6421/n1474 ) );
  FA_X1 \DP_OP_751_130_6421/U1085  ( .A(\DP_OP_751_130_6421/n1571 ), .B(
        \DP_OP_751_130_6421/n1510 ), .CI(\DP_OP_751_130_6421/n1570 ), .CO(
        \DP_OP_751_130_6421/n1471 ), .S(\DP_OP_751_130_6421/n1472 ) );
  FA_X1 \DP_OP_751_130_6421/U1084  ( .A(\DP_OP_751_130_6421/n1569 ), .B(
        \DP_OP_751_130_6421/n1509 ), .CI(\DP_OP_751_130_6421/n1568 ), .CO(
        \DP_OP_751_130_6421/n1469 ), .S(\DP_OP_751_130_6421/n1470 ) );
  FA_X1 \DP_OP_751_130_6421/U1083  ( .A(\DP_OP_751_130_6421/n1567 ), .B(
        \DP_OP_751_130_6421/n1508 ), .CI(\DP_OP_751_130_6421/n1566 ), .CO(
        \DP_OP_751_130_6421/n1467 ), .S(\DP_OP_751_130_6421/n1468 ) );
  FA_X1 \DP_OP_751_130_6421/U1082  ( .A(\DP_OP_751_130_6421/n1565 ), .B(
        \DP_OP_751_130_6421/n1507 ), .CI(\DP_OP_751_130_6421/n1564 ), .CO(
        \DP_OP_751_130_6421/n1465 ), .S(\DP_OP_751_130_6421/n1466 ) );
  FA_X1 \DP_OP_751_130_6421/U1081  ( .A(\DP_OP_751_130_6421/n1563 ), .B(
        \DP_OP_751_130_6421/n1506 ), .CI(\DP_OP_751_130_6421/n1562 ), .CO(
        \DP_OP_751_130_6421/n1463 ), .S(\DP_OP_751_130_6421/n1464 ) );
  FA_X1 \DP_OP_751_130_6421/U1080  ( .A(\DP_OP_751_130_6421/n1561 ), .B(
        \DP_OP_751_130_6421/n1505 ), .CI(\DP_OP_751_130_6421/n1560 ), .CO(
        \DP_OP_751_130_6421/n1461 ), .S(\DP_OP_751_130_6421/n1462 ) );
  FA_X1 \DP_OP_751_130_6421/U1079  ( .A(\DP_OP_751_130_6421/n1559 ), .B(
        \DP_OP_751_130_6421/n1504 ), .CI(\DP_OP_751_130_6421/n1558 ), .CO(
        \DP_OP_751_130_6421/n1459 ), .S(\DP_OP_751_130_6421/n1460 ) );
  FA_X1 \DP_OP_751_130_6421/U1078  ( .A(\DP_OP_751_130_6421/n1557 ), .B(
        \DP_OP_751_130_6421/n1503 ), .CI(\DP_OP_751_130_6421/n1556 ), .CO(
        \DP_OP_751_130_6421/n1457 ), .S(\DP_OP_751_130_6421/n1458 ) );
  FA_X1 \DP_OP_751_130_6421/U1077  ( .A(\DP_OP_751_130_6421/n1555 ), .B(
        \DP_OP_751_130_6421/n1502 ), .CI(\DP_OP_751_130_6421/n1554 ), .CO(
        \DP_OP_751_130_6421/n1455 ), .S(\DP_OP_751_130_6421/n1456 ) );
  FA_X1 \DP_OP_751_130_6421/U1076  ( .A(\DP_OP_751_130_6421/n1553 ), .B(
        \DP_OP_751_130_6421/n1501 ), .CI(\DP_OP_751_130_6421/n1552 ), .CO(
        \DP_OP_751_130_6421/n1453 ), .S(\DP_OP_751_130_6421/n1454 ) );
  FA_X1 \DP_OP_751_130_6421/U1075  ( .A(\DP_OP_751_130_6421/n1551 ), .B(
        \DP_OP_751_130_6421/n1500 ), .CI(\DP_OP_751_130_6421/n1550 ), .CO(
        \DP_OP_751_130_6421/n1451 ), .S(\DP_OP_751_130_6421/n1452 ) );
  FA_X1 \DP_OP_751_130_6421/U1074  ( .A(\DP_OP_751_130_6421/n1549 ), .B(
        \DP_OP_751_130_6421/n1499 ), .CI(\DP_OP_751_130_6421/n1548 ), .CO(
        \DP_OP_751_130_6421/n1449 ), .S(\DP_OP_751_130_6421/n1450 ) );
  FA_X1 \DP_OP_751_130_6421/U1073  ( .A(\DP_OP_751_130_6421/n1547 ), .B(
        \DP_OP_751_130_6421/n1498 ), .CI(\DP_OP_751_130_6421/n1546 ), .CO(
        \DP_OP_751_130_6421/n1447 ), .S(\DP_OP_751_130_6421/n1448 ) );
  FA_X1 \DP_OP_751_130_6421/U1072  ( .A(\DP_OP_751_130_6421/n1545 ), .B(
        \DP_OP_751_130_6421/n1497 ), .CI(\DP_OP_751_130_6421/n1544 ), .CO(
        \DP_OP_751_130_6421/n1445 ), .S(\DP_OP_751_130_6421/n1446 ) );
  FA_X1 \DP_OP_751_130_6421/U1071  ( .A(\DP_OP_751_130_6421/n1543 ), .B(
        \DP_OP_751_130_6421/n1496 ), .CI(\DP_OP_751_130_6421/n1542 ), .CO(
        \DP_OP_751_130_6421/n1443 ), .S(\DP_OP_751_130_6421/n1444 ) );
  FA_X1 \DP_OP_751_130_6421/U1070  ( .A(\DP_OP_751_130_6421/n1495 ), .B(
        \DP_OP_751_130_6421/n1541 ), .CI(\DP_OP_751_130_6421/n1540 ), .CO(
        \DP_OP_751_130_6421/n1441 ), .S(\DP_OP_751_130_6421/n1442 ) );
  FA_X1 \DP_OP_751_130_6421/U1069  ( .A(\DP_OP_751_130_6421/n1539 ), .B(
        \DP_OP_751_130_6421/n1494 ), .CI(\DP_OP_751_130_6421/n1538 ), .CO(
        \DP_OP_751_130_6421/n1439 ), .S(\DP_OP_751_130_6421/n1440 ) );
  FA_X1 \DP_OP_751_130_6421/U1068  ( .A(\DP_OP_751_130_6421/n1537 ), .B(
        \DP_OP_751_130_6421/n1493 ), .CI(\DP_OP_751_130_6421/n1536 ), .CO(
        \DP_OP_751_130_6421/n1437 ), .S(\DP_OP_751_130_6421/n1438 ) );
  FA_X1 \DP_OP_751_130_6421/U1067  ( .A(\DP_OP_751_130_6421/n1535 ), .B(
        \DP_OP_751_130_6421/n1492 ), .CI(\DP_OP_751_130_6421/n1534 ), .CO(
        \DP_OP_751_130_6421/n1435 ), .S(\DP_OP_751_130_6421/n1436 ) );
  FA_X1 \DP_OP_751_130_6421/U1066  ( .A(\DP_OP_751_130_6421/n1533 ), .B(
        \DP_OP_751_130_6421/n1491 ), .CI(\DP_OP_751_130_6421/n1532 ), .CO(
        \DP_OP_751_130_6421/n1433 ), .S(\DP_OP_751_130_6421/n1434 ) );
  FA_X1 \DP_OP_751_130_6421/U1064  ( .A(\DP_OP_751_130_6421/n1529 ), .B(
        \DP_OP_751_130_6421/n1489 ), .CI(\DP_OP_751_130_6421/n1528 ), .S(
        \DP_OP_751_130_6421/n1430 ) );
  FA_X1 \DP_OP_751_130_6421/U1018  ( .A(\DP_OP_751_130_6421/n1475 ), .B(
        \DP_OP_751_130_6421/n1411 ), .CI(\DP_OP_751_130_6421/n1474 ), .CO(
        \DP_OP_751_130_6421/n1375 ), .S(\DP_OP_751_130_6421/n1376 ) );
  FA_X1 \DP_OP_751_130_6421/U1017  ( .A(\DP_OP_751_130_6421/n1473 ), .B(
        \DP_OP_751_130_6421/n1410 ), .CI(\DP_OP_751_130_6421/n1472 ), .CO(
        \DP_OP_751_130_6421/n1373 ), .S(\DP_OP_751_130_6421/n1374 ) );
  FA_X1 \DP_OP_751_130_6421/U1016  ( .A(\DP_OP_751_130_6421/n1471 ), .B(
        \DP_OP_751_130_6421/n1409 ), .CI(\DP_OP_751_130_6421/n1470 ), .CO(
        \DP_OP_751_130_6421/n1371 ), .S(\DP_OP_751_130_6421/n1372 ) );
  FA_X1 \DP_OP_751_130_6421/U1015  ( .A(\DP_OP_751_130_6421/n1469 ), .B(
        \DP_OP_751_130_6421/n1408 ), .CI(\DP_OP_751_130_6421/n1468 ), .CO(
        \DP_OP_751_130_6421/n1369 ), .S(\DP_OP_751_130_6421/n1370 ) );
  FA_X1 \DP_OP_751_130_6421/U1014  ( .A(\DP_OP_751_130_6421/n1467 ), .B(
        \DP_OP_751_130_6421/n1407 ), .CI(\DP_OP_751_130_6421/n1466 ), .CO(
        \DP_OP_751_130_6421/n1367 ), .S(\DP_OP_751_130_6421/n1368 ) );
  FA_X1 \DP_OP_751_130_6421/U1013  ( .A(\DP_OP_751_130_6421/n1465 ), .B(
        \DP_OP_751_130_6421/n1406 ), .CI(\DP_OP_751_130_6421/n1464 ), .CO(
        \DP_OP_751_130_6421/n1365 ), .S(\DP_OP_751_130_6421/n1366 ) );
  FA_X1 \DP_OP_751_130_6421/U1012  ( .A(\DP_OP_751_130_6421/n1463 ), .B(
        \DP_OP_751_130_6421/n1405 ), .CI(\DP_OP_751_130_6421/n1462 ), .CO(
        \DP_OP_751_130_6421/n1363 ), .S(\DP_OP_751_130_6421/n1364 ) );
  FA_X1 \DP_OP_751_130_6421/U1011  ( .A(\DP_OP_751_130_6421/n1461 ), .B(
        \DP_OP_751_130_6421/n1404 ), .CI(\DP_OP_751_130_6421/n1460 ), .CO(
        \DP_OP_751_130_6421/n1361 ), .S(\DP_OP_751_130_6421/n1362 ) );
  FA_X1 \DP_OP_751_130_6421/U1010  ( .A(\DP_OP_751_130_6421/n1459 ), .B(
        \DP_OP_751_130_6421/n1403 ), .CI(\DP_OP_751_130_6421/n1458 ), .CO(
        \DP_OP_751_130_6421/n1359 ), .S(\DP_OP_751_130_6421/n1360 ) );
  FA_X1 \DP_OP_751_130_6421/U1009  ( .A(\DP_OP_751_130_6421/n1457 ), .B(
        \DP_OP_751_130_6421/n1402 ), .CI(\DP_OP_751_130_6421/n1456 ), .CO(
        \DP_OP_751_130_6421/n1357 ), .S(\DP_OP_751_130_6421/n1358 ) );
  FA_X1 \DP_OP_751_130_6421/U1008  ( .A(\DP_OP_751_130_6421/n1455 ), .B(
        \DP_OP_751_130_6421/n1401 ), .CI(\DP_OP_751_130_6421/n1454 ), .CO(
        \DP_OP_751_130_6421/n1355 ), .S(\DP_OP_751_130_6421/n1356 ) );
  FA_X1 \DP_OP_751_130_6421/U1007  ( .A(\DP_OP_751_130_6421/n1453 ), .B(
        \DP_OP_751_130_6421/n1400 ), .CI(\DP_OP_751_130_6421/n1452 ), .CO(
        \DP_OP_751_130_6421/n1353 ), .S(\DP_OP_751_130_6421/n1354 ) );
  FA_X1 \DP_OP_751_130_6421/U1006  ( .A(\DP_OP_751_130_6421/n1451 ), .B(
        \DP_OP_751_130_6421/n1399 ), .CI(\DP_OP_751_130_6421/n1450 ), .CO(
        \DP_OP_751_130_6421/n1351 ), .S(\DP_OP_751_130_6421/n1352 ) );
  FA_X1 \DP_OP_751_130_6421/U1005  ( .A(\DP_OP_751_130_6421/n1449 ), .B(
        \DP_OP_751_130_6421/n1398 ), .CI(\DP_OP_751_130_6421/n1448 ), .CO(
        \DP_OP_751_130_6421/n1349 ), .S(\DP_OP_751_130_6421/n1350 ) );
  FA_X1 \DP_OP_751_130_6421/U1004  ( .A(\DP_OP_751_130_6421/n1447 ), .B(
        \DP_OP_751_130_6421/n1397 ), .CI(\DP_OP_751_130_6421/n1446 ), .CO(
        \DP_OP_751_130_6421/n1347 ), .S(\DP_OP_751_130_6421/n1348 ) );
  FA_X1 \DP_OP_751_130_6421/U1003  ( .A(\DP_OP_751_130_6421/n1445 ), .B(
        \DP_OP_751_130_6421/n1396 ), .CI(\DP_OP_751_130_6421/n1444 ), .CO(
        \DP_OP_751_130_6421/n1345 ), .S(\DP_OP_751_130_6421/n1346 ) );
  FA_X1 \DP_OP_751_130_6421/U1002  ( .A(\DP_OP_751_130_6421/n1443 ), .B(
        \DP_OP_751_130_6421/n1395 ), .CI(\DP_OP_751_130_6421/n1442 ), .CO(
        \DP_OP_751_130_6421/n1343 ), .S(\DP_OP_751_130_6421/n1344 ) );
  FA_X1 \DP_OP_751_130_6421/U1001  ( .A(\DP_OP_751_130_6421/n1441 ), .B(
        \DP_OP_751_130_6421/n1394 ), .CI(\DP_OP_751_130_6421/n1440 ), .CO(
        \DP_OP_751_130_6421/n1341 ), .S(\DP_OP_751_130_6421/n1342 ) );
  FA_X1 \DP_OP_751_130_6421/U1000  ( .A(\DP_OP_751_130_6421/n1439 ), .B(
        \DP_OP_751_130_6421/n1393 ), .CI(\DP_OP_751_130_6421/n1438 ), .CO(
        \DP_OP_751_130_6421/n1339 ), .S(\DP_OP_751_130_6421/n1340 ) );
  FA_X1 \DP_OP_751_130_6421/U999  ( .A(\DP_OP_751_130_6421/n1437 ), .B(
        \DP_OP_751_130_6421/n1392 ), .CI(\DP_OP_751_130_6421/n1436 ), .CO(
        \DP_OP_751_130_6421/n1337 ), .S(\DP_OP_751_130_6421/n1338 ) );
  FA_X1 \DP_OP_751_130_6421/U998  ( .A(\DP_OP_751_130_6421/n1435 ), .B(
        \DP_OP_751_130_6421/n1391 ), .CI(\DP_OP_751_130_6421/n1434 ), .CO(
        \DP_OP_751_130_6421/n1335 ), .S(\DP_OP_751_130_6421/n1336 ) );
  FA_X1 \DP_OP_751_130_6421/U996  ( .A(\DP_OP_751_130_6421/n1431 ), .B(
        \DP_OP_751_130_6421/n1389 ), .CI(\DP_OP_751_130_6421/n1430 ), .S(
        \DP_OP_751_130_6421/n1332 ) );
  FA_X1 \DP_OP_751_130_6421/U949  ( .A(\DP_OP_751_130_6421/n1310 ), .B(n8055), 
        .CI(\DP_OP_751_130_6421/n1375 ), .CO(\DP_OP_751_130_6421/n1275 ), .S(
        \DP_OP_751_130_6421/n1276 ) );
  FA_X1 \DP_OP_751_130_6421/U948  ( .A(\DP_OP_751_130_6421/n1373 ), .B(
        \DP_OP_751_130_6421/n1309 ), .CI(\DP_OP_751_130_6421/n1372 ), .CO(
        \DP_OP_751_130_6421/n1273 ), .S(\DP_OP_751_130_6421/n1274 ) );
  FA_X1 \DP_OP_751_130_6421/U947  ( .A(\DP_OP_751_130_6421/n1371 ), .B(
        \DP_OP_751_130_6421/n1308 ), .CI(\DP_OP_751_130_6421/n1370 ), .CO(
        \DP_OP_751_130_6421/n1271 ), .S(\DP_OP_751_130_6421/n1272 ) );
  FA_X1 \DP_OP_751_130_6421/U946  ( .A(\DP_OP_751_130_6421/n1369 ), .B(
        \DP_OP_751_130_6421/n1307 ), .CI(\DP_OP_751_130_6421/n1368 ), .CO(
        \DP_OP_751_130_6421/n1269 ), .S(\DP_OP_751_130_6421/n1270 ) );
  FA_X1 \DP_OP_751_130_6421/U945  ( .A(\DP_OP_751_130_6421/n1367 ), .B(
        \DP_OP_751_130_6421/n1306 ), .CI(\DP_OP_751_130_6421/n1366 ), .CO(
        \DP_OP_751_130_6421/n1267 ), .S(\DP_OP_751_130_6421/n1268 ) );
  FA_X1 \DP_OP_751_130_6421/U944  ( .A(\DP_OP_751_130_6421/n1365 ), .B(
        \DP_OP_751_130_6421/n1305 ), .CI(\DP_OP_751_130_6421/n1364 ), .CO(
        \DP_OP_751_130_6421/n1265 ), .S(\DP_OP_751_130_6421/n1266 ) );
  FA_X1 \DP_OP_751_130_6421/U943  ( .A(\DP_OP_751_130_6421/n1363 ), .B(
        \DP_OP_751_130_6421/n1304 ), .CI(\DP_OP_751_130_6421/n1362 ), .CO(
        \DP_OP_751_130_6421/n1263 ), .S(\DP_OP_751_130_6421/n1264 ) );
  FA_X1 \DP_OP_751_130_6421/U942  ( .A(\DP_OP_751_130_6421/n1361 ), .B(
        \DP_OP_751_130_6421/n1303 ), .CI(\DP_OP_751_130_6421/n1360 ), .CO(
        \DP_OP_751_130_6421/n1261 ), .S(\DP_OP_751_130_6421/n1262 ) );
  FA_X1 \DP_OP_751_130_6421/U941  ( .A(\DP_OP_751_130_6421/n1359 ), .B(
        \DP_OP_751_130_6421/n1302 ), .CI(\DP_OP_751_130_6421/n1358 ), .CO(
        \DP_OP_751_130_6421/n1259 ), .S(\DP_OP_751_130_6421/n1260 ) );
  FA_X1 \DP_OP_751_130_6421/U940  ( .A(\DP_OP_751_130_6421/n1357 ), .B(
        \DP_OP_751_130_6421/n1301 ), .CI(\DP_OP_751_130_6421/n1356 ), .CO(
        \DP_OP_751_130_6421/n1257 ), .S(\DP_OP_751_130_6421/n1258 ) );
  FA_X1 \DP_OP_751_130_6421/U939  ( .A(\DP_OP_751_130_6421/n1355 ), .B(
        \DP_OP_751_130_6421/n1300 ), .CI(\DP_OP_751_130_6421/n1354 ), .CO(
        \DP_OP_751_130_6421/n1255 ), .S(\DP_OP_751_130_6421/n1256 ) );
  FA_X1 \DP_OP_751_130_6421/U938  ( .A(\DP_OP_751_130_6421/n1353 ), .B(
        \DP_OP_751_130_6421/n1299 ), .CI(\DP_OP_751_130_6421/n1352 ), .CO(
        \DP_OP_751_130_6421/n1253 ), .S(\DP_OP_751_130_6421/n1254 ) );
  FA_X1 \DP_OP_751_130_6421/U937  ( .A(\DP_OP_751_130_6421/n1351 ), .B(
        \DP_OP_751_130_6421/n1298 ), .CI(\DP_OP_751_130_6421/n1350 ), .CO(
        \DP_OP_751_130_6421/n1251 ), .S(\DP_OP_751_130_6421/n1252 ) );
  FA_X1 \DP_OP_751_130_6421/U936  ( .A(\DP_OP_751_130_6421/n1349 ), .B(
        \DP_OP_751_130_6421/n1297 ), .CI(\DP_OP_751_130_6421/n1348 ), .CO(
        \DP_OP_751_130_6421/n1249 ), .S(\DP_OP_751_130_6421/n1250 ) );
  FA_X1 \DP_OP_751_130_6421/U935  ( .A(\DP_OP_751_130_6421/n1347 ), .B(
        \DP_OP_751_130_6421/n1296 ), .CI(\DP_OP_751_130_6421/n1346 ), .CO(
        \DP_OP_751_130_6421/n1247 ), .S(\DP_OP_751_130_6421/n1248 ) );
  FA_X1 \DP_OP_751_130_6421/U934  ( .A(\DP_OP_751_130_6421/n1345 ), .B(
        \DP_OP_751_130_6421/n1295 ), .CI(\DP_OP_751_130_6421/n1344 ), .CO(
        \DP_OP_751_130_6421/n1245 ), .S(\DP_OP_751_130_6421/n1246 ) );
  FA_X1 \DP_OP_751_130_6421/U933  ( .A(\DP_OP_751_130_6421/n1343 ), .B(
        \DP_OP_751_130_6421/n1294 ), .CI(\DP_OP_751_130_6421/n1342 ), .CO(
        \DP_OP_751_130_6421/n1243 ), .S(\DP_OP_751_130_6421/n1244 ) );
  FA_X1 \DP_OP_751_130_6421/U932  ( .A(\DP_OP_751_130_6421/n1341 ), .B(
        \DP_OP_751_130_6421/n1293 ), .CI(\DP_OP_751_130_6421/n1340 ), .CO(
        \DP_OP_751_130_6421/n1241 ), .S(\DP_OP_751_130_6421/n1242 ) );
  FA_X1 \DP_OP_751_130_6421/U931  ( .A(\DP_OP_751_130_6421/n1339 ), .B(
        \DP_OP_751_130_6421/n1292 ), .CI(\DP_OP_751_130_6421/n1338 ), .CO(
        \DP_OP_751_130_6421/n1239 ), .S(\DP_OP_751_130_6421/n1240 ) );
  FA_X1 \DP_OP_751_130_6421/U930  ( .A(\DP_OP_751_130_6421/n1337 ), .B(
        \DP_OP_751_130_6421/n1291 ), .CI(\DP_OP_751_130_6421/n1336 ), .CO(
        \DP_OP_751_130_6421/n1237 ), .S(\DP_OP_751_130_6421/n1238 ) );
  FA_X1 \DP_OP_751_130_6421/U929  ( .A(\DP_OP_751_130_6421/n1335 ), .B(
        \DP_OP_751_130_6421/n1290 ), .CI(\DP_OP_751_130_6421/n1334 ), .CO(
        \DP_OP_751_130_6421/n1235 ), .S(\DP_OP_751_130_6421/n1236 ) );
  FA_X1 \DP_OP_751_130_6421/U928  ( .A(\DP_OP_751_130_6421/n1333 ), .B(
        \DP_OP_751_130_6421/n1289 ), .CI(\DP_OP_751_130_6421/n1332 ), .S(
        \DP_OP_751_130_6421/n1234 ) );
  FA_X1 \DP_OP_751_130_6421/U878  ( .A(\DP_OP_751_130_6421/n1271 ), .B(
        \DP_OP_751_130_6421/n1207 ), .CI(\DP_OP_751_130_6421/n1270 ), .CO(
        \DP_OP_751_130_6421/n1171 ), .S(\DP_OP_751_130_6421/n1172 ) );
  FA_X1 \DP_OP_751_130_6421/U877  ( .A(\DP_OP_751_130_6421/n1269 ), .B(
        \DP_OP_751_130_6421/n1206 ), .CI(\DP_OP_751_130_6421/n1268 ), .CO(
        \DP_OP_751_130_6421/n1169 ), .S(\DP_OP_751_130_6421/n1170 ) );
  FA_X1 \DP_OP_751_130_6421/U876  ( .A(\DP_OP_751_130_6421/n1267 ), .B(
        \DP_OP_751_130_6421/n1205 ), .CI(\DP_OP_751_130_6421/n1266 ), .CO(
        \DP_OP_751_130_6421/n1167 ), .S(\DP_OP_751_130_6421/n1168 ) );
  FA_X1 \DP_OP_751_130_6421/U875  ( .A(\DP_OP_751_130_6421/n1265 ), .B(
        \DP_OP_751_130_6421/n1204 ), .CI(\DP_OP_751_130_6421/n1264 ), .CO(
        \DP_OP_751_130_6421/n1165 ), .S(\DP_OP_751_130_6421/n1166 ) );
  FA_X1 \DP_OP_751_130_6421/U874  ( .A(\DP_OP_751_130_6421/n1263 ), .B(
        \DP_OP_751_130_6421/n1203 ), .CI(\DP_OP_751_130_6421/n1262 ), .CO(
        \DP_OP_751_130_6421/n1163 ), .S(\DP_OP_751_130_6421/n1164 ) );
  FA_X1 \DP_OP_751_130_6421/U873  ( .A(\DP_OP_751_130_6421/n1261 ), .B(
        \DP_OP_751_130_6421/n1202 ), .CI(\DP_OP_751_130_6421/n1260 ), .CO(
        \DP_OP_751_130_6421/n1161 ), .S(\DP_OP_751_130_6421/n1162 ) );
  FA_X1 \DP_OP_751_130_6421/U872  ( .A(\DP_OP_751_130_6421/n1259 ), .B(
        \DP_OP_751_130_6421/n1201 ), .CI(\DP_OP_751_130_6421/n1258 ), .CO(
        \DP_OP_751_130_6421/n1159 ), .S(\DP_OP_751_130_6421/n1160 ) );
  FA_X1 \DP_OP_751_130_6421/U871  ( .A(\DP_OP_751_130_6421/n1257 ), .B(
        \DP_OP_751_130_6421/n1200 ), .CI(\DP_OP_751_130_6421/n1256 ), .CO(
        \DP_OP_751_130_6421/n1157 ), .S(\DP_OP_751_130_6421/n1158 ) );
  FA_X1 \DP_OP_751_130_6421/U869  ( .A(\DP_OP_751_130_6421/n1253 ), .B(
        \DP_OP_751_130_6421/n1198 ), .CI(\DP_OP_751_130_6421/n1252 ), .CO(
        \DP_OP_751_130_6421/n1153 ), .S(\DP_OP_751_130_6421/n1154 ) );
  FA_X1 \DP_OP_751_130_6421/U868  ( .A(\DP_OP_751_130_6421/n1251 ), .B(
        \DP_OP_751_130_6421/n1197 ), .CI(\DP_OP_751_130_6421/n1250 ), .CO(
        \DP_OP_751_130_6421/n1151 ), .S(\DP_OP_751_130_6421/n1152 ) );
  FA_X1 \DP_OP_751_130_6421/U867  ( .A(\DP_OP_751_130_6421/n1249 ), .B(
        \DP_OP_751_130_6421/n1196 ), .CI(\DP_OP_751_130_6421/n1248 ), .CO(
        \DP_OP_751_130_6421/n1149 ), .S(\DP_OP_751_130_6421/n1150 ) );
  FA_X1 \DP_OP_751_130_6421/U866  ( .A(\DP_OP_751_130_6421/n1247 ), .B(
        \DP_OP_751_130_6421/n1195 ), .CI(\DP_OP_751_130_6421/n1246 ), .CO(
        \DP_OP_751_130_6421/n1147 ), .S(\DP_OP_751_130_6421/n1148 ) );
  FA_X1 \DP_OP_751_130_6421/U865  ( .A(\DP_OP_751_130_6421/n1245 ), .B(
        \DP_OP_751_130_6421/n1194 ), .CI(\DP_OP_751_130_6421/n1244 ), .CO(
        \DP_OP_751_130_6421/n1145 ), .S(\DP_OP_751_130_6421/n1146 ) );
  FA_X1 \DP_OP_751_130_6421/U864  ( .A(\DP_OP_751_130_6421/n1243 ), .B(
        \DP_OP_751_130_6421/n1193 ), .CI(\DP_OP_751_130_6421/n1242 ), .CO(
        \DP_OP_751_130_6421/n1143 ), .S(\DP_OP_751_130_6421/n1144 ) );
  FA_X1 \DP_OP_751_130_6421/U863  ( .A(\DP_OP_751_130_6421/n1241 ), .B(
        \DP_OP_751_130_6421/n1192 ), .CI(\DP_OP_751_130_6421/n1240 ), .CO(
        \DP_OP_751_130_6421/n1141 ), .S(\DP_OP_751_130_6421/n1142 ) );
  FA_X1 \DP_OP_751_130_6421/U862  ( .A(\DP_OP_751_130_6421/n1239 ), .B(
        \DP_OP_751_130_6421/n1191 ), .CI(\DP_OP_751_130_6421/n1238 ), .CO(
        \DP_OP_751_130_6421/n1139 ), .S(\DP_OP_751_130_6421/n1140 ) );
  FA_X1 \DP_OP_751_130_6421/U861  ( .A(\DP_OP_751_130_6421/n1237 ), .B(
        \DP_OP_751_130_6421/n1190 ), .CI(\DP_OP_751_130_6421/n1236 ), .CO(
        \DP_OP_751_130_6421/n1137 ), .S(\DP_OP_751_130_6421/n1138 ) );
  FA_X1 \DP_OP_751_130_6421/U860  ( .A(\DP_OP_751_130_6421/n1235 ), .B(
        \DP_OP_751_130_6421/n1189 ), .CI(\DP_OP_751_130_6421/n1234 ), .S(
        \DP_OP_751_130_6421/n1136 ) );
  FA_X1 \DP_OP_751_130_6421/U808  ( .A(\DP_OP_751_130_6421/n1169 ), .B(
        \DP_OP_751_130_6421/n1105 ), .CI(\DP_OP_751_130_6421/n1168 ), .CO(
        \DP_OP_751_130_6421/n1069 ), .S(\DP_OP_751_130_6421/n1070 ) );
  FA_X1 \DP_OP_751_130_6421/U807  ( .A(\DP_OP_751_130_6421/n1167 ), .B(
        \DP_OP_751_130_6421/n1104 ), .CI(\DP_OP_751_130_6421/n1166 ), .CO(
        \DP_OP_751_130_6421/n1067 ), .S(\DP_OP_751_130_6421/n1068 ) );
  FA_X1 \DP_OP_751_130_6421/U806  ( .A(\DP_OP_751_130_6421/n1165 ), .B(
        \DP_OP_751_130_6421/n1103 ), .CI(\DP_OP_751_130_6421/n1164 ), .CO(
        \DP_OP_751_130_6421/n1065 ), .S(\DP_OP_751_130_6421/n1066 ) );
  FA_X1 \DP_OP_751_130_6421/U805  ( .A(\DP_OP_751_130_6421/n1163 ), .B(
        \DP_OP_751_130_6421/n1102 ), .CI(\DP_OP_751_130_6421/n1162 ), .CO(
        \DP_OP_751_130_6421/n1063 ), .S(\DP_OP_751_130_6421/n1064 ) );
  FA_X1 \DP_OP_751_130_6421/U804  ( .A(\DP_OP_751_130_6421/n1161 ), .B(
        \DP_OP_751_130_6421/n1101 ), .CI(\DP_OP_751_130_6421/n1160 ), .CO(
        \DP_OP_751_130_6421/n1061 ), .S(\DP_OP_751_130_6421/n1062 ) );
  FA_X1 \DP_OP_751_130_6421/U803  ( .A(\DP_OP_751_130_6421/n1159 ), .B(
        \DP_OP_751_130_6421/n1100 ), .CI(\DP_OP_751_130_6421/n1158 ), .CO(
        \DP_OP_751_130_6421/n1059 ), .S(\DP_OP_751_130_6421/n1060 ) );
  FA_X1 \DP_OP_751_130_6421/U802  ( .A(\DP_OP_751_130_6421/n1157 ), .B(
        \DP_OP_751_130_6421/n1099 ), .CI(\DP_OP_751_130_6421/n1156 ), .CO(
        \DP_OP_751_130_6421/n1057 ), .S(\DP_OP_751_130_6421/n1058 ) );
  FA_X1 \DP_OP_751_130_6421/U801  ( .A(\DP_OP_751_130_6421/n1155 ), .B(
        \DP_OP_751_130_6421/n1098 ), .CI(\DP_OP_751_130_6421/n1154 ), .CO(
        \DP_OP_751_130_6421/n1055 ), .S(\DP_OP_751_130_6421/n1056 ) );
  FA_X1 \DP_OP_751_130_6421/U800  ( .A(\DP_OP_751_130_6421/n1153 ), .B(
        \DP_OP_751_130_6421/n1097 ), .CI(\DP_OP_751_130_6421/n1152 ), .CO(
        \DP_OP_751_130_6421/n1053 ), .S(\DP_OP_751_130_6421/n1054 ) );
  FA_X1 \DP_OP_751_130_6421/U799  ( .A(\DP_OP_751_130_6421/n1151 ), .B(
        \DP_OP_751_130_6421/n1096 ), .CI(\DP_OP_751_130_6421/n1150 ), .CO(
        \DP_OP_751_130_6421/n1051 ), .S(\DP_OP_751_130_6421/n1052 ) );
  FA_X1 \DP_OP_751_130_6421/U798  ( .A(\DP_OP_751_130_6421/n1149 ), .B(
        \DP_OP_751_130_6421/n1095 ), .CI(\DP_OP_751_130_6421/n1148 ), .CO(
        \DP_OP_751_130_6421/n1049 ), .S(\DP_OP_751_130_6421/n1050 ) );
  FA_X1 \DP_OP_751_130_6421/U797  ( .A(\DP_OP_751_130_6421/n1147 ), .B(
        \DP_OP_751_130_6421/n1094 ), .CI(\DP_OP_751_130_6421/n1146 ), .CO(
        \DP_OP_751_130_6421/n1047 ), .S(\DP_OP_751_130_6421/n1048 ) );
  FA_X1 \DP_OP_751_130_6421/U796  ( .A(\DP_OP_751_130_6421/n1145 ), .B(
        \DP_OP_751_130_6421/n1093 ), .CI(\DP_OP_751_130_6421/n1144 ), .CO(
        \DP_OP_751_130_6421/n1045 ), .S(\DP_OP_751_130_6421/n1046 ) );
  FA_X1 \DP_OP_751_130_6421/U795  ( .A(\DP_OP_751_130_6421/n1143 ), .B(
        \DP_OP_751_130_6421/n1092 ), .CI(\DP_OP_751_130_6421/n1142 ), .CO(
        \DP_OP_751_130_6421/n1043 ), .S(\DP_OP_751_130_6421/n1044 ) );
  FA_X1 \DP_OP_751_130_6421/U794  ( .A(\DP_OP_751_130_6421/n1141 ), .B(
        \DP_OP_751_130_6421/n1091 ), .CI(\DP_OP_751_130_6421/n1140 ), .CO(
        \DP_OP_751_130_6421/n1041 ), .S(\DP_OP_751_130_6421/n1042 ) );
  FA_X1 \DP_OP_751_130_6421/U793  ( .A(\DP_OP_751_130_6421/n1139 ), .B(
        \DP_OP_751_130_6421/n1090 ), .CI(\DP_OP_751_130_6421/n1138 ), .CO(
        \DP_OP_751_130_6421/n1039 ), .S(\DP_OP_751_130_6421/n1040 ) );
  FA_X1 \DP_OP_751_130_6421/U792  ( .A(\DP_OP_751_130_6421/n1137 ), .B(
        \DP_OP_751_130_6421/n1089 ), .CI(\DP_OP_751_130_6421/n1136 ), .S(
        \DP_OP_751_130_6421/n1038 ) );
  FA_X1 \DP_OP_751_130_6421/U738  ( .A(\DP_OP_751_130_6421/n1067 ), .B(
        \DP_OP_751_130_6421/n1003 ), .CI(\DP_OP_751_130_6421/n1066 ), .CO(
        \DP_OP_751_130_6421/n967 ), .S(\DP_OP_751_130_6421/n968 ) );
  FA_X1 \DP_OP_751_130_6421/U737  ( .A(\DP_OP_751_130_6421/n1065 ), .B(
        \DP_OP_751_130_6421/n1002 ), .CI(\DP_OP_751_130_6421/n1064 ), .CO(
        \DP_OP_751_130_6421/n965 ), .S(\DP_OP_751_130_6421/n966 ) );
  FA_X1 \DP_OP_751_130_6421/U736  ( .A(\DP_OP_751_130_6421/n1063 ), .B(
        \DP_OP_751_130_6421/n1001 ), .CI(\DP_OP_751_130_6421/n1062 ), .CO(
        \DP_OP_751_130_6421/n963 ), .S(\DP_OP_751_130_6421/n964 ) );
  FA_X1 \DP_OP_751_130_6421/U735  ( .A(\DP_OP_751_130_6421/n1061 ), .B(
        \DP_OP_751_130_6421/n1000 ), .CI(\DP_OP_751_130_6421/n1060 ), .CO(
        \DP_OP_751_130_6421/n961 ), .S(\DP_OP_751_130_6421/n962 ) );
  FA_X1 \DP_OP_751_130_6421/U734  ( .A(\DP_OP_751_130_6421/n1059 ), .B(
        \DP_OP_751_130_6421/n999 ), .CI(\DP_OP_751_130_6421/n1058 ), .CO(
        \DP_OP_751_130_6421/n959 ), .S(\DP_OP_751_130_6421/n960 ) );
  FA_X1 \DP_OP_751_130_6421/U733  ( .A(\DP_OP_751_130_6421/n1057 ), .B(
        \DP_OP_751_130_6421/n998 ), .CI(\DP_OP_751_130_6421/n1056 ), .CO(
        \DP_OP_751_130_6421/n957 ), .S(\DP_OP_751_130_6421/n958 ) );
  FA_X1 \DP_OP_751_130_6421/U732  ( .A(\DP_OP_751_130_6421/n1055 ), .B(
        \DP_OP_751_130_6421/n997 ), .CI(\DP_OP_751_130_6421/n1054 ), .CO(
        \DP_OP_751_130_6421/n955 ), .S(\DP_OP_751_130_6421/n956 ) );
  FA_X1 \DP_OP_751_130_6421/U731  ( .A(\DP_OP_751_130_6421/n1053 ), .B(
        \DP_OP_751_130_6421/n996 ), .CI(\DP_OP_751_130_6421/n1052 ), .CO(
        \DP_OP_751_130_6421/n953 ), .S(\DP_OP_751_130_6421/n954 ) );
  FA_X1 \DP_OP_751_130_6421/U730  ( .A(\DP_OP_751_130_6421/n1051 ), .B(
        \DP_OP_751_130_6421/n995 ), .CI(\DP_OP_751_130_6421/n1050 ), .CO(
        \DP_OP_751_130_6421/n951 ), .S(\DP_OP_751_130_6421/n952 ) );
  FA_X1 \DP_OP_751_130_6421/U729  ( .A(\DP_OP_751_130_6421/n1049 ), .B(
        \DP_OP_751_130_6421/n994 ), .CI(\DP_OP_751_130_6421/n1048 ), .CO(
        \DP_OP_751_130_6421/n949 ), .S(\DP_OP_751_130_6421/n950 ) );
  FA_X1 \DP_OP_751_130_6421/U728  ( .A(\DP_OP_751_130_6421/n1047 ), .B(
        \DP_OP_751_130_6421/n993 ), .CI(\DP_OP_751_130_6421/n1046 ), .CO(
        \DP_OP_751_130_6421/n947 ), .S(\DP_OP_751_130_6421/n948 ) );
  FA_X1 \DP_OP_751_130_6421/U727  ( .A(\DP_OP_751_130_6421/n1045 ), .B(
        \DP_OP_751_130_6421/n992 ), .CI(\DP_OP_751_130_6421/n1044 ), .CO(
        \DP_OP_751_130_6421/n945 ), .S(\DP_OP_751_130_6421/n946 ) );
  FA_X1 \DP_OP_751_130_6421/U726  ( .A(\DP_OP_751_130_6421/n1043 ), .B(
        \DP_OP_751_130_6421/n991 ), .CI(\DP_OP_751_130_6421/n1042 ), .CO(
        \DP_OP_751_130_6421/n943 ), .S(\DP_OP_751_130_6421/n944 ) );
  FA_X1 \DP_OP_751_130_6421/U725  ( .A(\DP_OP_751_130_6421/n1041 ), .B(
        \DP_OP_751_130_6421/n990 ), .CI(\DP_OP_751_130_6421/n1040 ), .CO(
        \DP_OP_751_130_6421/n941 ), .S(\DP_OP_751_130_6421/n942 ) );
  FA_X1 \DP_OP_751_130_6421/U724  ( .A(\DP_OP_751_130_6421/n1039 ), .B(
        \DP_OP_751_130_6421/n989 ), .CI(\DP_OP_751_130_6421/n1038 ), .S(
        \DP_OP_751_130_6421/n940 ) );
  FA_X1 \DP_OP_751_130_6421/U668  ( .A(\DP_OP_751_130_6421/n965 ), .B(
        \DP_OP_751_130_6421/n901 ), .CI(\DP_OP_751_130_6421/n964 ), .CO(
        \DP_OP_751_130_6421/n865 ), .S(\DP_OP_751_130_6421/n866 ) );
  FA_X1 \DP_OP_751_130_6421/U667  ( .A(\DP_OP_751_130_6421/n963 ), .B(
        \DP_OP_751_130_6421/n900 ), .CI(\DP_OP_751_130_6421/n962 ), .CO(
        \DP_OP_751_130_6421/n863 ), .S(\DP_OP_751_130_6421/n864 ) );
  FA_X1 \DP_OP_751_130_6421/U666  ( .A(\DP_OP_751_130_6421/n961 ), .B(
        \DP_OP_751_130_6421/n899 ), .CI(\DP_OP_751_130_6421/n960 ), .CO(
        \DP_OP_751_130_6421/n861 ), .S(\DP_OP_751_130_6421/n862 ) );
  FA_X1 \DP_OP_751_130_6421/U665  ( .A(\DP_OP_751_130_6421/n959 ), .B(
        \DP_OP_751_130_6421/n898 ), .CI(\DP_OP_751_130_6421/n958 ), .CO(
        \DP_OP_751_130_6421/n859 ), .S(\DP_OP_751_130_6421/n860 ) );
  FA_X1 \DP_OP_751_130_6421/U664  ( .A(\DP_OP_751_130_6421/n957 ), .B(
        \DP_OP_751_130_6421/n897 ), .CI(\DP_OP_751_130_6421/n956 ), .CO(
        \DP_OP_751_130_6421/n857 ), .S(\DP_OP_751_130_6421/n858 ) );
  FA_X1 \DP_OP_751_130_6421/U663  ( .A(\DP_OP_751_130_6421/n955 ), .B(
        \DP_OP_751_130_6421/n896 ), .CI(\DP_OP_751_130_6421/n954 ), .CO(
        \DP_OP_751_130_6421/n855 ), .S(\DP_OP_751_130_6421/n856 ) );
  FA_X1 \DP_OP_751_130_6421/U662  ( .A(\DP_OP_751_130_6421/n953 ), .B(
        \DP_OP_751_130_6421/n895 ), .CI(\DP_OP_751_130_6421/n952 ), .CO(
        \DP_OP_751_130_6421/n853 ), .S(\DP_OP_751_130_6421/n854 ) );
  FA_X1 \DP_OP_751_130_6421/U661  ( .A(\DP_OP_751_130_6421/n951 ), .B(
        \DP_OP_751_130_6421/n894 ), .CI(\DP_OP_751_130_6421/n950 ), .CO(
        \DP_OP_751_130_6421/n851 ), .S(\DP_OP_751_130_6421/n852 ) );
  FA_X1 \DP_OP_751_130_6421/U660  ( .A(\DP_OP_751_130_6421/n949 ), .B(
        \DP_OP_751_130_6421/n893 ), .CI(\DP_OP_751_130_6421/n948 ), .CO(
        \DP_OP_751_130_6421/n849 ), .S(\DP_OP_751_130_6421/n850 ) );
  FA_X1 \DP_OP_751_130_6421/U659  ( .A(\DP_OP_751_130_6421/n947 ), .B(
        \DP_OP_751_130_6421/n892 ), .CI(\DP_OP_751_130_6421/n946 ), .CO(
        \DP_OP_751_130_6421/n847 ), .S(\DP_OP_751_130_6421/n848 ) );
  FA_X1 \DP_OP_751_130_6421/U658  ( .A(\DP_OP_751_130_6421/n945 ), .B(
        \DP_OP_751_130_6421/n891 ), .CI(\DP_OP_751_130_6421/n944 ), .CO(
        \DP_OP_751_130_6421/n845 ), .S(\DP_OP_751_130_6421/n846 ) );
  FA_X1 \DP_OP_751_130_6421/U657  ( .A(\DP_OP_751_130_6421/n943 ), .B(
        \DP_OP_751_130_6421/n890 ), .CI(\DP_OP_751_130_6421/n942 ), .CO(
        \DP_OP_751_130_6421/n843 ), .S(\DP_OP_751_130_6421/n844 ) );
  FA_X1 \DP_OP_751_130_6421/U656  ( .A(\DP_OP_751_130_6421/n941 ), .B(
        \DP_OP_751_130_6421/n889 ), .CI(\DP_OP_751_130_6421/n940 ), .S(
        \DP_OP_751_130_6421/n842 ) );
  FA_X1 \DP_OP_751_130_6421/U598  ( .A(\DP_OP_751_130_6421/n863 ), .B(
        \DP_OP_751_130_6421/n799 ), .CI(\DP_OP_751_130_6421/n862 ), .CO(
        \DP_OP_751_130_6421/n763 ), .S(\DP_OP_751_130_6421/n764 ) );
  FA_X1 \DP_OP_751_130_6421/U597  ( .A(\DP_OP_751_130_6421/n861 ), .B(
        \DP_OP_751_130_6421/n798 ), .CI(\DP_OP_751_130_6421/n860 ), .CO(
        \DP_OP_751_130_6421/n761 ), .S(\DP_OP_751_130_6421/n762 ) );
  FA_X1 \DP_OP_751_130_6421/U596  ( .A(\DP_OP_751_130_6421/n859 ), .B(
        \DP_OP_751_130_6421/n797 ), .CI(\DP_OP_751_130_6421/n858 ), .CO(
        \DP_OP_751_130_6421/n759 ), .S(\DP_OP_751_130_6421/n760 ) );
  FA_X1 \DP_OP_751_130_6421/U595  ( .A(\DP_OP_751_130_6421/n857 ), .B(
        \DP_OP_751_130_6421/n796 ), .CI(\DP_OP_751_130_6421/n856 ), .CO(
        \DP_OP_751_130_6421/n757 ), .S(\DP_OP_751_130_6421/n758 ) );
  FA_X1 \DP_OP_751_130_6421/U594  ( .A(\DP_OP_751_130_6421/n855 ), .B(
        \DP_OP_751_130_6421/n795 ), .CI(\DP_OP_751_130_6421/n854 ), .CO(
        \DP_OP_751_130_6421/n755 ), .S(\DP_OP_751_130_6421/n756 ) );
  FA_X1 \DP_OP_751_130_6421/U593  ( .A(\DP_OP_751_130_6421/n853 ), .B(
        \DP_OP_751_130_6421/n794 ), .CI(\DP_OP_751_130_6421/n852 ), .CO(
        \DP_OP_751_130_6421/n753 ), .S(\DP_OP_751_130_6421/n754 ) );
  FA_X1 \DP_OP_751_130_6421/U592  ( .A(\DP_OP_751_130_6421/n851 ), .B(
        \DP_OP_751_130_6421/n793 ), .CI(\DP_OP_751_130_6421/n850 ), .CO(
        \DP_OP_751_130_6421/n751 ), .S(\DP_OP_751_130_6421/n752 ) );
  FA_X1 \DP_OP_751_130_6421/U591  ( .A(\DP_OP_751_130_6421/n849 ), .B(
        \DP_OP_751_130_6421/n792 ), .CI(\DP_OP_751_130_6421/n848 ), .CO(
        \DP_OP_751_130_6421/n749 ), .S(\DP_OP_751_130_6421/n750 ) );
  FA_X1 \DP_OP_751_130_6421/U590  ( .A(\DP_OP_751_130_6421/n847 ), .B(
        \DP_OP_751_130_6421/n791 ), .CI(\DP_OP_751_130_6421/n846 ), .CO(
        \DP_OP_751_130_6421/n747 ), .S(\DP_OP_751_130_6421/n748 ) );
  FA_X1 \DP_OP_751_130_6421/U589  ( .A(\DP_OP_751_130_6421/n845 ), .B(
        \DP_OP_751_130_6421/n790 ), .CI(\DP_OP_751_130_6421/n844 ), .CO(
        \DP_OP_751_130_6421/n745 ), .S(\DP_OP_751_130_6421/n746 ) );
  FA_X1 \DP_OP_751_130_6421/U528  ( .A(\DP_OP_751_130_6421/n761 ), .B(
        \DP_OP_751_130_6421/n697 ), .CI(\DP_OP_751_130_6421/n760 ), .CO(
        \DP_OP_751_130_6421/n661 ), .S(\DP_OP_751_130_6421/n662 ) );
  FA_X1 \DP_OP_751_130_6421/U527  ( .A(\DP_OP_751_130_6421/n759 ), .B(
        \DP_OP_751_130_6421/n696 ), .CI(\DP_OP_751_130_6421/n758 ), .CO(
        \DP_OP_751_130_6421/n659 ), .S(\DP_OP_751_130_6421/n660 ) );
  FA_X1 \DP_OP_751_130_6421/U526  ( .A(\DP_OP_751_130_6421/n757 ), .B(
        \DP_OP_751_130_6421/n695 ), .CI(\DP_OP_751_130_6421/n756 ), .CO(
        \DP_OP_751_130_6421/n657 ), .S(\DP_OP_751_130_6421/n658 ) );
  FA_X1 \DP_OP_751_130_6421/U525  ( .A(\DP_OP_751_130_6421/n755 ), .B(
        \DP_OP_751_130_6421/n694 ), .CI(\DP_OP_751_130_6421/n754 ), .CO(
        \DP_OP_751_130_6421/n655 ), .S(\DP_OP_751_130_6421/n656 ) );
  FA_X1 \DP_OP_751_130_6421/U524  ( .A(\DP_OP_751_130_6421/n753 ), .B(
        \DP_OP_751_130_6421/n693 ), .CI(\DP_OP_751_130_6421/n752 ), .CO(
        \DP_OP_751_130_6421/n653 ), .S(\DP_OP_751_130_6421/n654 ) );
  FA_X1 \DP_OP_751_130_6421/U523  ( .A(\DP_OP_751_130_6421/n751 ), .B(
        \DP_OP_751_130_6421/n692 ), .CI(\DP_OP_751_130_6421/n750 ), .CO(
        \DP_OP_751_130_6421/n651 ), .S(\DP_OP_751_130_6421/n652 ) );
  FA_X1 \DP_OP_751_130_6421/U522  ( .A(\DP_OP_751_130_6421/n749 ), .B(
        \DP_OP_751_130_6421/n691 ), .CI(\DP_OP_751_130_6421/n748 ), .CO(
        \DP_OP_751_130_6421/n649 ), .S(\DP_OP_751_130_6421/n650 ) );
  FA_X1 \DP_OP_751_130_6421/U521  ( .A(\DP_OP_751_130_6421/n747 ), .B(
        \DP_OP_751_130_6421/n690 ), .CI(\DP_OP_751_130_6421/n746 ), .CO(
        \DP_OP_751_130_6421/n647 ), .S(\DP_OP_751_130_6421/n648 ) );
  FA_X1 \DP_OP_751_130_6421/U520  ( .A(\DP_OP_751_130_6421/n745 ), .B(
        \DP_OP_751_130_6421/n689 ), .CI(\DP_OP_751_130_6421/n744 ), .S(
        \DP_OP_751_130_6421/n646 ) );
  FA_X1 \DP_OP_751_130_6421/U458  ( .A(\DP_OP_751_130_6421/n659 ), .B(
        \DP_OP_751_130_6421/n595 ), .CI(\DP_OP_751_130_6421/n658 ), .CO(
        \DP_OP_751_130_6421/n559 ), .S(\DP_OP_751_130_6421/n560 ) );
  FA_X1 \DP_OP_751_130_6421/U457  ( .A(\DP_OP_751_130_6421/n657 ), .B(
        \DP_OP_751_130_6421/n594 ), .CI(\DP_OP_751_130_6421/n656 ), .CO(
        \DP_OP_751_130_6421/n557 ), .S(\DP_OP_751_130_6421/n558 ) );
  FA_X1 \DP_OP_751_130_6421/U456  ( .A(\DP_OP_751_130_6421/n655 ), .B(
        \DP_OP_751_130_6421/n593 ), .CI(\DP_OP_751_130_6421/n654 ), .CO(
        \DP_OP_751_130_6421/n555 ), .S(\DP_OP_751_130_6421/n556 ) );
  FA_X1 \DP_OP_751_130_6421/U455  ( .A(\DP_OP_751_130_6421/n653 ), .B(
        \DP_OP_751_130_6421/n592 ), .CI(\DP_OP_751_130_6421/n652 ), .CO(
        \DP_OP_751_130_6421/n553 ), .S(\DP_OP_751_130_6421/n554 ) );
  FA_X1 \DP_OP_751_130_6421/U454  ( .A(\DP_OP_751_130_6421/n651 ), .B(
        \DP_OP_751_130_6421/n591 ), .CI(\DP_OP_751_130_6421/n650 ), .CO(
        \DP_OP_751_130_6421/n551 ), .S(\DP_OP_751_130_6421/n552 ) );
  FA_X1 \DP_OP_751_130_6421/U453  ( .A(\DP_OP_751_130_6421/n649 ), .B(
        \DP_OP_751_130_6421/n590 ), .CI(\DP_OP_751_130_6421/n648 ), .CO(
        \DP_OP_751_130_6421/n549 ), .S(\DP_OP_751_130_6421/n550 ) );
  FA_X1 \DP_OP_751_130_6421/U452  ( .A(\DP_OP_751_130_6421/n647 ), .B(
        \DP_OP_751_130_6421/n589 ), .CI(\DP_OP_751_130_6421/n646 ), .S(
        \DP_OP_751_130_6421/n548 ) );
  FA_X1 \DP_OP_751_130_6421/U388  ( .A(\DP_OP_751_130_6421/n557 ), .B(
        \DP_OP_751_130_6421/n493 ), .CI(\DP_OP_751_130_6421/n556 ), .CO(
        \DP_OP_751_130_6421/n457 ), .S(\DP_OP_751_130_6421/n458 ) );
  FA_X1 \DP_OP_751_130_6421/U386  ( .A(\DP_OP_751_130_6421/n553 ), .B(
        \DP_OP_751_130_6421/n491 ), .CI(\DP_OP_751_130_6421/n552 ), .CO(
        \DP_OP_751_130_6421/n453 ), .S(\DP_OP_751_130_6421/n454 ) );
  FA_X1 \DP_OP_751_130_6421/U385  ( .A(\DP_OP_751_130_6421/n551 ), .B(
        \DP_OP_751_130_6421/n490 ), .CI(\DP_OP_751_130_6421/n550 ), .CO(
        \DP_OP_751_130_6421/n451 ), .S(\DP_OP_751_130_6421/n452 ) );
  FA_X1 \DP_OP_751_130_6421/U384  ( .A(\DP_OP_751_130_6421/n549 ), .B(
        \DP_OP_751_130_6421/n489 ), .CI(\DP_OP_751_130_6421/n548 ), .S(
        \DP_OP_751_130_6421/n450 ) );
  FA_X1 \DP_OP_751_130_6421/U318  ( .A(\DP_OP_751_130_6421/n455 ), .B(
        \DP_OP_751_130_6421/n391 ), .CI(\DP_OP_751_130_6421/n454 ), .CO(
        \DP_OP_751_130_6421/n355 ), .S(\DP_OP_751_130_6421/n356 ) );
  FA_X1 \DP_OP_751_130_6421/U317  ( .A(\DP_OP_751_130_6421/n453 ), .B(
        \DP_OP_751_130_6421/n390 ), .CI(\DP_OP_751_130_6421/n452 ), .CO(
        \DP_OP_751_130_6421/n353 ), .S(\DP_OP_751_130_6421/n354 ) );
  FA_X1 \DP_OP_751_130_6421/U316  ( .A(\DP_OP_751_130_6421/n451 ), .B(
        \DP_OP_751_130_6421/n389 ), .CI(\DP_OP_751_130_6421/n450 ), .S(
        \DP_OP_751_130_6421/n352 ) );
  DFF_X2 \DataPath/WRF_CUhw/curr_addr_reg[31]  ( .D(n8257), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[31] ) );
  DFFS_X1 \IR_reg[27]  ( .D(n10259), .CK(CLK), .SN(n8463), .Q(n8285), .QN(
        IR[27]) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[2]  ( .D(n7684), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[2] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[3]  ( .D(n7683), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[3] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[4]  ( .D(n7682), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[4] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[5]  ( .D(n7681), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[5] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[6]  ( .D(n7680), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[6] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[7]  ( .D(n7679), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[7] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[8]  ( .D(n7678), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[8] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[9]  ( .D(n7677), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[9] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[10]  ( .D(n7676), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[10] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[11]  ( .D(n7675), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[11] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[12]  ( .D(n7674), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[12] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[13]  ( .D(n7673), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[13] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[14]  ( .D(n7672), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[14] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[15]  ( .D(n7671), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[15] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[16]  ( .D(n7670), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[16] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[17]  ( .D(n7669), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[17] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[18]  ( .D(n7668), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[18] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[23]  ( .D(n7667), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[23] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[19]  ( .D(n7666), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[19] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[20]  ( .D(n7665), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[20] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[24]  ( .D(n7664), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[24] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[21]  ( .D(n7663), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[21] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[25]  ( .D(n7662), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[25] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[22]  ( .D(n7661), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[22] ), .QN(n8048) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[26]  ( .D(n7660), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[26] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[27]  ( .D(n7659), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[27] ) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[28]  ( .D(n7658), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[28] ) );
  DFFR_X1 \IR_reg[9]  ( .D(n7139), .CK(CLK), .RN(n8464), .Q(IR[9]), .QN(n8101)
         );
  DFFR_X1 \IR_reg[6]  ( .D(n40), .CK(CLK), .RN(n8468), .Q(IR[6]), .QN(n8107)
         );
  DFFR_X1 \IR_reg[2]  ( .D(n36), .CK(CLK), .RN(n8458), .Q(IR[2]), .QN(n8196)
         );
  DFFR_X1 \IR_reg[14]  ( .D(n7138), .CK(CLK), .RN(n8468), .Q(n8134), .QN(n184)
         );
  DFFR_X1 \IR_reg[3]  ( .D(n37), .CK(CLK), .RN(n8462), .Q(IR[3]), .QN(n8097)
         );
  DFFR_X1 \IR_reg[5]  ( .D(n39), .CK(CLK), .RN(n8465), .Q(IR[5]), .QN(n8096)
         );
  DFFR_X1 \IR_reg[4]  ( .D(n38), .CK(CLK), .RN(n8461), .Q(IR[4]), .QN(n7975)
         );
  DFFR_X1 \IR_reg[22]  ( .D(n7130), .CK(CLK), .RN(n8457), .Q(n8175), .QN(n176)
         );
  DFFR_X1 \IR_reg[21]  ( .D(n7131), .CK(CLK), .RN(n8470), .Q(n8176), .QN(n177)
         );
  DFFR_X1 \IR_reg[20]  ( .D(n7132), .CK(CLK), .RN(n8464), .Q(n8177), .QN(n178)
         );
  DFFR_X1 \IR_reg[19]  ( .D(n7133), .CK(CLK), .RN(n8457), .Q(n8184), .QN(n179)
         );
  DFFR_X1 \IR_reg[18]  ( .D(n7134), .CK(CLK), .RN(n8469), .Q(n8179), .QN(n180)
         );
  DFFR_X1 \IR_reg[15]  ( .D(n7137), .CK(CLK), .RN(n8462), .Q(n8205), .QN(n183)
         );
  DFFR_X1 \IR_reg[12]  ( .D(n43), .CK(CLK), .RN(n8466), .Q(n8100), .QN(n185)
         );
  DFFR_X1 \IR_reg[11]  ( .D(n42), .CK(CLK), .RN(n8461), .Q(n8099), .QN(n186)
         );
  DFFR_X1 \IR_reg[7]  ( .D(n41), .CK(CLK), .RN(n8457), .Q(IR[7]), .QN(n8098)
         );
  DFFR_X1 \IR_reg[1]  ( .D(n35), .CK(CLK), .RN(n8462), .Q(IR[1]), .QN(n8094)
         );
  DFFR_X1 \IR_reg[0]  ( .D(n34), .CK(CLK), .RN(n8467), .Q(IR[0]), .QN(n8086)
         );
  DFFR_X1 \PC_reg[9]  ( .D(n7047), .CK(CLK), .RN(n8470), .Q(IRAM_ADDRESS[9]), 
        .QN(n208) );
  DFFR_X1 \PC_reg[5]  ( .D(n7051), .CK(CLK), .RN(n8467), .Q(IRAM_ADDRESS[5]), 
        .QN(\intadd_1/A[4] ) );
  DFFR_X1 \PC_reg[4]  ( .D(n7052), .CK(CLK), .RN(n8458), .Q(IRAM_ADDRESS[4]), 
        .QN(\intadd_1/A[3] ) );
  DFFR_X1 \PC_reg[8]  ( .D(n7048), .CK(CLK), .RN(n8466), .Q(IRAM_ADDRESS[8]), 
        .QN(n8169) );
  DFFR_X1 \PC_reg[3]  ( .D(n7053), .CK(CLK), .RN(n8460), .Q(IRAM_ADDRESS[3]), 
        .QN(n8133) );
  DFFR_X1 \PC_reg[11]  ( .D(n7045), .CK(CLK), .RN(n8469), .Q(IRAM_ADDRESS[11]), 
        .QN(\intadd_0/A[0] ) );
  DFFR_X1 \PC_reg[7]  ( .D(n7049), .CK(CLK), .RN(n8463), .Q(IRAM_ADDRESS[7]), 
        .QN(n210) );
  DFFR_X1 \PC_reg[2]  ( .D(n7054), .CK(CLK), .RN(n8470), .Q(IRAM_ADDRESS[2]), 
        .QN(\intadd_1/A[1] ) );
  DFFR_X1 \PC_reg[1]  ( .D(n7055), .CK(CLK), .RN(n8465), .Q(IRAM_ADDRESS[1]), 
        .QN(\intadd_1/A[0] ) );
  DFFR_X1 \PC_reg[17]  ( .D(n7039), .CK(CLK), .RN(n8461), .Q(IRAM_ADDRESS[17]), 
        .QN(n8181) );
  DFFR_X1 \PC_reg[20]  ( .D(n7036), .CK(CLK), .RN(n8458), .Q(IRAM_ADDRESS[20])
         );
  DFFR_X1 \PC_reg[15]  ( .D(n7041), .CK(CLK), .RN(n8459), .Q(IRAM_ADDRESS[15]), 
        .QN(n8125) );
  DFFR_X1 \PC_reg[12]  ( .D(n7044), .CK(CLK), .RN(n8463), .Q(IRAM_ADDRESS[12]), 
        .QN(n8128) );
  DFFR_X1 \PC_reg[13]  ( .D(n7043), .CK(CLK), .RN(n8462), .Q(IRAM_ADDRESS[13]), 
        .QN(n8127) );
  DFFR_X1 \PC_reg[19]  ( .D(n7037), .CK(CLK), .RN(n8460), .Q(IRAM_ADDRESS[19]), 
        .QN(n8180) );
  DFFR_X1 \PC_reg[14]  ( .D(n7042), .CK(CLK), .RN(n8468), .Q(IRAM_ADDRESS[14]), 
        .QN(n8126) );
  DFFR_X1 \PC_reg[26]  ( .D(n7030), .CK(CLK), .RN(n8469), .Q(IRAM_ADDRESS[26]), 
        .QN(n8103) );
  DFFR_X1 \PC_reg[27]  ( .D(n7029), .CK(CLK), .RN(n8469), .Q(IRAM_ADDRESS[27]), 
        .QN(n8185) );
  DFFR_X1 \PC_reg[28]  ( .D(n7028), .CK(CLK), .RN(n8464), .Q(IRAM_ADDRESS[28]), 
        .QN(n8178) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[15]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N61 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[15] ), .QN(n8224) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[4]  ( .D(n11557), .CK(CLK), .Q(n8166), .QN(\DECODEhw/i_tickcounter[4] ) );
  DFF_X1 \CU_I/CW_MEM_reg[MEM_EN]  ( .D(n7094), .CK(CLK), .Q(
        \CU_I/CW_MEM[MEM_EN] ), .QN(n8278) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[0]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N46 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[0] ), .QN(n8212) );
  DFF_X1 \DataPath/REG_B/Q_reg[4]  ( .D(n7075), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_B[4] ), .QN(n8209) );
  DFF_X1 \DataPath/REG_B/Q_reg[6]  ( .D(n7074), .CK(CLK), .Q(n8140), .QN(n481)
         );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[15]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N61 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[15] ), .QN(n8172) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_state_reg[0]  ( .D(n7058), .CK(CLK), 
        .Q(n8207), .QN(n877) );
  DFF_X1 \DataPath/RF/PUSH_ADDRGEN/curr_addr_reg[0]  ( .D(
        \DataPath/RF/PUSH_ADDRGEN/N46 ), .CK(CLK), .Q(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[0] ), .QN(n8210) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[27]  ( .D(n6829), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[123] ), .QN(n701) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[25]  ( .D(n6831), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[121] ), .QN(n699) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[24]  ( .D(n6832), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[120] ), .QN(n698) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[22]  ( .D(n6834), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[118] ), .QN(n696) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[9]  ( .D(n6847), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[105] ), .QN(n683) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[8]  ( .D(n6848), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[104] ), .QN(n682) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[27]  ( .D(n6925), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[219] ), .QN(n797) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[25]  ( .D(n6927), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[217] ), .QN(n795) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[24]  ( .D(n6928), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[216] ), .QN(n794) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[22]  ( .D(n6930), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[214] ), .QN(n792) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[9]  ( .D(n6943), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[201] ), .QN(n779) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[8]  ( .D(n6944), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[200] ), .QN(n778) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[27]  ( .D(n6893), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[187] ), .QN(n765) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[25]  ( .D(n6895), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[185] ), .QN(n763) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[24]  ( .D(n6896), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[184] ), .QN(n762) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[22]  ( .D(n6898), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[182] ), .QN(n760) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[10]  ( .D(n6910), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[170] ), .QN(n748) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[9]  ( .D(n6911), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[169] ), .QN(n747) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[8]  ( .D(n6912), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[168] ), .QN(n746) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[27]  ( .D(n6861), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[155] ), .QN(n733) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[25]  ( .D(n6863), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[153] ), .QN(n731) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[24]  ( .D(n6864), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[152] ), .QN(n730) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[22]  ( .D(n6866), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[150] ), .QN(n728) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[10]  ( .D(n6878), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[138] ), .QN(n716) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[9]  ( .D(n6879), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[137] ), .QN(n715) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[8]  ( .D(n6880), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[136] ), .QN(n714) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[27]  ( .D(n6957), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[251] ), .QN(n829) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[25]  ( .D(n6959), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[249] ), .QN(n827) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[24]  ( .D(n6960), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[248] ), .QN(n826) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[22]  ( .D(n6962), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[246] ), .QN(n824) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[9]  ( .D(n6975), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[233] ), .QN(n811) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[8]  ( .D(n6976), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[232] ), .QN(n810) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[27]  ( .D(n6797), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[91] ), .QN(n669) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[25]  ( .D(n6799), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[89] ), .QN(n667) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[24]  ( .D(n6800), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[88] ), .QN(n666) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[22]  ( .D(n6802), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[86] ), .QN(n664) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[9]  ( .D(n6815), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[73] ), .QN(n651) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[8]  ( .D(n6816), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[72] ), .QN(n650) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[27]  ( .D(n6765), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[59] ), .QN(n637) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[25]  ( .D(n6767), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[57] ), .QN(n635) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[24]  ( .D(n6768), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[56] ), .QN(n634) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[22]  ( .D(n6770), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[54] ), .QN(n632) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[10]  ( .D(n6782), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[42] ), .QN(n620) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[9]  ( .D(n6783), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[41] ), .QN(n619) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[8]  ( .D(n6784), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[40] ), .QN(n618) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[0]  ( .D(n6984), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[224] ), .QN(n802) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[0]  ( .D(n6952), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[192] ), .QN(n770) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[0]  ( .D(n6856), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[96] ), .QN(n674) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[0]  ( .D(n6824), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[64] ), .QN(n642) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[23]  ( .D(n6961), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[247] ), .QN(n825) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[7]  ( .D(n6977), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[231] ), .QN(n809) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[23]  ( .D(n6929), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[215] ), .QN(n793) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[7]  ( .D(n6945), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[199] ), .QN(n777) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[23]  ( .D(n6833), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[119] ), .QN(n697) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[7]  ( .D(n6849), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[103] ), .QN(n681) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[23]  ( .D(n6801), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[87] ), .QN(n665) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[7]  ( .D(n6817), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[71] ), .QN(n649) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[0]  ( .D(n6920), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[160] ), .QN(n738) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[0]  ( .D(n6888), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[128] ), .QN(n706) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[0]  ( .D(n6792), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[32] ), .QN(n610) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[23]  ( .D(n6897), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[183] ), .QN(n761) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[7]  ( .D(n6913), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[167] ), .QN(n745) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[23]  ( .D(n6865), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[151] ), .QN(n729) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[7]  ( .D(n6881), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[135] ), .QN(n713) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[23]  ( .D(n6769), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[55] ), .QN(n633) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[7]  ( .D(n6785), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[39] ), .QN(n617) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[3]  ( .D(n6981), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[227] ), .QN(n805) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[2]  ( .D(n6982), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[226] ), .QN(n804) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[1]  ( .D(n6983), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[225] ), .QN(n803) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[3]  ( .D(n6949), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[195] ), .QN(n773) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[2]  ( .D(n6950), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[194] ), .QN(n772) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[1]  ( .D(n6951), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[193] ), .QN(n771) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[3]  ( .D(n6853), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[99] ), .QN(n677) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[2]  ( .D(n6854), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[98] ), .QN(n676) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[1]  ( .D(n6855), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[97] ), .QN(n675) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[3]  ( .D(n6821), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[67] ), .QN(n645) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[2]  ( .D(n6822), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[66] ), .QN(n644) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[1]  ( .D(n6823), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[65] ), .QN(n643) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[6]  ( .D(n6978), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[230] ), .QN(n808) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[5]  ( .D(n6979), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[229] ), .QN(n807) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[6]  ( .D(n6946), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[198] ), .QN(n776) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[5]  ( .D(n6947), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[197] ), .QN(n775) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[6]  ( .D(n6850), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[102] ), .QN(n680) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[5]  ( .D(n6851), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[101] ), .QN(n679) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[6]  ( .D(n6818), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[70] ), .QN(n648) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[5]  ( .D(n6819), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[69] ), .QN(n647) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[13]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N59 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[13] ), .QN(n8195) );
  DFF_X1 \DataPath/RF/POP_ADDRGEN/curr_addr_reg[8]  ( .D(
        \DataPath/RF/POP_ADDRGEN/N54 ), .CK(CLK), .Q(
        \DataPath/RF/POP_ADDRGEN/curr_addr[8] ), .QN(n8194) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[3]  ( .D(n6917), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[163] ), .QN(n741) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[2]  ( .D(n6918), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[162] ), .QN(n740) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[1]  ( .D(n6919), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[161] ), .QN(n739) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[3]  ( .D(n6885), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[131] ), .QN(n709) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[2]  ( .D(n6886), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[130] ), .QN(n708) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[1]  ( .D(n6887), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[129] ), .QN(n707) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[3]  ( .D(n6789), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[35] ), .QN(n613) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[2]  ( .D(n6790), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[34] ), .QN(n612) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[1]  ( .D(n6791), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[33] ), .QN(n611) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[6]  ( .D(n6914), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[166] ), .QN(n744) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[5]  ( .D(n6915), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[165] ), .QN(n743) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[6]  ( .D(n6882), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[134] ), .QN(n712) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[5]  ( .D(n6883), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[133] ), .QN(n711) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[6]  ( .D(n6786), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[38] ), .QN(n616) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[5]  ( .D(n6787), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[37] ), .QN(n615) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_7/Q_reg[4]  ( .D(n6980), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[228] ), .QN(n806) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_6/Q_reg[4]  ( .D(n6948), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[196] ), .QN(n774) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_3/Q_reg[4]  ( .D(n6852), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[100] ), .QN(n678) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_2/Q_reg[4]  ( .D(n6820), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[68] ), .QN(n646) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_5/Q_reg[4]  ( .D(n6916), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[164] ), .QN(n742) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_4/Q_reg[4]  ( .D(n6884), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[132] ), .QN(n710) );
  DFF_X1 \DataPath/RF/BLOCK_GLOB_1/Q_reg[4]  ( .D(n6788), .CK(CLK), .Q(
        \DataPath/RF/bus_complete_win_data[36] ), .QN(n614) );
  DFF_X1 \DataPath/RF/SWP/Q_reg[0]  ( .D(n7063), .CK(CLK), .Q(
        \DataPath/RF/c_swin[0] ), .QN(n8117) );
  DFF_X1 \DataPath/RF/SWP/Q_reg[1]  ( .D(n7062), .CK(CLK), .Q(
        \DataPath/RF/c_swin[1] ), .QN(n835) );
  DFF_X1 \DataPath/RF/SWP/Q_reg[4]  ( .D(n7059), .CK(CLK), .Q(n8282), .QN(
        n8286) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[15]  ( .D(n2854), .CK(CLK), .Q(n8158), .QN(
        \DataPath/i_PIPLIN_IN1[15] ) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[12]  ( .D(n2857), .CK(CLK), .Q(n8159), .QN(
        \DataPath/i_PIPLIN_IN1[12] ) );
  DFF_X1 \DataPath/REG_IN1/Q_reg[11]  ( .D(n2858), .CK(CLK), .Q(n8160), .QN(
        \DataPath/i_PIPLIN_IN1[11] ) );
  DFF_X1 \DataPath/RF/SWP/Q_reg[3]  ( .D(n7060), .CK(CLK), .Q(
        \DataPath/RF/c_swin[3] ), .QN(n8272) );
  DFF_X1 \DataPath/RF/SWP/Q_reg[2]  ( .D(n7061), .CK(CLK), .Q(
        \DataPath/RF/c_swin[2] ), .QN(n836) );
  DFF_X1 \DataPath/REG_IN2/Q_reg[14]  ( .D(n7016), .CK(CLK), .Q(
        \DataPath/i_PIPLIN_IN2[14] ), .QN(n8204) );
  DFF_X1 \DECODEhw/HALF_ADDER_COUNTER/REG_TICK/Q_reg[2]  ( .D(n11554), .CK(CLK), .QN(\DECODEhw/i_tickcounter[2] ) );
  DFFS_X1 \IR_reg[29]  ( .D(n8255), .CK(CLK), .SN(n8469), .Q(n166), .QN(n8280)
         );
  DFFR_X1 \PC_reg[31]  ( .D(n7025), .CK(CLK), .RN(n8466), .Q(IRAM_ADDRESS[31]), 
        .QN(n7918) );
  DFFR_X1 \IR_reg[26]  ( .D(n7657), .CK(CLK), .RN(n8470), .Q(n172), .QN(n8090)
         );
  DFFS_X1 \IR_reg[31]  ( .D(n10256), .CK(CLK), .SN(n8465), .Q(n8115), .QN(
        IR[31]) );
  DFF_X2 \DataPath/RF/CWP/Q_reg[3]  ( .D(n7066), .CK(CLK), .Q(
        \DataPath/RF/c_win[3] ), .QN(n590) );
  DFF_X2 \CU_I/aluOpcode1_reg[2]  ( .D(n7088), .CK(CLK), .Q(i_ALU_OP[2]), .QN(
        n8084) );
  DFF_X2 \DataPath/RF/CWP/Q_reg[4]  ( .D(n7065), .CK(CLK), .Q(n7648), .QN(
        n8173) );
  DFF_X1 \DataPath/WRF_CUhw/curr_addr_reg[29]  ( .D(n8259), .CK(CLK), .Q(
        \DataPath/WRF_CUhw/curr_addr[29] ) );
  XNOR2_X1 U7545 ( .A(\DP_OP_751_130_6421/n559 ), .B(n7893), .ZN(
        \DP_OP_751_130_6421/n460 ) );
  AND2_X1 U7546 ( .A1(\DP_OP_751_130_6421/n764 ), .A2(
        \DP_OP_751_130_6421/n765 ), .ZN(n7708) );
  NAND2_X1 U7547 ( .A1(\DP_OP_751_130_6421/n1433 ), .A2(
        \DP_OP_751_130_6421/n1390 ), .ZN(n7897) );
  BUF_X1 U7548 ( .A(n8868), .Z(n8326) );
  BUF_X2 U7549 ( .A(n8863), .Z(n8319) );
  NOR2_X1 U7550 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[30] ), .ZN(
        n8075) );
  BUF_X2 U7551 ( .A(n8863), .Z(n8318) );
  BUF_X2 U7552 ( .A(n8868), .Z(n8327) );
  INV_X1 U7553 ( .A(n7737), .ZN(n8813) );
  BUF_X2 U7554 ( .A(n8869), .Z(n8330) );
  AND2_X1 U7555 ( .A1(n8860), .A2(n8859), .ZN(n8116) );
  CLKBUF_X3 U7556 ( .A(n7709), .Z(n8060) );
  INV_X1 U7557 ( .A(n10308), .ZN(n8478) );
  INV_X1 U7558 ( .A(n8274), .ZN(n8275) );
  INV_X2 U7559 ( .A(n9129), .ZN(n7705) );
  INV_X2 U7560 ( .A(n9121), .ZN(n9125) );
  INV_X2 U7561 ( .A(n9151), .ZN(n9157) );
  INV_X1 U7562 ( .A(n10289), .ZN(n11734) );
  BUF_X1 U7563 ( .A(n10258), .Z(n8299) );
  XNOR2_X1 U7564 ( .A(\DP_OP_751_130_6421/n458 ), .B(\DP_OP_751_130_6421/n459 ), .ZN(n7915) );
  XNOR2_X1 U7565 ( .A(\DP_OP_751_130_6421/n460 ), .B(\DP_OP_751_130_6421/n558 ), .ZN(n7921) );
  INV_X1 U7566 ( .A(n7708), .ZN(\DP_OP_751_130_6421/n78 ) );
  XNOR2_X1 U7567 ( .A(\DataPath/ALUhw/MULT/mux_out[1][7] ), .B(n7690), .ZN(
        n7191) );
  INV_X1 U7568 ( .A(n8060), .ZN(n7192) );
  AOI22_X1 U7569 ( .A1(n8060), .A2(\DataPath/ALUhw/MULT/mux_out[0][7] ), .B1(
        \DP_OP_751_130_6421/n1780 ), .B2(n7192), .ZN(n7193) );
  XOR2_X1 U7570 ( .A(n7191), .B(n7193), .Z(\DP_OP_751_130_6421/n1674 ) );
  NOR2_X1 U7571 ( .A1(n7193), .A2(n7191), .ZN(\DP_OP_751_130_6421/n1673 ) );
  AOI22_X1 U7572 ( .A1(n7775), .A2(n11682), .B1(n11680), .B2(n7792), .ZN(n7194) );
  INV_X1 U7573 ( .A(n7194), .ZN(n9411) );
  INV_X1 U7574 ( .A(n9909), .ZN(n7195) );
  OAI21_X1 U7575 ( .B1(n8315), .B2(n9911), .A(n7195), .ZN(n9915) );
  INV_X1 U7576 ( .A(\DP_OP_751_130_6421/n101 ), .ZN(n7196) );
  NOR2_X1 U7577 ( .A1(\DP_OP_751_130_6421/n100 ), .A2(n7196), .ZN(n7197) );
  XNOR2_X1 U7578 ( .A(n7197), .B(\DP_OP_751_130_6421/n102 ), .ZN(n7198) );
  AOI221_X1 U7579 ( .B1(n9777), .B2(n9770), .C1(n9778), .C2(n9770), .A(n9771), 
        .ZN(n7199) );
  XOR2_X1 U7580 ( .A(n9772), .B(n9775), .Z(n7200) );
  NOR2_X1 U7581 ( .A1(n7199), .A2(n7200), .ZN(n7201) );
  AOI211_X1 U7582 ( .C1(n7199), .C2(n7200), .A(n9786), .B(n7201), .ZN(n7202)
         );
  OAI21_X1 U7583 ( .B1(n9777), .B2(n9778), .A(n9770), .ZN(n7203) );
  NAND2_X1 U7584 ( .A1(n7200), .A2(n7203), .ZN(n7204) );
  OAI211_X1 U7585 ( .C1(n7200), .C2(n7203), .A(n9785), .B(n7204), .ZN(n7205)
         );
  NAND3_X1 U7586 ( .A1(n9774), .A2(\DP_OP_751_130_6421/n1107 ), .A3(n9992), 
        .ZN(n7206) );
  NAND3_X1 U7587 ( .A1(n7767), .A2(n9775), .A3(n9990), .ZN(n7207) );
  AOI21_X1 U7588 ( .B1(\DP_OP_751_130_6421/n1107 ), .B2(n9774), .A(n9850), 
        .ZN(n7208) );
  OAI21_X1 U7589 ( .B1(\DP_OP_751_130_6421/n1107 ), .B2(n9774), .A(n7208), 
        .ZN(n7209) );
  NAND4_X1 U7590 ( .A1(n7205), .A2(n7206), .A3(n7207), .A4(n7209), .ZN(n7210)
         );
  AOI211_X1 U7591 ( .C1(n10004), .C2(n7198), .A(n7202), .B(n7210), .ZN(n7211)
         );
  OAI22_X1 U7592 ( .A1(n9790), .A2(n9918), .B1(n9788), .B2(n9939), .ZN(n7212)
         );
  AOI22_X1 U7593 ( .A1(n10019), .A2(n10021), .B1(n10010), .B2(n11721), .ZN(
        n7213) );
  AOI22_X1 U7594 ( .A1(n7759), .A2(n10022), .B1(n10286), .B2(n10024), .ZN(
        n7214) );
  OAI211_X1 U7595 ( .C1(n9941), .C2(n9982), .A(n7213), .B(n7214), .ZN(n7215)
         );
  OAI22_X1 U7596 ( .A1(n9881), .A2(n9878), .B1(n10008), .B2(n10027), .ZN(n7216) );
  NOR3_X1 U7597 ( .A1(n7212), .A2(n7215), .A3(n7216), .ZN(n7217) );
  OAI222_X1 U7598 ( .A1(n11735), .A2(n7211), .B1(n11734), .B2(n516), .C1(n7217), .C2(n11730), .ZN(n7001) );
  INV_X1 U7599 ( .A(n8060), .ZN(n7218) );
  AOI22_X1 U7600 ( .A1(n8060), .A2(\DataPath/ALUhw/MULT/mux_out[0][6] ), .B1(
        \DP_OP_751_130_6421/n1781 ), .B2(n7218), .ZN(n7219) );
  XNOR2_X1 U7601 ( .A(\DataPath/ALUhw/MULT/mux_out[1][6] ), .B(n7690), .ZN(
        n7220) );
  NOR2_X1 U7602 ( .A1(n7219), .A2(n7220), .ZN(\DP_OP_751_130_6421/n1675 ) );
  XOR2_X1 U7603 ( .A(n7219), .B(n7220), .Z(\DP_OP_751_130_6421/n1676 ) );
  AOI22_X1 U7604 ( .A1(n9361), .A2(n11682), .B1(n11680), .B2(n7786), .ZN(n7221) );
  INV_X1 U7605 ( .A(n7221), .ZN(n9341) );
  NAND2_X1 U7606 ( .A1(n8066), .A2(\DP_OP_751_130_6421/n106 ), .ZN(n7222) );
  XNOR2_X1 U7607 ( .A(n7222), .B(\DP_OP_751_130_6421/n107 ), .ZN(n7223) );
  XNOR2_X1 U7608 ( .A(n9778), .B(n9776), .ZN(n7224) );
  INV_X1 U7609 ( .A(n9779), .ZN(n7225) );
  AOI22_X1 U7610 ( .A1(n9779), .A2(n9797), .B1(n9850), .B2(n7225), .ZN(n7226)
         );
  AOI221_X1 U7611 ( .B1(n9795), .B2(n7225), .C1(n9850), .C2(n9779), .A(n9780), 
        .ZN(n7227) );
  AOI21_X1 U7612 ( .B1(n9780), .B2(n7226), .A(n7227), .ZN(n7228) );
  INV_X1 U7613 ( .A(n9778), .ZN(n7229) );
  INV_X1 U7614 ( .A(n9777), .ZN(n7230) );
  OAI221_X1 U7615 ( .B1(n9778), .B2(n9777), .C1(n7229), .C2(n7230), .A(n9785), 
        .ZN(n7231) );
  OAI211_X1 U7616 ( .C1(n9786), .C2(n7224), .A(n7228), .B(n7231), .ZN(n7232)
         );
  AOI21_X1 U7617 ( .B1(n7223), .B2(n8337), .A(n7232), .ZN(n7233) );
  OAI22_X1 U7618 ( .A1(n9790), .A2(n9942), .B1(n10008), .B2(n10017), .ZN(n7234) );
  AOI22_X1 U7619 ( .A1(n10022), .A2(n10023), .B1(n10284), .B2(n9974), .ZN(
        n7235) );
  AOI22_X1 U7620 ( .A1(n9977), .A2(n10020), .B1(n7759), .B2(n11721), .ZN(n7236) );
  OAI211_X1 U7621 ( .C1(n9983), .C2(n9939), .A(n7235), .B(n7236), .ZN(n7237)
         );
  OAI22_X1 U7622 ( .A1(n9881), .A2(n10027), .B1(n9789), .B2(n9880), .ZN(n7238)
         );
  NOR3_X1 U7623 ( .A1(n7234), .A2(n7237), .A3(n7238), .ZN(n7239) );
  OAI222_X1 U7624 ( .A1(n11735), .A2(n7233), .B1(n11734), .B2(n515), .C1(n7239), .C2(n11730), .ZN(n7002) );
  AND2_X1 U7625 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[19] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N23 ) );
  AND2_X1 U7626 ( .A1(n8462), .A2(\DataPath/RF/internal_out1[29] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N33 ) );
  XNOR2_X1 U7627 ( .A(\DataPath/ALUhw/MULT/mux_out[1][15] ), .B(n7690), .ZN(
        n7240) );
  XOR2_X1 U7628 ( .A(\DataPath/ALUhw/MULT/mux_out[0][15] ), .B(n7974), .Z(
        n7241) );
  XOR2_X1 U7629 ( .A(n7240), .B(n7241), .Z(\DP_OP_751_130_6421/n1658 ) );
  NOR2_X1 U7630 ( .A1(n7241), .A2(n7240), .ZN(\DP_OP_751_130_6421/n1657 ) );
  AOI22_X1 U7631 ( .A1(\DataPath/i_PIPLIN_A[7] ), .A2(n8442), .B1(
        \DataPath/i_PIPLIN_IN1[7] ), .B2(n8443), .ZN(n7242) );
  INV_X1 U7632 ( .A(n7242), .ZN(n9151) );
  OAI22_X1 U7633 ( .A1(n7741), .A2(n9910), .B1(n8314), .B2(n8260), .ZN(n7243)
         );
  XNOR2_X1 U7634 ( .A(n8060), .B(n7243), .ZN(\DP_OP_751_130_6421/n159 ) );
  INV_X1 U7635 ( .A(n9137), .ZN(n7244) );
  INV_X1 U7636 ( .A(n8325), .ZN(n7245) );
  NAND3_X1 U7637 ( .A1(n9686), .A2(n11716), .A3(n10283), .ZN(n7246) );
  OAI21_X1 U7638 ( .B1(n9545), .B2(n7245), .A(n7246), .ZN(n7247) );
  AOI22_X1 U7639 ( .A1(n9687), .A2(n9196), .B1(n9691), .B2(n9078), .ZN(n7248)
         );
  OAI21_X1 U7640 ( .B1(n9633), .B2(n9543), .A(n7248), .ZN(n7249) );
  AOI211_X1 U7641 ( .C1(n9195), .C2(n7244), .A(n7247), .B(n7249), .ZN(n9940)
         );
  NAND2_X1 U7642 ( .A1(n8067), .A2(\DP_OP_751_130_6421/n114 ), .ZN(n7250) );
  XNOR2_X1 U7643 ( .A(n7250), .B(\DP_OP_751_130_6421/n115 ), .ZN(n7251) );
  OR2_X1 U7644 ( .A1(n9963), .A2(n9781), .ZN(n7252) );
  INV_X1 U7645 ( .A(n9782), .ZN(n7253) );
  AOI22_X1 U7646 ( .A1(n9782), .A2(n9803), .B1(n9990), .B2(n7253), .ZN(n7254)
         );
  INV_X1 U7647 ( .A(n9783), .ZN(n7255) );
  OAI221_X1 U7648 ( .B1(n9783), .B2(n9992), .C1(n7255), .C2(n9803), .A(n9784), 
        .ZN(n7256) );
  OAI21_X1 U7649 ( .B1(n7254), .B2(n9784), .A(n7256), .ZN(n7257) );
  AOI21_X1 U7650 ( .B1(n9785), .B2(n7252), .A(n7257), .ZN(n7258) );
  OAI21_X1 U7651 ( .B1(n9786), .B2(n7252), .A(n7258), .ZN(n7259) );
  AOI21_X1 U7652 ( .B1(n7251), .B2(n8337), .A(n7259), .ZN(n7260) );
  OAI22_X1 U7653 ( .A1(n9790), .A2(n9860), .B1(n9788), .B2(n9942), .ZN(n7261)
         );
  AOI22_X1 U7654 ( .A1(n9977), .A2(n10010), .B1(n9978), .B2(n11721), .ZN(n7262) );
  AOI22_X1 U7655 ( .A1(n10286), .A2(n10022), .B1(n10284), .B2(n9979), .ZN(
        n7263) );
  OAI211_X1 U7656 ( .C1(n9983), .C2(n9918), .A(n7262), .B(n7263), .ZN(n7264)
         );
  OAI22_X1 U7657 ( .A1(n9943), .A2(n9939), .B1(n9789), .B2(n9878), .ZN(n7265)
         );
  NOR3_X1 U7658 ( .A1(n7261), .A2(n7264), .A3(n7265), .ZN(n7266) );
  OAI222_X1 U7659 ( .A1(n11735), .A2(n7260), .B1(n11734), .B2(n514), .C1(n7266), .C2(n11730), .ZN(n7004) );
  AND2_X1 U7660 ( .A1(n8459), .A2(\DataPath/RF/internal_out2[29] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N33 ) );
  AND2_X1 U7661 ( .A1(n8470), .A2(\DataPath/RF/internal_out1[19] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N23 ) );
  AOI22_X1 U7662 ( .A1(n8084), .A2(n9889), .B1(i_ALU_OP[2]), .B2(n9966), .ZN(
        n7267) );
  INV_X1 U7663 ( .A(n7267), .ZN(n9285) );
  XOR2_X1 U7664 ( .A(\DataPath/ALUhw/MULT/mux_out[0][4] ), .B(n8060), .Z(n7268) );
  OAI22_X1 U7665 ( .A1(n8322), .A2(n8308), .B1(n8318), .B2(n8313), .ZN(n7269)
         );
  XNOR2_X1 U7666 ( .A(n7690), .B(n7269), .ZN(n7270) );
  NOR2_X1 U7667 ( .A1(n7268), .A2(n7270), .ZN(\DP_OP_751_130_6421/n1679 ) );
  XOR2_X1 U7668 ( .A(n7268), .B(n7270), .Z(\DP_OP_751_130_6421/n1680 ) );
  AOI21_X1 U7669 ( .B1(n7974), .B2(n8452), .A(n9064), .ZN(n7271) );
  INV_X1 U7670 ( .A(n7271), .ZN(n9065) );
  INV_X1 U7671 ( .A(n9497), .ZN(n7272) );
  OAI21_X1 U7672 ( .B1(n8302), .B2(n9007), .A(n7272), .ZN(n9075) );
  OAI21_X1 U7673 ( .B1(n181), .B2(n10153), .A(n10155), .ZN(n11672) );
  INV_X1 U7674 ( .A(n11732), .ZN(n7273) );
  INV_X1 U7675 ( .A(n9595), .ZN(n7274) );
  INV_X1 U7676 ( .A(n9341), .ZN(n7275) );
  NAND2_X1 U7677 ( .A1(n9143), .A2(n7275), .ZN(n7276) );
  AOI222_X1 U7678 ( .A1(n7273), .A2(n9681), .B1(n7274), .B2(n9045), .C1(n7276), 
        .C2(n9683), .ZN(n7277) );
  INV_X1 U7679 ( .A(n7786), .ZN(n7278) );
  OAI222_X1 U7680 ( .A1(n7278), .A2(n9018), .B1(n9157), .B2(n9281), .C1(n9138), 
        .C2(n9547), .ZN(n7279) );
  AOI21_X1 U7681 ( .B1(n9588), .B2(n9043), .A(n7279), .ZN(n7280) );
  OAI211_X1 U7682 ( .C1(n9592), .C2(n9139), .A(n7277), .B(n7280), .ZN(n9920)
         );
  INV_X1 U7683 ( .A(\DP_OP_751_130_6421/n117 ), .ZN(n7281) );
  NOR2_X1 U7684 ( .A1(\DP_OP_751_130_6421/n116 ), .A2(n7281), .ZN(n7282) );
  XNOR2_X1 U7685 ( .A(n7282), .B(\DP_OP_751_130_6421/n118 ), .ZN(n7283) );
  NOR3_X1 U7686 ( .A1(n7771), .A2(n9797), .A3(n9796), .ZN(n7284) );
  OAI22_X1 U7687 ( .A1(n9787), .A2(n9939), .B1(n9788), .B2(n9880), .ZN(n7285)
         );
  OAI22_X1 U7688 ( .A1(n9789), .A2(n10027), .B1(n9790), .B2(n9878), .ZN(n7286)
         );
  AOI22_X1 U7689 ( .A1(n11719), .A2(n10284), .B1(n11721), .B2(n10286), .ZN(
        n7287) );
  OAI21_X1 U7690 ( .B1(n9791), .B2(n9918), .A(n7287), .ZN(n7288) );
  OAI22_X1 U7691 ( .A1(n9941), .A2(n9860), .B1(n9983), .B2(n9942), .ZN(n7289)
         );
  NOR4_X1 U7692 ( .A1(n7285), .A2(n7286), .A3(n7288), .A4(n7289), .ZN(n7290)
         );
  NOR2_X1 U7693 ( .A1(n7799), .A2(\DP_OP_751_130_6421/n1311 ), .ZN(n7291) );
  AOI22_X1 U7694 ( .A1(n7799), .A2(\DP_OP_751_130_6421/n1311 ), .B1(n7291), 
        .B2(n9795), .ZN(n7292) );
  OAI21_X1 U7695 ( .B1(n7291), .B2(n9803), .A(n7292), .ZN(n7293) );
  XOR2_X1 U7696 ( .A(n7799), .B(n9792), .Z(n7294) );
  NAND2_X1 U7697 ( .A1(n9793), .A2(n7294), .ZN(n7295) );
  OAI211_X1 U7698 ( .C1(n9793), .C2(n7294), .A(n9958), .B(n7295), .ZN(n7296)
         );
  OAI211_X1 U7699 ( .C1(n7290), .C2(n9815), .A(n7293), .B(n7296), .ZN(n7297)
         );
  AOI211_X1 U7700 ( .C1(n8337), .C2(n7283), .A(n7284), .B(n7297), .ZN(n7298)
         );
  OAI22_X1 U7701 ( .A1(n513), .A2(n11734), .B1(n11735), .B2(n7298), .ZN(n7005)
         );
  AND2_X1 U7702 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[17] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N21 ) );
  AND2_X1 U7703 ( .A1(n8459), .A2(\DataPath/RF/internal_out1[18] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N22 ) );
  OAI21_X1 U7704 ( .B1(n182), .B2(n10153), .A(n10155), .ZN(n8822) );
  INV_X1 U7705 ( .A(n8325), .ZN(n7299) );
  NOR2_X1 U7706 ( .A1(n9495), .A2(n7299), .ZN(n7300) );
  OAI22_X1 U7707 ( .A1(n9538), .A2(n9201), .B1(n9498), .B2(n9633), .ZN(n7301)
         );
  AOI211_X1 U7708 ( .C1(n9691), .C2(n9075), .A(n7300), .B(n7301), .ZN(n7302)
         );
  OAI21_X1 U7709 ( .B1(n8085), .B2(n9199), .A(n9667), .ZN(n7303) );
  OAI211_X1 U7710 ( .C1(n9516), .C2(n11733), .A(n9686), .B(n7303), .ZN(n7304)
         );
  NAND2_X1 U7711 ( .A1(n7302), .A2(n7304), .ZN(n9211) );
  XOR2_X1 U7712 ( .A(\DP_OP_751_130_6421/n159 ), .B(\DP_OP_751_130_6421/n161 ), 
        .Z(n7305) );
  NAND3_X1 U7713 ( .A1(n7974), .A2(n8312), .A3(n9990), .ZN(n7306) );
  NAND3_X1 U7714 ( .A1(n7747), .A2(n9913), .A3(n9992), .ZN(n7307) );
  NOR3_X1 U7715 ( .A1(n9911), .A2(n8315), .A3(n11696), .ZN(n7308) );
  OAI221_X1 U7716 ( .B1(n7308), .B2(n10288), .C1(n7308), .C2(n9912), .A(n9909), 
        .ZN(n7309) );
  NAND3_X1 U7717 ( .A1(n7306), .A2(n7307), .A3(n7309), .ZN(n7310) );
  INV_X1 U7718 ( .A(n9914), .ZN(n7311) );
  OAI22_X1 U7719 ( .A1(n9916), .A2(n7311), .B1(n11696), .B2(n9915), .ZN(n7312)
         );
  AOI211_X1 U7720 ( .C1(n7305), .C2(n10004), .A(n7310), .B(n7312), .ZN(n7313)
         );
  OAI22_X1 U7721 ( .A1(n9917), .A2(n10027), .B1(n9919), .B2(n9918), .ZN(n7314)
         );
  AOI21_X1 U7722 ( .B1(n11698), .B2(n10021), .A(n7314), .ZN(n7315) );
  AOI22_X1 U7723 ( .A1(n9920), .A2(n10023), .B1(n10284), .B2(n9921), .ZN(n7316) );
  AOI22_X1 U7724 ( .A1(n9922), .A2(n10286), .B1(n7759), .B2(n9923), .ZN(n7317)
         );
  AOI22_X1 U7725 ( .A1(n9924), .A2(n10010), .B1(n10013), .B2(n9925), .ZN(n7318) );
  NAND4_X1 U7726 ( .A1(n7315), .A2(n7316), .A3(n7317), .A4(n7318), .ZN(n7319)
         );
  XNOR2_X1 U7727 ( .A(n7974), .B(n8312), .ZN(n7320) );
  OAI22_X1 U7728 ( .A1(n9953), .A2(n7320), .B1(n508), .B2(n11734), .ZN(n7321)
         );
  AOI21_X1 U7729 ( .B1(n10280), .B2(n7319), .A(n7321), .ZN(n7322) );
  OAI21_X1 U7730 ( .B1(n10032), .B2(n7313), .A(n7322), .ZN(n7012) );
  AND2_X1 U7731 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[18] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N22 ) );
  AND2_X1 U7732 ( .A1(n8466), .A2(\DataPath/RF/internal_out1[17] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N21 ) );
  OAI22_X1 U7733 ( .A1(n8321), .A2(n9783), .B1(n8318), .B2(n9796), .ZN(n7323)
         );
  XNOR2_X1 U7734 ( .A(n8059), .B(n7323), .ZN(n7324) );
  OAI22_X1 U7735 ( .A1(n8261), .A2(n8303), .B1(n7740), .B2(n9972), .ZN(n7325)
         );
  XOR2_X1 U7736 ( .A(n7974), .B(n7325), .Z(n7326) );
  NOR2_X1 U7737 ( .A1(n7324), .A2(n7326), .ZN(\DP_OP_751_130_6421/n1659 ) );
  XOR2_X1 U7738 ( .A(n7324), .B(n7326), .Z(\DP_OP_751_130_6421/n1660 ) );
  OAI21_X1 U7739 ( .B1(\DP_OP_751_130_6421/n1255 ), .B2(
        \DP_OP_751_130_6421/n1199 ), .A(\DP_OP_751_130_6421/n1254 ), .ZN(n7931) );
  INV_X1 U7740 ( .A(n9286), .ZN(n7327) );
  AOI21_X1 U7741 ( .B1(n9285), .B2(n11722), .A(n7327), .ZN(n9412) );
  AND4_X1 U7742 ( .A1(n8090), .A2(n7720), .A3(n7992), .A4(n8246), .ZN(n8242)
         );
  OAI21_X1 U7743 ( .B1(n9928), .B2(n9926), .A(n9927), .ZN(n7328) );
  INV_X1 U7744 ( .A(n9951), .ZN(n7329) );
  AOI222_X1 U7745 ( .A1(n9929), .A2(n7328), .B1(n9929), .B2(n9932), .C1(n7328), 
        .C2(n7329), .ZN(n9234) );
  INV_X1 U7746 ( .A(n9088), .ZN(n7330) );
  AOI21_X1 U7747 ( .B1(n7970), .B2(n8084), .A(n7330), .ZN(n9911) );
  INV_X1 U7748 ( .A(n9590), .ZN(n7331) );
  INV_X1 U7749 ( .A(n9589), .ZN(n7332) );
  AOI222_X1 U7750 ( .A1(n7331), .A2(n7332), .B1(n9591), .B2(n9683), .C1(n9588), 
        .C2(n8325), .ZN(n7333) );
  OAI21_X1 U7751 ( .B1(n9592), .B2(n9593), .A(n9220), .ZN(n7334) );
  AOI22_X1 U7752 ( .A1(n9687), .A2(n9597), .B1(n9594), .B2(n7334), .ZN(n7335)
         );
  OAI211_X1 U7753 ( .C1(n9595), .C2(n9596), .A(n7333), .B(n7335), .ZN(n10024)
         );
  XOR2_X1 U7754 ( .A(n10186), .B(IRAM_ADDRESS[20]), .Z(n7336) );
  XNOR2_X1 U7755 ( .A(n10152), .B(n7336), .ZN(n7337) );
  AOI22_X1 U7756 ( .A1(n10266), .A2(IRAM_ADDRESS[20]), .B1(i_RD1[20]), .B2(
        n10267), .ZN(n7338) );
  OAI21_X1 U7757 ( .B1(n11678), .B2(n7337), .A(n7338), .ZN(n7036) );
  AOI22_X1 U7758 ( .A1(n10286), .A2(n9979), .B1(n9978), .B2(n11719), .ZN(n7339) );
  AOI22_X1 U7759 ( .A1(n10020), .A2(n9920), .B1(n10013), .B2(n9924), .ZN(n7340) );
  OAI211_X1 U7760 ( .C1(n9940), .C2(n9880), .A(n7339), .B(n7340), .ZN(n7341)
         );
  AOI22_X1 U7761 ( .A1(n9176), .A2(n10021), .B1(n7759), .B2(n9211), .ZN(n7342)
         );
  OAI21_X1 U7762 ( .B1(n9982), .B2(n9798), .A(n7342), .ZN(n7343) );
  NOR2_X1 U7763 ( .A1(n9878), .A2(n9787), .ZN(n7344) );
  NOR3_X1 U7764 ( .A1(n7344), .A2(n7341), .A3(n7343), .ZN(n7345) );
  NAND2_X1 U7765 ( .A1(DRAM_ADDRESS[5]), .A2(n7764), .ZN(n7346) );
  NAND2_X1 U7766 ( .A1(n8057), .A2(n7792), .ZN(n7347) );
  NAND2_X1 U7767 ( .A1(n9850), .A2(n7347), .ZN(n7348) );
  OAI221_X1 U7768 ( .B1(n7347), .B2(n9992), .C1(n8057), .C2(n7792), .A(n7348), 
        .ZN(n7349) );
  AOI21_X1 U7769 ( .B1(n9100), .B2(n9809), .A(n9135), .ZN(n7350) );
  OAI21_X1 U7770 ( .B1(n9100), .B2(n9809), .A(n7350), .ZN(n7351) );
  OAI211_X1 U7771 ( .C1(n9100), .C2(n9811), .A(n10278), .B(n9123), .ZN(n7352)
         );
  NAND3_X1 U7772 ( .A1(n8445), .A2(n9125), .A3(n9990), .ZN(n7353) );
  NAND4_X1 U7773 ( .A1(n7349), .A2(n7351), .A3(n7352), .A4(n7353), .ZN(n7354)
         );
  NAND2_X1 U7774 ( .A1(n8073), .A2(\DP_OP_751_130_6421/n144 ), .ZN(n7355) );
  XNOR2_X1 U7775 ( .A(n7355), .B(\DP_OP_751_130_6421/n145 ), .ZN(n7356) );
  OAI221_X1 U7776 ( .B1(n7354), .B2(n7356), .C1(n7354), .C2(n8337), .A(n10279), 
        .ZN(n7357) );
  OAI211_X1 U7777 ( .C1(n7345), .C2(n11730), .A(n7346), .B(n7357), .ZN(n7010)
         );
  AND2_X1 U7778 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[15] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N19 ) );
  AND2_X1 U7779 ( .A1(n8464), .A2(\DataPath/RF/internal_out1[16] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N20 ) );
  OAI22_X1 U7780 ( .A1(\DataPath/RF/c_win[1] ), .A2(n8272), .B1(n589), .B2(
        n8282), .ZN(n7358) );
  NOR3_X1 U7781 ( .A1(n8236), .A2(n8250), .A3(n7358), .ZN(n8235) );
  OAI22_X1 U7782 ( .A1(n8321), .A2(n8305), .B1(n8317), .B2(n8308), .ZN(n7359)
         );
  XNOR2_X1 U7783 ( .A(n8059), .B(n7359), .ZN(n7360) );
  XOR2_X1 U7784 ( .A(\DataPath/ALUhw/MULT/mux_out[0][5] ), .B(n8060), .Z(n7361) );
  XOR2_X1 U7785 ( .A(n7360), .B(n7361), .Z(\DP_OP_751_130_6421/n1678 ) );
  NOR2_X1 U7786 ( .A1(n7360), .A2(n7361), .ZN(\DP_OP_751_130_6421/n1677 ) );
  AOI22_X1 U7787 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[19] ), .B1(
        n7945), .B2(n7935), .ZN(n7362) );
  INV_X1 U7788 ( .A(n7362), .ZN(n7848) );
  OAI21_X1 U7789 ( .B1(n180), .B2(n10153), .A(n10155), .ZN(n8826) );
  NAND3_X1 U7790 ( .A1(IR[1]), .A2(n8802), .A3(n8803), .ZN(\intadd_1/B[0] ) );
  OAI21_X1 U7791 ( .B1(n10299), .B2(n9324), .A(n9329), .ZN(n9427) );
  INV_X1 U7792 ( .A(\DP_OP_751_130_6421/n1208 ), .ZN(n7363) );
  INV_X1 U7793 ( .A(\DP_OP_751_130_6421/n1209 ), .ZN(n7364) );
  OAI21_X1 U7794 ( .B1(\DP_OP_751_130_6421/n1209 ), .B2(
        \DP_OP_751_130_6421/n1208 ), .A(\DP_OP_751_130_6421/n1273 ), .ZN(n7365) );
  OAI21_X1 U7795 ( .B1(n7363), .B2(n7364), .A(n7365), .ZN(
        \DP_OP_751_130_6421/n1173 ) );
  NAND3_X1 U7796 ( .A1(\DP_OP_751_130_6421/n393 ), .A2(n9992), .A3(n7775), 
        .ZN(n7366) );
  NAND3_X1 U7797 ( .A1(n9826), .A2(n9824), .A3(n9990), .ZN(n7367) );
  INV_X1 U7798 ( .A(n9825), .ZN(n7368) );
  OAI221_X1 U7799 ( .B1(n9821), .B2(n9822), .C1(n9821), .C2(n9823), .A(n7368), 
        .ZN(n7369) );
  AOI21_X1 U7800 ( .B1(n9823), .B2(n9819), .A(n9820), .ZN(n7370) );
  OAI21_X1 U7801 ( .B1(n9823), .B2(n9819), .A(n7370), .ZN(n7371) );
  NAND4_X1 U7802 ( .A1(n7366), .A2(n7367), .A3(n7369), .A4(n7371), .ZN(n7859)
         );
  NAND2_X1 U7803 ( .A1(n11716), .A2(n10285), .ZN(n7372) );
  INV_X1 U7804 ( .A(n9686), .ZN(n7373) );
  INV_X1 U7805 ( .A(n8325), .ZN(n7374) );
  OAI222_X1 U7806 ( .A1(n7372), .A2(n7373), .B1(n9139), .B2(n9221), .C1(n7374), 
        .C2(n9475), .ZN(n7375) );
  NOR2_X1 U7807 ( .A1(n9137), .A2(n9081), .ZN(n7376) );
  AOI21_X1 U7808 ( .B1(n9224), .B2(n9687), .A(n7376), .ZN(n7377) );
  OAI21_X1 U7809 ( .B1(n9477), .B2(n9633), .A(n7377), .ZN(n7378) );
  AOI211_X1 U7810 ( .C1(n9691), .C2(n9084), .A(n7375), .B(n7378), .ZN(n9787)
         );
  AOI22_X2 U7811 ( .A1(n7692), .A2(\DataPath/i_PIPLIN_A[9] ), .B1(n8443), .B2(
        \DataPath/i_PIPLIN_IN1[9] ), .ZN(n9951) );
  INV_X1 U7812 ( .A(n8306), .ZN(n7379) );
  NOR2_X1 U7813 ( .A1(n9080), .A2(n7379), .ZN(n9095) );
  INV_X1 U7814 ( .A(IR[31]), .ZN(n7380) );
  NOR3_X1 U7815 ( .A1(n8492), .A2(n7969), .A3(n7380), .ZN(n10136) );
  INV_X1 U7816 ( .A(n11617), .ZN(n7381) );
  NOR4_X1 U7817 ( .A1(IR[4]), .A2(n8097), .A3(IR[5]), .A4(n7381), .ZN(n10240)
         );
  OR2_X1 U7818 ( .A1(n8827), .A2(n7928), .ZN(n7382) );
  INV_X1 U7819 ( .A(n8824), .ZN(n7383) );
  OAI221_X1 U7820 ( .B1(n8824), .B2(n7382), .C1(n7383), .C2(n8823), .A(n10149), 
        .ZN(n7384) );
  AOI22_X1 U7821 ( .A1(n10266), .A2(IRAM_ADDRESS[17]), .B1(i_RD1[17]), .B2(
        n10267), .ZN(n7385) );
  OAI21_X1 U7822 ( .B1(n11678), .B2(n7384), .A(n7385), .ZN(n7039) );
  INV_X1 U7823 ( .A(n9914), .ZN(n7386) );
  NAND2_X1 U7824 ( .A1(n9090), .A2(n7386), .ZN(n7387) );
  XNOR2_X1 U7825 ( .A(n11695), .B(n7387), .ZN(n7388) );
  INV_X1 U7826 ( .A(\DP_OP_751_130_6421/n155 ), .ZN(n7389) );
  NOR2_X1 U7827 ( .A1(\DP_OP_751_130_6421/n154 ), .A2(n7389), .ZN(n7390) );
  XNOR2_X1 U7828 ( .A(n9069), .B(n8309), .ZN(n7391) );
  NAND3_X1 U7829 ( .A1(n9069), .A2(n8309), .A3(n9990), .ZN(n7392) );
  NAND3_X1 U7830 ( .A1(n7860), .A2(n9992), .A3(n9070), .ZN(n7393) );
  OAI211_X1 U7831 ( .C1(n9850), .C2(n7391), .A(n7392), .B(n7393), .ZN(n7394)
         );
  XNOR2_X1 U7832 ( .A(n7390), .B(\DP_OP_751_130_6421/n158 ), .ZN(n7395) );
  AOI21_X1 U7833 ( .B1(n7395), .B2(n8337), .A(n7394), .ZN(n7396) );
  OAI221_X1 U7834 ( .B1(n11697), .B2(n10282), .C1(n11697), .C2(n11695), .A(
        n9072), .ZN(n7397) );
  OAI211_X1 U7835 ( .C1(n9916), .C2(n7388), .A(n7396), .B(n7397), .ZN(n7398)
         );
  OAI22_X1 U7836 ( .A1(n9917), .A2(n9878), .B1(n9938), .B2(n10017), .ZN(n7399)
         );
  AOI21_X1 U7837 ( .B1(n10013), .B2(n9921), .A(n7399), .ZN(n7400) );
  AOI22_X1 U7838 ( .A1(n9922), .A2(n9978), .B1(n10284), .B2(n9079), .ZN(n7401)
         );
  AOI22_X1 U7839 ( .A1(n9920), .A2(n7759), .B1(n10010), .B2(n9923), .ZN(n7402)
         );
  AOI22_X1 U7840 ( .A1(n10021), .A2(n9924), .B1(n10020), .B2(n11698), .ZN(
        n7403) );
  NAND4_X1 U7841 ( .A1(n7400), .A2(n7401), .A3(n7402), .A4(n7403), .ZN(n7404)
         );
  AOI222_X1 U7842 ( .A1(n7398), .A2(n10281), .B1(DRAM_ADDRESS[2]), .B2(n7764), 
        .C1(n7404), .C2(n10280), .ZN(n2165) );
  AND2_X1 U7843 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[16] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N20 ) );
  AND2_X1 U7844 ( .A1(n8466), .A2(\DataPath/RF/internal_out1[15] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N19 ) );
  OAI22_X1 U7845 ( .A1(n8858), .A2(n9277), .B1(n8974), .B2(n9460), .ZN(n7405)
         );
  XNOR2_X1 U7846 ( .A(n7880), .B(n7405), .ZN(\DP_OP_751_130_6421/n1725 ) );
  AOI22_X1 U7847 ( .A1(\DataPath/RF/c_swin[2] ), .A2(n589), .B1(n836), .B2(
        \DataPath/RF/c_win[2] ), .ZN(n7406) );
  OAI21_X1 U7848 ( .B1(n8282), .B2(n8173), .A(n7406), .ZN(n7989) );
  INV_X1 U7849 ( .A(n10327), .ZN(n7407) );
  INV_X1 U7850 ( .A(n10318), .ZN(n7408) );
  INV_X1 U7851 ( .A(n10319), .ZN(n7409) );
  INV_X1 U7852 ( .A(n10320), .ZN(n7410) );
  OAI221_X1 U7853 ( .B1(n7410), .B2(n10322), .C1(n7410), .C2(n10820), .A(
        n10321), .ZN(n7411) );
  OAI221_X1 U7854 ( .B1(n7409), .B2(n10324), .C1(n7409), .C2(n7411), .A(n10323), .ZN(n7412) );
  OAI221_X1 U7855 ( .B1(n7408), .B2(n10326), .C1(n7408), .C2(n7412), .A(n10325), .ZN(n7413) );
  OAI221_X1 U7856 ( .B1(n7407), .B2(n10328), .C1(n7407), .C2(n7413), .A(n10329), .ZN(n7414) );
  NAND2_X1 U7857 ( .A1(n10330), .A2(n7414), .ZN(n10349) );
  OR2_X1 U7858 ( .A1(\DP_OP_751_130_6421/n458 ), .A2(\DP_OP_751_130_6421/n459 ), .ZN(n7914) );
  AOI22_X1 U7859 ( .A1(n8042), .A2(n7848), .B1(n7649), .B2(n7847), .ZN(n7415)
         );
  INV_X1 U7860 ( .A(n8078), .ZN(n7416) );
  OAI21_X1 U7861 ( .B1(n8077), .B2(n7416), .A(n8047), .ZN(n7417) );
  OAI211_X1 U7862 ( .C1(n8046), .C2(n8079), .A(n7415), .B(n7417), .ZN(n7808)
         );
  NAND3_X1 U7863 ( .A1(IR[5]), .A2(n8802), .A3(n8803), .ZN(\intadd_1/B[4] ) );
  NOR3_X1 U7864 ( .A1(n7726), .A2(n11735), .A3(n7748), .ZN(n7418) );
  NAND3_X1 U7865 ( .A1(\DP_OP_751_130_6421/n61 ), .A2(n7823), .A3(n7418), .ZN(
        n7822) );
  NOR2_X1 U7866 ( .A1(n8330), .A2(n9910), .ZN(n7419) );
  XOR2_X1 U7867 ( .A(\DP_OP_751_130_6421/n1681 ), .B(n7419), .Z(
        \DP_OP_751_130_6421/n1582 ) );
  NOR2_X1 U7868 ( .A1(n8330), .A2(n9910), .ZN(n7420) );
  MUX2_X1 U7869 ( .A(n8057), .B(\DP_OP_751_130_6421/n1681 ), .S(n7420), .Z(
        \DP_OP_751_130_6421/n1581 ) );
  INV_X1 U7870 ( .A(n7705), .ZN(n7421) );
  NOR2_X1 U7871 ( .A1(n9124), .A2(n7421), .ZN(n9155) );
  INV_X1 U7872 ( .A(n9086), .ZN(n7422) );
  AOI21_X1 U7873 ( .B1(i_ALU_OP[2]), .B2(n9806), .A(n7422), .ZN(n9692) );
  INV_X1 U7874 ( .A(n9105), .ZN(n7423) );
  AOI21_X1 U7875 ( .B1(n9125), .B2(i_ALU_OP[2]), .A(n7423), .ZN(n9408) );
  NAND2_X1 U7876 ( .A1(n8818), .A2(n10188), .ZN(n7424) );
  NAND3_X1 U7877 ( .A1(n7424), .A2(\intadd_0/n16 ), .A3(n8093), .ZN(n8254) );
  NOR2_X1 U7878 ( .A1(n7940), .A2(n8148), .ZN(n7425) );
  AOI21_X1 U7879 ( .B1(n7940), .B2(\DataPath/i_PIPLIN_IN2[15] ), .A(n7425), 
        .ZN(n7767) );
  NAND3_X1 U7880 ( .A1(n11716), .A2(n9691), .A3(n10283), .ZN(n7426) );
  NAND2_X1 U7881 ( .A1(n8325), .A2(n9194), .ZN(n7427) );
  OAI211_X1 U7882 ( .C1(n9220), .C2(n9545), .A(n7426), .B(n7427), .ZN(n7428)
         );
  AOI21_X1 U7883 ( .B1(n9195), .B2(n9226), .A(n7428), .ZN(n7429) );
  NAND2_X1 U7884 ( .A1(n9686), .A2(n9196), .ZN(n7430) );
  OAI211_X1 U7885 ( .C1(n9538), .C2(n9540), .A(n7429), .B(n7430), .ZN(n10014)
         );
  NAND2_X1 U7886 ( .A1(n10232), .A2(n10066), .ZN(n7431) );
  NOR2_X1 U7887 ( .A1(n172), .A2(n165), .ZN(n7432) );
  NOR3_X1 U7888 ( .A1(n7432), .A2(n10140), .A3(n8287), .ZN(n7433) );
  AOI211_X1 U7889 ( .C1(n8287), .C2(n7431), .A(n7433), .B(n10136), .ZN(n10297)
         );
  INV_X1 U7890 ( .A(i_RD1[8]), .ZN(n7434) );
  XOR2_X1 U7891 ( .A(n10194), .B(n8169), .Z(n7435) );
  NAND2_X1 U7892 ( .A1(n7894), .A2(n10195), .ZN(n7436) );
  OAI22_X1 U7893 ( .A1(n7436), .A2(n10196), .B1(n7894), .B2(n7435), .ZN(n7437)
         );
  OAI222_X1 U7894 ( .A1(n7434), .A2(n7750), .B1(n7437), .B2(n11678), .C1(
        n10210), .C2(n8169), .ZN(n7048) );
  NAND2_X1 U7895 ( .A1(\DP_OP_751_130_6421/n151 ), .A2(
        \DP_OP_751_130_6421/n152 ), .ZN(n7438) );
  XNOR2_X1 U7896 ( .A(n7438), .B(\DP_OP_751_130_6421/n153 ), .ZN(n7439) );
  INV_X1 U7897 ( .A(n9095), .ZN(n7440) );
  NAND2_X1 U7898 ( .A1(n9094), .A2(n7440), .ZN(n7441) );
  AOI21_X1 U7899 ( .B1(n11697), .B2(n7441), .A(n11696), .ZN(n7442) );
  NOR2_X1 U7900 ( .A1(n7442), .A2(n10288), .ZN(n7443) );
  INV_X1 U7901 ( .A(n9093), .ZN(n7444) );
  NOR2_X1 U7902 ( .A1(n11695), .A2(n9914), .ZN(n7445) );
  AOI21_X1 U7903 ( .B1(n7445), .B2(n9090), .A(n7444), .ZN(n7446) );
  NAND2_X1 U7904 ( .A1(n11697), .A2(n7442), .ZN(n7447) );
  NOR2_X1 U7905 ( .A1(n7446), .A2(n7441), .ZN(n7448) );
  AOI221_X1 U7906 ( .B1(n7446), .B2(n7441), .C1(n7448), .C2(n7447), .A(n7443), 
        .ZN(n7449) );
  NOR3_X1 U7907 ( .A1(n7770), .A2(n8305), .A3(n9797), .ZN(n7450) );
  AOI211_X1 U7908 ( .C1(n7439), .C2(n8337), .A(n7449), .B(n7450), .ZN(n7451)
         );
  NOR3_X1 U7909 ( .A1(n9795), .A2(n9085), .A3(n7690), .ZN(n7452) );
  XNOR2_X1 U7910 ( .A(n8059), .B(n8306), .ZN(n7453) );
  AOI21_X1 U7911 ( .B1(n7453), .B2(n9803), .A(n7452), .ZN(n7454) );
  NAND2_X1 U7912 ( .A1(n7451), .A2(n7454), .ZN(n7455) );
  AOI22_X1 U7913 ( .A1(n9923), .A2(n10021), .B1(n7759), .B2(n9176), .ZN(n7456)
         );
  INV_X1 U7914 ( .A(n9920), .ZN(n7457) );
  OAI22_X1 U7915 ( .A1(n9919), .A2(n9939), .B1(n9880), .B2(n7457), .ZN(n7458)
         );
  INV_X1 U7916 ( .A(n9924), .ZN(n7459) );
  OAI22_X1 U7917 ( .A1(n9938), .A2(n10027), .B1(n9918), .B2(n7459), .ZN(n7460)
         );
  AOI211_X1 U7918 ( .C1(n10284), .C2(n11698), .A(n7458), .B(n7460), .ZN(n7461)
         );
  AOI22_X1 U7919 ( .A1(n10286), .A2(n9947), .B1(n9922), .B2(n10023), .ZN(n7462) );
  NAND3_X1 U7920 ( .A1(n7456), .A2(n7461), .A3(n7462), .ZN(n7463) );
  AOI222_X1 U7921 ( .A1(n7455), .A2(n10281), .B1(n7764), .B2(DRAM_ADDRESS[3]), 
        .C1(n7463), .C2(n10280), .ZN(n2133) );
  AND2_X1 U7922 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[13] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N17 ) );
  AND2_X1 U7923 ( .A1(n8462), .A2(\DataPath/RF/internal_out1[14] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N18 ) );
  OAI22_X1 U7924 ( .A1(n8261), .A2(n8428), .B1(n7740), .B2(n9904), .ZN(n7464)
         );
  XNOR2_X1 U7925 ( .A(n8060), .B(n7464), .ZN(\DP_OP_751_130_6421/n1730 ) );
  OAI21_X1 U7926 ( .B1(\DataPath/WRF_CUhw/curr_addr[21] ), .B2(n7776), .A(
        n8047), .ZN(n8046) );
  NAND2_X1 U7927 ( .A1(n9453), .A2(n9449), .ZN(n7465) );
  OAI21_X1 U7928 ( .B1(n11729), .B2(n11728), .A(n10276), .ZN(n7466) );
  OAI221_X1 U7929 ( .B1(n7465), .B2(n9450), .C1(n7465), .C2(n7466), .A(n9452), 
        .ZN(n9359) );
  NAND2_X1 U7930 ( .A1(n8021), .A2(n8033), .ZN(n7467) );
  NAND2_X1 U7931 ( .A1(n7651), .A2(n8035), .ZN(n7468) );
  OAI211_X1 U7932 ( .C1(n8037), .C2(n8032), .A(n7467), .B(n7468), .ZN(n8017)
         );
  INV_X1 U7933 ( .A(\DP_OP_751_130_6421/n902 ), .ZN(n7469) );
  INV_X1 U7934 ( .A(n8061), .ZN(n7470) );
  OAI21_X1 U7935 ( .B1(n8061), .B2(\DP_OP_751_130_6421/n902 ), .A(
        \DP_OP_751_130_6421/n967 ), .ZN(n7471) );
  OAI21_X1 U7936 ( .B1(n7469), .B2(n7470), .A(n7471), .ZN(
        \DP_OP_751_130_6421/n867 ) );
  INV_X1 U7937 ( .A(\DP_OP_751_130_6421/n597 ), .ZN(n7472) );
  NAND2_X1 U7938 ( .A1(n9528), .A2(n9609), .ZN(n7473) );
  OAI221_X1 U7939 ( .B1(n9528), .B2(\DP_OP_751_130_6421/n597 ), .C1(n9609), 
        .C2(n7472), .A(n7473), .ZN(n8926) );
  NOR2_X1 U7940 ( .A1(n7745), .A2(n8315), .ZN(n7474) );
  XOR2_X1 U7941 ( .A(\DP_OP_751_130_6421/n1477 ), .B(n7474), .Z(
        \DP_OP_751_130_6421/n1378 ) );
  NOR2_X1 U7942 ( .A1(n7745), .A2(n8315), .ZN(n7475) );
  MUX2_X1 U7943 ( .A(\DP_OP_751_130_6421/n1413 ), .B(
        \DP_OP_751_130_6421/n1477 ), .S(n7475), .Z(\DP_OP_751_130_6421/n1377 )
         );
  OAI21_X1 U7944 ( .B1(\DP_OP_751_130_6421/n1069 ), .B2(
        \DP_OP_751_130_6421/n1004 ), .A(\DP_OP_751_130_6421/n1005 ), .ZN(n7476) );
  OAI21_X1 U7945 ( .B1(n7477), .B2(n7478), .A(n7476), .ZN(
        \DP_OP_751_130_6421/n969 ) );
  INV_X1 U7946 ( .A(\DP_OP_751_130_6421/n1069 ), .ZN(n7477) );
  INV_X1 U7947 ( .A(\DP_OP_751_130_6421/n1004 ), .ZN(n7478) );
  INV_X1 U7948 ( .A(n9809), .ZN(n7479) );
  AOI21_X1 U7949 ( .B1(n9126), .B2(n9125), .A(n7479), .ZN(n9153) );
  AOI22_X1 U7950 ( .A1(\DataPath/i_PIPLIN_A[13] ), .A2(n7692), .B1(
        \DataPath/i_PIPLIN_IN1[13] ), .B2(n8443), .ZN(n7480) );
  INV_X1 U7951 ( .A(n7480), .ZN(n9966) );
  AOI22_X1 U7952 ( .A1(n9691), .A2(n9087), .B1(n8325), .B2(n9692), .ZN(n7481)
         );
  NOR2_X1 U7953 ( .A1(n9137), .A2(n9330), .ZN(n7482) );
  INV_X1 U7954 ( .A(n9685), .ZN(n7483) );
  INV_X1 U7955 ( .A(n9682), .ZN(n7484) );
  OAI22_X1 U7956 ( .A1(n9140), .A2(n7483), .B1(n9139), .B2(n7484), .ZN(n7485)
         );
  AOI211_X1 U7957 ( .C1(n9683), .C2(n9689), .A(n7482), .B(n7485), .ZN(n7486)
         );
  OAI211_X1 U7958 ( .C1(n9633), .C2(n9324), .A(n7481), .B(n7486), .ZN(n11719)
         );
  AND3_X1 U7959 ( .A1(n8242), .A2(n8238), .A3(n11635), .ZN(n7487) );
  OAI21_X1 U7960 ( .B1(n877), .B2(n7487), .A(n11660), .ZN(n11666) );
  INV_X1 U7961 ( .A(\DataPath/RF/PUSH_ADDRGEN/curr_addr[15] ), .ZN(n7488) );
  NOR2_X1 U7962 ( .A1(n10821), .A2(n7488), .ZN(n11846) );
  NAND2_X1 U7963 ( .A1(IR[2]), .A2(n10063), .ZN(n7489) );
  OAI22_X1 U7964 ( .A1(n11830), .A2(n10217), .B1(n10045), .B2(n7489), .ZN(
        n7490) );
  NOR3_X1 U7965 ( .A1(n10057), .A2(n10051), .A3(n7490), .ZN(n10242) );
  XOR2_X1 U7966 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[20] ), .Z(n7491)
         );
  OAI21_X1 U7967 ( .B1(\DP_OP_1091J1_126_6973/n13 ), .B2(n7491), .A(n10822), 
        .ZN(n7492) );
  AOI21_X1 U7968 ( .B1(\DP_OP_1091J1_126_6973/n13 ), .B2(n7491), .A(n7492), 
        .ZN(DRAMRF_ADDRESS[20]) );
  AOI21_X1 U7969 ( .B1(n8825), .B2(n8029), .A(n8030), .ZN(n7493) );
  INV_X1 U7970 ( .A(n7493), .ZN(n10152) );
  INV_X1 U7971 ( .A(n11678), .ZN(n7494) );
  XOR2_X1 U7972 ( .A(n10157), .B(IRAM_ADDRESS[30]), .Z(n7495) );
  AOI222_X1 U7973 ( .A1(n7494), .A2(n7495), .B1(i_RD1[30]), .B2(n10267), .C1(
        n10266), .C2(IRAM_ADDRESS[30]), .ZN(n8256) );
  AND2_X1 U7974 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[14] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N18 ) );
  AND2_X1 U7975 ( .A1(n8468), .A2(\DataPath/RF/internal_out1[13] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N17 ) );
  XNOR2_X1 U7976 ( .A(\DataPath/ALUhw/MULT/mux_out[2][31] ), .B(n8057), .ZN(
        n7496) );
  NAND2_X1 U7977 ( .A1(\DP_OP_751_130_6421/n1692 ), .A2(n7933), .ZN(n7497) );
  XNOR2_X1 U7978 ( .A(n7497), .B(n7496), .ZN(n7903) );
  AOI22_X1 U7979 ( .A1(n8275), .A2(n8272), .B1(n589), .B2(n8282), .ZN(n7498)
         );
  INV_X1 U7980 ( .A(n7498), .ZN(n8250) );
  NAND2_X1 U7981 ( .A1(n10331), .A2(n10338), .ZN(n7499) );
  OAI21_X1 U7982 ( .B1(n7499), .B2(n10334), .A(n10335), .ZN(n10337) );
  INV_X1 U7983 ( .A(n8077), .ZN(n7500) );
  NAND3_X1 U7984 ( .A1(n8076), .A2(n8048), .A3(n7500), .ZN(n8047) );
  OAI21_X1 U7985 ( .B1(n10299), .B2(n9290), .A(n9291), .ZN(n9393) );
  OAI21_X1 U7986 ( .B1(n7975), .B2(n7736), .A(\intadd_1/A[3] ), .ZN(
        \intadd_1/n17 ) );
  INV_X1 U7987 ( .A(n8026), .ZN(n7501) );
  NAND2_X1 U7988 ( .A1(n8022), .A2(n7501), .ZN(n8012) );
  NOR2_X1 U7989 ( .A1(n7949), .A2(\DP_OP_751_130_6421/n355 ), .ZN(n7502) );
  AOI211_X1 U7990 ( .C1(n7949), .C2(\DP_OP_751_130_6421/n355 ), .A(
        \DP_OP_751_130_6421/n354 ), .B(n7502), .ZN(\DP_OP_751_130_6421/n60 )
         );
  INV_X1 U7991 ( .A(\DP_OP_751_130_6421/n392 ), .ZN(n7503) );
  INV_X1 U7992 ( .A(\DP_OP_751_130_6421/n393 ), .ZN(n7504) );
  OAI21_X1 U7993 ( .B1(\DP_OP_751_130_6421/n393 ), .B2(
        \DP_OP_751_130_6421/n392 ), .A(\DP_OP_751_130_6421/n457 ), .ZN(n7505)
         );
  OAI21_X1 U7994 ( .B1(n7503), .B2(n7504), .A(n7505), .ZN(
        \DP_OP_751_130_6421/n357 ) );
  AOI211_X1 U7995 ( .C1(n11720), .C2(n9913), .A(n11685), .B(n9040), .ZN(n9317)
         );
  INV_X1 U7996 ( .A(n8059), .ZN(n7506) );
  OAI22_X1 U7997 ( .A1(n7740), .A2(n8311), .B1(n8261), .B2(n8308), .ZN(n7507)
         );
  XOR2_X1 U7998 ( .A(n8060), .B(n7507), .Z(n7508) );
  NOR2_X1 U7999 ( .A1(n7506), .A2(n7508), .ZN(\DP_OP_751_130_6421/n1686 ) );
  XNOR2_X1 U8000 ( .A(n8059), .B(n7508), .ZN(\DP_OP_751_130_6421/n1684 ) );
  AOI22_X1 U8001 ( .A1(\DataPath/i_PIPLIN_A[4] ), .A2(n7732), .B1(
        \DataPath/i_PIPLIN_IN1[4] ), .B2(n8443), .ZN(n7509) );
  INV_X1 U8002 ( .A(n7509), .ZN(n9099) );
  NOR3_X1 U8003 ( .A1(n380), .A2(DATA_SIZE[1]), .A3(n10733), .ZN(n7510) );
  OAI21_X1 U8004 ( .B1(n11616), .B2(n217), .A(n7510), .ZN(n10783) );
  INV_X1 U8005 ( .A(n10148), .ZN(n7511) );
  AND3_X1 U8006 ( .A1(n10151), .A2(n8824), .A3(n7511), .ZN(n8029) );
  OAI21_X1 U8007 ( .B1(\DP_OP_751_130_6421/n495 ), .B2(
        \DP_OP_751_130_6421/n494 ), .A(\DP_OP_751_130_6421/n559 ), .ZN(n7512)
         );
  OAI21_X1 U8008 ( .B1(n7513), .B2(n7514), .A(n7512), .ZN(
        \DP_OP_751_130_6421/n459 ) );
  INV_X1 U8009 ( .A(\DP_OP_751_130_6421/n494 ), .ZN(n7513) );
  INV_X1 U8010 ( .A(\DP_OP_751_130_6421/n495 ), .ZN(n7514) );
  AOI22_X1 U8011 ( .A1(n7738), .A2(\DataPath/i_PIPLIN_IN2[8] ), .B1(
        \DataPath/i_PIPLIN_B[8] ), .B2(n8455), .ZN(n7515) );
  INV_X1 U8012 ( .A(n7515), .ZN(n9182) );
  INV_X1 U8013 ( .A(n9966), .ZN(n7516) );
  OAI21_X1 U8014 ( .B1(n9237), .B2(n7516), .A(n9768), .ZN(n9961) );
  NOR2_X1 U8015 ( .A1(n7940), .A2(n8149), .ZN(n7517) );
  AOI21_X1 U8016 ( .B1(n7940), .B2(\DataPath/i_PIPLIN_IN2[17] ), .A(n7517), 
        .ZN(n8449) );
  AOI22_X1 U8017 ( .A1(n9075), .A2(n9683), .B1(n9198), .B2(n9024), .ZN(n7518)
         );
  INV_X1 U8018 ( .A(n9547), .ZN(n7519) );
  AOI22_X1 U8019 ( .A1(n9687), .A2(n9496), .B1(n9500), .B2(n7519), .ZN(n7520)
         );
  OAI211_X1 U8020 ( .C1(n9019), .C2(n9498), .A(n7518), .B(n7520), .ZN(n7521)
         );
  AOI21_X1 U8021 ( .B1(n9516), .B2(n9031), .A(n7521), .ZN(n7522) );
  OAI21_X1 U8022 ( .B1(n8308), .B2(n9049), .A(n7522), .ZN(n9921) );
  NAND2_X1 U8023 ( .A1(n8093), .A2(\intadd_0/n17 ), .ZN(n7523) );
  OAI211_X1 U8024 ( .C1(n8254), .C2(n8818), .A(\intadd_0/n14 ), .B(n7523), 
        .ZN(n8253) );
  XOR2_X1 U8025 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[18] ), .Z(n7524)
         );
  OAI21_X1 U8026 ( .B1(\DP_OP_1091J1_126_6973/n15 ), .B2(n7524), .A(n10822), 
        .ZN(n7525) );
  AOI21_X1 U8027 ( .B1(\DP_OP_1091J1_126_6973/n15 ), .B2(n7524), .A(n7525), 
        .ZN(DRAMRF_ADDRESS[18]) );
  XOR2_X1 U8028 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[21] ), .Z(n7526)
         );
  OAI21_X1 U8029 ( .B1(n7776), .B2(\DataPath/WRF_CUhw/curr_addr[20] ), .A(
        \DP_OP_1091J1_126_6973/n13 ), .ZN(n7527) );
  NAND2_X1 U8030 ( .A1(n7527), .A2(n8079), .ZN(n7528) );
  OAI21_X1 U8031 ( .B1(n7526), .B2(n7528), .A(n10822), .ZN(n7529) );
  AOI21_X1 U8032 ( .B1(n7526), .B2(n7528), .A(n7529), .ZN(DRAMRF_ADDRESS[21])
         );
  AOI222_X1 U8033 ( .A1(n11643), .A2(n7648), .B1(n11645), .B2(
        \DataPath/RF/c_win[3] ), .C1(\DataPath/RF/c_win[0] ), .C2(n11644), 
        .ZN(n7530) );
  NOR2_X1 U8034 ( .A1(RST), .A2(n7530), .ZN(n7065) );
  INV_X1 U8035 ( .A(IR[1]), .ZN(n7531) );
  NAND2_X1 U8036 ( .A1(n7969), .A2(n8287), .ZN(n7532) );
  NAND2_X1 U8037 ( .A1(n10232), .A2(n7532), .ZN(n7533) );
  AOI22_X1 U8038 ( .A1(n10060), .A2(n10059), .B1(n10219), .B2(n7533), .ZN(
        n7534) );
  OAI222_X1 U8039 ( .A1(n11620), .A2(n10058), .B1(n11828), .B2(n8084), .C1(
        n11830), .C2(n7534), .ZN(n7535) );
  AOI21_X1 U8040 ( .B1(n10057), .B2(n7531), .A(n7535), .ZN(n7536) );
  NAND3_X1 U8041 ( .A1(n10061), .A2(n8196), .A3(n10063), .ZN(n7537) );
  NAND2_X1 U8042 ( .A1(n7536), .A2(n7537), .ZN(n7088) );
  NOR2_X1 U8043 ( .A1(n166), .A2(n8294), .ZN(n7538) );
  AOI21_X1 U8044 ( .B1(IRAM_DATA[29]), .B2(n10258), .A(n7538), .ZN(n8255) );
  NAND2_X1 U8045 ( .A1(n8072), .A2(\DP_OP_751_130_6421/n136 ), .ZN(n7539) );
  XNOR2_X1 U8046 ( .A(n7539), .B(\DP_OP_751_130_6421/n137 ), .ZN(n7540) );
  XOR2_X1 U8047 ( .A(n9158), .B(n7786), .Z(n7541) );
  OAI21_X1 U8048 ( .B1(n9150), .B2(n11713), .A(n9149), .ZN(n7542) );
  OAI21_X1 U8049 ( .B1(n7541), .B2(n7542), .A(n9810), .ZN(n7543) );
  AOI21_X1 U8050 ( .B1(n7541), .B2(n7542), .A(n7543), .ZN(n7544) );
  NAND2_X1 U8051 ( .A1(n9149), .A2(n9152), .ZN(n7545) );
  OAI21_X1 U8052 ( .B1(n7541), .B2(n7545), .A(n10278), .ZN(n7546) );
  AOI21_X1 U8053 ( .B1(n7541), .B2(n7545), .A(n7546), .ZN(n7547) );
  AOI211_X1 U8054 ( .C1(n7540), .C2(n8337), .A(n7544), .B(n7547), .ZN(n7548)
         );
  NAND2_X1 U8055 ( .A1(\DP_OP_751_130_6421/n1515 ), .A2(n7786), .ZN(n7549) );
  NAND2_X1 U8056 ( .A1(n9850), .A2(n7549), .ZN(n7550) );
  OAI221_X1 U8057 ( .B1(n7549), .B2(n9992), .C1(\DP_OP_751_130_6421/n1515 ), 
        .C2(n7786), .A(n7550), .ZN(n7551) );
  NAND3_X1 U8058 ( .A1(n8446), .A2(n9990), .A3(n9157), .ZN(n7552) );
  NAND3_X1 U8059 ( .A1(n7548), .A2(n7551), .A3(n7552), .ZN(n7553) );
  AOI22_X1 U8060 ( .A1(n9974), .A2(n10286), .B1(n7759), .B2(n11719), .ZN(n7554) );
  AOI22_X1 U8061 ( .A1(n9211), .A2(n10021), .B1(n9920), .B2(n10013), .ZN(n7555) );
  AOI22_X1 U8062 ( .A1(n9947), .A2(n10010), .B1(n10284), .B2(n9176), .ZN(n7556) );
  AOI22_X1 U8063 ( .A1(n9946), .A2(n9978), .B1(n10023), .B2(n9979), .ZN(n7557)
         );
  NAND2_X1 U8064 ( .A1(n7556), .A2(n7557), .ZN(n7558) );
  AOI21_X1 U8065 ( .B1(n9922), .B2(n10020), .A(n7558), .ZN(n7559) );
  NAND3_X1 U8066 ( .A1(n7554), .A2(n7555), .A3(n7559), .ZN(n7560) );
  AOI222_X1 U8067 ( .A1(n7553), .A2(n10281), .B1(n7764), .B2(DRAM_ADDRESS[7]), 
        .C1(n7560), .C2(n10280), .ZN(n2011) );
  AOI22_X1 U8068 ( .A1(IRAM_ADDRESS[23]), .A2(n10266), .B1(n10267), .B2(
        i_RD1[23]), .ZN(n7561) );
  INV_X1 U8069 ( .A(\intadd_2/n33 ), .ZN(n7562) );
  OAI21_X1 U8070 ( .B1(\intadd_2/n22 ), .B2(n7562), .A(\intadd_2/n23 ), .ZN(
        n7563) );
  INV_X1 U8071 ( .A(\intadd_2/n18 ), .ZN(n7564) );
  NOR2_X1 U8072 ( .A1(\intadd_2/n17 ), .A2(n7564), .ZN(n7565) );
  NAND2_X1 U8073 ( .A1(n7565), .A2(n7563), .ZN(n7566) );
  OAI211_X1 U8074 ( .C1(n7565), .C2(n7563), .A(n7566), .B(n8421), .ZN(n7567)
         );
  NAND2_X1 U8075 ( .A1(n7561), .A2(n7567), .ZN(n7033) );
  AND2_X1 U8076 ( .A1(n8458), .A2(\DataPath/RF/internal_out2[30] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N34 ) );
  AND2_X1 U8077 ( .A1(n8470), .A2(\DataPath/RF/internal_out2[28] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N32 ) );
  AND2_X1 U8078 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[27] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N31 ) );
  AND2_X1 U8079 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[26] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N30 ) );
  AND2_X1 U8080 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[25] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N29 ) );
  AND2_X1 U8081 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[24] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N28 ) );
  AND2_X1 U8082 ( .A1(n8463), .A2(\DataPath/RF/internal_out2[23] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N27 ) );
  AND2_X1 U8083 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[22] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N26 ) );
  AND2_X1 U8084 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[21] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N25 ) );
  AND2_X1 U8085 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[20] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N24 ) );
  AND2_X1 U8086 ( .A1(n8465), .A2(\DataPath/RF/internal_out2[11] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N15 ) );
  AND2_X1 U8087 ( .A1(n8468), .A2(\DataPath/RF/internal_out2[10] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N14 ) );
  AND2_X1 U8088 ( .A1(n8466), .A2(\DataPath/RF/internal_out2[9] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N13 ) );
  AND2_X1 U8089 ( .A1(n8458), .A2(\DataPath/RF/internal_out2[8] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N12 ) );
  AND2_X1 U8090 ( .A1(n8465), .A2(\DataPath/RF/internal_out2[7] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N11 ) );
  AND2_X1 U8091 ( .A1(n8464), .A2(\DataPath/RF/internal_out2[6] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N10 ) );
  AND2_X1 U8092 ( .A1(n8467), .A2(\DataPath/RF/internal_out2[5] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N9 ) );
  AND2_X1 U8093 ( .A1(n8464), .A2(\DataPath/RF/internal_out2[4] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N8 ) );
  AND2_X1 U8094 ( .A1(n8468), .A2(\DataPath/RF/internal_out2[3] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N7 ) );
  AND2_X1 U8095 ( .A1(n8461), .A2(\DataPath/RF/internal_out2[2] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N6 ) );
  AND2_X1 U8096 ( .A1(n8462), .A2(\DataPath/RF/internal_out2[1] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N5 ) );
  AND2_X1 U8097 ( .A1(n8457), .A2(\DataPath/RF/internal_out2[0] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N4 ) );
  AND2_X1 U8098 ( .A1(n8469), .A2(\DataPath/RF/internal_out1[12] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N16 ) );
  AND2_X1 U8099 ( .A1(n8469), .A2(\DataPath/RF/internal_out1[31] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N35 ) );
  OAI22_X1 U8100 ( .A1(n7740), .A2(n8428), .B1(n9608), .B2(n8261), .ZN(n7929)
         );
  OAI22_X1 U8101 ( .A1(n8321), .A2(n9796), .B1(n8317), .B2(n8941), .ZN(n7568)
         );
  XNOR2_X1 U8102 ( .A(n7690), .B(n7568), .ZN(n7569) );
  XOR2_X1 U8103 ( .A(\DataPath/ALUhw/MULT/mux_out[0][13] ), .B(n7974), .Z(
        n7570) );
  XOR2_X1 U8104 ( .A(n7569), .B(n7570), .Z(\DP_OP_751_130_6421/n1662 ) );
  NOR2_X1 U8105 ( .A1(n7569), .A2(n7570), .ZN(\DP_OP_751_130_6421/n1661 ) );
  INV_X1 U8106 ( .A(\DP_OP_751_130_6421/n291 ), .ZN(n7571) );
  NAND2_X1 U8107 ( .A1(n9377), .A2(n9824), .ZN(n7572) );
  OAI221_X1 U8108 ( .B1(n9377), .B2(\DP_OP_751_130_6421/n291 ), .C1(n9824), 
        .C2(n7571), .A(n7572), .ZN(n7573) );
  OAI22_X1 U8109 ( .A1(n8316), .A2(n7573), .B1(n8311), .B2(n8942), .ZN(
        \DataPath/ALUhw/MULT/mux_out[15][31] ) );
  INV_X1 U8110 ( .A(n10333), .ZN(n7574) );
  AOI221_X1 U8111 ( .B1(n10331), .B2(n7574), .C1(n10334), .C2(n7574), .A(
        n10332), .ZN(n7575) );
  AOI221_X1 U8112 ( .B1(n7575), .B2(n10315), .C1(n10316), .C2(n10315), .A(
        n10311), .ZN(n7576) );
  NOR2_X1 U8113 ( .A1(n7576), .A2(n10317), .ZN(n10353) );
  INV_X1 U8114 ( .A(n11846), .ZN(n7577) );
  NAND3_X1 U8115 ( .A1(n10293), .A2(DRAMRF_READY), .A3(n7577), .ZN(n7982) );
  NOR3_X1 U8116 ( .A1(n7736), .A2(n7975), .A3(\intadd_1/A[3] ), .ZN(
        \intadd_1/n16 ) );
  NOR2_X1 U8117 ( .A1(IRAM_ADDRESS[29]), .A2(IRAM_ADDRESS[28]), .ZN(n7578) );
  NAND2_X1 U8118 ( .A1(n10175), .A2(n7578), .ZN(n7962) );
  INV_X1 U8119 ( .A(\DP_OP_751_130_6421/n495 ), .ZN(n7579) );
  NAND2_X1 U8120 ( .A1(n9517), .A2(n9847), .ZN(n7580) );
  OAI221_X1 U8121 ( .B1(n9517), .B2(\DP_OP_751_130_6421/n495 ), .C1(n9847), 
        .C2(n7579), .A(n7580), .ZN(n8930) );
  OAI21_X1 U8122 ( .B1(n10299), .B2(n9498), .A(n9298), .ZN(n7581) );
  INV_X1 U8123 ( .A(n7581), .ZN(n9503) );
  INV_X1 U8124 ( .A(\DP_OP_751_130_6421/n800 ), .ZN(n7582) );
  INV_X1 U8125 ( .A(n8062), .ZN(n7583) );
  OAI21_X1 U8126 ( .B1(n8062), .B2(\DP_OP_751_130_6421/n800 ), .A(
        \DP_OP_751_130_6421/n865 ), .ZN(n7584) );
  OAI21_X1 U8127 ( .B1(n7582), .B2(n7583), .A(n7584), .ZN(
        \DP_OP_751_130_6421/n765 ) );
  INV_X1 U8128 ( .A(n9082), .ZN(n7585) );
  AOI21_X1 U8129 ( .B1(i_ALU_OP[2]), .B2(n7693), .A(n7585), .ZN(n9225) );
  OAI22_X1 U8130 ( .A1(n7740), .A2(n8308), .B1(n8260), .B2(n8305), .ZN(n7586)
         );
  XNOR2_X1 U8131 ( .A(n8060), .B(n7586), .ZN(n7587) );
  AND2_X1 U8132 ( .A1(n7587), .A2(\DP_OP_751_130_6421/n1686 ), .ZN(
        \DP_OP_751_130_6421/n1681 ) );
  XOR2_X1 U8133 ( .A(n7587), .B(\DP_OP_751_130_6421/n1686 ), .Z(
        \DP_OP_751_130_6421/n1682 ) );
  AOI211_X1 U8134 ( .C1(n11720), .C2(n9085), .A(n9006), .B(n11685), .ZN(n7588)
         );
  INV_X1 U8135 ( .A(n7588), .ZN(n9476) );
  INV_X1 U8136 ( .A(IRAM_ADDRESS[19]), .ZN(n7589) );
  NAND2_X1 U8137 ( .A1(n10151), .A2(n8831), .ZN(n7590) );
  OAI22_X1 U8138 ( .A1(n10150), .A2(n7589), .B1(n10146), .B2(n7590), .ZN(n8030) );
  INV_X1 U8139 ( .A(\DP_OP_751_130_6421/n698 ), .ZN(n7591) );
  INV_X1 U8140 ( .A(n7782), .ZN(n7592) );
  OAI21_X1 U8141 ( .B1(n7782), .B2(\DP_OP_751_130_6421/n698 ), .A(
        \DP_OP_751_130_6421/n763 ), .ZN(n7593) );
  OAI21_X1 U8142 ( .B1(n7591), .B2(n7592), .A(n7593), .ZN(
        \DP_OP_751_130_6421/n663 ) );
  XNOR2_X1 U8143 ( .A(n7633), .B(\DP_OP_751_130_6421/n357 ), .ZN(n7594) );
  NAND2_X1 U8144 ( .A1(n7881), .A2(n7821), .ZN(n7595) );
  XNOR2_X1 U8145 ( .A(n7595), .B(n7594), .ZN(\DataPath/ALUhw/i_Q_EXTENDED[61] ) );
  INV_X1 U8146 ( .A(n9782), .ZN(n7596) );
  NOR2_X1 U8147 ( .A1(n9239), .A2(n7596), .ZN(n9963) );
  INV_X1 U8148 ( .A(n9669), .ZN(n7597) );
  AOI22_X1 U8149 ( .A1(n9025), .A2(n9415), .B1(n9024), .B2(n7597), .ZN(n7598)
         );
  INV_X1 U8150 ( .A(n9104), .ZN(n7599) );
  AOI22_X1 U8151 ( .A1(n7792), .A2(n8981), .B1(n7775), .B2(n8980), .ZN(n7600)
         );
  OAI21_X1 U8152 ( .B1(n7599), .B2(n9411), .A(n9683), .ZN(n7601) );
  AND2_X1 U8153 ( .A1(n7601), .A2(n7600), .ZN(n7602) );
  OAI211_X1 U8154 ( .C1(n9019), .C2(n9671), .A(n7598), .B(n7602), .ZN(n9924)
         );
  INV_X1 U8155 ( .A(n10239), .ZN(n7603) );
  NAND3_X1 U8156 ( .A1(IR[2]), .A2(IR[1]), .A3(n7603), .ZN(n10243) );
  XOR2_X1 U8157 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[17] ), .Z(n7604)
         );
  OAI21_X1 U8158 ( .B1(n7704), .B2(n7604), .A(n10822), .ZN(n7605) );
  AOI21_X1 U8159 ( .B1(n7704), .B2(n7604), .A(n7605), .ZN(DRAMRF_ADDRESS[17])
         );
  AOI21_X1 U8160 ( .B1(n7936), .B2(\DP_OP_1091J1_126_6973/n15 ), .A(n7935), 
        .ZN(n7606) );
  XNOR2_X1 U8161 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[19] ), .ZN(n7607) );
  OAI21_X1 U8162 ( .B1(n7606), .B2(n7607), .A(n10822), .ZN(n7608) );
  AOI21_X1 U8163 ( .B1(n7606), .B2(n7607), .A(n7608), .ZN(DRAMRF_ADDRESS[19])
         );
  XOR2_X1 U8164 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[22] ), .Z(n7609)
         );
  INV_X1 U8165 ( .A(n8079), .ZN(n7610) );
  AOI21_X1 U8166 ( .B1(\DP_OP_1091J1_126_6973/n13 ), .B2(n8044), .A(n7610), 
        .ZN(n7611) );
  NOR2_X1 U8167 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[21] ), .ZN(
        n7612) );
  OAI21_X1 U8168 ( .B1(n7611), .B2(n7612), .A(n8078), .ZN(n7613) );
  OAI21_X1 U8169 ( .B1(n7609), .B2(n7613), .A(n10822), .ZN(n7614) );
  AOI21_X1 U8170 ( .B1(n7609), .B2(n7613), .A(n7614), .ZN(DRAMRF_ADDRESS[22])
         );
  XOR2_X1 U8171 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[28] ), .Z(n7615)
         );
  OAI21_X1 U8172 ( .B1(\DP_OP_1091J1_126_6973/n5 ), .B2(n7615), .A(n10822), 
        .ZN(n7616) );
  AOI21_X1 U8173 ( .B1(\DP_OP_1091J1_126_6973/n5 ), .B2(n7615), .A(n7616), 
        .ZN(DRAMRF_ADDRESS[28]) );
  INV_X1 U8174 ( .A(n10822), .ZN(n7617) );
  NOR2_X1 U8175 ( .A1(n8028), .A2(n7617), .ZN(DRAMRF_ADDRESS[30]) );
  AND2_X1 U8176 ( .A1(\C620/DATA2_31 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[31])
         );
  NOR2_X1 U8177 ( .A1(n7907), .A2(n8145), .ZN(n7618) );
  AOI21_X1 U8178 ( .B1(n7907), .B2(\DataPath/i_PIPLIN_IN2[11] ), .A(n7618), 
        .ZN(n7771) );
  AOI22_X1 U8179 ( .A1(n7940), .A2(\DataPath/i_PIPLIN_IN2[14] ), .B1(
        \DataPath/i_PIPLIN_B[14] ), .B2(n8455), .ZN(n7619) );
  INV_X1 U8180 ( .A(n7619), .ZN(n9780) );
  AOI222_X1 U8181 ( .A1(n11643), .A2(\DataPath/RF/c_win[2] ), .B1(n11644), 
        .B2(\DataPath/RF/c_win[3] ), .C1(n11645), .C2(\DataPath/RF/c_win[1] ), 
        .ZN(n7620) );
  NOR2_X1 U8182 ( .A1(RST), .A2(n7620), .ZN(n7067) );
  NOR2_X1 U8183 ( .A1(n7695), .A2(n8253), .ZN(n7621) );
  XOR2_X1 U8184 ( .A(n10187), .B(n7621), .Z(n7622) );
  AOI22_X1 U8185 ( .A1(n10266), .A2(IRAM_ADDRESS[16]), .B1(i_RD1[16]), .B2(
        n10267), .ZN(n7623) );
  OAI21_X1 U8186 ( .B1(n11678), .B2(n7622), .A(n7623), .ZN(n7040) );
  INV_X1 U8187 ( .A(n10217), .ZN(n7624) );
  AOI211_X1 U8188 ( .C1(IR[31]), .C2(n10234), .A(n10218), .B(n7624), .ZN(n7625) );
  INV_X1 U8189 ( .A(n8287), .ZN(n7626) );
  OAI222_X1 U8190 ( .A1(n7626), .A2(n8090), .B1(n7626), .B2(n10219), .C1(
        n10303), .C2(n8287), .ZN(n7627) );
  OAI211_X1 U8191 ( .C1(n10221), .C2(n10220), .A(n7625), .B(n7627), .ZN(
        \CU_I/CW[UNSIGNED_ID] ) );
  AND2_X1 U8192 ( .A1(n8469), .A2(\DataPath/RF/internal_out2[12] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N16 ) );
  AND2_X1 U8193 ( .A1(n8464), .A2(\DataPath/RF/internal_out1[30] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N34 ) );
  AND2_X1 U8194 ( .A1(n8459), .A2(\DataPath/RF/internal_out1[28] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N32 ) );
  AND2_X1 U8195 ( .A1(n8460), .A2(\DataPath/RF/internal_out1[27] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N31 ) );
  AND2_X1 U8196 ( .A1(n8465), .A2(\DataPath/RF/internal_out1[26] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N30 ) );
  AND2_X1 U8197 ( .A1(n8468), .A2(\DataPath/RF/internal_out1[25] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N29 ) );
  AND2_X1 U8198 ( .A1(n8459), .A2(\DataPath/RF/internal_out1[24] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N28 ) );
  AND2_X1 U8199 ( .A1(n8468), .A2(\DataPath/RF/internal_out1[23] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N27 ) );
  AND2_X1 U8200 ( .A1(n8459), .A2(\DataPath/RF/internal_out1[22] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N26 ) );
  AND2_X1 U8201 ( .A1(n8458), .A2(\DataPath/RF/internal_out1[21] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N25 ) );
  AND2_X1 U8202 ( .A1(n8469), .A2(\DataPath/RF/internal_out1[20] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N24 ) );
  AND2_X1 U8203 ( .A1(n8460), .A2(\DataPath/RF/internal_out1[11] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N15 ) );
  AND2_X1 U8204 ( .A1(n8461), .A2(\DataPath/RF/internal_out1[10] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N14 ) );
  AND2_X1 U8205 ( .A1(n8458), .A2(\DataPath/RF/internal_out1[9] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N13 ) );
  AND2_X1 U8206 ( .A1(n8467), .A2(\DataPath/RF/internal_out1[8] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N12 ) );
  AND2_X1 U8207 ( .A1(n8461), .A2(\DataPath/RF/internal_out1[7] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N11 ) );
  AND2_X1 U8208 ( .A1(n8457), .A2(\DataPath/RF/internal_out1[6] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N10 ) );
  AND2_X1 U8209 ( .A1(n8463), .A2(\DataPath/RF/internal_out1[5] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N9 ) );
  AND2_X1 U8210 ( .A1(n8461), .A2(\DataPath/RF/internal_out1[4] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N8 ) );
  AND2_X1 U8211 ( .A1(n8465), .A2(\DataPath/RF/internal_out1[3] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N7 ) );
  AND2_X1 U8212 ( .A1(n8462), .A2(\DataPath/RF/internal_out1[2] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N6 ) );
  AND2_X1 U8213 ( .A1(n8463), .A2(\DataPath/RF/internal_out1[1] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N5 ) );
  AND2_X1 U8214 ( .A1(n8468), .A2(\DataPath/RF/internal_out1[0] ), .ZN(
        \DataPath/RF/RDPORT0_OUTLATCH/N4 ) );
  AND2_X1 U8215 ( .A1(n8465), .A2(\DataPath/RF/internal_out2[31] ), .ZN(
        \DataPath/RF/RDPORT1_OUTLATCH/N35 ) );
  CLKBUF_X3 U8216 ( .A(n465), .Z(n7731) );
  INV_X1 U8217 ( .A(n465), .ZN(n8443) );
  BUF_X2 U8218 ( .A(n465), .Z(n7732) );
  BUF_X1 U8219 ( .A(\DP_OP_751_130_6421/n64 ), .Z(n7628) );
  BUF_X1 U8220 ( .A(\DP_OP_751_130_6421/n72 ), .Z(n7629) );
  INV_X1 U8221 ( .A(n8116), .ZN(n7630) );
  BUF_X2 U8222 ( .A(\DP_OP_751_130_6421/n1719 ), .Z(n8058) );
  BUF_X4 U8223 ( .A(n8058), .Z(n7690) );
  NOR2_X1 U8224 ( .A1(n7631), .A2(n7632), .ZN(n7817) );
  XOR2_X1 U8225 ( .A(n7802), .B(n7827), .Z(n7631) );
  OR2_X1 U8226 ( .A1(n7804), .A2(\DP_OP_751_130_6421/n60 ), .ZN(n7632) );
  BUF_X1 U8227 ( .A(\DP_OP_751_130_6421/n356 ), .Z(n7633) );
  INV_X1 U8228 ( .A(n9516), .ZN(n7634) );
  INV_X1 U8229 ( .A(n7709), .ZN(n7635) );
  OR2_X2 U8230 ( .A1(n7709), .A2(n9062), .ZN(n8858) );
  BUF_X1 U8231 ( .A(n8819), .Z(n7636) );
  CLKBUF_X3 U8232 ( .A(\DP_OP_751_130_6421/n1515 ), .Z(n8056) );
  INV_X1 U8233 ( .A(n7709), .ZN(\DP_OP_751_130_6421/n1752 ) );
  OAI21_X1 U8234 ( .B1(n7630), .B2(\DP_OP_751_130_6421/n1752 ), .A(n8862), 
        .ZN(n7637) );
  INV_X2 U8235 ( .A(n7768), .ZN(n8321) );
  BUF_X1 U8236 ( .A(n8593), .Z(n7638) );
  OAI21_X1 U8237 ( .B1(n8572), .B2(i_RD1[8]), .A(n8558), .ZN(n7639) );
  OR2_X1 U8238 ( .A1(n8625), .A2(i_RD1[4]), .ZN(n7640) );
  BUF_X1 U8239 ( .A(\DP_OP_751_130_6421/n79 ), .Z(n7641) );
  BUF_X1 U8240 ( .A(\DP_OP_751_130_6421/n82 ), .Z(n7642) );
  BUF_X1 U8241 ( .A(\DP_OP_751_130_6421/n90 ), .Z(n7643) );
  NAND2_X1 U8242 ( .A1(n7736), .A2(n8811), .ZN(n10210) );
  AND2_X1 U8243 ( .A1(n7644), .A2(n7645), .ZN(n8708) );
  NOR4_X1 U8244 ( .A1(n8697), .A2(n8717), .A3(n8696), .A4(n8745), .ZN(n7644)
         );
  AND2_X1 U8245 ( .A1(n8780), .A2(n8728), .ZN(n7645) );
  AND2_X2 U8246 ( .A1(n8799), .A2(n8001), .ZN(n8000) );
  BUF_X1 U8247 ( .A(n8718), .Z(n7646) );
  BUF_X1 U8248 ( .A(n10092), .Z(n7647) );
  AND3_X1 U8249 ( .A1(n7996), .A2(n7998), .A3(IR[0]), .ZN(n10211) );
  INV_X2 U8250 ( .A(n8084), .ZN(n8452) );
  INV_X2 U8251 ( .A(n9774), .ZN(n9775) );
  INV_X2 U8252 ( .A(n8058), .ZN(n7770) );
  BUF_X2 U8253 ( .A(n8858), .Z(n7741) );
  INV_X2 U8254 ( .A(n9711), .ZN(n7693) );
  BUF_X2 U8255 ( .A(n7709), .Z(n7880) );
  AND2_X4 U8256 ( .A1(n8845), .A2(n8844), .ZN(n9161) );
  INV_X2 U8257 ( .A(n9794), .ZN(n9796) );
  BUF_X2 U8258 ( .A(n9910), .Z(n8315) );
  NAND2_X2 U8259 ( .A1(\DataPath/i_PIPLIN_A[16] ), .A2(n7692), .ZN(n9250) );
  INV_X2 U8260 ( .A(n9327), .ZN(n8301) );
  AND2_X1 U8261 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[17] ), .ZN(
        n7649) );
  NAND2_X2 U8262 ( .A1(n10210), .A2(n8812), .ZN(n11678) );
  OR2_X2 U8263 ( .A1(n8285), .A2(n172), .ZN(n10232) );
  INV_X2 U8264 ( .A(n9782), .ZN(n9783) );
  BUF_X4 U8265 ( .A(\DP_OP_751_130_6421/n1617 ), .Z(n8057) );
  BUF_X2 U8266 ( .A(n8858), .Z(n7740) );
  OR3_X2 U8267 ( .A1(n10270), .A2(n10291), .A3(n8521), .ZN(n7721) );
  AND2_X1 U8268 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[5] ), .ZN(n7650) );
  NOR2_X1 U8269 ( .A1(n165), .A2(n167), .ZN(n10041) );
  BUF_X2 U8270 ( .A(n10041), .Z(n7720) );
  AND2_X4 U8271 ( .A1(\CU_I/CW_MEM[MEM_EN] ), .A2(n10300), .ZN(n11835) );
  INV_X2 U8272 ( .A(n7749), .ZN(n8302) );
  NAND2_X2 U8273 ( .A1(\DataPath/i_PIPLIN_A[24] ), .A2(n8442), .ZN(n9527) );
  XNOR2_X1 U8274 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[31] ), .ZN(n7651) );
  XOR2_X1 U8275 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[29] ), .Z(n7652)
         );
  OR2_X1 U8276 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[17] ), .ZN(n7653) );
  NAND2_X2 U8277 ( .A1(\DataPath/i_PIPLIN_A[29] ), .A2(n7732), .ZN(n9826) );
  XNOR2_X1 U8278 ( .A(\DataPath/ALUhw/MULT/mux_out[15][31] ), .B(
        \DP_OP_751_130_6421/n291 ), .ZN(n7654) );
  BUF_X1 U8279 ( .A(n10004), .Z(n8337) );
  OR2_X1 U8280 ( .A1(n11734), .A2(n528), .ZN(n7655) );
  INV_X2 U8281 ( .A(n9889), .ZN(n9904) );
  NOR2_X2 U8282 ( .A1(n10273), .A2(n178), .ZN(i_ADD_RS2[4]) );
  INV_X1 U8283 ( .A(n7712), .ZN(\DP_OP_1091J1_126_6973/n17 ) );
  AOI21_X1 U8284 ( .B1(\DP_OP_1091J1_126_6973/n18 ), .B2(n7713), .A(n7714), 
        .ZN(n7712) );
  OAI21_X2 U8285 ( .B1(n8446), .B2(n9130), .A(n7796), .ZN(n8872) );
  NAND2_X1 U8286 ( .A1(n9002), .A2(n9016), .ZN(n7656) );
  NAND2_X2 U8287 ( .A1(n10108), .A2(n10271), .ZN(n8295) );
  INV_X1 U8290 ( .A(n7126), .ZN(n7657) );
  AND2_X1 U8291 ( .A1(DRAMRF_ADDRESS[28]), .A2(n8468), .ZN(n7658) );
  AND2_X1 U8292 ( .A1(DRAMRF_ADDRESS[27]), .A2(n8470), .ZN(n7659) );
  AND2_X1 U8293 ( .A1(DRAMRF_ADDRESS[26]), .A2(n8466), .ZN(n7660) );
  AND2_X1 U8294 ( .A1(DRAMRF_ADDRESS[22]), .A2(n8457), .ZN(n7661) );
  AND2_X1 U8295 ( .A1(DRAMRF_ADDRESS[25]), .A2(n8460), .ZN(n7662) );
  AND2_X1 U8296 ( .A1(DRAMRF_ADDRESS[21]), .A2(n8461), .ZN(n7663) );
  AND2_X1 U8297 ( .A1(DRAMRF_ADDRESS[24]), .A2(n8470), .ZN(n7664) );
  AND2_X1 U8298 ( .A1(DRAMRF_ADDRESS[20]), .A2(n8462), .ZN(n7665) );
  AND2_X1 U8299 ( .A1(DRAMRF_ADDRESS[19]), .A2(n8467), .ZN(n7666) );
  AND2_X1 U8300 ( .A1(DRAMRF_ADDRESS[23]), .A2(n8470), .ZN(n7667) );
  AND2_X1 U8301 ( .A1(DRAMRF_ADDRESS[18]), .A2(n8457), .ZN(n7668) );
  AND2_X1 U8302 ( .A1(DRAMRF_ADDRESS[17]), .A2(n8459), .ZN(n7669) );
  AND2_X1 U8303 ( .A1(DRAMRF_ADDRESS[16]), .A2(n8458), .ZN(n7670) );
  AND2_X1 U8304 ( .A1(DRAMRF_ADDRESS[15]), .A2(n8465), .ZN(n7671) );
  AND2_X1 U8305 ( .A1(DRAMRF_ADDRESS[14]), .A2(n8463), .ZN(n7672) );
  AND2_X1 U8306 ( .A1(DRAMRF_ADDRESS[13]), .A2(n8459), .ZN(n7673) );
  AND2_X1 U8307 ( .A1(DRAMRF_ADDRESS[12]), .A2(n8458), .ZN(n7674) );
  AND2_X1 U8308 ( .A1(DRAMRF_ADDRESS[11]), .A2(n8470), .ZN(n7675) );
  AND2_X1 U8309 ( .A1(DRAMRF_ADDRESS[10]), .A2(n8460), .ZN(n7676) );
  AND2_X1 U8310 ( .A1(DRAMRF_ADDRESS[9]), .A2(n8459), .ZN(n7677) );
  AND2_X1 U8311 ( .A1(DRAMRF_ADDRESS[8]), .A2(n8466), .ZN(n7678) );
  AND2_X1 U8312 ( .A1(DRAMRF_ADDRESS[7]), .A2(n8467), .ZN(n7679) );
  AND2_X1 U8313 ( .A1(DRAMRF_ADDRESS[6]), .A2(n8462), .ZN(n7680) );
  AND2_X1 U8314 ( .A1(DRAMRF_ADDRESS[5]), .A2(n8462), .ZN(n7681) );
  AND2_X1 U8315 ( .A1(DRAMRF_ADDRESS[4]), .A2(n8462), .ZN(n7682) );
  AND2_X1 U8316 ( .A1(DRAMRF_ADDRESS[3]), .A2(n8462), .ZN(n7683) );
  AND2_X1 U8317 ( .A1(DRAMRF_ADDRESS[2]), .A2(n8462), .ZN(n7684) );
  INV_X1 U8318 ( .A(n7688), .ZN(n7685) );
  BUF_X1 U8319 ( .A(n8317), .Z(n7686) );
  BUF_X1 U8320 ( .A(n8329), .Z(n7687) );
  BUF_X1 U8321 ( .A(n8869), .Z(n8329) );
  OAI21_X1 U8322 ( .B1(\DP_OP_751_130_6421/n1433 ), .B2(
        \DP_OP_751_130_6421/n1390 ), .A(n7899), .ZN(n7898) );
  AOI21_X1 U8323 ( .B1(\intadd_2/CO ), .B2(n10180), .A(n7891), .ZN(n10177) );
  NOR2_X2 U8324 ( .A1(n10273), .A2(n180), .ZN(i_ADD_RS2[2]) );
  BUF_X1 U8325 ( .A(n8974), .Z(n8261) );
  BUF_X2 U8326 ( .A(n8863), .Z(n8317) );
  AND2_X1 U8327 ( .A1(n8867), .A2(n8866), .ZN(n7688) );
  NAND2_X1 U8328 ( .A1(n9002), .A2(n9016), .ZN(n7689) );
  OR2_X2 U8329 ( .A1(\DP_OP_751_130_6421/n1752 ), .A2(n7727), .ZN(n9002) );
  AND2_X1 U8330 ( .A1(\DP_OP_751_130_6421/n1697 ), .A2(
        \DP_OP_751_130_6421/n1727 ), .ZN(\DP_OP_751_130_6421/n1637 ) );
  INV_X1 U8331 ( .A(n9846), .ZN(n7691) );
  INV_X2 U8332 ( .A(n8444), .ZN(n7692) );
  INV_X1 U8333 ( .A(n8444), .ZN(n8442) );
  XOR2_X1 U8334 ( .A(\DP_OP_751_130_6421/n1697 ), .B(
        \DP_OP_751_130_6421/n1727 ), .Z(\DP_OP_751_130_6421/n1638 ) );
  CLKBUF_X3 U8335 ( .A(n8974), .Z(n8260) );
  XOR2_X1 U8336 ( .A(\DP_OP_751_130_6421/n1004 ), .B(
        \DP_OP_751_130_6421/n1005 ), .Z(n7694) );
  XOR2_X1 U8337 ( .A(\DP_OP_751_130_6421/n1069 ), .B(n7694), .Z(
        \DP_OP_751_130_6421/n970 ) );
  OAI21_X1 U8338 ( .B1(n8159), .B2(n7732), .A(n8841), .ZN(n9782) );
  MUX2_X2 U8339 ( .A(n9678), .B(n8049), .S(\DP_OP_751_130_6421/n1617 ), .Z(
        n8868) );
  AND2_X2 U8340 ( .A1(n7731), .A2(\DataPath/i_PIPLIN_A[26] ), .ZN(n9516) );
  BUF_X1 U8341 ( .A(n8252), .Z(n7695) );
  BUF_X1 U8342 ( .A(\intadd_1/CO ), .Z(n7696) );
  BUF_X1 U8343 ( .A(n10200), .Z(n7697) );
  INV_X2 U8344 ( .A(n9991), .ZN(n10005) );
  BUF_X2 U8345 ( .A(n8868), .Z(n7734) );
  AND2_X2 U8346 ( .A1(n7731), .A2(\DataPath/i_PIPLIN_A[19] ), .ZN(n9711) );
  BUF_X1 U8347 ( .A(n8801), .Z(n7698) );
  AOI21_X1 U8348 ( .B1(\DP_OP_1091J1_126_6973/n5 ), .B2(n8022), .A(n8021), 
        .ZN(n7699) );
  XOR2_X1 U8349 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[27] ), .Z(n7700)
         );
  XOR2_X1 U8350 ( .A(\DP_OP_1091J1_126_6973/n6 ), .B(n7700), .Z(
        \C620/DATA2_27 ) );
  NAND2_X1 U8351 ( .A1(\DP_OP_1091J1_126_6973/n6 ), .A2(n7776), .ZN(n7701) );
  NAND2_X1 U8352 ( .A1(\DP_OP_1091J1_126_6973/n6 ), .A2(
        \DataPath/WRF_CUhw/curr_addr[27] ), .ZN(n7702) );
  NAND2_X1 U8353 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[27] ), .ZN(
        n7703) );
  NAND3_X2 U8354 ( .A1(n7701), .A2(n7702), .A3(n7703), .ZN(
        \DP_OP_1091J1_126_6973/n5 ) );
  BUF_X1 U8355 ( .A(\DP_OP_1091J1_126_6973/n16 ), .Z(n7704) );
  AOI21_X1 U8356 ( .B1(\DP_OP_1091J1_126_6973/n5 ), .B2(n8022), .A(n8021), 
        .ZN(n8016) );
  XNOR2_X1 U8357 ( .A(n7802), .B(n7827), .ZN(n7706) );
  NOR2_X1 U8358 ( .A1(\DP_OP_751_130_6421/n356 ), .A2(
        \DP_OP_751_130_6421/n357 ), .ZN(n7707) );
  XOR2_X1 U8359 ( .A(\DP_OP_751_130_6421/n1696 ), .B(
        \DP_OP_751_130_6421/n1726 ), .Z(\DP_OP_751_130_6421/n1636 ) );
  NAND2_X2 U8360 ( .A1(n8847), .A2(n8846), .ZN(n9129) );
  MUX2_X1 U8361 ( .A(n7710), .B(n7711), .S(n8087), .Z(n7709) );
  OAI21_X2 U8362 ( .B1(n8162), .B2(n7731), .A(n8843), .ZN(n9230) );
  BUF_X1 U8363 ( .A(\DP_OP_751_130_6421/n164 ), .Z(n7892) );
  XNOR2_X1 U8364 ( .A(n7628), .B(n7883), .ZN(\DataPath/ALUhw/i_Q_EXTENDED[60] ) );
  OR2_X1 U8365 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[15] ), .ZN(n7713) );
  AND2_X1 U8366 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[15] ), .ZN(
        n7714) );
  OR2_X1 U8367 ( .A1(n7735), .A2(n7715), .ZN(\intadd_1/n26 ) );
  OR2_X1 U8368 ( .A1(IR[2]), .A2(IRAM_ADDRESS[2]), .ZN(n7715) );
  AOI21_X1 U8369 ( .B1(n8768), .B2(n8767), .A(n8766), .ZN(n7716) );
  AOI22_X1 U8370 ( .A1(n8605), .A2(i_RD1[1]), .B1(n7718), .B2(i_RD1[2]), .ZN(
        n7717) );
  AOI21_X1 U8371 ( .B1(n10091), .B2(n8456), .A(n8584), .ZN(n7718) );
  BUF_X1 U8372 ( .A(\intadd_1/n17 ), .Z(n7719) );
  OR3_X1 U8373 ( .A1(n10270), .A2(n10291), .A3(n8521), .ZN(n8705) );
  BUF_X1 U8374 ( .A(i_S2), .Z(n7738) );
  XNOR2_X1 U8375 ( .A(\DP_OP_751_130_6421/n73 ), .B(n7958), .ZN(
        \DataPath/ALUhw/i_Q_EXTENDED[55] ) );
  INV_X1 U8376 ( .A(n7965), .ZN(\DP_OP_751_130_6421/n66 ) );
  NAND2_X1 U8377 ( .A1(\DP_OP_751_130_6421/n1255 ), .A2(
        \DP_OP_751_130_6421/n1199 ), .ZN(n7930) );
  XOR2_X1 U8378 ( .A(\DP_OP_751_130_6421/n555 ), .B(\DP_OP_751_130_6421/n492 ), 
        .Z(n7722) );
  XOR2_X1 U8379 ( .A(\DP_OP_751_130_6421/n554 ), .B(n7722), .Z(
        \DP_OP_751_130_6421/n456 ) );
  NAND2_X1 U8380 ( .A1(\DP_OP_751_130_6421/n554 ), .A2(
        \DP_OP_751_130_6421/n555 ), .ZN(n7723) );
  NAND2_X1 U8381 ( .A1(\DP_OP_751_130_6421/n554 ), .A2(
        \DP_OP_751_130_6421/n492 ), .ZN(n7724) );
  NAND2_X1 U8382 ( .A1(\DP_OP_751_130_6421/n555 ), .A2(
        \DP_OP_751_130_6421/n492 ), .ZN(n7725) );
  NAND3_X1 U8383 ( .A1(n7723), .A2(n7724), .A3(n7725), .ZN(
        \DP_OP_751_130_6421/n455 ) );
  XNOR2_X1 U8384 ( .A(\DP_OP_751_130_6421/n355 ), .B(n7949), .ZN(n7726) );
  BUF_X1 U8385 ( .A(n9071), .Z(n7727) );
  NAND2_X1 U8386 ( .A1(n10041), .A2(n8280), .ZN(n10216) );
  CLKBUF_X1 U8387 ( .A(n9062), .Z(n7970) );
  CLKBUF_X1 U8388 ( .A(n7880), .Z(n7974) );
  OAI22_X1 U8389 ( .A1(n8858), .A2(n9460), .B1(n8974), .B2(n8300), .ZN(n7910)
         );
  CLKBUF_X1 U8390 ( .A(n8049), .Z(n7937) );
  AND2_X1 U8391 ( .A1(n7824), .A2(\DP_OP_751_130_6421/n1724 ), .ZN(
        \DP_OP_751_130_6421/n1631 ) );
  CLKBUF_X3 U8392 ( .A(n8058), .Z(n8059) );
  AND2_X1 U8393 ( .A1(\DP_OP_751_130_6421/n1693 ), .A2(n7884), .ZN(
        \DP_OP_751_130_6421/n1629 ) );
  OR2_X1 U8394 ( .A1(n8260), .A2(n9904), .ZN(n7728) );
  OR2_X1 U8395 ( .A1(n9026), .A2(n8974), .ZN(n7729) );
  OAI21_X2 U8396 ( .B1(n8143), .B2(n8453), .A(n8870), .ZN(
        \DP_OP_751_130_6421/n1515 ) );
  BUF_X2 U8397 ( .A(n8873), .Z(n8331) );
  OAI21_X2 U8398 ( .B1(n8449), .B2(n9735), .A(n8907), .ZN(n8908) );
  OAI21_X2 U8399 ( .B1(n7767), .B2(n9755), .A(n8900), .ZN(n8901) );
  OAI21_X2 U8400 ( .B1(n8448), .B2(n9780), .A(n8894), .ZN(n8895) );
  OAI21_X2 U8401 ( .B1(n8890), .B2(\DP_OP_751_130_6421/n1311 ), .A(n8889), 
        .ZN(n8891) );
  BUF_X4 U8402 ( .A(n8454), .Z(n7907) );
  BUF_X2 U8403 ( .A(n8878), .Z(n8333) );
  NOR2_X1 U8404 ( .A1(\DP_OP_751_130_6421/n460 ), .A2(
        \DP_OP_751_130_6421/n558 ), .ZN(n7730) );
  INV_X2 U8405 ( .A(n9099), .ZN(n9806) );
  BUF_X1 U8406 ( .A(n8868), .Z(n7733) );
  BUF_X1 U8407 ( .A(n8821), .Z(n7735) );
  BUF_X2 U8408 ( .A(n8821), .Z(n7736) );
  BUF_X2 U8409 ( .A(n8821), .Z(n7737) );
  NAND2_X1 U8410 ( .A1(n7996), .A2(n7998), .ZN(n8821) );
  BUF_X2 U8411 ( .A(n8087), .Z(n7739) );
  AND2_X1 U8412 ( .A1(n7706), .A2(n8014), .ZN(n7814) );
  XNOR2_X1 U8413 ( .A(n7916), .B(n7915), .ZN(\DataPath/ALUhw/i_Q_EXTENDED[59] ) );
  AND2_X1 U8414 ( .A1(n8709), .A2(n8119), .ZN(n7794) );
  NOR2_X1 U8415 ( .A1(n7752), .A2(n8743), .ZN(n7864) );
  NAND2_X1 U8416 ( .A1(n7856), .A2(i_RD2[31]), .ZN(n8685) );
  NOR2_X2 U8417 ( .A1(n10356), .A2(n10355), .ZN(n8353) );
  NOR2_X2 U8418 ( .A1(n10356), .A2(n10355), .ZN(n8354) );
  NOR2_X2 U8419 ( .A1(n10359), .A2(n10357), .ZN(n8351) );
  NOR2_X2 U8420 ( .A1(n10359), .A2(n10354), .ZN(n8348) );
  NOR2_X2 U8421 ( .A1(n10359), .A2(n10357), .ZN(n8350) );
  NOR2_X2 U8422 ( .A1(n10357), .A2(n10356), .ZN(n8356) );
  NOR2_X2 U8423 ( .A1(n10358), .A2(n10342), .ZN(n8344) );
  NOR2_X2 U8424 ( .A1(n10357), .A2(n10356), .ZN(n8357) );
  NOR2_X2 U8425 ( .A1(n10359), .A2(n10358), .ZN(n8358) );
  NOR2_X2 U8426 ( .A1(n10358), .A2(n10342), .ZN(n8343) );
  NOR2_X2 U8427 ( .A1(n10359), .A2(n10354), .ZN(n8349) );
  NOR2_X2 U8428 ( .A1(n10355), .A2(n10342), .ZN(n8342) );
  NOR2_X2 U8429 ( .A1(n10354), .A2(n10341), .ZN(n8340) );
  NOR2_X2 U8430 ( .A1(n10354), .A2(n10342), .ZN(n8345) );
  NOR2_X2 U8431 ( .A1(n10354), .A2(n10342), .ZN(n8346) );
  AOI22_X1 U8432 ( .A1(\DP_OP_751_130_6421/n1171 ), .A2(n7924), .B1(
        \DP_OP_751_130_6421/n1106 ), .B2(\DP_OP_751_130_6421/n1107 ), .ZN(
        n7923) );
  INV_X2 U8433 ( .A(n10886), .ZN(n10885) );
  INV_X2 U8434 ( .A(n10891), .ZN(n10890) );
  INV_X2 U8435 ( .A(n10897), .ZN(n10896) );
  NOR2_X2 U8436 ( .A1(n10273), .A2(n182), .ZN(i_ADD_RS2[0]) );
  INV_X2 U8437 ( .A(n10997), .ZN(n10994) );
  AND2_X2 U8438 ( .A1(n8470), .A2(n11329), .ZN(n11330) );
  INV_X2 U8439 ( .A(n10949), .ZN(n10948) );
  INV_X2 U8440 ( .A(n11037), .ZN(n11035) );
  AND2_X2 U8441 ( .A1(n8470), .A2(n11335), .ZN(n11336) );
  OAI222_X4 U8442 ( .A1(n11345), .A2(n11102), .B1(n11194), .B2(n8271), .C1(
        n11346), .C2(n11640), .ZN(n11066) );
  NAND2_X1 U8443 ( .A1(n8700), .A2(n8684), .ZN(n10072) );
  AND2_X1 U8444 ( .A1(n8494), .A2(n8456), .ZN(n7855) );
  XNOR2_X1 U8445 ( .A(\DP_OP_751_130_6421/n1106 ), .B(
        \DP_OP_751_130_6421/n1107 ), .ZN(n7925) );
  OR2_X1 U8446 ( .A1(\DP_OP_751_130_6421/n1106 ), .A2(
        \DP_OP_751_130_6421/n1107 ), .ZN(n7924) );
  BUF_X1 U8447 ( .A(n8892), .Z(n7760) );
  BUF_X1 U8448 ( .A(n8902), .Z(n7763) );
  BUF_X1 U8449 ( .A(n8909), .Z(n7758) );
  INV_X2 U8450 ( .A(n10999), .ZN(n11003) );
  BUF_X2 U8451 ( .A(n8883), .Z(n7742) );
  BUF_X1 U8452 ( .A(n10011), .Z(n7759) );
  AND2_X2 U8453 ( .A1(n11841), .A2(\DataPath/RF/c_swin[0] ), .ZN(n8183) );
  INV_X1 U8454 ( .A(i_SEL_CMPB), .ZN(n8456) );
  AOI222_X1 U8455 ( .A1(\DataPath/RF/c_swin[2] ), .A2(n11658), .B1(n8281), 
        .B2(n11656), .C1(\DataPath/RF/c_swin[3] ), .C2(n11657), .ZN(n11655) );
  INV_X2 U8456 ( .A(n7767), .ZN(\DP_OP_751_130_6421/n1107 ) );
  BUF_X1 U8457 ( .A(n8896), .Z(n7765) );
  BUF_X2 U8458 ( .A(n8872), .Z(n7743) );
  BUF_X2 U8459 ( .A(n8884), .Z(n7744) );
  BUF_X2 U8460 ( .A(n8879), .Z(n7745) );
  BUF_X1 U8461 ( .A(n9678), .Z(n7942) );
  BUF_X2 U8462 ( .A(n8873), .Z(n7746) );
  INV_X1 U8463 ( .A(n7880), .ZN(n7747) );
  OR2_X1 U8464 ( .A1(n8031), .A2(n7773), .ZN(n8026) );
  NOR2_X1 U8465 ( .A1(i_BUSY_WINDOW), .A2(n7986), .ZN(n8801) );
  NOR2_X1 U8466 ( .A1(n7773), .A2(n8075), .ZN(n8037) );
  OAI21_X1 U8467 ( .B1(n8189), .B2(n7907), .A(n8939), .ZN(
        \DP_OP_751_130_6421/n291 ) );
  OAI21_X2 U8468 ( .B1(n8156), .B2(n7907), .A(n8924), .ZN(
        \DP_OP_751_130_6421/n597 ) );
  CLKBUF_X1 U8469 ( .A(n9151), .Z(n7786) );
  INV_X1 U8470 ( .A(n10245), .ZN(n10099) );
  XNOR2_X1 U8471 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[11] ), .ZN(n7871) );
  OR2_X1 U8472 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[19] ), .ZN(n7945) );
  OR2_X1 U8473 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[12] ), .ZN(n7957) );
  AND2_X1 U8474 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[12] ), .ZN(
        n7956) );
  INV_X1 U8475 ( .A(n9607), .ZN(n9608) );
  OR2_X1 U8476 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[28] ), .ZN(n8022) );
  AND2_X1 U8477 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[22] ), .ZN(
        n8077) );
  OR2_X1 U8478 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[5] ), .ZN(n8045)
         );
  XNOR2_X1 U8479 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[4] ), .ZN(n7886)
         );
  NAND2_X1 U8480 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[29] ), .ZN(
        n8036) );
  AND2_X1 U8481 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[28] ), .ZN(
        n8021) );
  OR2_X1 U8482 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[20] ), .ZN(n8044) );
  XNOR2_X1 U8483 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[16] ), .ZN(n7904) );
  AND2_X2 U8484 ( .A1(n8840), .A2(n8839), .ZN(n8303) );
  XNOR2_X1 U8485 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[14] ), .ZN(n7971) );
  OR2_X1 U8486 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[18] ), .ZN(n7936) );
  XNOR2_X1 U8487 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[12] ), .ZN(n7955) );
  AND2_X1 U8488 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[13] ), .ZN(
        n8082) );
  AND2_X1 U8489 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[18] ), .ZN(
        n7935) );
  AND2_X2 U8490 ( .A1(n7732), .A2(\DataPath/i_PIPLIN_A[23] ), .ZN(n9607) );
  AND2_X1 U8491 ( .A1(\DataPath/i_PIPLIN_A[22] ), .A2(n8442), .ZN(n11723) );
  BUF_X4 U8492 ( .A(n8282), .Z(n8281) );
  NAND2_X1 U8493 ( .A1(n10822), .A2(n8462), .ZN(n8051) );
  AND2_X1 U8494 ( .A1(\DataPath/i_PIPLIN_A[20] ), .A2(n7692), .ZN(n9327) );
  AND2_X2 U8495 ( .A1(\DataPath/i_PIPLIN_A[28] ), .A2(n8442), .ZN(n9689) );
  INV_X1 U8496 ( .A(n8337), .ZN(n7748) );
  INV_X1 U8497 ( .A(n9246), .ZN(n7749) );
  NAND3_X1 U8498 ( .A1(n7987), .A2(n7720), .A3(n8115), .ZN(n7986) );
  NOR2_X1 U8499 ( .A1(IR[27]), .A2(n8090), .ZN(n10059) );
  NAND2_X1 U8500 ( .A1(n7832), .A2(n7837), .ZN(\intadd_2/n33 ) );
  NAND2_X1 U8501 ( .A1(n10152), .A2(n7838), .ZN(n7832) );
  NAND2_X1 U8502 ( .A1(n7928), .A2(n8824), .ZN(n10149) );
  BUF_X1 U8503 ( .A(n8825), .Z(n7928) );
  BUF_X1 U8504 ( .A(n10191), .Z(n7917) );
  AND2_X1 U8505 ( .A1(\intadd_2/n9 ), .A2(n7830), .ZN(n7829) );
  BUF_X1 U8506 ( .A(n10197), .Z(n7894) );
  NAND2_X1 U8507 ( .A1(n7833), .A2(n7836), .ZN(n7830) );
  AND2_X1 U8508 ( .A1(n8164), .A2(n7834), .ZN(n7833) );
  NAND2_X1 U8509 ( .A1(n7835), .A2(n7837), .ZN(n7834) );
  OR2_X1 U8510 ( .A1(n10163), .A2(IRAM_ADDRESS[26]), .ZN(n7919) );
  INV_X1 U8511 ( .A(n7838), .ZN(n7835) );
  INV_X1 U8512 ( .A(n7837), .ZN(n7836) );
  OR2_X1 U8513 ( .A1(n10186), .A2(IRAM_ADDRESS[20]), .ZN(n7838) );
  NAND2_X1 U8514 ( .A1(n10186), .A2(IRAM_ADDRESS[20]), .ZN(n7837) );
  AND2_X1 U8515 ( .A1(n10175), .A2(IRAM_ADDRESS[25]), .ZN(n7891) );
  INV_X1 U8516 ( .A(n10267), .ZN(n7750) );
  INV_X1 U8517 ( .A(n11678), .ZN(n8421) );
  OR2_X1 U8518 ( .A1(n10196), .A2(n8814), .ZN(n7943) );
  AND2_X1 U8519 ( .A1(n8808), .A2(n210), .ZN(n7793) );
  OR2_X1 U8520 ( .A1(\intadd_0/B[4] ), .A2(n7636), .ZN(n10155) );
  INV_X1 U8521 ( .A(n10210), .ZN(n10266) );
  AND2_X1 U8522 ( .A1(n10198), .A2(IRAM_ADDRESS[7]), .ZN(n7922) );
  NAND2_X1 U8523 ( .A1(n7997), .A2(n8000), .ZN(n8803) );
  AOI21_X1 U8524 ( .B1(n8000), .B2(n7999), .A(n11667), .ZN(n7998) );
  XNOR2_X1 U8525 ( .A(\DP_OP_751_130_6421/n66 ), .B(n7921), .ZN(
        \DataPath/ALUhw/i_Q_EXTENDED[58] ) );
  XNOR2_X1 U8526 ( .A(n7892), .B(n7967), .ZN(\DataPath/ALUhw/i_Q_EXTENDED[57] ) );
  AOI21_X1 U8527 ( .B1(n7699), .B2(n8027), .A(n8009), .ZN(n8028) );
  NAND2_X1 U8528 ( .A1(n8790), .A2(n10231), .ZN(n8001) );
  AOI21_X1 U8529 ( .B1(\DP_OP_1091J1_126_6973/n5 ), .B2(n8018), .A(n8017), 
        .ZN(n8019) );
  AND2_X1 U8530 ( .A1(\C620/DATA2_27 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[27])
         );
  AND2_X1 U8531 ( .A1(\C620/DATA2_26 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[26])
         );
  AOI21_X1 U8532 ( .B1(n9386), .B2(n10281), .A(n8013), .ZN(n8003) );
  XNOR2_X1 U8533 ( .A(n7953), .B(\DP_OP_751_130_6421/n165 ), .ZN(
        \DataPath/ALUhw/i_Q_EXTENDED[54] ) );
  INV_X1 U8534 ( .A(n8230), .ZN(n7751) );
  INV_X1 U8535 ( .A(n7846), .ZN(\DP_OP_1091J1_126_6973/n13 ) );
  AOI21_X1 U8536 ( .B1(\DP_OP_1091J1_126_6973/n15 ), .B2(n7849), .A(n7848), 
        .ZN(n7846) );
  INV_X1 U8537 ( .A(n7807), .ZN(\DP_OP_1091J1_126_6973/n15 ) );
  AOI21_X1 U8538 ( .B1(n7864), .B2(n7868), .A(n7863), .ZN(n7861) );
  AND2_X1 U8539 ( .A1(n7869), .A2(n7866), .ZN(n7865) );
  OAI21_X1 U8540 ( .B1(n7639), .B2(n8733), .A(n8736), .ZN(n7868) );
  AOI21_X1 U8541 ( .B1(n7704), .B2(n7653), .A(n7649), .ZN(n7807) );
  INV_X1 U8542 ( .A(n8737), .ZN(n7869) );
  OAI21_X1 U8543 ( .B1(n8740), .B2(n8743), .A(n8742), .ZN(n7863) );
  AND2_X1 U8544 ( .A1(n8741), .A2(n8734), .ZN(n7867) );
  INV_X1 U8545 ( .A(n8743), .ZN(n7866) );
  AND2_X1 U8546 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  XNOR2_X1 U8547 ( .A(\DP_OP_1091J1_126_6973/n17 ), .B(n7904), .ZN(
        \C620/DATA2_16 ) );
  AND2_X1 U8548 ( .A1(n8727), .A2(i_RD1[5]), .ZN(n7876) );
  NAND2_X1 U8549 ( .A1(n8572), .A2(i_RD1[8]), .ZN(n8733) );
  INV_X1 U8550 ( .A(n8741), .ZN(n7752) );
  INV_X2 U8551 ( .A(n11839), .ZN(n7753) );
  XNOR2_X1 U8552 ( .A(\DP_OP_1091J1_126_6973/n19 ), .B(n7971), .ZN(
        \C620/DATA2_14 ) );
  AND2_X1 U8553 ( .A1(n8802), .A2(IR[3]), .ZN(n8006) );
  XNOR2_X1 U8554 ( .A(\DP_OP_751_130_6421/n358 ), .B(\DP_OP_751_130_6421/n456 ), .ZN(n7883) );
  OR2_X1 U8555 ( .A1(i_HAZARD_SIG_CU), .A2(n8483), .ZN(n11667) );
  XNOR2_X1 U8556 ( .A(\DP_OP_751_130_6421/n560 ), .B(\DP_OP_751_130_6421/n561 ), .ZN(n7967) );
  XNOR2_X1 U8557 ( .A(\DP_OP_751_130_6421/n457 ), .B(n7800), .ZN(
        \DP_OP_751_130_6421/n358 ) );
  NAND2_X1 U8558 ( .A1(n7788), .A2(n7787), .ZN(\DP_OP_751_130_6421/n561 ) );
  XNOR2_X1 U8559 ( .A(\DP_OP_1091J1_126_6973/n21 ), .B(n7955), .ZN(
        \C620/DATA2_12 ) );
  NAND2_X1 U8560 ( .A1(\DP_OP_751_130_6421/n661 ), .A2(n7789), .ZN(n7788) );
  XNOR2_X1 U8561 ( .A(\DP_OP_751_130_6421/n662 ), .B(\DP_OP_751_130_6421/n663 ), .ZN(n7958) );
  XNOR2_X1 U8562 ( .A(\DP_OP_751_130_6421/n661 ), .B(n7790), .ZN(
        \DP_OP_751_130_6421/n562 ) );
  XNOR2_X1 U8563 ( .A(\DP_OP_751_130_6421/n664 ), .B(\DP_OP_751_130_6421/n762 ), .ZN(n7953) );
  XNOR2_X1 U8564 ( .A(\DP_OP_1091J1_126_6973/n22 ), .B(n7871), .ZN(
        \C620/DATA2_11 ) );
  NAND2_X1 U8565 ( .A1(\DP_OP_751_130_6421/n664 ), .A2(
        \DP_OP_751_130_6421/n762 ), .ZN(n7950) );
  XNOR2_X1 U8566 ( .A(\DP_OP_751_130_6421/n763 ), .B(n7801), .ZN(
        \DP_OP_751_130_6421/n664 ) );
  XNOR2_X1 U8567 ( .A(\DP_OP_751_130_6421/n865 ), .B(n7909), .ZN(
        \DP_OP_751_130_6421/n766 ) );
  NAND2_X1 U8568 ( .A1(n7931), .A2(n7930), .ZN(\DP_OP_751_130_6421/n1155 ) );
  XNOR2_X1 U8569 ( .A(\DP_OP_751_130_6421/n967 ), .B(n7784), .ZN(
        \DP_OP_751_130_6421/n868 ) );
  NAND2_X1 U8570 ( .A1(n9839), .A2(n9840), .ZN(n7902) );
  BUF_X1 U8571 ( .A(n11158), .Z(n8389) );
  BUF_X1 U8572 ( .A(n10930), .Z(n8368) );
  BUF_X1 U8573 ( .A(n11739), .Z(n8430) );
  BUF_X1 U8574 ( .A(n11742), .Z(n8431) );
  BUF_X1 U8575 ( .A(n11755), .Z(n8433) );
  BUF_X1 U8576 ( .A(n11045), .Z(n8379) );
  BUF_X1 U8577 ( .A(n11821), .Z(n8439) );
  BUF_X1 U8578 ( .A(n10867), .Z(n8361) );
  BUF_X1 U8579 ( .A(n11171), .Z(n8395) );
  INV_X1 U8580 ( .A(n7923), .ZN(\DP_OP_751_130_6421/n1071 ) );
  BUF_X1 U8581 ( .A(n11801), .Z(n8438) );
  AND2_X2 U8582 ( .A1(n8470), .A2(n11377), .ZN(n11404) );
  INV_X2 U8583 ( .A(n11413), .ZN(n8409) );
  BUF_X1 U8584 ( .A(n11771), .Z(n8435) );
  INV_X2 U8585 ( .A(n11200), .ZN(n11199) );
  XNOR2_X1 U8586 ( .A(\DP_OP_751_130_6421/n1171 ), .B(n7925), .ZN(
        \DP_OP_751_130_6421/n1072 ) );
  INV_X2 U8587 ( .A(n10955), .ZN(n8266) );
  INV_X2 U8588 ( .A(n11235), .ZN(n11234) );
  INV_X2 U8589 ( .A(n11105), .ZN(n11104) );
  INV_X2 U8590 ( .A(n11117), .ZN(n11116) );
  INV_X1 U8591 ( .A(n10880), .ZN(n10879) );
  INV_X2 U8592 ( .A(n11351), .ZN(n11350) );
  BUF_X1 U8593 ( .A(n10863), .Z(n8359) );
  INV_X2 U8594 ( .A(n10907), .ZN(n10906) );
  INV_X2 U8595 ( .A(n11101), .ZN(n11100) );
  INV_X2 U8596 ( .A(n11598), .ZN(n8420) );
  AND2_X2 U8597 ( .A1(n8470), .A2(n11362), .ZN(n11364) );
  INV_X2 U8598 ( .A(n11344), .ZN(n11343) );
  AND2_X1 U8599 ( .A1(n8462), .A2(n11802), .ZN(n11800) );
  AND2_X2 U8600 ( .A1(n8462), .A2(n11759), .ZN(n11770) );
  AND2_X2 U8601 ( .A1(n8468), .A2(n11159), .ZN(n11160) );
  AND2_X2 U8602 ( .A1(n8467), .A2(n11154), .ZN(n11155) );
  INV_X2 U8603 ( .A(n11153), .ZN(n11151) );
  INV_X2 U8604 ( .A(n11114), .ZN(n11113) );
  NAND2_X1 U8605 ( .A1(n7898), .A2(n7897), .ZN(\DP_OP_751_130_6421/n1333 ) );
  AND2_X2 U8606 ( .A1(n8467), .A2(n11094), .ZN(n11097) );
  INV_X2 U8607 ( .A(n11065), .ZN(n11064) );
  AND2_X2 U8608 ( .A1(n8467), .A2(n11059), .ZN(n11060) );
  AND2_X2 U8609 ( .A1(n8464), .A2(n10939), .ZN(n10940) );
  AND2_X2 U8610 ( .A1(n8467), .A2(n11056), .ZN(n11057) );
  AND2_X2 U8611 ( .A1(n8467), .A2(n11052), .ZN(n11053) );
  AND2_X2 U8612 ( .A1(n8464), .A2(n10942), .ZN(n10943) );
  AND2_X2 U8613 ( .A1(n8466), .A2(n11049), .ZN(n11050) );
  AND2_X2 U8614 ( .A1(n8466), .A2(n11048), .ZN(n11046) );
  AND2_X2 U8615 ( .A1(n8465), .A2(n11043), .ZN(n11041) );
  INV_X2 U8616 ( .A(n10952), .ZN(n7754) );
  AND2_X2 U8617 ( .A1(n8464), .A2(n10973), .ZN(n10977) );
  INV_X2 U8618 ( .A(n10987), .ZN(n7755) );
  AND2_X2 U8619 ( .A1(n8469), .A2(n10864), .ZN(n10862) );
  INV_X2 U8620 ( .A(n10874), .ZN(n10872) );
  AND2_X2 U8621 ( .A1(n8469), .A2(n11307), .ZN(n11308) );
  INV_X2 U8622 ( .A(n11271), .ZN(n11269) );
  INV_X2 U8623 ( .A(n11225), .ZN(n11224) );
  INV_X2 U8624 ( .A(n10914), .ZN(n10913) );
  INV_X2 U8625 ( .A(n10902), .ZN(n10901) );
  AND2_X2 U8626 ( .A1(n8468), .A2(n11165), .ZN(n11166) );
  INV_X2 U8627 ( .A(n11193), .ZN(n11190) );
  XNOR2_X1 U8628 ( .A(\DP_OP_751_130_6421/n1273 ), .B(n7791), .ZN(
        \DP_OP_751_130_6421/n1174 ) );
  AND2_X2 U8629 ( .A1(n8468), .A2(n11168), .ZN(n11169) );
  AND2_X2 U8630 ( .A1(n8468), .A2(n11173), .ZN(n11186) );
  XNOR2_X1 U8631 ( .A(\DP_OP_1091J1_126_6973/n29 ), .B(n7886), .ZN(
        \C620/DATA2_4 ) );
  AND2_X1 U8632 ( .A1(n10271), .A2(i_RF2), .ZN(n7839) );
  NAND2_X1 U8633 ( .A1(n7896), .A2(n7895), .ZN(\DP_OP_751_130_6421/n1431 ) );
  OR2_X1 U8634 ( .A1(\DP_OP_751_130_6421/n1682 ), .A2(
        \DP_OP_751_130_6421/n1683 ), .ZN(\DP_OP_751_130_6421/n151 ) );
  XNOR2_X1 U8635 ( .A(\DP_OP_751_130_6421/n902 ), .B(n8061), .ZN(n7784) );
  INV_X1 U8636 ( .A(n10295), .ZN(n10934) );
  OR4_X1 U8637 ( .A1(n9553), .A2(n9552), .A3(n9551), .A4(n9550), .ZN(n10018)
         );
  NAND2_X1 U8638 ( .A1(\DP_OP_751_130_6421/n1490 ), .A2(
        \DP_OP_751_130_6421/n1531 ), .ZN(n7895) );
  OAI21_X1 U8639 ( .B1(\DP_OP_751_130_6421/n1490 ), .B2(
        \DP_OP_751_130_6421/n1531 ), .A(\DP_OP_751_130_6421/n1530 ), .ZN(n7896) );
  BUF_X1 U8640 ( .A(n11073), .Z(n7779) );
  XNOR2_X1 U8641 ( .A(\DP_OP_751_130_6421/n596 ), .B(\DP_OP_751_130_6421/n597 ), .ZN(n7790) );
  INV_X1 U8642 ( .A(n8183), .ZN(n8437) );
  BUF_X1 U8643 ( .A(n11110), .Z(n7778) );
  NOR2_X1 U8644 ( .A1(n11735), .A2(n7748), .ZN(n7841) );
  NAND2_X1 U8645 ( .A1(\DP_OP_751_130_6421/n596 ), .A2(
        \DP_OP_751_130_6421/n597 ), .ZN(n7787) );
  OR2_X1 U8646 ( .A1(\DP_OP_751_130_6421/n596 ), .A2(\DP_OP_751_130_6421/n597 ), .ZN(n7789) );
  BUF_X1 U8647 ( .A(n11084), .Z(n7780) );
  BUF_X1 U8648 ( .A(n11081), .Z(n7781) );
  AND2_X1 U8649 ( .A1(\DP_OP_751_130_6421/n1696 ), .A2(
        \DP_OP_751_130_6421/n1726 ), .ZN(\DP_OP_751_130_6421/n1635 ) );
  XNOR2_X1 U8650 ( .A(\DP_OP_751_130_6421/n290 ), .B(\DP_OP_751_130_6421/n291 ), .ZN(n7949) );
  BUF_X2 U8651 ( .A(n11419), .Z(n8410) );
  INV_X4 U8652 ( .A(n11419), .ZN(n7756) );
  OR2_X1 U8653 ( .A1(\DP_OP_751_130_6421/n290 ), .A2(\DP_OP_751_130_6421/n291 ), .ZN(n7948) );
  AND2_X1 U8654 ( .A1(\DP_OP_751_130_6421/n290 ), .A2(
        \DP_OP_751_130_6421/n291 ), .ZN(n7947) );
  INV_X1 U8655 ( .A(n7934), .ZN(n7933) );
  AND2_X1 U8656 ( .A1(\DP_OP_751_130_6421/n1730 ), .A2(
        \DP_OP_751_130_6421/n1700 ), .ZN(\DP_OP_751_130_6421/n1643 ) );
  XNOR2_X1 U8657 ( .A(\DP_OP_751_130_6421/n698 ), .B(n7782), .ZN(n7801) );
  XNOR2_X1 U8658 ( .A(\DP_OP_751_130_6421/n392 ), .B(\DP_OP_751_130_6421/n393 ), .ZN(n7800) );
  INV_X1 U8659 ( .A(n8456), .ZN(n7856) );
  XNOR2_X1 U8660 ( .A(\DP_OP_751_130_6421/n800 ), .B(n8062), .ZN(n7909) );
  AND2_X1 U8661 ( .A1(n7847), .A2(n7653), .ZN(n7809) );
  OR2_X1 U8662 ( .A1(n11735), .A2(n7748), .ZN(n8004) );
  INV_X1 U8663 ( .A(n7885), .ZN(n7884) );
  INV_X1 U8664 ( .A(n10101), .ZN(i_ADD_WS1[2]) );
  BUF_X2 U8665 ( .A(n11836), .Z(n7757) );
  NOR2_X2 U8666 ( .A1(n835), .A2(n8054), .ZN(n11419) );
  NOR2_X1 U8667 ( .A1(n8010), .A2(n8023), .ZN(n8008) );
  BUF_X2 U8668 ( .A(n11237), .Z(n7761) );
  BUF_X2 U8669 ( .A(n11119), .Z(n7762) );
  AND2_X1 U8670 ( .A1(n8042), .A2(n7849), .ZN(n7847) );
  AND3_X1 U8671 ( .A1(n8239), .A2(n8240), .A3(n7981), .ZN(n7980) );
  BUF_X2 U8672 ( .A(n10289), .Z(n7764) );
  INV_X2 U8673 ( .A(n8449), .ZN(\DP_OP_751_130_6421/n1005 ) );
  INV_X1 U8674 ( .A(n7740), .ZN(n9017) );
  OR2_X1 U8675 ( .A1(n8974), .A2(n9826), .ZN(n7908) );
  NOR2_X1 U8676 ( .A1(n8026), .A2(n8011), .ZN(n8010) );
  AND2_X1 U8677 ( .A1(n8024), .A2(n8025), .ZN(n8023) );
  INV_X1 U8678 ( .A(n8032), .ZN(n8015) );
  AND2_X1 U8679 ( .A1(n8033), .A2(n8022), .ZN(n8018) );
  NOR2_X1 U8680 ( .A1(n8046), .A2(n8043), .ZN(n8042) );
  INV_X1 U8681 ( .A(\DataPath/ALUhw/MULT/mux_out[0][0] ), .ZN(n7766) );
  INV_X1 U8682 ( .A(n8864), .ZN(n7768) );
  BUF_X2 U8683 ( .A(n10290), .Z(n7769) );
  INV_X1 U8684 ( .A(n7860), .ZN(n9069) );
  BUF_X1 U8685 ( .A(\DP_OP_751_130_6421/n699 ), .Z(n7782) );
  OR2_X1 U8686 ( .A1(\DP_OP_751_130_6421/n1719 ), .A2(n9802), .ZN(n8049) );
  NAND2_X2 U8687 ( .A1(n8886), .A2(n8885), .ZN(\DP_OP_751_130_6421/n1209 ) );
  AND2_X1 U8688 ( .A1(n8036), .A2(n8031), .ZN(n8027) );
  AND2_X1 U8689 ( .A1(n7992), .A2(n7991), .ZN(n7990) );
  OR2_X1 U8690 ( .A1(n8858), .A2(n8300), .ZN(n7870) );
  AND2_X1 U8691 ( .A1(n7945), .A2(n7936), .ZN(n7849) );
  INV_X1 U8692 ( .A(n8116), .ZN(\DP_OP_751_130_6421/n1719 ) );
  INV_X1 U8693 ( .A(n7798), .ZN(n7772) );
  OAI21_X1 U8694 ( .B1(n8075), .B2(n8036), .A(n8038), .ZN(n8035) );
  INV_X1 U8695 ( .A(n8021), .ZN(n8011) );
  INV_X1 U8696 ( .A(\DP_OP_751_130_6421/n1515 ), .ZN(n8446) );
  BUF_X1 U8697 ( .A(n9794), .Z(n7799) );
  INV_X1 U8698 ( .A(n10231), .ZN(n7999) );
  BUF_X1 U8699 ( .A(n9121), .Z(n7792) );
  INV_X2 U8700 ( .A(n9966), .ZN(n9972) );
  INV_X1 U8701 ( .A(n8044), .ZN(n8043) );
  AND2_X1 U8702 ( .A1(n8090), .A2(n7720), .ZN(n7991) );
  INV_X1 U8703 ( .A(n8036), .ZN(n8034) );
  INV_X1 U8704 ( .A(n8074), .ZN(n8031) );
  INV_X2 U8705 ( .A(n11457), .ZN(n11458) );
  NAND2_X2 U8706 ( .A1(n8460), .A2(n11478), .ZN(n11510) );
  INV_X2 U8707 ( .A(n11461), .ZN(n11462) );
  INV_X1 U8708 ( .A(n9516), .ZN(n9277) );
  INV_X2 U8709 ( .A(n11469), .ZN(n11470) );
  NAND2_X2 U8710 ( .A1(n8460), .A2(n11473), .ZN(n11474) );
  INV_X1 U8711 ( .A(n8039), .ZN(n7773) );
  INV_X2 U8712 ( .A(n11465), .ZN(n11466) );
  AND2_X1 U8713 ( .A1(n7994), .A2(n8478), .ZN(n7993) );
  AND2_X2 U8714 ( .A1(n8857), .A2(n8856), .ZN(n9910) );
  AND2_X2 U8715 ( .A1(n8855), .A2(n8854), .ZN(n8311) );
  NAND2_X2 U8716 ( .A1(n8460), .A2(n11453), .ZN(n11454) );
  AND2_X2 U8717 ( .A1(n8853), .A2(n8852), .ZN(n8308) );
  AND2_X2 U8718 ( .A1(n8851), .A2(n8850), .ZN(n8305) );
  AND2_X1 U8719 ( .A1(DRAMRF_READY), .A2(n8292), .ZN(n8291) );
  INV_X1 U8720 ( .A(n9250), .ZN(n7774) );
  INV_X1 U8721 ( .A(n9826), .ZN(n7775) );
  BUF_X4 U8722 ( .A(\DP_OP_1091J1_126_6973/n72 ), .Z(n7776) );
  NAND2_X2 U8723 ( .A1(n470), .A2(n471), .ZN(n10822) );
  BUF_X1 U8724 ( .A(IR[27]), .Z(n7969) );
  OR2_X1 U8725 ( .A1(n8117), .A2(\DataPath/RF/c_win[3] ), .ZN(n8247) );
  INV_X2 U8726 ( .A(i_DATAMEM_RM), .ZN(n11616) );
  INV_X2 U8727 ( .A(DRAMRF_READY), .ZN(n11840) );
  BUF_X1 U8728 ( .A(n10926), .Z(n8365) );
  BUF_X1 U8729 ( .A(n10917), .Z(n8362) );
  BUF_X1 U8730 ( .A(n11738), .Z(n8429) );
  OAI211_X2 U8731 ( .C1(n10249), .C2(n182), .A(n10248), .B(n10247), .ZN(
        i_ADD_WS1[0]) );
  INV_X1 U8732 ( .A(n10018), .ZN(n7777) );
  AOI22_X2 U8733 ( .A1(n11419), .A2(n11282), .B1(n11489), .B2(n7756), .ZN(
        n11384) );
  AOI22_X2 U8734 ( .A1(n11419), .A2(n11277), .B1(n11484), .B2(n7756), .ZN(
        n11380) );
  NOR2_X2 U8735 ( .A1(n10359), .A2(n10358), .ZN(n8113) );
  NOR2_X2 U8736 ( .A1(DATA_SIZE[0]), .A2(n381), .ZN(n10800) );
  NOR2_X2 U8737 ( .A1(n10341), .A2(n10355), .ZN(n8112) );
  NOR2_X2 U8738 ( .A1(n10356), .A2(n10358), .ZN(n8111) );
  NOR3_X2 U8739 ( .A1(i_ADD_WB[3]), .A2(n8102), .A3(n8192), .ZN(n10932) );
  NOR3_X2 U8740 ( .A1(n8168), .A2(n10703), .A3(n10694), .ZN(n10737) );
  NOR2_X2 U8741 ( .A1(n10341), .A2(n10355), .ZN(n8110) );
  NOR3_X2 U8742 ( .A1(n508), .A2(n10703), .A3(n10694), .ZN(n10736) );
  BUF_X2 U8743 ( .A(n11405), .Z(n8407) );
  BUF_X2 U8744 ( .A(n11365), .Z(n8406) );
  OAI22_X2 U8745 ( .A1(n11415), .A2(n11758), .B1(n7756), .B2(n11757), .ZN(
        n11316) );
  OAI22_X2 U8746 ( .A1(n11415), .A2(n11773), .B1(n7756), .B2(n11772), .ZN(
        n11318) );
  XNOR2_X1 U8747 ( .A(\DP_OP_751_130_6421/n494 ), .B(\DP_OP_751_130_6421/n495 ), .ZN(n7893) );
  OAI21_X1 U8748 ( .B1(n8154), .B2(n7907), .A(n8917), .ZN(
        \DP_OP_751_130_6421/n699 ) );
  BUF_X1 U8749 ( .A(n11044), .Z(n8378) );
  BUF_X1 U8750 ( .A(n10945), .Z(n8372) );
  BUF_X1 U8751 ( .A(n11157), .Z(n8388) );
  NOR4_X2 U8752 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n9144), .ZN(n9788)
         );
  AOI22_X2 U8753 ( .A1(n7762), .A2(n11281), .B1(n11488), .B2(n11102), .ZN(
        n11078) );
  AOI22_X2 U8754 ( .A1(n7761), .A2(n11283), .B1(n11490), .B2(n11211), .ZN(
        n11229) );
  AOI22_X2 U8755 ( .A1(n7762), .A2(n11290), .B1(n11497), .B2(n11102), .ZN(
        n11085) );
  NOR4_X4 U8756 ( .A1(n9483), .A2(n9482), .A3(n9481), .A4(n9480), .ZN(n9879)
         );
  NAND2_X2 U8757 ( .A1(n8960), .A2(n8959), .ZN(n9850) );
  OAI22_X2 U8758 ( .A1(n7756), .A2(n11276), .B1(n11483), .B2(n8410), .ZN(
        n11379) );
  XNOR2_X1 U8759 ( .A(\DP_OP_751_130_6421/n1208 ), .B(
        \DP_OP_751_130_6421/n1209 ), .ZN(n7791) );
  NOR2_X2 U8760 ( .A1(n10355), .A2(n10342), .ZN(n8109) );
  NOR2_X2 U8761 ( .A1(n10354), .A2(n10341), .ZN(n8108) );
  NOR3_X4 U8762 ( .A1(i_ADD_WB[4]), .A2(i_ADD_WB[3]), .A3(n8192), .ZN(n11476)
         );
  OAI22_X2 U8763 ( .A1(n11640), .A2(n11758), .B1(n11211), .B2(n11757), .ZN(
        n11162) );
  NOR2_X2 U8764 ( .A1(n10356), .A2(n10358), .ZN(n8089) );
  AOI22_X2 U8765 ( .A1(n8410), .A2(n11301), .B1(n11508), .B2(n7756), .ZN(
        n11402) );
  AOI22_X2 U8766 ( .A1(n8410), .A2(n11284), .B1(n11491), .B2(n7756), .ZN(
        n11386) );
  AOI221_X2 U8767 ( .B1(n507), .B2(n10693), .C1(n10692), .C2(n10693), .A(
        n11616), .ZN(n10738) );
  NOR2_X2 U8768 ( .A1(n10760), .A2(n10761), .ZN(n10779) );
  NOR2_X2 U8769 ( .A1(n9589), .A2(n11733), .ZN(n9683) );
  AOI211_X2 U8770 ( .C1(n9687), .C2(n9639), .A(n9638), .B(n9637), .ZN(n10008)
         );
  OAI22_X2 U8771 ( .A1(n8450), .A2(n11773), .B1(n8436), .B2(n11772), .ZN(
        n11802) );
  INV_X1 U8772 ( .A(n8183), .ZN(n8436) );
  NOR2_X2 U8773 ( .A1(n8338), .A2(n11646), .ZN(n10815) );
  OAI22_X2 U8774 ( .A1(n11415), .A2(n11322), .B1(n7756), .B2(n11321), .ZN(
        n11323) );
  NOR2_X2 U8775 ( .A1(i_DATAMEM_RM), .A2(n10703), .ZN(n10790) );
  OAI22_X2 U8776 ( .A1(n8271), .A2(n11737), .B1(n11102), .B2(n11736), .ZN(
        n11039) );
  OAI21_X2 U8777 ( .B1(n8187), .B2(n7907), .A(n8932), .ZN(
        \DP_OP_751_130_6421/n393 ) );
  AOI22_X2 U8778 ( .A1(n8410), .A2(n11275), .B1(n11482), .B2(n7756), .ZN(
        n11423) );
  AOI22_X2 U8779 ( .A1(n8410), .A2(n11274), .B1(n11481), .B2(n7756), .ZN(
        n11422) );
  XNOR2_X1 U8780 ( .A(n7783), .B(n7770), .ZN(n7824) );
  OAI22_X1 U8781 ( .A1(n7689), .A2(n9277), .B1(n7637), .B2(n9846), .ZN(n7783)
         );
  XNOR2_X1 U8782 ( .A(\DataPath/ALUhw/MULT/mux_out[1][19] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1703 ) );
  BUF_X1 U8783 ( .A(n9002), .Z(n7785) );
  XNOR2_X1 U8784 ( .A(\DataPath/ALUhw/MULT/mux_out[1][16] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1706 ) );
  AND2_X1 U8785 ( .A1(\DP_OP_751_130_6421/n356 ), .A2(
        \DP_OP_751_130_6421/n357 ), .ZN(n7819) );
  XNOR2_X1 U8786 ( .A(\DataPath/ALUhw/MULT/mux_out[1][24] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1698 ) );
  XNOR2_X1 U8787 ( .A(\DataPath/ALUhw/MULT/mux_out[1][17] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1705 ) );
  NOR2_X1 U8788 ( .A1(n8807), .A2(n7793), .ZN(n10197) );
  NAND3_X1 U8789 ( .A1(n8708), .A2(n8710), .A3(n7794), .ZN(n10105) );
  XNOR2_X1 U8790 ( .A(n7795), .B(\DP_OP_751_130_6421/n1700 ), .ZN(
        \DP_OP_751_130_6421/n1644 ) );
  XNOR2_X1 U8791 ( .A(\DataPath/ALUhw/MULT/mux_out[1][22] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1700 ) );
  INV_X1 U8792 ( .A(\DP_OP_751_130_6421/n1730 ), .ZN(n7795) );
  XNOR2_X1 U8793 ( .A(\DataPath/ALUhw/MULT/mux_out[1][25] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1697 ) );
  XNOR2_X1 U8794 ( .A(\DataPath/ALUhw/MULT/mux_out[1][26] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1696 ) );
  AOI21_X1 U8795 ( .B1(n7798), .B2(n9130), .A(n7797), .ZN(n7796) );
  NOR2_X1 U8796 ( .A1(\DP_OP_751_130_6421/n1515 ), .A2(
        \DP_OP_751_130_6421/n1617 ), .ZN(n7797) );
  INV_X1 U8797 ( .A(n8445), .ZN(n7798) );
  XNOR2_X1 U8798 ( .A(\DataPath/ALUhw/MULT/mux_out[2][27] ), .B(n7772), .ZN(
        \DP_OP_751_130_6421/n1593 ) );
  INV_X1 U8799 ( .A(n7739), .ZN(n8454) );
  INV_X1 U8800 ( .A(n7721), .ZN(n8495) );
  XNOR2_X1 U8801 ( .A(\DataPath/ALUhw/MULT/mux_out[2][28] ), .B(n7772), .ZN(
        \DP_OP_751_130_6421/n1592 ) );
  XNOR2_X1 U8802 ( .A(n7803), .B(\DP_OP_751_130_6421/n352 ), .ZN(n7802) );
  XNOR2_X1 U8803 ( .A(\DP_OP_751_130_6421/n353 ), .B(n7654), .ZN(n7803) );
  NAND2_X1 U8804 ( .A1(n10281), .A2(n8337), .ZN(n7804) );
  AND2_X1 U8805 ( .A1(\DP_OP_751_130_6421/n61 ), .A2(n7805), .ZN(n8005) );
  INV_X1 U8806 ( .A(\DP_OP_751_130_6421/n60 ), .ZN(n7805) );
  INV_X1 U8807 ( .A(n7806), .ZN(\DP_OP_1091J1_126_6973/n10 ) );
  AOI21_X1 U8808 ( .B1(\DP_OP_1091J1_126_6973/n16 ), .B2(n7809), .A(n7808), 
        .ZN(n7806) );
  NOR2_X1 U8809 ( .A1(n7810), .A2(n7706), .ZN(n7812) );
  NAND2_X1 U8810 ( .A1(\DP_OP_751_130_6421/n61 ), .A2(n7841), .ZN(n7810) );
  NAND4_X1 U8811 ( .A1(n7815), .A2(n7842), .A3(n7813), .A4(n7811), .ZN(n6985)
         );
  NAND2_X1 U8812 ( .A1(n7850), .A2(n7812), .ZN(n7811) );
  NAND2_X1 U8813 ( .A1(n7814), .A2(n10281), .ZN(n7813) );
  AOI21_X1 U8814 ( .B1(\DP_OP_751_130_6421/n62 ), .B2(n7817), .A(n7816), .ZN(
        n7815) );
  NOR2_X1 U8815 ( .A1(n7840), .A2(n11735), .ZN(n7816) );
  OAI21_X1 U8816 ( .B1(n7821), .B2(n7707), .A(n7818), .ZN(
        \DP_OP_751_130_6421/n62 ) );
  AOI21_X1 U8817 ( .B1(n7826), .B2(n7820), .A(n7819), .ZN(n7818) );
  INV_X1 U8818 ( .A(n7881), .ZN(n7820) );
  NAND2_X1 U8819 ( .A1(n7882), .A2(\DP_OP_751_130_6421/n64 ), .ZN(n7821) );
  OAI21_X1 U8820 ( .B1(n7822), .B2(n7706), .A(n7655), .ZN(n7851) );
  INV_X1 U8821 ( .A(\DP_OP_751_130_6421/n354 ), .ZN(n7823) );
  NAND2_X1 U8822 ( .A1(n7726), .A2(\DP_OP_751_130_6421/n354 ), .ZN(
        \DP_OP_751_130_6421/n61 ) );
  XNOR2_X1 U8823 ( .A(n7824), .B(n7877), .ZN(\DP_OP_751_130_6421/n1632 ) );
  AOI21_X1 U8824 ( .B1(n7966), .B2(\DP_OP_751_130_6421/n164 ), .A(n7963), .ZN(
        n7965) );
  NAND2_X1 U8825 ( .A1(n7825), .A2(\DP_OP_751_130_6421/n71 ), .ZN(
        \DP_OP_751_130_6421/n164 ) );
  NAND2_X1 U8826 ( .A1(\DP_OP_751_130_6421/n72 ), .A2(n8070), .ZN(n7825) );
  OR2_X1 U8827 ( .A1(\DP_OP_751_130_6421/n562 ), .A2(\DP_OP_751_130_6421/n660 ), .ZN(n8070) );
  NAND2_X1 U8828 ( .A1(n7960), .A2(n7959), .ZN(\DP_OP_751_130_6421/n72 ) );
  OR2_X1 U8829 ( .A1(\DP_OP_751_130_6421/n356 ), .A2(\DP_OP_751_130_6421/n357 ), .ZN(n7826) );
  AOI21_X1 U8830 ( .B1(\DP_OP_751_130_6421/n355 ), .B2(n7948), .A(n7947), .ZN(
        n7827) );
  NOR2_X1 U8831 ( .A1(n7828), .A2(n7857), .ZN(\DP_OP_751_130_6421/n1633 ) );
  XNOR2_X1 U8832 ( .A(n7858), .B(n8059), .ZN(n7857) );
  INV_X1 U8833 ( .A(\DP_OP_751_130_6421/n1725 ), .ZN(n7828) );
  NAND2_X1 U8834 ( .A1(n10152), .A2(n7833), .ZN(n7831) );
  NAND2_X1 U8835 ( .A1(n7831), .A2(n7829), .ZN(\intadd_2/CO ) );
  INV_X1 U8836 ( .A(n10270), .ZN(n10272) );
  OR2_X2 U8837 ( .A1(n8819), .A2(n10245), .ZN(n10270) );
  NAND2_X1 U8838 ( .A1(n10272), .A2(n7839), .ZN(n10273) );
  INV_X1 U8839 ( .A(n9371), .ZN(n7840) );
  INV_X1 U8840 ( .A(n7851), .ZN(n7842) );
  NAND2_X1 U8841 ( .A1(n7914), .A2(n7916), .ZN(n7913) );
  OAI21_X1 U8842 ( .B1(n7965), .B2(n7730), .A(n7920), .ZN(n7916) );
  NAND2_X1 U8843 ( .A1(n7844), .A2(n7843), .ZN(n6987) );
  AOI21_X1 U8844 ( .B1(n7859), .B2(n10279), .A(n7902), .ZN(n7843) );
  NAND2_X1 U8845 ( .A1(\DataPath/ALUhw/i_Q_EXTENDED[61] ), .A2(n7845), .ZN(
        n7844) );
  NOR2_X1 U8846 ( .A1(n10032), .A2(n7748), .ZN(n7845) );
  INV_X1 U8847 ( .A(\DP_OP_751_130_6421/n62 ), .ZN(n7850) );
  NAND2_X1 U8848 ( .A1(n7853), .A2(n7852), .ZN(n8688) );
  NAND2_X1 U8849 ( .A1(n8495), .A2(n7855), .ZN(n7852) );
  INV_X1 U8850 ( .A(n7854), .ZN(n7853) );
  OAI21_X1 U8851 ( .B1(n8684), .B2(n7856), .A(n8685), .ZN(n7854) );
  NAND2_X2 U8852 ( .A1(n8495), .A2(n8494), .ZN(n8700) );
  INV_X1 U8853 ( .A(n8688), .ZN(n8686) );
  XNOR2_X1 U8854 ( .A(\DP_OP_751_130_6421/n1725 ), .B(n7857), .ZN(
        \DP_OP_751_130_6421/n1634 ) );
  OAI22_X1 U8855 ( .A1(n9527), .A2(n7637), .B1(n7689), .B2(n9846), .ZN(n7858)
         );
  CLKBUF_X1 U8856 ( .A(n7727), .Z(n7860) );
  INV_X1 U8857 ( .A(n8864), .ZN(n8320) );
  NAND2_X1 U8858 ( .A1(n9002), .A2(n9016), .ZN(n8864) );
  NAND2_X1 U8859 ( .A1(n7862), .A2(n7861), .ZN(n8748) );
  NAND3_X1 U8860 ( .A1(n8735), .A2(n7865), .A3(n7867), .ZN(n7862) );
  NAND2_X1 U8861 ( .A1(n7870), .A2(n7908), .ZN(n7938) );
  INV_X1 U8862 ( .A(n7872), .ZN(\DP_OP_1091J1_126_6973/n20 ) );
  AOI21_X1 U8863 ( .B1(\DP_OP_1091J1_126_6973/n21 ), .B2(n7957), .A(n7956), 
        .ZN(n7872) );
  OAI21_X1 U8864 ( .B1(n7875), .B2(n7874), .A(n7873), .ZN(
        \DP_OP_1091J1_126_6973/n21 ) );
  NAND2_X1 U8865 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[11] ), .ZN(
        n7873) );
  NOR2_X1 U8866 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[11] ), .ZN(
        n7874) );
  INV_X1 U8867 ( .A(\DP_OP_1091J1_126_6973/n22 ), .ZN(n7875) );
  AOI21_X1 U8868 ( .B1(n8729), .B2(n8728), .A(n7876), .ZN(n8732) );
  INV_X1 U8869 ( .A(\DP_OP_751_130_6421/n1724 ), .ZN(n7877) );
  NAND2_X1 U8870 ( .A1(n7879), .A2(n7878), .ZN(n7027) );
  NAND2_X1 U8871 ( .A1(n10267), .A2(i_RD1[29]), .ZN(n7878) );
  NAND2_X1 U8872 ( .A1(n10161), .A2(n7750), .ZN(n7879) );
  XNOR2_X1 U8873 ( .A(\DP_OP_751_130_6421/n1693 ), .B(n7885), .ZN(
        \DP_OP_751_130_6421/n1630 ) );
  XNOR2_X1 U8874 ( .A(n7938), .B(n7747), .ZN(n7885) );
  XNOR2_X1 U8875 ( .A(\DataPath/ALUhw/MULT/mux_out[1][29] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1693 ) );
  NAND2_X1 U8876 ( .A1(\DP_OP_751_130_6421/n358 ), .A2(
        \DP_OP_751_130_6421/n456 ), .ZN(n7881) );
  OR2_X1 U8877 ( .A1(\DP_OP_751_130_6421/n358 ), .A2(\DP_OP_751_130_6421/n456 ), .ZN(n7882) );
  INV_X1 U8878 ( .A(n7887), .ZN(\DP_OP_1091J1_126_6973/n27 ) );
  AOI21_X1 U8879 ( .B1(\DP_OP_1091J1_126_6973/n28 ), .B2(n8045), .A(n7650), 
        .ZN(n7887) );
  NAND2_X1 U8880 ( .A1(n7889), .A2(n7888), .ZN(\DP_OP_1091J1_126_6973/n28 ) );
  NAND2_X1 U8881 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[4] ), .ZN(
        n7888) );
  NAND2_X1 U8882 ( .A1(\DP_OP_1091J1_126_6973/n29 ), .A2(n7890), .ZN(n7889) );
  OR2_X1 U8883 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[4] ), .ZN(n7890)
         );
  XNOR2_X1 U8884 ( .A(\DP_OP_751_130_6421/n843 ), .B(\DP_OP_751_130_6421/n789 ), .ZN(n7964) );
  XNOR2_X1 U8885 ( .A(n7964), .B(\DP_OP_751_130_6421/n842 ), .ZN(
        \DP_OP_751_130_6421/n744 ) );
  OAI21_X2 U8886 ( .B1(n8142), .B2(n8453), .A(n8865), .ZN(
        \DP_OP_751_130_6421/n1617 ) );
  XNOR2_X1 U8887 ( .A(n7901), .B(n7899), .ZN(\DP_OP_751_130_6421/n1334 ) );
  XNOR2_X1 U8888 ( .A(n7900), .B(\DP_OP_751_130_6421/n1530 ), .ZN(n7899) );
  XNOR2_X1 U8889 ( .A(\DP_OP_751_130_6421/n1490 ), .B(
        \DP_OP_751_130_6421/n1531 ), .ZN(n7900) );
  XNOR2_X1 U8890 ( .A(\DP_OP_751_130_6421/n1433 ), .B(
        \DP_OP_751_130_6421/n1390 ), .ZN(n7901) );
  XNOR2_X1 U8891 ( .A(\DataPath/ALUhw/MULT/mux_out[1][23] ), .B(n7770), .ZN(
        \DP_OP_751_130_6421/n1699 ) );
  XNOR2_X1 U8892 ( .A(\DP_OP_751_130_6421/n1626 ), .B(n7903), .ZN(
        \DP_OP_751_130_6421/n1528 ) );
  OAI21_X1 U8893 ( .B1(n7712), .B2(n7906), .A(n7905), .ZN(
        \DP_OP_1091J1_126_6973/n16 ) );
  NAND2_X1 U8894 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[16] ), .ZN(
        n7905) );
  NOR2_X1 U8895 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[16] ), .ZN(
        n7906) );
  INV_X1 U8896 ( .A(n7739), .ZN(n8453) );
  OAI21_X1 U8897 ( .B1(n7740), .B2(n9826), .A(n7729), .ZN(n7944) );
  XNOR2_X1 U8898 ( .A(n7910), .B(n7880), .ZN(\DP_OP_751_130_6421/n1724 ) );
  NAND2_X1 U8899 ( .A1(n7911), .A2(n8227), .ZN(n8226) );
  NAND2_X1 U8900 ( .A1(n7716), .A2(n7751), .ZN(n7911) );
  NOR2_X1 U8901 ( .A1(n10216), .A2(n8244), .ZN(n10224) );
  NAND2_X1 U8902 ( .A1(n172), .A2(IR[27]), .ZN(n8244) );
  NOR2_X1 U8903 ( .A1(IR[31]), .A2(n8280), .ZN(n10226) );
  NAND2_X1 U8904 ( .A1(n7913), .A2(n7912), .ZN(\DP_OP_751_130_6421/n64 ) );
  NAND2_X1 U8905 ( .A1(\DP_OP_751_130_6421/n458 ), .A2(
        \DP_OP_751_130_6421/n459 ), .ZN(n7912) );
  OAI22_X1 U8906 ( .A1(n10261), .A2(n7962), .B1(n10260), .B2(n8050), .ZN(
        n10157) );
  XNOR2_X1 U8907 ( .A(n10265), .B(n7918), .ZN(n10269) );
  NAND2_X1 U8908 ( .A1(n8050), .A2(n7919), .ZN(n10158) );
  NAND2_X1 U8909 ( .A1(\DP_OP_751_130_6421/n460 ), .A2(
        \DP_OP_751_130_6421/n558 ), .ZN(n7920) );
  INV_X1 U8910 ( .A(n8454), .ZN(n8455) );
  NOR2_X1 U8911 ( .A1(n10200), .A2(n7922), .ZN(n8807) );
  XNOR2_X1 U8912 ( .A(n7926), .B(n8060), .ZN(\DP_OP_751_130_6421/n1735 ) );
  OAI22_X1 U8913 ( .A1(n7740), .A2(n9250), .B1(n8260), .B2(n10005), .ZN(n7926)
         );
  XNOR2_X1 U8914 ( .A(n7927), .B(n8060), .ZN(\DP_OP_751_130_6421/n1734 ) );
  OAI22_X1 U8915 ( .A1(n7740), .A2(n10005), .B1(n8260), .B2(n9246), .ZN(n7927)
         );
  XNOR2_X1 U8916 ( .A(n7929), .B(n7880), .ZN(\DP_OP_751_130_6421/n1729 ) );
  XNOR2_X1 U8917 ( .A(n7932), .B(\DP_OP_751_130_6421/n1254 ), .ZN(
        \DP_OP_751_130_6421/n1156 ) );
  XNOR2_X1 U8918 ( .A(\DP_OP_751_130_6421/n1255 ), .B(
        \DP_OP_751_130_6421/n1199 ), .ZN(n7932) );
  XNOR2_X1 U8919 ( .A(\DP_OP_751_130_6421/n1692 ), .B(n7934), .ZN(
        \DP_OP_751_130_6421/n1628 ) );
  XNOR2_X1 U8920 ( .A(n7944), .B(n7747), .ZN(n7934) );
  NOR2_X1 U8921 ( .A1(n10261), .A2(n7962), .ZN(n10264) );
  BUF_X1 U8922 ( .A(\intadd_1/n25 ), .Z(n7939) );
  BUF_X2 U8923 ( .A(n7907), .Z(n7940) );
  XNOR2_X1 U8924 ( .A(n7941), .B(n8060), .ZN(\DP_OP_751_130_6421/n1732 ) );
  OAI22_X1 U8925 ( .A1(n7740), .A2(n7693), .B1(n8260), .B2(n8301), .ZN(n7941)
         );
  AOI21_X1 U8926 ( .B1(n10197), .B2(n10195), .A(n7943), .ZN(n8816) );
  XNOR2_X1 U8927 ( .A(n7946), .B(n7880), .ZN(\DP_OP_751_130_6421/n1731 ) );
  OAI21_X1 U8928 ( .B1(n7740), .B2(n8301), .A(n7728), .ZN(n7946) );
  NAND2_X1 U8929 ( .A1(n7951), .A2(n7950), .ZN(\DP_OP_751_130_6421/n73 ) );
  NAND2_X1 U8930 ( .A1(\DP_OP_751_130_6421/n165 ), .A2(n7952), .ZN(n7951) );
  OR2_X1 U8931 ( .A1(\DP_OP_751_130_6421/n664 ), .A2(\DP_OP_751_130_6421/n762 ), .ZN(n7952) );
  BUF_X1 U8932 ( .A(n10226), .Z(n7954) );
  AOI21_X1 U8933 ( .B1(\DP_OP_1091J1_126_6973/n20 ), .B2(n8041), .A(n8082), 
        .ZN(n8040) );
  NAND2_X1 U8934 ( .A1(\DP_OP_751_130_6421/n662 ), .A2(
        \DP_OP_751_130_6421/n663 ), .ZN(n7959) );
  NAND2_X1 U8935 ( .A1(\DP_OP_751_130_6421/n73 ), .A2(n7961), .ZN(n7960) );
  OR2_X1 U8936 ( .A1(\DP_OP_751_130_6421/n662 ), .A2(\DP_OP_751_130_6421/n663 ), .ZN(n7961) );
  AND2_X1 U8937 ( .A1(\DP_OP_751_130_6421/n560 ), .A2(
        \DP_OP_751_130_6421/n561 ), .ZN(n7963) );
  OR2_X1 U8938 ( .A1(\DP_OP_751_130_6421/n560 ), .A2(\DP_OP_751_130_6421/n561 ), .ZN(n7966) );
  XNOR2_X1 U8939 ( .A(n7968), .B(n8060), .ZN(\DP_OP_751_130_6421/n1733 ) );
  OAI22_X1 U8940 ( .A1(n7693), .A2(n8260), .B1(n7740), .B2(n9246), .ZN(n7968)
         );
  OAI21_X1 U8941 ( .B1(n8040), .B2(n7973), .A(n7972), .ZN(
        \DP_OP_1091J1_126_6973/n18 ) );
  NAND2_X1 U8942 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[14] ), .ZN(
        n7972) );
  NOR2_X1 U8943 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[14] ), .ZN(
        n7973) );
  XNOR2_X1 U8944 ( .A(n7976), .B(n8076), .ZN(\DP_OP_1091J1_126_6973/n37 ) );
  OAI211_X1 U8945 ( .C1(n7982), .C2(n7980), .A(n7978), .B(n7977), .ZN(n7976)
         );
  NAND2_X1 U8946 ( .A1(n11647), .A2(n7993), .ZN(n7977) );
  NAND2_X1 U8947 ( .A1(n7979), .A2(n8291), .ZN(n7978) );
  NAND2_X1 U8948 ( .A1(n11647), .A2(n8478), .ZN(n7979) );
  NAND2_X1 U8949 ( .A1(n8801), .A2(n10304), .ZN(n11647) );
  OR2_X1 U8950 ( .A1(n8243), .A2(n8241), .ZN(n7981) );
  NAND2_X1 U8951 ( .A1(n11633), .A2(n10801), .ZN(n8239) );
  NAND2_X1 U8952 ( .A1(n7988), .A2(n8290), .ZN(n11633) );
  NOR2_X1 U8953 ( .A1(n7985), .A2(n7983), .ZN(n10304) );
  NAND2_X1 U8954 ( .A1(n7984), .A2(n8235), .ZN(n7983) );
  INV_X1 U8955 ( .A(n8248), .ZN(n7984) );
  OAI21_X1 U8956 ( .B1(n7648), .B2(n835), .A(n8247), .ZN(n7985) );
  AND4_X1 U8957 ( .A1(n8280), .A2(IR[27]), .A3(n8167), .A4(n172), .ZN(n7987)
         );
  NOR2_X1 U8958 ( .A1(n7989), .A2(n10307), .ZN(n7988) );
  NOR2_X1 U8959 ( .A1(n8285), .A2(n166), .ZN(n7992) );
  AND2_X1 U8960 ( .A1(\DP_OP_1091J1_126_6973/n72 ), .A2(DRAMRF_READY), .ZN(
        n7994) );
  NAND2_X1 U8961 ( .A1(n7995), .A2(n8000), .ZN(n7996) );
  INV_X1 U8962 ( .A(n8791), .ZN(n7995) );
  NAND2_X1 U8963 ( .A1(n8791), .A2(n10231), .ZN(n7997) );
  XNOR2_X1 U8964 ( .A(n8016), .B(n7652), .ZN(\C620/DATA2_29 ) );
  NAND2_X1 U8965 ( .A1(n8015), .A2(n7699), .ZN(n8020) );
  OAI21_X1 U8966 ( .B1(n8002), .B2(n8004), .A(n8003), .ZN(n6986) );
  XNOR2_X1 U8967 ( .A(\DP_OP_751_130_6421/n62 ), .B(n8005), .ZN(n8002) );
  NAND2_X1 U8968 ( .A1(n8803), .A2(n8006), .ZN(\intadd_1/B[2] ) );
  OAI21_X1 U8969 ( .B1(n8007), .B2(n8012), .A(n8008), .ZN(n8009) );
  INV_X1 U8970 ( .A(\DP_OP_1091J1_126_6973/n5 ), .ZN(n8007) );
  OAI22_X1 U8971 ( .A1(n9404), .A2(n11730), .B1(n11734), .B2(n527), .ZN(n8013)
         );
  NOR2_X1 U8972 ( .A1(\DP_OP_751_130_6421/n61 ), .A2(n7748), .ZN(n8014) );
  NAND2_X1 U8973 ( .A1(n8020), .A2(n8019), .ZN(\C620/DATA2_31 ) );
  NOR2_X1 U8974 ( .A1(n8028), .A2(n8051), .ZN(n8258) );
  NAND2_X1 U8975 ( .A1(n8036), .A2(n8074), .ZN(n8024) );
  OAI21_X1 U8976 ( .B1(n8034), .B2(n8039), .A(n8031), .ZN(n8025) );
  OR2_X1 U8977 ( .A1(n7651), .A2(n8035), .ZN(n8032) );
  AND2_X1 U8978 ( .A1(n8037), .A2(n7651), .ZN(n8033) );
  AND2_X1 U8979 ( .A1(n8171), .A2(\C620/DATA2_31 ), .ZN(n8257) );
  NAND2_X1 U8980 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[30] ), .ZN(
        n8038) );
  OR2_X1 U8981 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[29] ), .ZN(n8039) );
  INV_X1 U8982 ( .A(n8040), .ZN(\DP_OP_1091J1_126_6973/n19 ) );
  OR2_X1 U8983 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[13] ), .ZN(n8041) );
  BUF_X1 U8984 ( .A(n10159), .Z(n8050) );
  OAI21_X1 U8985 ( .B1(n8141), .B2(i_S2), .A(n8861), .ZN(n9071) );
  AND2_X1 U8986 ( .A1(\C620/DATA2_29 ), .A2(n8171), .ZN(n8259) );
  AND2_X1 U8987 ( .A1(\C620/DATA2_29 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[29])
         );
  INV_X1 U8988 ( .A(n10309), .ZN(n8052) );
  INV_X1 U8989 ( .A(n8243), .ZN(n8053) );
  OAI211_X1 U8990 ( .C1(n8243), .C2(n8241), .A(n8240), .B(n8239), .ZN(n8054)
         );
  OR2_X1 U8991 ( .A1(n8242), .A2(n8484), .ZN(n8240) );
  INV_X1 U8992 ( .A(n8054), .ZN(n11841) );
  INV_X1 U8993 ( .A(\DP_OP_751_130_6421/n106 ), .ZN(\DP_OP_751_130_6421/n104 )
         );
  INV_X1 U8994 ( .A(\DP_OP_751_130_6421/n114 ), .ZN(\DP_OP_751_130_6421/n112 )
         );
  INV_X1 U8995 ( .A(\DP_OP_751_130_6421/n122 ), .ZN(\DP_OP_751_130_6421/n120 )
         );
  INV_X1 U8996 ( .A(\DP_OP_751_130_6421/n124 ), .ZN(\DP_OP_751_130_6421/n123 )
         );
  INV_X1 U8997 ( .A(\DP_OP_751_130_6421/n128 ), .ZN(\DP_OP_751_130_6421/n126 )
         );
  INV_X1 U8998 ( .A(\DP_OP_751_130_6421/n136 ), .ZN(\DP_OP_751_130_6421/n134 )
         );
  INV_X1 U8999 ( .A(\DP_OP_751_130_6421/n144 ), .ZN(\DP_OP_751_130_6421/n142 )
         );
  INV_X1 U9000 ( .A(\DP_OP_751_130_6421/n152 ), .ZN(\DP_OP_751_130_6421/n150 )
         );
  INV_X1 U9001 ( .A(\DP_OP_751_130_6421/n163 ), .ZN(\DP_OP_751_130_6421/n161 )
         );
  INV_X1 U9002 ( .A(\DP_OP_751_130_6421/n74 ), .ZN(\DP_OP_751_130_6421/n165 )
         );
  INV_X1 U9003 ( .A(\DP_OP_751_130_6421/n80 ), .ZN(\DP_OP_751_130_6421/n169 )
         );
  INV_X1 U9004 ( .A(\DP_OP_751_130_6421/n88 ), .ZN(\DP_OP_751_130_6421/n171 )
         );
  INV_X1 U9005 ( .A(\DP_OP_751_130_6421/n96 ), .ZN(\DP_OP_751_130_6421/n173 )
         );
  INV_X1 U9006 ( .A(\DataPath/ALUhw/MULT/mux_out[0][31] ), .ZN(
        \DP_OP_751_130_6421/n1756 ) );
  INV_X1 U9007 ( .A(\DP_OP_751_130_6421/n108 ), .ZN(\DP_OP_751_130_6421/n176 )
         );
  INV_X1 U9008 ( .A(\DataPath/ALUhw/MULT/mux_out[0][26] ), .ZN(
        \DP_OP_751_130_6421/n1761 ) );
  INV_X1 U9009 ( .A(\DataPath/ALUhw/MULT/mux_out[0][25] ), .ZN(
        \DP_OP_751_130_6421/n1762 ) );
  INV_X1 U9010 ( .A(\DataPath/ALUhw/MULT/mux_out[0][24] ), .ZN(
        \DP_OP_751_130_6421/n1763 ) );
  INV_X1 U9011 ( .A(\DataPath/ALUhw/MULT/mux_out[0][16] ), .ZN(
        \DP_OP_751_130_6421/n1771 ) );
  INV_X1 U9012 ( .A(\DataPath/ALUhw/MULT/mux_out[0][12] ), .ZN(
        \DP_OP_751_130_6421/n1775 ) );
  INV_X1 U9013 ( .A(\DataPath/ALUhw/MULT/mux_out[0][11] ), .ZN(
        \DP_OP_751_130_6421/n1776 ) );
  INV_X1 U9014 ( .A(\DataPath/ALUhw/MULT/mux_out[0][10] ), .ZN(
        \DP_OP_751_130_6421/n1777 ) );
  INV_X1 U9015 ( .A(\DataPath/ALUhw/MULT/mux_out[0][9] ), .ZN(
        \DP_OP_751_130_6421/n1778 ) );
  INV_X1 U9016 ( .A(\DataPath/ALUhw/MULT/mux_out[0][8] ), .ZN(
        \DP_OP_751_130_6421/n1779 ) );
  INV_X1 U9017 ( .A(\DataPath/ALUhw/MULT/mux_out[0][7] ), .ZN(
        \DP_OP_751_130_6421/n1780 ) );
  INV_X1 U9018 ( .A(\DataPath/ALUhw/MULT/mux_out[0][6] ), .ZN(
        \DP_OP_751_130_6421/n1781 ) );
  INV_X1 U9019 ( .A(\DP_OP_751_130_6421/n130 ), .ZN(\DP_OP_751_130_6421/n181 )
         );
  INV_X1 U9020 ( .A(\DP_OP_751_130_6421/n138 ), .ZN(\DP_OP_751_130_6421/n183 )
         );
  INV_X1 U9021 ( .A(\DP_OP_751_130_6421/n146 ), .ZN(\DP_OP_751_130_6421/n185 )
         );
  INV_X1 U9022 ( .A(\DP_OP_751_130_6421/n86 ), .ZN(\DP_OP_751_130_6421/n84 )
         );
  INV_X1 U9023 ( .A(\DP_OP_751_130_6421/n94 ), .ZN(\DP_OP_751_130_6421/n92 )
         );
  INV_X1 U9024 ( .A(\DP_OP_751_130_6421/n99 ), .ZN(\DP_OP_751_130_6421/n98 )
         );
  AOI21_X1 U9025 ( .B1(n8065), .B2(\DP_OP_751_130_6421/n129 ), .A(
        \DP_OP_751_130_6421/n126 ), .ZN(\DP_OP_751_130_6421/n124 ) );
  OAI21_X1 U9026 ( .B1(\DP_OP_751_130_6421/n100 ), .B2(
        \DP_OP_751_130_6421/n102 ), .A(\DP_OP_751_130_6421/n101 ), .ZN(
        \DP_OP_751_130_6421/n99 ) );
  OAI21_X1 U9027 ( .B1(\DP_OP_751_130_6421/n130 ), .B2(
        \DP_OP_751_130_6421/n132 ), .A(\DP_OP_751_130_6421/n131 ), .ZN(
        \DP_OP_751_130_6421/n129 ) );
  OAI21_X1 U9028 ( .B1(\DP_OP_751_130_6421/n116 ), .B2(
        \DP_OP_751_130_6421/n118 ), .A(\DP_OP_751_130_6421/n117 ), .ZN(
        \DP_OP_751_130_6421/n115 ) );
  OAI21_X1 U9029 ( .B1(\DP_OP_751_130_6421/n80 ), .B2(\DP_OP_751_130_6421/n82 ), .A(\DP_OP_751_130_6421/n81 ), .ZN(\DP_OP_751_130_6421/n79 ) );
  XOR2_X1 U9030 ( .A(\DP_OP_751_130_6421/n6 ), .B(n7642), .Z(
        \DataPath/ALUhw/i_Q_EXTENDED[52] ) );
  XNOR2_X1 U9031 ( .A(\DP_OP_751_130_6421/n87 ), .B(\DP_OP_751_130_6421/n7 ), 
        .ZN(\DataPath/ALUhw/i_Q_EXTENDED[51] ) );
  XOR2_X1 U9032 ( .A(\DP_OP_751_130_6421/n18 ), .B(\DP_OP_751_130_6421/n132 ), 
        .Z(\DataPath/ALUhw/i_Q_EXTENDED[40] ) );
  AOI21_X1 U9033 ( .B1(n8064), .B2(\DP_OP_751_130_6421/n79 ), .A(n7708), .ZN(
        \DP_OP_751_130_6421/n74 ) );
  XNOR2_X1 U9034 ( .A(\DP_OP_751_130_6421/n5 ), .B(n7641), .ZN(
        \DataPath/ALUhw/i_Q_EXTENDED[53] ) );
  XNOR2_X1 U9035 ( .A(\DP_OP_751_130_6421/n17 ), .B(\DP_OP_751_130_6421/n129 ), 
        .ZN(\DataPath/ALUhw/i_Q_EXTENDED[41] ) );
  NAND2_X1 U9036 ( .A1(\DP_OP_751_130_6421/n1753 ), .A2(n7747), .ZN(
        \DP_OP_751_130_6421/n163 ) );
  OAI21_X1 U9037 ( .B1(\DP_OP_751_130_6421/n108 ), .B2(
        \DP_OP_751_130_6421/n110 ), .A(\DP_OP_751_130_6421/n109 ), .ZN(
        \DP_OP_751_130_6421/n107 ) );
  XOR2_X1 U9038 ( .A(\DP_OP_751_130_6421/n13 ), .B(\DP_OP_751_130_6421/n110 ), 
        .Z(\DataPath/ALUhw/i_Q_EXTENDED[45] ) );
  AND2_X1 U9039 ( .A1(n8063), .A2(\DP_OP_751_130_6421/n163 ), .ZN(
        \DataPath/ALUhw/i_Q_EXTENDED[32] ) );
  OR2_X1 U9040 ( .A1(\DP_OP_751_130_6421/n1753 ), .A2(n7747), .ZN(n8063) );
  OR2_X1 U9041 ( .A1(\DP_OP_751_130_6421/n764 ), .A2(\DP_OP_751_130_6421/n765 ), .ZN(n8064) );
  OR2_X1 U9042 ( .A1(\DP_OP_751_130_6421/n1072 ), .A2(
        \DP_OP_751_130_6421/n1170 ), .ZN(n8066) );
  OR2_X1 U9043 ( .A1(\DP_OP_751_130_6421/n1174 ), .A2(
        \DP_OP_751_130_6421/n1272 ), .ZN(n8067) );
  OR2_X1 U9044 ( .A1(\DP_OP_751_130_6421/n1276 ), .A2(
        \DP_OP_751_130_6421/n1374 ), .ZN(n8071) );
  OR2_X1 U9045 ( .A1(\DP_OP_751_130_6421/n1376 ), .A2(
        \DP_OP_751_130_6421/n1377 ), .ZN(n8065) );
  OR2_X1 U9046 ( .A1(\DP_OP_751_130_6421/n1478 ), .A2(
        \DP_OP_751_130_6421/n1479 ), .ZN(n8072) );
  NOR2_X1 U9047 ( .A1(\DP_OP_751_130_6421/n1684 ), .A2(
        \DP_OP_751_130_6421/n1685 ), .ZN(\DP_OP_751_130_6421/n154 ) );
  OR2_X1 U9048 ( .A1(\DP_OP_751_130_6421/n1580 ), .A2(
        \DP_OP_751_130_6421/n1581 ), .ZN(n8073) );
  AOI21_X1 U9049 ( .B1(n8067), .B2(\DP_OP_751_130_6421/n115 ), .A(
        \DP_OP_751_130_6421/n112 ), .ZN(\DP_OP_751_130_6421/n110 ) );
  AOI21_X1 U9050 ( .B1(n8066), .B2(\DP_OP_751_130_6421/n107 ), .A(
        \DP_OP_751_130_6421/n104 ), .ZN(\DP_OP_751_130_6421/n102 ) );
  OAI21_X1 U9051 ( .B1(\DP_OP_751_130_6421/n98 ), .B2(\DP_OP_751_130_6421/n96 ), .A(\DP_OP_751_130_6421/n97 ), .ZN(\DP_OP_751_130_6421/n95 ) );
  OR2_X1 U9052 ( .A1(\DP_OP_751_130_6421/n968 ), .A2(\DP_OP_751_130_6421/n969 ), .ZN(n8069) );
  AOI21_X1 U9053 ( .B1(\DP_OP_751_130_6421/n95 ), .B2(n8069), .A(
        \DP_OP_751_130_6421/n92 ), .ZN(\DP_OP_751_130_6421/n90 ) );
  OAI21_X1 U9054 ( .B1(\DP_OP_751_130_6421/n90 ), .B2(\DP_OP_751_130_6421/n88 ), .A(\DP_OP_751_130_6421/n89 ), .ZN(\DP_OP_751_130_6421/n87 ) );
  OR2_X1 U9055 ( .A1(\DP_OP_751_130_6421/n866 ), .A2(\DP_OP_751_130_6421/n867 ), .ZN(n8068) );
  AOI21_X1 U9056 ( .B1(\DP_OP_751_130_6421/n87 ), .B2(n8068), .A(
        \DP_OP_751_130_6421/n84 ), .ZN(\DP_OP_751_130_6421/n82 ) );
  BUF_X1 U9057 ( .A(\DP_OP_751_130_6421/n801 ), .Z(n8062) );
  BUF_X1 U9058 ( .A(\DP_OP_751_130_6421/n903 ), .Z(n8061) );
  BUF_X1 U9059 ( .A(\DP_OP_751_130_6421/n1311 ), .Z(n8055) );
  INV_X1 U9060 ( .A(\DP_OP_1091J1_126_6973/n72 ), .ZN(n8076) );
  XNOR2_X1 U9061 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[30] ), .ZN(n8074) );
  NAND2_X1 U9062 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[21] ), .ZN(
        n8078) );
  NAND2_X1 U9063 ( .A1(n7776), .A2(\DataPath/WRF_CUhw/curr_addr[20] ), .ZN(
        n8079) );
  XOR2_X1 U9064 ( .A(\DP_OP_1091J1_126_6973/n18 ), .B(n8080), .Z(
        \C620/DATA2_15 ) );
  XOR2_X1 U9065 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[15] ), .Z(n8080)
         );
  XOR2_X1 U9066 ( .A(\DP_OP_1091J1_126_6973/n28 ), .B(n8081), .Z(
        \C620/DATA2_5 ) );
  XOR2_X1 U9067 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[5] ), .Z(n8081)
         );
  XOR2_X1 U9068 ( .A(\DP_OP_1091J1_126_6973/n20 ), .B(n8083), .Z(
        \C620/DATA2_13 ) );
  XOR2_X1 U9069 ( .A(n7776), .B(\DataPath/WRF_CUhw/curr_addr[13] ), .Z(n8083)
         );
  AND2_X1 U9070 ( .A1(n8052), .A2(n8478), .ZN(n10295) );
  BUF_X1 U9071 ( .A(n11196), .Z(n8397) );
  INV_X1 U9072 ( .A(n11358), .ZN(n11357) );
  BUF_X1 U9073 ( .A(n11000), .Z(n8375) );
  BUF_X1 U9074 ( .A(n11309), .Z(n8399) );
  BUF_X1 U9075 ( .A(n11306), .Z(n8398) );
  BUF_X1 U9076 ( .A(n11312), .Z(n8400) );
  BUF_X1 U9077 ( .A(n11320), .Z(n8402) );
  BUF_X1 U9078 ( .A(n11315), .Z(n8401) );
  BUF_X1 U9079 ( .A(n11325), .Z(n8403) );
  BUF_X1 U9080 ( .A(n10946), .Z(n8373) );
  BUF_X1 U9081 ( .A(n10927), .Z(n8366) );
  BUF_X1 U9082 ( .A(n10918), .Z(n8363) );
  NAND2_X2 U9083 ( .A1(n11841), .A2(n8281), .ZN(n10999) );
  NOR2_X1 U9084 ( .A1(RST), .A2(n8360), .ZN(n10867) );
  NOR2_X1 U9085 ( .A1(RST), .A2(n8434), .ZN(n11755) );
  NOR2_X1 U9086 ( .A1(RST), .A2(n8432), .ZN(n11742) );
  NOR2_X1 U9087 ( .A1(RST), .A2(n8440), .ZN(n11821) );
  NOR2_X1 U9088 ( .A1(RST), .A2(n8429), .ZN(n11739) );
  OR2_X1 U9089 ( .A1(n11840), .A2(n10801), .ZN(n11662) );
  BUF_X1 U9090 ( .A(n10292), .Z(n8294) );
  NOR2_X2 U9091 ( .A1(n10266), .A2(n8812), .ZN(n10267) );
  NOR2_X1 U9092 ( .A1(n11667), .A2(n8138), .ZN(n10292) );
  INV_X1 U9093 ( .A(n11667), .ZN(n8802) );
  INV_X1 U9094 ( .A(n8246), .ZN(n2872) );
  BUF_X1 U9095 ( .A(n8295), .Z(n8296) );
  INV_X1 U9096 ( .A(n11210), .ZN(n11209) );
  INV_X1 U9097 ( .A(n11222), .ZN(n11221) );
  BUF_X1 U9098 ( .A(n11051), .Z(n8381) );
  BUF_X1 U9099 ( .A(n11161), .Z(n8390) );
  BUF_X1 U9100 ( .A(n11187), .Z(n8396) );
  BUF_X1 U9101 ( .A(n11054), .Z(n8382) );
  BUF_X1 U9102 ( .A(n11058), .Z(n8383) );
  BUF_X1 U9103 ( .A(n11047), .Z(n8380) );
  BUF_X1 U9104 ( .A(n11170), .Z(n8393) );
  BUF_X1 U9105 ( .A(n11042), .Z(n8377) );
  BUF_X1 U9106 ( .A(n10978), .Z(n8374) );
  BUF_X1 U9107 ( .A(n11098), .Z(n8386) );
  BUF_X1 U9108 ( .A(n11061), .Z(n8384) );
  BUF_X1 U9109 ( .A(n11167), .Z(n8392) );
  BUF_X1 U9110 ( .A(n11069), .Z(n8385) );
  BUF_X1 U9111 ( .A(n10923), .Z(n8364) );
  BUF_X1 U9112 ( .A(n11164), .Z(n8391) );
  INV_X1 U9113 ( .A(n11372), .ZN(n11371) );
  BUF_X1 U9114 ( .A(n11040), .Z(n8376) );
  BUF_X1 U9115 ( .A(n10938), .Z(n8369) );
  INV_X1 U9116 ( .A(n7754), .ZN(n8262) );
  INV_X1 U9117 ( .A(n7755), .ZN(n8267) );
  BUF_X1 U9118 ( .A(n11331), .Z(n8404) );
  BUF_X1 U9119 ( .A(n11337), .Z(n8405) );
  INV_X1 U9120 ( .A(n8266), .ZN(n8264) );
  AND2_X1 U9121 ( .A1(n8468), .A2(n11305), .ZN(n11303) );
  INV_X1 U9122 ( .A(n11830), .ZN(n10300) );
  AND2_X1 U9123 ( .A1(n8469), .A2(n11310), .ZN(n11311) );
  AND2_X1 U9124 ( .A1(n8470), .A2(n11318), .ZN(n11319) );
  AND2_X1 U9125 ( .A1(n8469), .A2(n11316), .ZN(n11314) );
  INV_X1 U9126 ( .A(n8420), .ZN(n8418) );
  AND2_X1 U9127 ( .A1(n8470), .A2(n11323), .ZN(n11324) );
  AND2_X1 U9128 ( .A1(n8462), .A2(n11797), .ZN(n11752) );
  AND2_X1 U9129 ( .A1(n8463), .A2(n11763), .ZN(n11820) );
  AND2_X1 U9130 ( .A1(n8465), .A2(n11769), .ZN(n11803) );
  AND2_X1 U9131 ( .A1(n8463), .A2(n11782), .ZN(n11812) );
  AND2_X1 U9132 ( .A1(n8463), .A2(n11762), .ZN(n11819) );
  AND2_X1 U9133 ( .A1(n8463), .A2(n11764), .ZN(n11823) );
  INV_X1 U9134 ( .A(n11723), .ZN(n8428) );
  INV_X1 U9135 ( .A(n406), .ZN(n8447) );
  OR2_X1 U9136 ( .A1(n7736), .A2(n183), .ZN(\intadd_0/B[4] ) );
  NOR2_X1 U9137 ( .A1(n10273), .A2(n181), .ZN(i_ADD_RS2[1]) );
  AND2_X1 U9138 ( .A1(n8782), .A2(n8689), .ZN(n8779) );
  AND3_X2 U9139 ( .A1(n8788), .A2(n10059), .A3(n10041), .ZN(n10245) );
  AND2_X1 U9140 ( .A1(IR[31]), .A2(n166), .ZN(n8788) );
  INV_X1 U9141 ( .A(i_BUSY_WINDOW), .ZN(n8243) );
  BUF_X1 U9142 ( .A(n11156), .Z(n8387) );
  BUF_X1 U9143 ( .A(n10941), .Z(n8370) );
  BUF_X1 U9144 ( .A(n10944), .Z(n8371) );
  AND2_X1 U9145 ( .A1(n8464), .A2(n10936), .ZN(n10937) );
  AND2_X1 U9146 ( .A1(n8467), .A2(n11066), .ZN(n11068) );
  AND2_X1 U9147 ( .A1(n8470), .A2(n10921), .ZN(n10922) );
  AND2_X1 U9148 ( .A1(n8468), .A2(n11162), .ZN(n11163) );
  AND2_X1 U9149 ( .A1(n8464), .A2(n11039), .ZN(n11038) );
  INV_X1 U9150 ( .A(n8266), .ZN(n8265) );
  NOR2_X1 U9151 ( .A1(RST), .A2(n8394), .ZN(n11171) );
  BUF_X1 U9152 ( .A(n11836), .Z(n8441) );
  NOR2_X1 U9153 ( .A1(RST), .A2(n11835), .ZN(n11836) );
  NOR2_X1 U9154 ( .A1(RST), .A2(n8378), .ZN(n11045) );
  INV_X2 U9155 ( .A(n11119), .ZN(n11102) );
  AND2_X1 U9156 ( .A1(n8462), .A2(n10962), .ZN(n11014) );
  AND2_X1 U9157 ( .A1(n8463), .A2(n10981), .ZN(n11006) );
  AND2_X1 U9158 ( .A1(n8463), .A2(n10956), .ZN(n11004) );
  AND2_X1 U9159 ( .A1(n8464), .A2(n10960), .ZN(n11011) );
  AND2_X1 U9160 ( .A1(n8464), .A2(n10989), .ZN(n11010) );
  AND2_X1 U9161 ( .A1(n8463), .A2(n10957), .ZN(n11007) );
  AND2_X1 U9162 ( .A1(n8464), .A2(n10959), .ZN(n11009) );
  NOR2_X1 U9163 ( .A1(RST), .A2(n8388), .ZN(n11158) );
  INV_X2 U9164 ( .A(n11237), .ZN(n11211) );
  AND2_X1 U9165 ( .A1(n8464), .A2(n10958), .ZN(n11008) );
  AND2_X1 U9166 ( .A1(n8466), .A2(n10972), .ZN(n11028) );
  AND2_X1 U9167 ( .A1(n8462), .A2(n10995), .ZN(n11036) );
  AND2_X1 U9168 ( .A1(n8461), .A2(n10966), .ZN(n11020) );
  AND2_X1 U9169 ( .A1(n8460), .A2(n10970), .ZN(n11025) );
  INV_X1 U9170 ( .A(n11838), .ZN(n11679) );
  NOR2_X1 U9171 ( .A1(RST), .A2(n11802), .ZN(n11801) );
  AND2_X1 U9172 ( .A1(n8457), .A2(n11767), .ZN(n11794) );
  AND2_X1 U9173 ( .A1(n8463), .A2(n11792), .ZN(n11750) );
  AND2_X1 U9174 ( .A1(n8464), .A2(n11768), .ZN(n11796) );
  AND2_X1 U9175 ( .A1(n8462), .A2(n11790), .ZN(n11749) );
  AND2_X1 U9176 ( .A1(n8462), .A2(n11765), .ZN(n11791) );
  AND2_X1 U9177 ( .A1(n8458), .A2(n11798), .ZN(n11753) );
  AND2_X1 U9178 ( .A1(n8460), .A2(n11799), .ZN(n11754) );
  OAI22_X1 U9179 ( .A1(n8450), .A2(n11333), .B1(n8436), .B2(n11332), .ZN(
        n10868) );
  AND2_X1 U9180 ( .A1(n8469), .A2(n11766), .ZN(n11793) );
  OAI22_X1 U9181 ( .A1(n8450), .A2(n11741), .B1(n8436), .B2(n11740), .ZN(
        n11743) );
  OAI22_X1 U9182 ( .A1(n8450), .A2(n11322), .B1(n8437), .B2(n11321), .ZN(
        n11822) );
  AND2_X1 U9183 ( .A1(n8470), .A2(n11774), .ZN(n11804) );
  AND2_X1 U9184 ( .A1(n8464), .A2(n11775), .ZN(n11805) );
  AND2_X1 U9185 ( .A1(n8463), .A2(n11780), .ZN(n11810) );
  AND2_X1 U9186 ( .A1(n8459), .A2(n11779), .ZN(n11809) );
  AND2_X1 U9187 ( .A1(n8462), .A2(n11787), .ZN(n11746) );
  AND2_X1 U9188 ( .A1(n8463), .A2(n11786), .ZN(n11818) );
  AND2_X1 U9189 ( .A1(n8461), .A2(n11776), .ZN(n11806) );
  AND2_X1 U9190 ( .A1(n8462), .A2(n11788), .ZN(n11747) );
  AND2_X1 U9191 ( .A1(n8463), .A2(n11761), .ZN(n11816) );
  AND2_X1 U9192 ( .A1(n8463), .A2(n11783), .ZN(n11814) );
  AND2_X1 U9193 ( .A1(n8468), .A2(n11778), .ZN(n11808) );
  AND2_X1 U9194 ( .A1(n8467), .A2(n11777), .ZN(n11807) );
  AND2_X1 U9195 ( .A1(n8463), .A2(n11784), .ZN(n11815) );
  AND2_X1 U9196 ( .A1(n8462), .A2(n11789), .ZN(n11748) );
  AND2_X1 U9197 ( .A1(n8463), .A2(n11785), .ZN(n11817) );
  AND2_X1 U9198 ( .A1(n8463), .A2(n11760), .ZN(n11813) );
  AND2_X1 U9199 ( .A1(n8463), .A2(n11781), .ZN(n11811) );
  INV_X1 U9200 ( .A(n10095), .ZN(i_ADD_WS1[4]) );
  NAND2_X1 U9201 ( .A1(n8246), .A2(n8470), .ZN(n11830) );
  INV_X1 U9202 ( .A(n11731), .ZN(n9667) );
  INV_X1 U9203 ( .A(n11733), .ZN(n11731) );
  INV_X1 U9204 ( .A(n7771), .ZN(\DP_OP_751_130_6421/n1311 ) );
  NAND2_X1 U9205 ( .A1(n8493), .A2(n10226), .ZN(n10271) );
  OR2_X1 U9206 ( .A1(IR[31]), .A2(n166), .ZN(n10067) );
  NAND2_X1 U9207 ( .A1(n8491), .A2(n8490), .ZN(n8819) );
  INV_X1 U9208 ( .A(n11838), .ZN(n8426) );
  INV_X1 U9209 ( .A(n11838), .ZN(n8427) );
  NOR2_X1 U9210 ( .A1(RST), .A2(n11195), .ZN(n11196) );
  INV_X1 U9211 ( .A(n7755), .ZN(n8268) );
  INV_X1 U9212 ( .A(n7754), .ZN(n8263) );
  NOR2_X1 U9213 ( .A1(RST), .A2(n8269), .ZN(n11000) );
  NOR2_X1 U9214 ( .A1(RST), .A2(n8367), .ZN(n10930) );
  NOR2_X1 U9215 ( .A1(RST), .A2(n11318), .ZN(n11320) );
  NOR2_X1 U9216 ( .A1(RST), .A2(n11316), .ZN(n11315) );
  NOR2_X1 U9217 ( .A1(n8272), .A2(n8054), .ZN(n11119) );
  INV_X1 U9218 ( .A(n8420), .ZN(n8419) );
  NOR2_X1 U9219 ( .A1(RST), .A2(n11323), .ZN(n11325) );
  AND2_X1 U9220 ( .A1(n8463), .A2(n10980), .ZN(n11005) );
  AND2_X1 U9221 ( .A1(n8461), .A2(n10992), .ZN(n11030) );
  AND2_X1 U9222 ( .A1(n8464), .A2(n10961), .ZN(n11012) );
  AND2_X1 U9223 ( .A1(n8464), .A2(n10982), .ZN(n11013) );
  AND2_X1 U9224 ( .A1(n8462), .A2(n10993), .ZN(n11032) );
  AND2_X1 U9225 ( .A1(n8467), .A2(n10985), .ZN(n11029) );
  NOR2_X1 U9226 ( .A1(RST), .A2(n8372), .ZN(n10946) );
  NOR2_X1 U9227 ( .A1(RST), .A2(n8365), .ZN(n10927) );
  NOR2_X1 U9228 ( .A1(RST), .A2(n8362), .ZN(n10918) );
  AND2_X1 U9229 ( .A1(n8461), .A2(n10971), .ZN(n11027) );
  AND2_X1 U9230 ( .A1(n8459), .A2(n10984), .ZN(n11026) );
  AND2_X1 U9231 ( .A1(n8458), .A2(n10974), .ZN(n11031) );
  NOR2_X1 U9232 ( .A1(RST), .A2(n11759), .ZN(n11771) );
  NOR2_X1 U9233 ( .A1(RST), .A2(n10864), .ZN(n10863) );
  AND2_X1 U9234 ( .A1(n8469), .A2(n10964), .ZN(n11016) );
  AND2_X1 U9235 ( .A1(n8466), .A2(n10963), .ZN(n11015) );
  AND2_X1 U9236 ( .A1(n8459), .A2(n10965), .ZN(n11017) );
  AND2_X1 U9237 ( .A1(n8465), .A2(n10967), .ZN(n11021) );
  AND2_X1 U9238 ( .A1(n8458), .A2(n10990), .ZN(n11018) );
  AND2_X1 U9239 ( .A1(n8457), .A2(n10983), .ZN(n11023) );
  AND2_X1 U9240 ( .A1(n8470), .A2(n10969), .ZN(n11024) );
  AND2_X1 U9241 ( .A1(n8460), .A2(n10968), .ZN(n11022) );
  AND2_X1 U9242 ( .A1(n8464), .A2(n10991), .ZN(n11019) );
  AND2_X1 U9243 ( .A1(n8468), .A2(n10975), .ZN(n11033) );
  AND2_X1 U9244 ( .A1(n8464), .A2(n10976), .ZN(n11034) );
  AND2_X1 U9245 ( .A1(n8466), .A2(n11795), .ZN(n11751) );
  NOR2_X2 U9246 ( .A1(n10915), .A2(n11665), .ZN(n10802) );
  INV_X1 U9247 ( .A(n11661), .ZN(n11665) );
  OAI22_X1 U9248 ( .A1(n8450), .A2(n11737), .B1(n11736), .B2(n8437), .ZN(
        n11738) );
  NOR2_X2 U9249 ( .A1(n11662), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[15] ), 
        .ZN(n10915) );
  INV_X1 U9250 ( .A(n8295), .ZN(n10248) );
  INV_X1 U9251 ( .A(n10281), .ZN(n11735) );
  NOR2_X1 U9252 ( .A1(n10273), .A2(n179), .ZN(i_ADD_RS2[3]) );
  INV_X1 U9253 ( .A(n8779), .ZN(n8717) );
  INV_X1 U9254 ( .A(n11846), .ZN(n9270) );
  OR2_X1 U9255 ( .A1(n7648), .A2(n8286), .ZN(n8290) );
  OR2_X1 U9256 ( .A1(IR[31]), .A2(n8484), .ZN(n8241) );
  INV_X1 U9257 ( .A(n11626), .ZN(n11828) );
  NOR2_X1 U9258 ( .A1(RST), .A2(n11048), .ZN(n11047) );
  NOR2_X1 U9259 ( .A1(RST), .A2(n11168), .ZN(n11170) );
  NOR2_X1 U9260 ( .A1(RST), .A2(n11043), .ZN(n11042) );
  NOR2_X1 U9261 ( .A1(RST), .A2(n11094), .ZN(n11098) );
  NOR2_X1 U9262 ( .A1(RST), .A2(n11059), .ZN(n11061) );
  NOR2_X1 U9263 ( .A1(RST), .A2(n11165), .ZN(n11167) );
  NOR2_X1 U9264 ( .A1(RST), .A2(n11066), .ZN(n11069) );
  NOR2_X1 U9265 ( .A1(RST), .A2(n10921), .ZN(n10923) );
  OAI22_X1 U9266 ( .A1(n8293), .A2(n11741), .B1(n11740), .B2(n10999), .ZN(
        n10921) );
  NOR2_X1 U9267 ( .A1(RST), .A2(n11162), .ZN(n11164) );
  AND2_X1 U9268 ( .A1(n8466), .A2(n11093), .ZN(n11148) );
  AND2_X1 U9269 ( .A1(n8465), .A2(n11095), .ZN(n11150) );
  AND2_X1 U9270 ( .A1(n8461), .A2(n11181), .ZN(n11261) );
  AND2_X1 U9271 ( .A1(n8464), .A2(n11232), .ZN(n11259) );
  AND2_X1 U9272 ( .A1(n8465), .A2(n11111), .ZN(n11145) );
  AND2_X1 U9273 ( .A1(n8465), .A2(n11096), .ZN(n11152) );
  NOR2_X1 U9274 ( .A1(RST), .A2(n11039), .ZN(n11040) );
  NOR2_X1 U9275 ( .A1(RST), .A2(n10936), .ZN(n10938) );
  NOR2_X1 U9276 ( .A1(RST), .A2(n11329), .ZN(n11331) );
  NOR2_X1 U9277 ( .A1(RST), .A2(n11335), .ZN(n11337) );
  AND2_X1 U9278 ( .A1(n8469), .A2(n11388), .ZN(n11435) );
  NOR2_X1 U9279 ( .A1(RST), .A2(n11307), .ZN(n11309) );
  NOR2_X1 U9280 ( .A1(RST), .A2(n11305), .ZN(n11306) );
  AND2_X1 U9281 ( .A1(n8464), .A2(n11180), .ZN(n11255) );
  AND2_X1 U9282 ( .A1(n8466), .A2(n11179), .ZN(n11253) );
  AND2_X1 U9283 ( .A1(n8467), .A2(n11182), .ZN(n11263) );
  AND2_X1 U9284 ( .A1(n8467), .A2(n11227), .ZN(n11244) );
  AND2_X1 U9285 ( .A1(n8468), .A2(n11219), .ZN(n11268) );
  AND2_X1 U9286 ( .A1(n8467), .A2(n11177), .ZN(n11246) );
  AND2_X1 U9287 ( .A1(n8467), .A2(n11189), .ZN(n11242) );
  AND2_X1 U9288 ( .A1(n8469), .A2(n11399), .ZN(n11447) );
  AND2_X1 U9289 ( .A1(n8469), .A2(n11403), .ZN(n11597) );
  NOR2_X1 U9290 ( .A1(RST), .A2(n11310), .ZN(n11312) );
  OAI22_X1 U9291 ( .A1(n11415), .A2(n11745), .B1(n7756), .B2(n11744), .ZN(
        n11310) );
  AND2_X1 U9292 ( .A1(n8469), .A2(n11382), .ZN(n11429) );
  AND2_X1 U9293 ( .A1(n8469), .A2(n11401), .ZN(n11449) );
  AND2_X1 U9294 ( .A1(n8468), .A2(n11394), .ZN(n11442) );
  AND2_X1 U9295 ( .A1(n8468), .A2(n11400), .ZN(n11448) );
  AND2_X1 U9296 ( .A1(n8469), .A2(n11395), .ZN(n11443) );
  AND2_X1 U9297 ( .A1(n8466), .A2(n11055), .ZN(n11144) );
  AND2_X1 U9298 ( .A1(n8465), .A2(n11083), .ZN(n11136) );
  AND2_X1 U9299 ( .A1(n8465), .A2(n11067), .ZN(n11149) );
  AND2_X1 U9300 ( .A1(n8468), .A2(n11410), .ZN(n11438) );
  AND2_X1 U9301 ( .A1(n8470), .A2(n11397), .ZN(n11445) );
  AND2_X1 U9302 ( .A1(n8469), .A2(n11387), .ZN(n11434) );
  AND2_X1 U9303 ( .A1(n8467), .A2(n11174), .ZN(n11238) );
  AND2_X1 U9304 ( .A1(n8468), .A2(n11191), .ZN(n11270) );
  AND2_X1 U9305 ( .A1(n8467), .A2(n11175), .ZN(n11241) );
  AND2_X1 U9306 ( .A1(n8467), .A2(n11203), .ZN(n11240) );
  AND2_X1 U9307 ( .A1(n8460), .A2(n11178), .ZN(n11250) );
  AND2_X1 U9308 ( .A1(n8467), .A2(n11176), .ZN(n11243) );
  AND2_X1 U9309 ( .A1(n8468), .A2(n11183), .ZN(n11265) );
  AND2_X1 U9310 ( .A1(n8461), .A2(n11205), .ZN(n11254) );
  AND2_X1 U9311 ( .A1(n8467), .A2(n11213), .ZN(n11239) );
  AND2_X1 U9312 ( .A1(n8465), .A2(n11230), .ZN(n11256) );
  AND2_X1 U9313 ( .A1(n8468), .A2(n11184), .ZN(n11266) );
  AND2_X1 U9314 ( .A1(n8467), .A2(n11204), .ZN(n11247) );
  AND2_X1 U9315 ( .A1(n8462), .A2(n11231), .ZN(n11258) );
  AND2_X1 U9316 ( .A1(n8467), .A2(n11228), .ZN(n11248) );
  AND2_X1 U9317 ( .A1(n8468), .A2(n11207), .ZN(n11264) );
  AND2_X1 U9318 ( .A1(n8468), .A2(n11185), .ZN(n11267) );
  AND2_X1 U9319 ( .A1(n8467), .A2(n11214), .ZN(n11245) );
  AND2_X1 U9320 ( .A1(n8467), .A2(n11218), .ZN(n11260) );
  OAI22_X1 U9321 ( .A1(n11640), .A2(n11741), .B1(n11211), .B2(n11740), .ZN(
        n11157) );
  NOR2_X1 U9322 ( .A1(n836), .A2(n8054), .ZN(n11237) );
  INV_X1 U9323 ( .A(\DataPath/RF/c_win[3] ), .ZN(n8293) );
  AOI22_X1 U9324 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[4] ), 
        .B1(n10935), .B2(n10934), .ZN(n11772) );
  BUF_X2 U9325 ( .A(n10868), .Z(n8360) );
  BUF_X2 U9326 ( .A(n11756), .Z(n8434) );
  OAI22_X1 U9327 ( .A1(n8173), .A2(n11745), .B1(n8437), .B2(n11744), .ZN(
        n11756) );
  AOI22_X1 U9328 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[2] ), 
        .B1(n10925), .B2(n10934), .ZN(n11744) );
  BUF_X2 U9329 ( .A(n11743), .Z(n8432) );
  AOI22_X1 U9330 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[1] ), 
        .B1(n10920), .B2(n10934), .ZN(n11740) );
  BUF_X2 U9331 ( .A(n11822), .Z(n8440) );
  INV_X1 U9332 ( .A(n10280), .ZN(n11730) );
  AND2_X1 U9333 ( .A1(n10281), .A2(n10287), .ZN(n10280) );
  BUF_X1 U9334 ( .A(n8916), .Z(n8336) );
  NAND2_X1 U9335 ( .A1(n10292), .A2(IRAM_READY), .ZN(n8811) );
  BUF_X1 U9336 ( .A(n11463), .Z(n8413) );
  BUF_X1 U9337 ( .A(n11467), .Z(n8414) );
  BUF_X1 U9338 ( .A(n11511), .Z(n8417) );
  BUF_X1 U9339 ( .A(n11471), .Z(n8415) );
  BUF_X1 U9340 ( .A(n11459), .Z(n8412) );
  BUF_X1 U9341 ( .A(n11455), .Z(n8411) );
  BUF_X1 U9342 ( .A(n11475), .Z(n8416) );
  BUF_X1 U9343 ( .A(n10816), .Z(n8338) );
  INV_X1 U9344 ( .A(n11839), .ZN(n8422) );
  INV_X1 U9345 ( .A(n11839), .ZN(n8423) );
  INV_X1 U9346 ( .A(n11839), .ZN(n8424) );
  NOR2_X1 U9347 ( .A1(RST), .A2(n11154), .ZN(n11156) );
  NOR2_X1 U9348 ( .A1(RST), .A2(n11049), .ZN(n11051) );
  NOR2_X1 U9349 ( .A1(RST), .A2(n11159), .ZN(n11161) );
  NOR2_X1 U9350 ( .A1(RST), .A2(n11173), .ZN(n11187) );
  NOR2_X1 U9351 ( .A1(RST), .A2(n11052), .ZN(n11054) );
  NOR2_X1 U9352 ( .A1(RST), .A2(n11056), .ZN(n11058) );
  NOR2_X1 U9353 ( .A1(RST), .A2(n10973), .ZN(n10978) );
  NOR2_X1 U9354 ( .A1(RST), .A2(n10939), .ZN(n10941) );
  NOR2_X1 U9355 ( .A1(RST), .A2(n10942), .ZN(n10944) );
  OAI22_X1 U9356 ( .A1(n11640), .A2(n11773), .B1(n11211), .B2(n11772), .ZN(
        n11165) );
  AND2_X1 U9357 ( .A1(n8466), .A2(n11088), .ZN(n11141) );
  AND2_X1 U9358 ( .A1(n8466), .A2(n11087), .ZN(n11140) );
  AND2_X1 U9359 ( .A1(n8465), .A2(n11077), .ZN(n11128) );
  AND2_X1 U9360 ( .A1(n8466), .A2(n11082), .ZN(n11133) );
  AND2_X1 U9361 ( .A1(n8465), .A2(n11109), .ZN(n11134) );
  NOR2_X1 U9362 ( .A1(RST), .A2(n11377), .ZN(n11405) );
  NOR2_X1 U9363 ( .A1(RST), .A2(n11362), .ZN(n11365) );
  AND2_X1 U9364 ( .A1(n8469), .A2(n11383), .ZN(n11430) );
  OAI22_X1 U9365 ( .A1(n11415), .A2(n11741), .B1(n7756), .B2(n11740), .ZN(
        n11307) );
  OAI22_X1 U9366 ( .A1(n11415), .A2(n11737), .B1(n11736), .B2(n7756), .ZN(
        n11305) );
  AND2_X1 U9367 ( .A1(n8459), .A2(n11217), .ZN(n11257) );
  OAI22_X1 U9368 ( .A1(n11640), .A2(n11327), .B1(n11211), .B2(n11326), .ZN(
        n11172) );
  INV_X1 U9369 ( .A(n10693), .ZN(n10795) );
  AND2_X1 U9370 ( .A1(n8469), .A2(n11411), .ZN(n11451) );
  AND2_X1 U9371 ( .A1(n8469), .A2(n11390), .ZN(n11437) );
  AND2_X1 U9372 ( .A1(n8469), .A2(n11392), .ZN(n11440) );
  AND2_X1 U9373 ( .A1(n8469), .A2(n11389), .ZN(n11436) );
  AND2_X1 U9374 ( .A1(n8470), .A2(n11398), .ZN(n11446) );
  AND2_X1 U9375 ( .A1(n8469), .A2(n11385), .ZN(n11432) );
  AND2_X1 U9376 ( .A1(n8470), .A2(n11396), .ZN(n11444) );
  AND2_X1 U9377 ( .A1(n8466), .A2(n11079), .ZN(n11130) );
  AND2_X1 U9378 ( .A1(n8466), .A2(n11092), .ZN(n11147) );
  AND2_X1 U9379 ( .A1(n8465), .A2(n11107), .ZN(n11123) );
  AND2_X1 U9380 ( .A1(n8465), .A2(n11072), .ZN(n11121) );
  AND2_X1 U9381 ( .A1(n8466), .A2(n11080), .ZN(n11131) );
  AND2_X1 U9382 ( .A1(n8466), .A2(n11089), .ZN(n11142) );
  AND2_X1 U9383 ( .A1(n8464), .A2(n11076), .ZN(n11126) );
  AND2_X1 U9384 ( .A1(n8465), .A2(n11108), .ZN(n11127) );
  AND2_X1 U9385 ( .A1(n8465), .A2(n11086), .ZN(n11139) );
  AND2_X1 U9386 ( .A1(n8465), .A2(n11090), .ZN(n11143) );
  AND2_X1 U9387 ( .A1(n8465), .A2(n11091), .ZN(n11146) );
  AND2_X1 U9388 ( .A1(n8465), .A2(n11071), .ZN(n11120) );
  AND2_X1 U9389 ( .A1(n8464), .A2(n11074), .ZN(n11124) );
  OAI22_X1 U9390 ( .A1(n8271), .A2(n11745), .B1(n11744), .B2(n11102), .ZN(
        n11044) );
  AND2_X1 U9391 ( .A1(n8464), .A2(n11075), .ZN(n11125) );
  AND2_X1 U9392 ( .A1(n8458), .A2(n11206), .ZN(n11262) );
  AND2_X1 U9393 ( .A1(n8470), .A2(n11378), .ZN(n11420) );
  AND2_X1 U9394 ( .A1(n8470), .A2(n11391), .ZN(n11439) );
  AND2_X1 U9395 ( .A1(n8470), .A2(n11381), .ZN(n11428) );
  AND2_X1 U9396 ( .A1(n8465), .A2(n11216), .ZN(n11252) );
  AND2_X1 U9397 ( .A1(n8457), .A2(n11215), .ZN(n11251) );
  INV_X1 U9398 ( .A(n8275), .ZN(n11640) );
  OAI22_X1 U9399 ( .A1(n8293), .A2(n11333), .B1(n11332), .B2(n10999), .ZN(
        n10945) );
  OAI22_X1 U9400 ( .A1(n8293), .A2(n11745), .B1(n11744), .B2(n10999), .ZN(
        n10926) );
  OAI22_X1 U9401 ( .A1(n8293), .A2(n11737), .B1(n11736), .B2(n10999), .ZN(
        n10917) );
  INV_X2 U9402 ( .A(n8409), .ZN(n8408) );
  AOI22_X1 U9403 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[9] ), 
        .B1(n10876), .B2(n10934), .ZN(n11345) );
  AOI22_X1 U9404 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[3] ), 
        .B1(n10929), .B2(n10934), .ZN(n11757) );
  OAI22_X1 U9405 ( .A1(n8450), .A2(n11327), .B1(n8436), .B2(n11326), .ZN(
        n10864) );
  AOI22_X1 U9406 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[6] ), 
        .B1(n10843), .B2(n10934), .ZN(n11326) );
  NAND2_X1 U9407 ( .A1(n8460), .A2(n11513), .ZN(n11838) );
  INV_X1 U9408 ( .A(n11070), .ZN(n11355) );
  AOI22_X1 U9409 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[12] ), 
        .B1(n10893), .B2(n10934), .ZN(n11366) );
  AND2_X1 U9410 ( .A1(n10910), .A2(n11468), .ZN(n11369) );
  INV_X1 U9411 ( .A(n11359), .ZN(n11202) );
  NOR2_X1 U9412 ( .A1(i_ADD_WB[4]), .A2(n10870), .ZN(n10910) );
  INV_X1 U9413 ( .A(n10836), .ZN(n11505) );
  INV_X1 U9414 ( .A(n10835), .ZN(n11504) );
  INV_X1 U9415 ( .A(n10833), .ZN(n11502) );
  INV_X1 U9416 ( .A(n10837), .ZN(n11506) );
  INV_X1 U9417 ( .A(n10831), .ZN(n11500) );
  INV_X1 U9418 ( .A(n10832), .ZN(n11501) );
  INV_X1 U9419 ( .A(n10839), .ZN(n11508) );
  INV_X1 U9420 ( .A(n10840), .ZN(n11509) );
  AOI22_X1 U9421 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[7] ), 
        .B1(n10866), .B2(n10934), .ZN(n11332) );
  INV_X1 U9422 ( .A(n10834), .ZN(n11503) );
  INV_X1 U9423 ( .A(n10838), .ZN(n11507) );
  AOI22_X1 U9424 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[5] ), 
        .B1(n10828), .B2(n10934), .ZN(n11321) );
  INV_X1 U9425 ( .A(n7648), .ZN(n8450) );
  INV_X1 U9426 ( .A(n10844), .ZN(n11479) );
  INV_X1 U9427 ( .A(n10860), .ZN(n11495) );
  INV_X1 U9428 ( .A(n10845), .ZN(n11480) );
  INV_X1 U9429 ( .A(n10850), .ZN(n11485) );
  INV_X1 U9430 ( .A(n10849), .ZN(n11484) );
  INV_X1 U9431 ( .A(n10841), .ZN(n11512) );
  INV_X1 U9432 ( .A(n10826), .ZN(n11497) );
  INV_X1 U9433 ( .A(n10852), .ZN(n11487) );
  INV_X1 U9434 ( .A(n10858), .ZN(n11493) );
  INV_X1 U9435 ( .A(n10846), .ZN(n11481) );
  INV_X1 U9436 ( .A(n10829), .ZN(n11498) );
  INV_X1 U9437 ( .A(n10856), .ZN(n11491) );
  INV_X1 U9438 ( .A(n10854), .ZN(n11489) );
  INV_X1 U9439 ( .A(n10859), .ZN(n11494) );
  INV_X1 U9440 ( .A(n10848), .ZN(n11483) );
  INV_X1 U9441 ( .A(n10847), .ZN(n11482) );
  INV_X1 U9442 ( .A(n10855), .ZN(n11490) );
  INV_X1 U9443 ( .A(n10830), .ZN(n11499) );
  INV_X1 U9444 ( .A(n10861), .ZN(n11496) );
  INV_X1 U9445 ( .A(n10857), .ZN(n11492) );
  INV_X1 U9446 ( .A(n10853), .ZN(n11488) );
  INV_X1 U9447 ( .A(n10851), .ZN(n11486) );
  BUF_X1 U9448 ( .A(i_S3), .Z(n8451) );
  OAI211_X1 U9449 ( .C1(n10249), .C2(n181), .A(n10248), .B(n10103), .ZN(
        i_ADD_WS1[1]) );
  NOR2_X1 U9450 ( .A1(n566), .A2(n11567), .ZN(n11568) );
  NOR2_X1 U9451 ( .A1(n564), .A2(n11564), .ZN(n11565) );
  NOR2_X1 U9452 ( .A1(n562), .A2(n11561), .ZN(n11562) );
  INV_X1 U9453 ( .A(n10279), .ZN(n10032) );
  AND2_X1 U9454 ( .A1(n7769), .A2(n8105), .ZN(n10281) );
  NOR2_X1 U9455 ( .A1(n11830), .A2(n8191), .ZN(n10290) );
  INV_X1 U9456 ( .A(n9589), .ZN(n9686) );
  NAND2_X1 U9457 ( .A1(n10155), .A2(n10154), .ZN(n10175) );
  INV_X1 U9458 ( .A(n8130), .ZN(n8287) );
  NAND2_X1 U9459 ( .A1(DRAM_ISSUE), .A2(n8245), .ZN(n8246) );
  AOI21_X1 U9460 ( .B1(DRAM_READNOTWRITE), .B2(n8277), .A(n8278), .ZN(
        DRAM_ISSUE) );
  AND2_X1 U9461 ( .A1(\DataPath/RF/POP_ADDRGEN/curr_state[1] ), .A2(n877), 
        .ZN(n8484) );
  INV_X1 U9462 ( .A(n10104), .ZN(n10119) );
  NOR2_X1 U9463 ( .A1(RST), .A2(n11222), .ZN(n11220) );
  NOR2_X1 U9464 ( .A1(RST), .A2(n11210), .ZN(n11208) );
  OAI22_X1 U9465 ( .A1(n8271), .A2(n11333), .B1(n11332), .B2(n11102), .ZN(
        n11059) );
  AND2_X1 U9466 ( .A1(n8466), .A2(n11078), .ZN(n11129) );
  NOR2_X1 U9467 ( .A1(RST), .A2(n11372), .ZN(n11370) );
  OAI22_X1 U9468 ( .A1(n8293), .A2(n11773), .B1(n11772), .B2(n10999), .ZN(
        n10936) );
  AND2_X1 U9469 ( .A1(n8468), .A2(n11379), .ZN(n11424) );
  AND2_X1 U9470 ( .A1(n8470), .A2(n11386), .ZN(n11433) );
  AND2_X1 U9471 ( .A1(n8470), .A2(n11380), .ZN(n11425) );
  AND2_X1 U9472 ( .A1(n8470), .A2(n11384), .ZN(n11431) );
  BUF_X2 U9473 ( .A(n11001), .Z(n8269) );
  OAI222_X1 U9474 ( .A1(n10999), .A2(n10998), .B1(n11407), .B2(n8271), .C1(
        n11406), .C2(n8293), .ZN(n11001) );
  BUF_X2 U9475 ( .A(n10931), .Z(n8367) );
  OAI22_X1 U9476 ( .A1(n8293), .A2(n11758), .B1(n11757), .B2(n10999), .ZN(
        n10931) );
  BUF_X2 U9477 ( .A(n11172), .Z(n8394) );
  AND2_X1 U9478 ( .A1(n8466), .A2(n7778), .ZN(n11135) );
  AND2_X1 U9479 ( .A1(n8465), .A2(n7779), .ZN(n11122) );
  AND2_X1 U9480 ( .A1(n8466), .A2(n7780), .ZN(n11137) );
  AND2_X1 U9481 ( .A1(n8466), .A2(n7781), .ZN(n11132) );
  AND2_X1 U9482 ( .A1(n8466), .A2(n11085), .ZN(n11138) );
  AND2_X1 U9483 ( .A1(n8470), .A2(n11402), .ZN(n11450) );
  INV_X1 U9484 ( .A(\DataPath/RF/c_win[0] ), .ZN(n11415) );
  AND2_X1 U9485 ( .A1(n8459), .A2(n11229), .ZN(n11249) );
  INV_X1 U9486 ( .A(n10998), .ZN(n11409) );
  AOI22_X1 U9487 ( .A1(n10295), .A2(n8195), .B1(n10898), .B2(n10934), .ZN(
        n11373) );
  INV_X1 U9488 ( .A(n11194), .ZN(n11348) );
  AOI22_X1 U9489 ( .A1(n10295), .A2(n8194), .B1(n10869), .B2(n10934), .ZN(
        n11341) );
  BUF_X1 U9490 ( .A(n589), .Z(n8271) );
  OAI22_X1 U9491 ( .A1(n10295), .A2(n10908), .B1(n10916), .B2(n8172), .ZN(
        n11418) );
  NAND3_X1 U9492 ( .A1(\CU_I/CW_ID[ID_EN] ), .A2(n8246), .A3(n8457), .ZN(
        n11839) );
  AOI22_X1 U9493 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[11] ), 
        .B1(n10888), .B2(n10934), .ZN(n11361) );
  NOR2_X1 U9494 ( .A1(n8102), .A2(n10870), .ZN(n10909) );
  NAND2_X1 U9495 ( .A1(i_ADD_WB[3]), .A2(i_WF), .ZN(n10870) );
  OAI22_X1 U9496 ( .A1(\DataPath/RF/POP_ADDRGEN/curr_addr[0] ), .A2(n10916), 
        .B1(n10295), .B2(n11660), .ZN(n11736) );
  AOI21_X1 U9497 ( .B1(n7954), .B2(n8135), .A(n10245), .ZN(n10102) );
  NOR2_X1 U9498 ( .A1(n576), .A2(n11582), .ZN(n11583) );
  NOR2_X1 U9499 ( .A1(n574), .A2(n11579), .ZN(n11580) );
  NOR2_X1 U9500 ( .A1(n572), .A2(n11576), .ZN(n11577) );
  NOR2_X1 U9501 ( .A1(n570), .A2(n11573), .ZN(n11574) );
  NOR2_X1 U9502 ( .A1(n568), .A2(n11570), .ZN(n11571) );
  NOR2_X1 U9503 ( .A1(n560), .A2(n11558), .ZN(n11559) );
  NOR2_X1 U9504 ( .A1(n558), .A2(n11555), .ZN(n11556) );
  NOR2_X2 U9505 ( .A1(n8803), .A2(n8811), .ZN(n10258) );
  AND4_X1 U9506 ( .A1(n9570), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(n8121)
         );
  INV_X1 U9507 ( .A(n10020), .ZN(n9918) );
  NOR2_X1 U9508 ( .A1(n7769), .A2(RST), .ZN(n10289) );
  AND2_X1 U9509 ( .A1(n8943), .A2(n8958), .ZN(n9992) );
  AND2_X1 U9510 ( .A1(n9067), .A2(n9017), .ZN(n10020) );
  INV_X1 U9511 ( .A(n9942), .ZN(n10021) );
  AND2_X1 U9512 ( .A1(n9017), .A2(n9068), .ZN(n10023) );
  INV_X1 U9513 ( .A(n9593), .ZN(n9691) );
  NAND2_X1 U9514 ( .A1(n8819), .A2(n8497), .ZN(n10108) );
  AND2_X1 U9515 ( .A1(\DataPath/RF/c_win[3] ), .A2(n8272), .ZN(n8288) );
  NOR2_X1 U9516 ( .A1(\DataPath/RF/PUSH_ADDRGEN/curr_state[0] ), .A2(n849), 
        .ZN(n10308) );
  NOR2_X1 U9517 ( .A1(n471), .A2(n470), .ZN(\DP_OP_1091J1_126_6973/n72 ) );
  NOR2_X1 U9518 ( .A1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[15] ), .A2(n10821), 
        .ZN(n10816) );
  NOR2_X1 U9519 ( .A1(n8246), .A2(RST), .ZN(n11626) );
  NOR2_X1 U9520 ( .A1(n11839), .A2(n10109), .ZN(n10104) );
  INV_X2 U9521 ( .A(n11838), .ZN(n8425) );
  OAI22_X1 U9522 ( .A1(n8271), .A2(n11758), .B1(n11757), .B2(n11102), .ZN(
        n11048) );
  OAI22_X1 U9523 ( .A1(n11640), .A2(n11322), .B1(n11211), .B2(n11321), .ZN(
        n11168) );
  OAI22_X1 U9524 ( .A1(n8271), .A2(n11741), .B1(n11740), .B2(n11102), .ZN(
        n11043) );
  NOR2_X1 U9525 ( .A1(RST), .A2(n8268), .ZN(n10986) );
  NOR2_X1 U9526 ( .A1(RST), .A2(n8263), .ZN(n10951) );
  OAI22_X1 U9527 ( .A1(n11415), .A2(n11327), .B1(n7756), .B2(n11326), .ZN(
        n11329) );
  OAI22_X1 U9528 ( .A1(n11415), .A2(n11333), .B1(n7756), .B2(n11332), .ZN(
        n11335) );
  AOI211_X1 U9529 ( .C1(n11355), .C2(\DataPath/RF/c_win[3] ), .A(RST), .B(
        n10953), .ZN(n10955) );
  INV_X1 U9530 ( .A(n10777), .ZN(n10785) );
  INV_X1 U9531 ( .A(n10800), .ZN(n10703) );
  AOI22_X1 U9532 ( .A1(n7762), .A2(n11287), .B1(n11494), .B2(n11102), .ZN(
        n11110) );
  AOI22_X1 U9533 ( .A1(n7762), .A2(n11274), .B1(n11481), .B2(n11102), .ZN(
        n11073) );
  AOI22_X1 U9534 ( .A1(n7762), .A2(n11289), .B1(n11496), .B2(n11102), .ZN(
        n11084) );
  AOI22_X1 U9535 ( .A1(n7762), .A2(n11284), .B1(n11491), .B2(n11102), .ZN(
        n11081) );
  AOI211_X1 U9536 ( .C1(n8410), .C2(n11418), .A(RST), .B(n11417), .ZN(n11598)
         );
  AOI211_X1 U9537 ( .C1(n8410), .C2(n11409), .A(RST), .B(n11408), .ZN(n11413)
         );
  OAI22_X1 U9538 ( .A1(n10934), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[14] ), 
        .B1(n10904), .B2(n10295), .ZN(n10998) );
  NOR3_X1 U9539 ( .A1(n537), .A2(i_ADD_WB[1]), .A3(i_ADD_WB[2]), .ZN(n11477)
         );
  NOR3_X1 U9540 ( .A1(i_ADD_WB[0]), .A2(n539), .A3(i_ADD_WB[1]), .ZN(n11464)
         );
  NOR3_X1 U9541 ( .A1(i_ADD_WB[2]), .A2(n8170), .A3(n537), .ZN(n11468) );
  INV_X1 U9542 ( .A(n11546), .ZN(n11298) );
  INV_X1 U9543 ( .A(n11545), .ZN(n11297) );
  INV_X1 U9544 ( .A(n11543), .ZN(n11295) );
  INV_X1 U9545 ( .A(n11547), .ZN(n11299) );
  INV_X1 U9546 ( .A(n11541), .ZN(n11293) );
  INV_X1 U9547 ( .A(n11542), .ZN(n11294) );
  INV_X1 U9548 ( .A(n11549), .ZN(n11301) );
  INV_X1 U9549 ( .A(n11550), .ZN(n11302) );
  INV_X1 U9550 ( .A(n11544), .ZN(n11296) );
  INV_X1 U9551 ( .A(n11548), .ZN(n11300) );
  NOR3_X1 U9552 ( .A1(n539), .A2(n537), .A3(i_ADD_WB[1]), .ZN(n11460) );
  NOR3_X1 U9553 ( .A1(i_ADD_WB[0]), .A2(n8170), .A3(n539), .ZN(n11456) );
  NOR3_X1 U9554 ( .A1(i_ADD_WB[2]), .A2(i_ADD_WB[0]), .A3(n8170), .ZN(n11472)
         );
  INV_X1 U9555 ( .A(n11520), .ZN(n11272) );
  INV_X1 U9556 ( .A(n11536), .ZN(n11288) );
  INV_X1 U9557 ( .A(n11521), .ZN(n11273) );
  INV_X1 U9558 ( .A(n11526), .ZN(n11278) );
  INV_X1 U9559 ( .A(n11525), .ZN(n11277) );
  INV_X1 U9560 ( .A(n11551), .ZN(n11304) );
  INV_X1 U9561 ( .A(n11538), .ZN(n11290) );
  INV_X1 U9562 ( .A(n11528), .ZN(n11280) );
  INV_X1 U9563 ( .A(n11534), .ZN(n11286) );
  INV_X1 U9564 ( .A(n11522), .ZN(n11274) );
  INV_X1 U9565 ( .A(n11539), .ZN(n11291) );
  INV_X1 U9566 ( .A(n11532), .ZN(n11284) );
  INV_X1 U9567 ( .A(n11530), .ZN(n11282) );
  INV_X1 U9568 ( .A(n11535), .ZN(n11287) );
  INV_X1 U9569 ( .A(n11524), .ZN(n11276) );
  INV_X1 U9570 ( .A(n11523), .ZN(n11275) );
  INV_X1 U9571 ( .A(n11531), .ZN(n11283) );
  INV_X1 U9572 ( .A(n11540), .ZN(n11292) );
  INV_X1 U9573 ( .A(n11537), .ZN(n11289) );
  INV_X1 U9574 ( .A(n11533), .ZN(n11285) );
  INV_X1 U9575 ( .A(n11529), .ZN(n11281) );
  INV_X1 U9576 ( .A(n11527), .ZN(n11279) );
  NOR2_X1 U9577 ( .A1(n466), .A2(n11513), .ZN(\DECODEhw/i_WR1 ) );
  NAND2_X1 U9578 ( .A1(\CU_I/CW_ID[ID_EN] ), .A2(n8246), .ZN(n11513) );
  NOR2_X1 U9579 ( .A1(n578), .A2(n11585), .ZN(n11586) );
  INV_X1 U9580 ( .A(n10292), .ZN(n10257) );
  INV_X1 U9581 ( .A(n10284), .ZN(n9982) );
  AND2_X1 U9582 ( .A1(n10281), .A2(n9815), .ZN(n10279) );
  INV_X1 U9583 ( .A(n10287), .ZN(n9815) );
  INV_X1 U9584 ( .A(n10010), .ZN(n9880) );
  INV_X1 U9585 ( .A(n9939), .ZN(n10013) );
  INV_X1 U9586 ( .A(n10023), .ZN(n9878) );
  INV_X1 U9587 ( .A(n9978), .ZN(n10027) );
  INV_X1 U9588 ( .A(n9958), .ZN(n9935) );
  AND2_X1 U9589 ( .A1(i_ALU_OP[0]), .A2(i_ALU_OP[1]), .ZN(n10287) );
  INV_X1 U9590 ( .A(n10286), .ZN(n10017) );
  OR2_X1 U9591 ( .A1(n7688), .A2(n7690), .ZN(n9589) );
  NOR2_X1 U9592 ( .A1(n8182), .A2(i_ALU_OP[1]), .ZN(n10004) );
  AND4_X1 U9593 ( .A1(n10297), .A2(n8488), .A3(n10216), .A4(n10067), .ZN(n8138) );
  OR2_X1 U9594 ( .A1(RST), .A2(i_RF1), .ZN(\DataPath/RF/RDPORT0_OUTLATCH/N3 )
         );
  OR2_X1 U9595 ( .A1(RST), .A2(i_RF2), .ZN(\DataPath/RF/RDPORT1_OUTLATCH/N3 )
         );
  INV_X1 U9596 ( .A(RST), .ZN(n8461) );
  AND2_X1 U9597 ( .A1(n8244), .A2(n8489), .ZN(n10141) );
  BUF_X1 U9598 ( .A(n10678), .Z(n8352) );
  BUF_X1 U9599 ( .A(n10681), .Z(n8355) );
  OR2_X1 U9600 ( .A1(n10353), .A2(n10352), .ZN(n10356) );
  BUF_X1 U9601 ( .A(n10670), .Z(n8341) );
  BUF_X1 U9602 ( .A(n10669), .Z(n8339) );
  NOR2_X1 U9603 ( .A1(n10357), .A2(n10341), .ZN(n10669) );
  BUF_X1 U9604 ( .A(n10666), .Z(n8347) );
  NOR2_X1 U9605 ( .A1(n10357), .A2(n10342), .ZN(n10666) );
  NAND2_X1 U9606 ( .A1(n10335), .A2(n10336), .ZN(n10357) );
  OR2_X1 U9607 ( .A1(n10351), .A2(n10349), .ZN(n10342) );
  NAND2_X1 U9608 ( .A1(n10934), .A2(n10818), .ZN(n10314) );
  INV_X1 U9609 ( .A(RST), .ZN(n8459) );
  INV_X1 U9610 ( .A(RST), .ZN(n8458) );
  NAND3_X1 U9611 ( .A1(n11468), .A2(n11476), .A3(n8457), .ZN(n11471) );
  NAND3_X1 U9612 ( .A1(n11456), .A2(n11476), .A3(n8457), .ZN(n11459) );
  NAND3_X1 U9613 ( .A1(n11460), .A2(n11476), .A3(n8457), .ZN(n11463) );
  NAND3_X1 U9614 ( .A1(n11464), .A2(n11476), .A3(n8457), .ZN(n11467) );
  NAND3_X1 U9615 ( .A1(n11452), .A2(n11476), .A3(n8457), .ZN(n11455) );
  NAND3_X1 U9616 ( .A1(n11472), .A2(n11476), .A3(n8457), .ZN(n11475) );
  NAND3_X1 U9617 ( .A1(n11477), .A2(n11476), .A3(n8457), .ZN(n11511) );
  NOR2_X1 U9618 ( .A1(RST), .A2(n11358), .ZN(n11356) );
  INV_X1 U9619 ( .A(n10760), .ZN(n10791) );
  NOR2_X1 U9620 ( .A1(n10754), .A2(n10732), .ZN(n10777) );
  NAND2_X1 U9621 ( .A1(n10731), .A2(n10780), .ZN(n10754) );
  NOR2_X1 U9622 ( .A1(n11616), .A2(n10755), .ZN(n10760) );
  NOR2_X1 U9623 ( .A1(n10797), .A2(n10691), .ZN(n10741) );
  NOR2_X1 U9624 ( .A1(DATA_SIZE[1]), .A2(n10795), .ZN(n10797) );
  INV_X1 U9625 ( .A(RST), .ZN(n8466) );
  INV_X1 U9626 ( .A(RST), .ZN(n8465) );
  INV_X1 U9627 ( .A(RST), .ZN(n8469) );
  AOI22_X1 U9628 ( .A1(n8410), .A2(n11279), .B1(n11486), .B2(n7756), .ZN(
        n11381) );
  AOI22_X1 U9629 ( .A1(n8410), .A2(n11297), .B1(n11504), .B2(n7756), .ZN(
        n11398) );
  AOI22_X1 U9630 ( .A1(n8410), .A2(n11295), .B1(n11502), .B2(n7756), .ZN(
        n11396) );
  AOI22_X1 U9631 ( .A1(n8410), .A2(n11283), .B1(n11490), .B2(n7756), .ZN(
        n11385) );
  AOI22_X1 U9632 ( .A1(n8410), .A2(n11288), .B1(n11495), .B2(n7756), .ZN(
        n11390) );
  INV_X1 U9633 ( .A(RST), .ZN(n8470) );
  NOR2_X1 U9634 ( .A1(RST), .A2(n10880), .ZN(n10878) );
  INV_X1 U9635 ( .A(RST), .ZN(n8468) );
  INV_X1 U9636 ( .A(RST), .ZN(n8467) );
  AOI22_X1 U9637 ( .A1(n8410), .A2(n11302), .B1(n11509), .B2(n7756), .ZN(
        n11411) );
  NOR2_X1 U9638 ( .A1(RST), .A2(n8408), .ZN(n11412) );
  INV_X1 U9639 ( .A(RST), .ZN(n8457) );
  INV_X1 U9640 ( .A(RST), .ZN(n8460) );
  INV_X1 U9641 ( .A(RST), .ZN(n8464) );
  INV_X1 U9642 ( .A(RST), .ZN(n8463) );
  NOR3_X1 U9643 ( .A1(n539), .A2(n537), .A3(n8170), .ZN(n11452) );
  INV_X1 U9644 ( .A(n10097), .ZN(i_ADD_WS1[3]) );
  INV_X1 U9645 ( .A(n9460), .ZN(n9459) );
  AND2_X1 U9646 ( .A1(n7732), .A2(\DataPath/i_PIPLIN_A[31] ), .ZN(n9361) );
  INV_X1 U9647 ( .A(n9631), .ZN(n9026) );
  AND2_X1 U9648 ( .A1(n7732), .A2(\DataPath/i_PIPLIN_A[30] ), .ZN(n9631) );
  BUF_X1 U9649 ( .A(n8308), .Z(n8309) );
  INV_X1 U9650 ( .A(\DP_OP_751_130_6421/n393 ), .ZN(n9824) );
  INV_X1 U9651 ( .A(\DP_OP_751_130_6421/n597 ), .ZN(n9847) );
  BUF_X1 U9652 ( .A(n8305), .Z(n8307) );
  XNOR2_X1 U9653 ( .A(\DP_OP_751_130_6421/n801 ), .B(n9646), .ZN(n8923) );
  INV_X1 U9654 ( .A(n7782), .ZN(n9609) );
  XNOR2_X1 U9655 ( .A(\DP_OP_751_130_6421/n903 ), .B(n9660), .ZN(n8916) );
  OAI21_X1 U9656 ( .B1(n8131), .B2(n7907), .A(n8910), .ZN(
        \DP_OP_751_130_6421/n801 ) );
  OAI21_X1 U9657 ( .B1(n8151), .B2(n7940), .A(n8903), .ZN(
        \DP_OP_751_130_6421/n903 ) );
  BUF_X1 U9658 ( .A(n9951), .Z(n8304) );
  INV_X1 U9659 ( .A(\DP_OP_751_130_6421/n1209 ), .ZN(n8448) );
  AND2_X1 U9660 ( .A1(n7732), .A2(\DataPath/i_PIPLIN_A[21] ), .ZN(n9889) );
  BUF_X1 U9661 ( .A(n8884), .Z(n8335) );
  BUF_X1 U9662 ( .A(n8869), .Z(n8328) );
  BUF_X1 U9663 ( .A(n8872), .Z(n8332) );
  INV_X1 U9664 ( .A(\DP_OP_751_130_6421/n1617 ), .ZN(n8445) );
  INV_X1 U9665 ( .A(i_NPC_SEL), .ZN(n8812) );
  OR2_X2 U9666 ( .A1(n7736), .A2(n8820), .ZN(n10153) );
  NOR2_X1 U9667 ( .A1(n10270), .A2(n177), .ZN(i_ADD_RS1[0]) );
  NOR2_X1 U9668 ( .A1(n10270), .A2(n174), .ZN(i_ADD_RS1[3]) );
  NOR2_X1 U9669 ( .A1(n10270), .A2(n175), .ZN(i_ADD_RS1[2]) );
  NOR2_X1 U9670 ( .A1(n10270), .A2(n176), .ZN(i_ADD_RS1[1]) );
  NOR2_X1 U9671 ( .A1(n10270), .A2(n173), .ZN(i_ADD_RS1[4]) );
  NOR2_X1 U9672 ( .A1(n10220), .A2(n10232), .ZN(n10291) );
  INV_X1 U9673 ( .A(RST), .ZN(n8462) );
  INV_X1 U9674 ( .A(DRAM_READY), .ZN(n8245) );
  AOI211_X4 U9675 ( .C1(n8275), .C2(n11202), .A(RST), .B(n11201), .ZN(n11210)
         );
  AOI211_X4 U9676 ( .C1(\DataPath/RF/c_win[1] ), .C2(n11369), .A(RST), .B(
        n11212), .ZN(n11222) );
  AOI211_X4 U9677 ( .C1(n7762), .C2(n11341), .A(RST), .B(n11062), .ZN(n11065)
         );
  AOI211_X4 U9678 ( .C1(n7762), .C2(n11373), .A(RST), .B(n11106), .ZN(n11114)
         );
  AOI211_X4 U9679 ( .C1(n7761), .C2(n11409), .A(RST), .B(n11226), .ZN(n11235)
         );
  AOI211_X4 U9680 ( .C1(n7761), .C2(n11341), .A(RST), .B(n11188), .ZN(n11193)
         );
  AOI211_X4 U9681 ( .C1(n7762), .C2(n11418), .A(RST), .B(n11118), .ZN(n11153)
         );
  AOI211_X4 U9682 ( .C1(n7762), .C2(n11409), .A(RST), .B(n11115), .ZN(n11117)
         );
  AOI211_X4 U9683 ( .C1(n7761), .C2(n11418), .A(RST), .B(n11236), .ZN(n11271)
         );
  AOI211_X4 U9684 ( .C1(n7761), .C2(n11373), .A(RST), .B(n11223), .ZN(n11225)
         );
  AOI211_X4 U9685 ( .C1(\DataPath/RF/c_win[1] ), .C2(n11355), .A(RST), .B(
        n11197), .ZN(n11200) );
  AOI211_X4 U9686 ( .C1(n11369), .C2(\DataPath/RF/c_win[2] ), .A(RST), .B(
        n11103), .ZN(n11105) );
  AOI211_X4 U9687 ( .C1(n11202), .C2(\DataPath/RF/c_win[2] ), .A(RST), .B(
        n11099), .ZN(n11101) );
  OAI222_X4 U9688 ( .A1(n11345), .A2(n11211), .B1(n11346), .B2(n11415), .C1(
        n11640), .C2(n11194), .ZN(n11195) );
  AOI211_X4 U9689 ( .C1(\DataPath/RF/c_win[0] ), .C2(n11369), .A(RST), .B(
        n11368), .ZN(n11372) );
  AOI211_X4 U9690 ( .C1(\DataPath/RF/c_win[0] ), .C2(n11355), .A(RST), .B(
        n11354), .ZN(n11358) );
  AOI211_X1 U9691 ( .C1(n11348), .C2(\DataPath/RF/c_win[3] ), .A(RST), .B(
        n10950), .ZN(n10952) );
  AOI211_X1 U9692 ( .C1(n11369), .C2(\DataPath/RF/c_win[3] ), .A(RST), .B(
        n10979), .ZN(n10987) );
  AOI211_X4 U9693 ( .C1(n8410), .C2(n11341), .A(RST), .B(n11340), .ZN(n11344)
         );
  AOI211_X4 U9694 ( .C1(n8183), .C2(n11341), .A(RST), .B(n10871), .ZN(n10874)
         );
  AOI211_X4 U9695 ( .C1(n8183), .C2(n11373), .A(RST), .B(n10899), .ZN(n10902)
         );
  AOI211_X4 U9696 ( .C1(\DataPath/RF/c_win[0] ), .C2(n11348), .A(RST), .B(
        n11347), .ZN(n11351) );
  AOI211_X4 U9697 ( .C1(n8183), .C2(n11418), .A(RST), .B(n10912), .ZN(n10914)
         );
  AOI211_X4 U9698 ( .C1(n8183), .C2(n11409), .A(RST), .B(n10905), .ZN(n10907)
         );
  AOI221_X4 U9699 ( .B1(n8410), .B2(n11292), .C1(n7756), .C2(n11499), .A(RST), 
        .ZN(n11441) );
  AOI22_X2 U9700 ( .A1(n11419), .A2(n11278), .B1(n11485), .B2(n7756), .ZN(
        n11426) );
  AOI22_X2 U9701 ( .A1(n11419), .A2(n11273), .B1(n11480), .B2(n7756), .ZN(
        n11421) );
  AOI211_X4 U9702 ( .C1(n11003), .C2(n11373), .A(RST), .B(n10988), .ZN(n10997)
         );
  AOI211_X4 U9703 ( .C1(n7648), .C2(n11348), .A(RST), .B(n10877), .ZN(n10880)
         );
  AOI211_X4 U9704 ( .C1(n11003), .C2(n11341), .A(RST), .B(n10947), .ZN(n10949)
         );
  AOI211_X4 U9705 ( .C1(n11003), .C2(n11418), .A(RST), .B(n11002), .ZN(n11037)
         );
  AOI211_X4 U9706 ( .C1(n7648), .C2(n11355), .A(RST), .B(n10883), .ZN(n10886)
         );
  AOI211_X4 U9707 ( .C1(n7648), .C2(n11369), .A(RST), .B(n10894), .ZN(n10897)
         );
  AOI211_X4 U9708 ( .C1(n7648), .C2(n11202), .A(RST), .B(n10889), .ZN(n10891)
         );
  NOR3_X1 U9709 ( .A1(i_ADD_WB[1]), .A2(i_ADD_WB[0]), .A3(i_ADD_WB[2]), .ZN(
        n10911) );
  NOR2_X1 U9710 ( .A1(n10295), .A2(n11661), .ZN(n10916) );
  OAI21_X1 U9711 ( .B1(\DataPath/RF/POP_ADDRGEN/curr_state[1] ), .B2(n877), 
        .A(n10801), .ZN(n11661) );
  NAND2_X1 U9712 ( .A1(\DataPath/RF/POP_ADDRGEN/curr_state[1] ), .A2(n877), 
        .ZN(n10801) );
  NOR2_X2 U9713 ( .A1(n8957), .A2(n8956), .ZN(n9990) );
  NOR2_X2 U9714 ( .A1(n7942), .A2(n9667), .ZN(n9687) );
  NOR2_X2 U9715 ( .A1(n7785), .A2(n9088), .ZN(n10286) );
  NOR2_X2 U9716 ( .A1(n9054), .A2(n9069), .ZN(n10010) );
  NOR2_X2 U9717 ( .A1(n9053), .A2(n9052), .ZN(n10284) );
  AOI21_X2 U9718 ( .B1(n8969), .B2(n8968), .A(n8260), .ZN(n9978) );
  OAI21_X2 U9719 ( .B1(n8132), .B2(n7907), .A(n8928), .ZN(
        \DP_OP_751_130_6421/n495 ) );
  INV_X2 U9720 ( .A(n9230), .ZN(n8941) );
  INV_X2 U9721 ( .A(n8447), .ZN(\DP_OP_751_130_6421/n1413 ) );
  AND4_X2 U9722 ( .A1(n8678), .A2(n8771), .A3(n8677), .A4(n8776), .ZN(n8119)
         );
  AOI211_X1 U9723 ( .C1(n10236), .C2(n8115), .A(n10235), .B(n10234), .ZN(
        n10237) );
  AOI21_X1 U9724 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(n10238) );
  NOR2_X1 U9725 ( .A1(n10137), .A2(n11667), .ZN(n10274) );
  AOI211_X1 U9726 ( .C1(n10141), .C2(n10138), .A(n10136), .B(n10143), .ZN(
        n10137) );
  NOR2_X1 U9727 ( .A1(n10301), .A2(n10138), .ZN(\CU_I/CW[DATA_SIZE][0] ) );
  NOR2_X1 U9728 ( .A1(n10301), .A2(n10139), .ZN(\CU_I/CW[DATA_SIZE][1] ) );
  NAND2_X1 U9729 ( .A1(n10145), .A2(n10144), .ZN(\CU_I/CW[MUXB_SEL] ) );
  INV_X1 U9730 ( .A(n10143), .ZN(n10145) );
  NAND2_X1 U9731 ( .A1(n10215), .A2(n10214), .ZN(\CU_I/CW[NPC_SEL] ) );
  INV_X1 U9732 ( .A(n7990), .ZN(n10215) );
  OAI211_X1 U9733 ( .C1(n172), .C2(n10228), .A(n10230), .B(n10227), .ZN(
        \CU_I/CW[SEL_CMPB] ) );
  AOI211_X1 U9734 ( .C1(n7954), .C2(n10225), .A(n10224), .B(n10245), .ZN(
        n10227) );
  INV_X1 U9735 ( .A(\CU_I/CW[DRAM_WE] ), .ZN(n10229) );
  NOR2_X1 U9736 ( .A1(n10142), .A2(n10144), .ZN(\CU_I/CW[DRAM_WE] ) );
  NAND2_X1 U9737 ( .A1(n10141), .A2(n10140), .ZN(n10144) );
  INV_X1 U9738 ( .A(n10296), .ZN(n10142) );
  AOI21_X1 U9739 ( .B1(n10141), .B2(n8477), .A(n10143), .ZN(n10296) );
  NAND4_X1 U9740 ( .A1(n8476), .A2(n8475), .A3(n8800), .A4(n8474), .ZN(n10143)
         );
  NOR2_X1 U9741 ( .A1(n8244), .A2(IR[31]), .ZN(n8473) );
  AOI21_X1 U9742 ( .B1(n10233), .B2(n10066), .A(n10303), .ZN(n8475) );
  INV_X1 U9743 ( .A(n10067), .ZN(n10233) );
  OR2_X1 U9744 ( .A1(n8496), .A2(n165), .ZN(n8476) );
  NOR2_X1 U9745 ( .A1(n10048), .A2(n8280), .ZN(n8477) );
  AOI21_X1 U9746 ( .B1(n10223), .B2(n10222), .A(n10231), .ZN(n10230) );
  OAI22_X1 U9747 ( .A1(n11838), .A2(n8209), .B1(n11839), .B2(n10112), .ZN(
        n7075) );
  INV_X1 U9748 ( .A(i_RD2[4]), .ZN(n10112) );
  AOI22_X1 U9749 ( .A1(n10104), .A2(n8205), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_IN1[15] ), .ZN(n2854) );
  AOI22_X1 U9750 ( .A1(n10104), .A2(n8100), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_IN1[12] ), .ZN(n2857) );
  AOI22_X1 U9751 ( .A1(n10104), .A2(n8099), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_IN1[11] ), .ZN(n2858) );
  INV_X1 U9752 ( .A(\CU_I/CW_ID[UNSIGNED_ID] ), .ZN(n10298) );
  AOI22_X1 U9753 ( .A1(n10089), .A2(n7753), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_IN2[7] ), .ZN(n2389) );
  OAI211_X1 U9754 ( .C1(n10056), .C2(n10243), .A(n10055), .B(n10054), .ZN(
        n7086) );
  AOI22_X1 U9755 ( .A1(n10053), .A2(n10052), .B1(i_ALU_OP[4]), .B2(n11626), 
        .ZN(n10054) );
  INV_X1 U9756 ( .A(n8244), .ZN(n10052) );
  INV_X1 U9757 ( .A(n10051), .ZN(n10055) );
  AOI22_X1 U9758 ( .A1(i_ADD_WS1[1]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_WRB1[1] ), .ZN(n2869) );
  OAI211_X1 U9759 ( .C1(n8105), .C2(n11828), .A(n10037), .B(n10036), .ZN(n7082) );
  OAI21_X1 U9760 ( .B1(n10218), .B2(n10035), .A(n10300), .ZN(n10036) );
  INV_X1 U9761 ( .A(n10066), .ZN(n10236) );
  NOR3_X1 U9762 ( .A1(n10066), .A2(n8115), .A3(n166), .ZN(n10218) );
  OAI211_X1 U9763 ( .C1(n7975), .C2(n10034), .A(n10040), .B(n11623), .ZN(
        n10037) );
  INV_X1 U9764 ( .A(n11622), .ZN(n10034) );
  AOI22_X1 U9765 ( .A1(i_ADD_WS1[3]), .A2(n7753), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_WRB1[3] ), .ZN(n2867) );
  AOI22_X1 U9766 ( .A1(i_ADD_WS1[4]), .A2(n7753), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_WRB1[4] ), .ZN(n2866) );
  OAI22_X1 U9767 ( .A1(n10121), .A2(n11839), .B1(n497), .B2(n11838), .ZN(n7021) );
  INV_X1 U9768 ( .A(n10120), .ZN(n10121) );
  OAI22_X1 U9769 ( .A1(n10131), .A2(n11839), .B1(n11838), .B2(n8204), .ZN(
        n7016) );
  INV_X1 U9770 ( .A(n10130), .ZN(n10131) );
  OAI222_X1 U9771 ( .A1(n10239), .A2(n11621), .B1(n11828), .B2(n8198), .C1(
        n8090), .C2(n11619), .ZN(n7084) );
  OR2_X1 U9772 ( .A1(n11830), .A2(n8800), .ZN(n11619) );
  NAND2_X1 U9773 ( .A1(n8472), .A2(n8471), .ZN(n8800) );
  NAND2_X1 U9774 ( .A1(n8795), .A2(n10066), .ZN(n8472) );
  OAI211_X1 U9775 ( .C1(n11828), .C2(n222), .A(n10071), .B(n10070), .ZN(n7085)
         );
  OAI22_X1 U9776 ( .A1(n172), .A2(n10067), .B1(n10066), .B2(n166), .ZN(n10068)
         );
  INV_X1 U9777 ( .A(n10065), .ZN(n10069) );
  OAI211_X1 U9778 ( .C1(n10064), .C2(n10063), .A(n8196), .B(n10062), .ZN(
        n10071) );
  INV_X1 U9779 ( .A(n11618), .ZN(n10062) );
  NOR2_X1 U9780 ( .A1(n11620), .A2(IR[4]), .ZN(n10064) );
  OAI22_X1 U9781 ( .A1(n10114), .A2(n11839), .B1(n11838), .B2(n8221), .ZN(
        n7024) );
  INV_X1 U9782 ( .A(n10113), .ZN(n10114) );
  OAI211_X1 U9783 ( .C1(n11828), .C2(n8095), .A(n10050), .B(n10049), .ZN(n7087) );
  AOI21_X1 U9784 ( .B1(n10053), .B2(n10048), .A(n10047), .ZN(n10049) );
  NOR3_X1 U9785 ( .A1(n11830), .A2(n10232), .A3(n10228), .ZN(n10047) );
  INV_X1 U9786 ( .A(n10060), .ZN(n10228) );
  INV_X1 U9787 ( .A(n10138), .ZN(n10048) );
  OAI21_X1 U9788 ( .B1(IR[1]), .B2(n10061), .A(n10046), .ZN(n10050) );
  AOI211_X1 U9789 ( .C1(n10045), .C2(IR[1]), .A(n8196), .B(n11620), .ZN(n10046) );
  OAI211_X1 U9790 ( .C1(n11838), .C2(n8211), .A(n10119), .B(n10118), .ZN(n7022) );
  NAND2_X1 U9791 ( .A1(n10117), .A2(n7753), .ZN(n10118) );
  NAND2_X1 U9792 ( .A1(n8238), .A2(n8242), .ZN(n11634) );
  OR2_X1 U9793 ( .A1(n8243), .A2(IR[31]), .ZN(n8238) );
  OAI22_X1 U9794 ( .A1(n10119), .A2(n8094), .B1(n8214), .B2(n11838), .ZN(n7118) );
  OAI22_X1 U9795 ( .A1(n10119), .A2(n8086), .B1(n8213), .B2(n11838), .ZN(n7119) );
  OAI22_X1 U9796 ( .A1(n10119), .A2(n8107), .B1(n8218), .B2(n11838), .ZN(n7113) );
  OAI22_X1 U9797 ( .A1(n10119), .A2(n8096), .B1(n8217), .B2(n11838), .ZN(n7114) );
  OAI22_X1 U9798 ( .A1(n10119), .A2(n7975), .B1(n8216), .B2(n11838), .ZN(n7115) );
  OAI22_X1 U9799 ( .A1(n10119), .A2(n8101), .B1(n8220), .B2(n11838), .ZN(n7111) );
  OAI22_X1 U9800 ( .A1(n10119), .A2(n8098), .B1(n8219), .B2(n11838), .ZN(n7112) );
  OAI22_X1 U9801 ( .A1(n10119), .A2(n8097), .B1(n8215), .B2(n11838), .ZN(n7116) );
  INV_X1 U9802 ( .A(n10056), .ZN(n10061) );
  NAND2_X1 U9803 ( .A1(n10040), .A2(IR[0]), .ZN(n11620) );
  AND2_X1 U9804 ( .A1(\C620/DATA2_2 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[2]) );
  INV_X1 U9805 ( .A(n10290), .ZN(n11694) );
  OAI211_X1 U9806 ( .C1(n10044), .C2(n10056), .A(n10242), .B(n10043), .ZN(
        n7089) );
  AOI21_X1 U9807 ( .B1(n11626), .B2(i_ALU_OP[1]), .A(n10053), .ZN(n10043) );
  NOR2_X1 U9808 ( .A1(n11830), .A2(n10220), .ZN(n10053) );
  NAND2_X1 U9809 ( .A1(n10039), .A2(IR[5]), .ZN(n10056) );
  OAI211_X1 U9810 ( .C1(n8086), .C2(n8094), .A(n10040), .B(IR[2]), .ZN(n10044)
         );
  OAI211_X1 U9811 ( .C1(n10244), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n7090) );
  AOI22_X1 U9812 ( .A1(n10300), .A2(n10291), .B1(i_ALU_OP[0]), .B2(n11626), 
        .ZN(n10241) );
  NOR2_X1 U9813 ( .A1(n10042), .A2(n8094), .ZN(n10063) );
  NAND2_X1 U9814 ( .A1(n10060), .A2(n10138), .ZN(n10217) );
  NOR2_X1 U9815 ( .A1(n10058), .A2(n10042), .ZN(n10051) );
  INV_X1 U9816 ( .A(n10040), .ZN(n10042) );
  NAND2_X1 U9817 ( .A1(n10240), .A2(n11622), .ZN(n10058) );
  NOR3_X1 U9818 ( .A1(n10045), .A2(n8196), .A3(n10239), .ZN(n10057) );
  NAND2_X1 U9819 ( .A1(n10039), .A2(n8096), .ZN(n10045) );
  NOR3_X1 U9820 ( .A1(n10038), .A2(IR[4]), .A3(IR[3]), .ZN(n10039) );
  INV_X1 U9821 ( .A(n11617), .ZN(n10038) );
  NAND2_X1 U9822 ( .A1(n10040), .A2(n8086), .ZN(n10239) );
  NOR2_X1 U9823 ( .A1(n11830), .A2(n10098), .ZN(n10040) );
  INV_X1 U9824 ( .A(n10240), .ZN(n10244) );
  AOI22_X1 U9825 ( .A1(n10090), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[5] ), .ZN(n2392) );
  AOI22_X1 U9826 ( .A1(i_ADD_WS1[0]), .A2(n8423), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_WRB1[0] ), .ZN(n2870) );
  AOI22_X1 U9827 ( .A1(n10087), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[11] ), .ZN(n2383) );
  AOI22_X1 U9828 ( .A1(n10086), .A2(n7753), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_IN2[16] ), .ZN(n2377) );
  AOI22_X1 U9829 ( .A1(n10104), .A2(n8134), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN1[14] ), .ZN(n2855) );
  AOI22_X1 U9830 ( .A1(i_ADD_WS1[2]), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_WRB1[2] ), .ZN(n2868) );
  AOI22_X1 U9831 ( .A1(n10080), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[23] ), .ZN(n2362) );
  AOI22_X1 U9832 ( .A1(n10078), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[25] ), .ZN(n2358) );
  AOI22_X1 U9833 ( .A1(n10079), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[24] ), .ZN(n2360) );
  AOI22_X1 U9834 ( .A1(n10084), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[18] ), .ZN(n2373) );
  AOI22_X1 U9835 ( .A1(n10072), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[31] ), .ZN(n2346) );
  AOI22_X1 U9836 ( .A1(n10081), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[22] ), .ZN(n2364) );
  AOI22_X1 U9837 ( .A1(n10073), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[30] ), .ZN(n2348) );
  AOI22_X1 U9838 ( .A1(n10074), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[29] ), .ZN(n2350) );
  AOI22_X1 U9839 ( .A1(n10088), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[9] ), .ZN(n2386) );
  AOI22_X1 U9840 ( .A1(n10075), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[28] ), .ZN(n2352) );
  AOI22_X1 U9841 ( .A1(n10076), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[27] ), .ZN(n2354) );
  AOI22_X1 U9842 ( .A1(n10085), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[17] ), .ZN(n2375) );
  AOI22_X1 U9843 ( .A1(n10077), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[26] ), .ZN(n2356) );
  AOI22_X1 U9844 ( .A1(n10083), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[19] ), .ZN(n2371) );
  AOI22_X1 U9845 ( .A1(n10082), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[21] ), .ZN(n2366) );
  AOI22_X1 U9846 ( .A1(n10104), .A2(IR[8]), .B1(\DataPath/i_PIPLIN_IN1[8] ), 
        .B2(n8425), .ZN(n2861) );
  AOI22_X1 U9847 ( .A1(n10104), .A2(IR[13]), .B1(\DataPath/i_PIPLIN_IN1[13] ), 
        .B2(n8425), .ZN(n2856) );
  AOI22_X1 U9848 ( .A1(n10104), .A2(IR[10]), .B1(\DataPath/i_PIPLIN_IN1[10] ), 
        .B2(n8425), .ZN(n2859) );
  AND2_X1 U9849 ( .A1(\C620/DATA2_3 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[3]) );
  INV_X1 U9850 ( .A(n10133), .ZN(n7015) );
  AOI22_X1 U9851 ( .A1(n10132), .A2(n7753), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_IN2[15] ), .ZN(n10133) );
  INV_X1 U9852 ( .A(n10135), .ZN(n7014) );
  AOI22_X1 U9853 ( .A1(n10134), .A2(n8424), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_IN2[20] ), .ZN(n10135) );
  INV_X1 U9854 ( .A(n10125), .ZN(n7019) );
  AOI22_X1 U9855 ( .A1(n10124), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[10] ), .ZN(n10125) );
  INV_X1 U9856 ( .A(n10123), .ZN(n7020) );
  AOI22_X1 U9857 ( .A1(n10122), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[8] ), .ZN(n10123) );
  INV_X1 U9858 ( .A(n10116), .ZN(n7023) );
  AOI22_X1 U9859 ( .A1(n10115), .A2(n8424), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[3] ), .ZN(n10116) );
  INV_X1 U9860 ( .A(n10127), .ZN(n7018) );
  AOI22_X1 U9861 ( .A1(n10126), .A2(n8422), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[12] ), .ZN(n10127) );
  INV_X1 U9862 ( .A(n10129), .ZN(n7017) );
  AOI22_X1 U9863 ( .A1(n10128), .A2(n8423), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[13] ), .ZN(n10129) );
  INV_X1 U9864 ( .A(n10111), .ZN(n7117) );
  AOI22_X1 U9865 ( .A1(n10110), .A2(n7753), .B1(\DataPath/i_PIPLIN_IN1[2] ), 
        .B2(n8425), .ZN(n10111) );
  OAI21_X1 U9866 ( .B1(n10109), .B2(n8196), .A(n10108), .ZN(n10110) );
  INV_X1 U9867 ( .A(n10291), .ZN(n10109) );
  AND2_X1 U9868 ( .A1(\C620/DATA2_4 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[4]) );
  AND2_X1 U9869 ( .A1(\C620/DATA2_5 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[5]) );
  AND2_X1 U9870 ( .A1(\C620/DATA2_6 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[6]) );
  AND2_X1 U9871 ( .A1(\C620/DATA2_7 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[7]) );
  OAI22_X1 U9872 ( .A1(n10093), .A2(n11839), .B1(n8197), .B2(n11838), .ZN(n102) );
  AND2_X1 U9873 ( .A1(\C620/DATA2_8 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[8]) );
  OAI21_X1 U9874 ( .B1(n506), .B2(n11838), .A(n10107), .ZN(n7120) );
  AND2_X1 U9875 ( .A1(\C620/DATA2_9 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[9]) );
  OAI211_X1 U9876 ( .C1(n9136), .C2(n9135), .A(n9134), .B(n9133), .ZN(n11709)
         );
  NAND2_X1 U9877 ( .A1(\DataPath/ALUhw/i_Q_EXTENDED[38] ), .A2(n8337), .ZN(
        n9134) );
  INV_X1 U9878 ( .A(n9810), .ZN(n9135) );
  NAND2_X1 U9879 ( .A1(n9128), .A2(n9127), .ZN(n9150) );
  INV_X1 U9880 ( .A(n9153), .ZN(n9128) );
  NAND2_X1 U9881 ( .A1(n9149), .A2(n9148), .ZN(n11713) );
  INV_X1 U9882 ( .A(n9155), .ZN(n9149) );
  AOI222_X1 U9883 ( .A1(n11719), .A2(n10023), .B1(n9920), .B2(n10284), .C1(
        n9923), .C2(n10013), .ZN(n11704) );
  AOI22_X1 U9884 ( .A1(n9946), .A2(n10286), .B1(n9978), .B2(n9979), .ZN(n11705) );
  AOI22_X1 U9885 ( .A1(n9947), .A2(n10011), .B1(n10020), .B2(n9176), .ZN(
        n11706) );
  AOI22_X1 U9886 ( .A1(n9922), .A2(n10021), .B1(n10010), .B2(n9211), .ZN(
        n11707) );
  NOR2_X1 U9887 ( .A1(n9909), .A2(n9912), .ZN(n9914) );
  NAND2_X1 U9888 ( .A1(n9091), .A2(n9093), .ZN(n11695) );
  AND2_X1 U9889 ( .A1(n9915), .A2(n9090), .ZN(n10282) );
  NAND2_X1 U9890 ( .A1(n9089), .A2(n9090), .ZN(n9909) );
  OAI211_X1 U9891 ( .C1(n9063), .C2(n7970), .A(n9061), .B(n9060), .ZN(n11691)
         );
  OAI211_X1 U9892 ( .C1(n9803), .C2(n9072), .A(n8315), .B(n7970), .ZN(n9060)
         );
  INV_X1 U9893 ( .A(n11696), .ZN(n9072) );
  NAND2_X1 U9894 ( .A1(n9958), .A2(n8084), .ZN(n11696) );
  NAND2_X1 U9895 ( .A1(n9059), .A2(n10287), .ZN(n9061) );
  NAND4_X1 U9896 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), .ZN(n9059)
         );
  AOI22_X1 U9897 ( .A1(n9925), .A2(n10284), .B1(n11698), .B2(n10010), .ZN(
        n9055) );
  OAI211_X1 U9898 ( .C1(n8311), .C2(n9049), .A(n9048), .B(n9047), .ZN(n9925)
         );
  AOI22_X1 U9899 ( .A1(n9046), .A2(n10283), .B1(n9045), .B2(n9195), .ZN(n9047)
         );
  OAI21_X1 U9900 ( .B1(n9538), .B2(n11681), .A(n9670), .ZN(n9046) );
  AOI21_X1 U9901 ( .B1(n9043), .B2(n9194), .A(n9042), .ZN(n9048) );
  OAI22_X1 U9902 ( .A1(n9630), .A2(n9041), .B1(n9317), .B2(n9547), .ZN(n9042)
         );
  INV_X1 U9903 ( .A(n9078), .ZN(n9041) );
  AOI22_X1 U9904 ( .A1(n9079), .A2(n10021), .B1(n10023), .B2(n9923), .ZN(n9056) );
  INV_X1 U9905 ( .A(n9798), .ZN(n9923) );
  INV_X1 U9906 ( .A(n9919), .ZN(n9079) );
  NOR3_X1 U9907 ( .A1(n9014), .A2(n9013), .A3(n9012), .ZN(n9919) );
  OAI22_X1 U9908 ( .A1(n9011), .A2(n9081), .B1(n7942), .B2(n9474), .ZN(n9012)
         );
  AOI21_X1 U9909 ( .B1(n9010), .B2(n9281), .A(n8305), .ZN(n9013) );
  OAI21_X1 U9910 ( .B1(n9477), .B2(n9019), .A(n9009), .ZN(n9014) );
  AOI22_X1 U9911 ( .A1(n9025), .A2(n9476), .B1(n9683), .B2(n9084), .ZN(n9009)
         );
  AOI21_X1 U9912 ( .B1(n7759), .B2(n9924), .A(n9004), .ZN(n9057) );
  OAI22_X1 U9913 ( .A1(n9003), .A2(n9939), .B1(n9917), .B2(n10017), .ZN(n9004)
         );
  INV_X1 U9914 ( .A(n9176), .ZN(n9917) );
  AOI211_X1 U9915 ( .C1(n9170), .C2(n9043), .A(n8987), .B(n8986), .ZN(n9003)
         );
  OAI211_X1 U9916 ( .C1(n9011), .C2(n9167), .A(n8985), .B(n8984), .ZN(n8986)
         );
  NAND2_X1 U9917 ( .A1(n9028), .A2(n8991), .ZN(n8984) );
  OAI21_X1 U9918 ( .B1(n7774), .B2(n9559), .A(n9683), .ZN(n8985) );
  OAI22_X1 U9919 ( .A1(n9538), .A2(n9557), .B1(n9527), .B2(n9670), .ZN(n8987)
         );
  AOI22_X1 U9920 ( .A1(n9921), .A2(n10020), .B1(n9978), .B2(n9920), .ZN(n9058)
         );
  INV_X1 U9921 ( .A(n8981), .ZN(n9049) );
  AOI21_X1 U9922 ( .B1(n8315), .B2(n9990), .A(n8961), .ZN(n9063) );
  AOI21_X1 U9923 ( .B1(n9850), .B2(n9935), .A(n9910), .ZN(n8961) );
  OAI211_X1 U9924 ( .C1(n9916), .C2(n9912), .A(n8945), .B(n8944), .ZN(n11692)
         );
  AOI21_X1 U9925 ( .B1(\DataPath/ALUhw/MULT/mux_out[0][0] ), .B2(n9992), .A(
        i_SEL_ALU_SETCMP), .ZN(n8944) );
  NAND2_X1 U9926 ( .A1(\DataPath/ALUhw/i_Q_EXTENDED[32] ), .A2(n8337), .ZN(
        n8945) );
  NAND2_X1 U9927 ( .A1(n9911), .A2(n8315), .ZN(n9912) );
  INV_X1 U9928 ( .A(n10288), .ZN(n9916) );
  AND2_X1 U9929 ( .A1(n9958), .A2(n8452), .ZN(n10288) );
  AND2_X1 U9930 ( .A1(\C620/DATA2_10 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[10])
         );
  AOI211_X1 U9931 ( .C1(\DataPath/ALUhw/i_Q_EXTENDED[40] ), .C2(n10004), .A(
        n9189), .B(n9188), .ZN(n11714) );
  OAI21_X1 U9932 ( .B1(n9187), .B2(n9815), .A(n9186), .ZN(n9188) );
  NOR3_X1 U9933 ( .A1(n9181), .A2(n9180), .A3(n9179), .ZN(n9187) );
  OAI211_X1 U9934 ( .C1(n9983), .C2(n9878), .A(n9178), .B(n9177), .ZN(n9179)
         );
  AOI22_X1 U9935 ( .A1(n9211), .A2(n10020), .B1(n10013), .B2(n9176), .ZN(n9177) );
  AOI22_X1 U9936 ( .A1(n11719), .A2(n10010), .B1(n9977), .B2(n10286), .ZN(
        n9178) );
  OAI22_X1 U9937 ( .A1(n9791), .A2(n9860), .B1(n9940), .B2(n9982), .ZN(n9180)
         );
  OAI22_X1 U9938 ( .A1(n9788), .A2(n10027), .B1(n9787), .B2(n9942), .ZN(n9181)
         );
  AOI211_X1 U9939 ( .C1(n9928), .C2(n9166), .A(n9935), .B(n9165), .ZN(n9189)
         );
  NOR3_X1 U9940 ( .A1(n9928), .A2(n9926), .A3(n9164), .ZN(n9165) );
  INV_X1 U9941 ( .A(n9927), .ZN(n9164) );
  XNOR2_X1 U9942 ( .A(n9162), .B(n9161), .ZN(n9166) );
  OAI21_X1 U9943 ( .B1(n9957), .B2(n10032), .A(n9956), .ZN(n7007) );
  AOI21_X1 U9944 ( .B1(n10280), .B2(n9955), .A(n9954), .ZN(n9956) );
  OAI22_X1 U9945 ( .A1(n9953), .A2(n9952), .B1(n8206), .B2(n11734), .ZN(n9954)
         );
  INV_X1 U9946 ( .A(n10007), .ZN(n9953) );
  AOI22_X1 U9947 ( .A1(n9947), .A2(n10020), .B1(n10010), .B2(n9979), .ZN(n9948) );
  AOI211_X1 U9948 ( .C1(n7759), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9949)
         );
  OAI22_X1 U9949 ( .A1(n9943), .A2(n9942), .B1(n9941), .B2(n10027), .ZN(n9944)
         );
  OAI22_X1 U9950 ( .A1(n9940), .A2(n9939), .B1(n9938), .B2(n9982), .ZN(n9945)
         );
  INV_X1 U9951 ( .A(n9211), .ZN(n9938) );
  INV_X1 U9952 ( .A(n9983), .ZN(n9946) );
  AOI22_X1 U9953 ( .A1(n9974), .A2(n10023), .B1(n10286), .B2(n10014), .ZN(
        n9950) );
  AOI21_X1 U9954 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[41] ), .B2(n8337), .A(
        n9937), .ZN(n9957) );
  OAI211_X1 U9955 ( .C1(n9936), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9937)
         );
  XNOR2_X1 U9956 ( .A(n9931), .B(n9930), .ZN(n9936) );
  XNOR2_X1 U9957 ( .A(n9929), .B(n9951), .ZN(n9930) );
  AOI21_X1 U9958 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(n9931) );
  OAI22_X1 U9959 ( .A1(n9818), .A2(n11735), .B1(n509), .B2(n11734), .ZN(n7011)
         );
  AOI21_X1 U9960 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[36] ), .B2(n8337), .A(
        n9817), .ZN(n9818) );
  OAI211_X1 U9961 ( .C1(n9816), .C2(n9815), .A(n9814), .B(n9813), .ZN(n9817)
         );
  OAI21_X1 U9962 ( .B1(n9812), .B2(n9811), .A(n9810), .ZN(n9813) );
  NOR2_X1 U9963 ( .A1(n9098), .A2(n9935), .ZN(n9810) );
  INV_X1 U9964 ( .A(n9154), .ZN(n9098) );
  INV_X1 U9965 ( .A(n9809), .ZN(n9812) );
  AOI21_X1 U9966 ( .B1(n10278), .B2(n9805), .A(n9804), .ZN(n9807) );
  AOI21_X1 U9967 ( .B1(n10278), .B2(n9801), .A(n9800), .ZN(n9808) );
  NOR2_X1 U9968 ( .A1(n9154), .A2(n9935), .ZN(n10278) );
  AOI211_X1 U9969 ( .C1(n10021), .C2(n9920), .A(n11703), .B(n9799), .ZN(n9816)
         );
  NOR2_X1 U9970 ( .A1(n9798), .A2(n9918), .ZN(n9799) );
  NOR2_X1 U9971 ( .A1(n9037), .A2(n9036), .ZN(n9798) );
  NAND4_X1 U9972 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(n9036)
         );
  NAND2_X1 U9973 ( .A1(n9031), .A2(n9631), .ZN(n9032) );
  OAI21_X1 U9974 ( .B1(n11723), .B2(n9627), .A(n9683), .ZN(n9033) );
  AOI22_X1 U9975 ( .A1(n9028), .A2(n9129), .B1(n9687), .B2(n9027), .ZN(n9034)
         );
  INV_X1 U9976 ( .A(n9391), .ZN(n9027) );
  INV_X1 U9977 ( .A(n9281), .ZN(n9028) );
  AOI22_X1 U9978 ( .A1(n9025), .A2(n9390), .B1(n9024), .B2(n9023), .ZN(n9035)
         );
  INV_X1 U9979 ( .A(n9634), .ZN(n9023) );
  OAI22_X1 U9980 ( .A1(n9019), .A2(n9290), .B1(n7705), .B2(n9018), .ZN(n9037)
         );
  NAND2_X1 U9981 ( .A1(n10013), .A2(n11698), .ZN(n11699) );
  NAND4_X1 U9982 ( .A1(n8955), .A2(n8954), .A3(n8953), .A4(n8952), .ZN(n11698)
         );
  OAI21_X1 U9983 ( .B1(n9087), .B2(n9685), .A(n9683), .ZN(n8952) );
  AOI22_X1 U9984 ( .A1(n9099), .A2(n8981), .B1(n8980), .B2(n9689), .ZN(n8953)
         );
  AOI22_X1 U9985 ( .A1(n9025), .A2(n9682), .B1(n9024), .B2(n9680), .ZN(n8954)
         );
  NAND2_X1 U9986 ( .A1(n9043), .A2(n9684), .ZN(n8955) );
  AOI22_X1 U9987 ( .A1(n10010), .A2(n9176), .B1(n10284), .B2(n9924), .ZN(
        n11700) );
  OR2_X1 U9988 ( .A1(n9031), .A2(n9687), .ZN(n8980) );
  NOR2_X1 U9989 ( .A1(n9670), .A2(i_ALU_OP[2]), .ZN(n9031) );
  NAND2_X1 U9990 ( .A1(n9018), .A2(n9281), .ZN(n8981) );
  INV_X1 U9991 ( .A(n9547), .ZN(n9025) );
  NAND4_X1 U9992 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(n9176)
         );
  OAI21_X1 U9993 ( .B1(n8997), .B2(n9559), .A(n9691), .ZN(n8998) );
  NOR2_X1 U9994 ( .A1(n9250), .A2(n9667), .ZN(n8997) );
  NAND2_X1 U9995 ( .A1(n8996), .A2(n8325), .ZN(n8999) );
  INV_X1 U9996 ( .A(n9305), .ZN(n8996) );
  OAI21_X1 U9997 ( .B1(n9564), .B2(n8085), .A(n9667), .ZN(n8993) );
  NAND2_X1 U9998 ( .A1(n9527), .A2(n11731), .ZN(n8990) );
  AOI22_X1 U9999 ( .A1(n10023), .A2(n9211), .B1(n7759), .B2(n9922), .ZN(n11701) );
  INV_X1 U10000 ( .A(n9940), .ZN(n9922) );
  NAND2_X1 U10001 ( .A1(n9548), .A2(n9039), .ZN(n9078) );
  NAND2_X1 U10002 ( .A1(n8979), .A2(n9991), .ZN(n9039) );
  AOI22_X1 U10003 ( .A1(n10286), .A2(n11719), .B1(n9978), .B2(n9947), .ZN(
        n11702) );
  INV_X1 U10004 ( .A(n9787), .ZN(n9947) );
  INV_X1 U10005 ( .A(n9019), .ZN(n9043) );
  OR2_X1 U10006 ( .A1(n9137), .A2(n8085), .ZN(n9019) );
  NAND2_X1 U10007 ( .A1(n9681), .A2(n8452), .ZN(n9018) );
  NAND2_X1 U10008 ( .A1(n8970), .A2(n9011), .ZN(n9045) );
  INV_X1 U10009 ( .A(n9024), .ZN(n9011) );
  NOR2_X1 U10010 ( .A1(n9593), .A2(n8948), .ZN(n9024) );
  NOR2_X1 U10011 ( .A1(n8084), .A2(i_ALU_OP[4]), .ZN(n8948) );
  NAND2_X1 U10012 ( .A1(n9687), .A2(n11718), .ZN(n8970) );
  AND2_X1 U10013 ( .A1(\C620/DATA2_11 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[11])
         );
  AOI21_X1 U10014 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[42] ), .B2(n8337), .A(
        n9219), .ZN(n11715) );
  OAI211_X1 U10015 ( .C1(n9218), .C2(n9935), .A(n9217), .B(n9216), .ZN(n9219)
         );
  OAI21_X1 U10016 ( .B1(n9215), .B2(n9214), .A(n10287), .ZN(n9216) );
  OAI211_X1 U10017 ( .C1(n9983), .C2(n9880), .A(n9213), .B(n9212), .ZN(n9214)
         );
  AOI22_X1 U10018 ( .A1(n9979), .A2(n10021), .B1(n9211), .B2(n10013), .ZN(
        n9212) );
  AOI22_X1 U10019 ( .A1(n11719), .A2(n10020), .B1(n9977), .B2(n10023), .ZN(
        n9213) );
  OAI211_X1 U10020 ( .C1(n9787), .C2(n9982), .A(n9210), .B(n9209), .ZN(n9215)
         );
  AOI22_X1 U10021 ( .A1(n10014), .A2(n9978), .B1(n10286), .B2(n10019), .ZN(
        n9209) );
  NAND2_X1 U10022 ( .A1(n9974), .A2(n7759), .ZN(n9210) );
  XNOR2_X1 U10023 ( .A(n9234), .B(n9190), .ZN(n9218) );
  XNOR2_X1 U10024 ( .A(n9231), .B(n9230), .ZN(n9190) );
  AND2_X1 U10025 ( .A1(\C620/DATA2_12 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[12])
         );
  INV_X1 U10026 ( .A(n9979), .ZN(n9791) );
  NAND2_X1 U10027 ( .A1(n9479), .A2(n9008), .ZN(n9084) );
  NAND2_X1 U10028 ( .A1(n8979), .A2(n9711), .ZN(n9008) );
  INV_X1 U10029 ( .A(n9225), .ZN(n9081) );
  NAND2_X1 U10030 ( .A1(n10258), .A2(IRAM_DATA[9]), .ZN(n11600) );
  NAND2_X1 U10031 ( .A1(n10258), .A2(IRAM_DATA[2]), .ZN(n11852) );
  NAND2_X1 U10032 ( .A1(n10258), .A2(IRAM_DATA[6]), .ZN(n11851) );
  NAND2_X1 U10033 ( .A1(n10258), .A2(IRAM_DATA[25]), .ZN(n11612) );
  NAND2_X1 U10034 ( .A1(n10258), .A2(IRAM_DATA[14]), .ZN(n11601) );
  NAND2_X1 U10035 ( .A1(n10258), .A2(IRAM_DATA[23]), .ZN(n11610) );
  NAND2_X1 U10036 ( .A1(n10258), .A2(IRAM_DATA[24]), .ZN(n11611) );
  AOI22_X1 U10037 ( .A1(n10258), .A2(IRAM_DATA[31]), .B1(IR[31]), .B2(n10257), 
        .ZN(n10256) );
  OAI21_X1 U10038 ( .B1(n8294), .B2(n8097), .A(n10253), .ZN(n37) );
  NAND2_X1 U10039 ( .A1(n10258), .A2(IRAM_DATA[3]), .ZN(n10253) );
  INV_X1 U10040 ( .A(n11719), .ZN(n9943) );
  NOR2_X1 U10041 ( .A1(n9007), .A2(n8301), .ZN(n9087) );
  OR2_X1 U10042 ( .A1(n8452), .A2(n11681), .ZN(n9007) );
  AND2_X1 U10043 ( .A1(\C620/DATA2_13 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[13])
         );
  AOI211_X1 U10044 ( .C1(n8177), .C2(n10102), .A(n10094), .B(n8296), .ZN(
        n10095) );
  AOI211_X1 U10045 ( .C1(n8184), .C2(n10102), .A(n10096), .B(n8297), .ZN(
        n10097) );
  AOI22_X1 U10046 ( .A1(n10246), .A2(n8099), .B1(n10245), .B2(n8176), .ZN(
        n10247) );
  AOI211_X1 U10047 ( .C1(n8179), .C2(n10102), .A(n10100), .B(n8295), .ZN(
        n10101) );
  AOI22_X1 U10048 ( .A1(n10246), .A2(n8100), .B1(n10245), .B2(n8175), .ZN(
        n10103) );
  INV_X1 U10049 ( .A(n10102), .ZN(n10249) );
  OAI211_X1 U10050 ( .C1(n9988), .C2(n10032), .A(n9987), .B(n9986), .ZN(n7003)
         );
  OAI21_X1 U10051 ( .B1(n9985), .B2(n9984), .A(n10280), .ZN(n9986) );
  OAI211_X1 U10052 ( .C1(n9983), .C2(n9982), .A(n9981), .B(n9980), .ZN(n9984)
         );
  AOI22_X1 U10053 ( .A1(n9979), .A2(n10013), .B1(n10022), .B2(n9978), .ZN(
        n9980) );
  OAI211_X1 U10054 ( .C1(n9140), .C2(n9666), .A(n8161), .B(n9110), .ZN(n9979)
         );
  OR2_X1 U10055 ( .A1(n9633), .A2(n9671), .ZN(n9110) );
  NAND2_X1 U10056 ( .A1(n9408), .A2(n8325), .ZN(n9106) );
  OR2_X1 U10057 ( .A1(n9593), .A2(n9104), .ZN(n9107) );
  NAND2_X1 U10058 ( .A1(n8979), .A2(n9889), .ZN(n9104) );
  NAND2_X1 U10059 ( .A1(n9687), .A2(n9415), .ZN(n9108) );
  NAND2_X1 U10060 ( .A1(n9103), .A2(n9686), .ZN(n9109) );
  OAI21_X1 U10061 ( .B1(n9669), .B2(n9102), .A(n9101), .ZN(n9103) );
  INV_X1 U10062 ( .A(n9674), .ZN(n9101) );
  AOI22_X1 U10063 ( .A1(n11721), .A2(n10023), .B1(n10021), .B2(n9977), .ZN(
        n9981) );
  NAND2_X1 U10064 ( .A1(n9976), .A2(n9975), .ZN(n9985) );
  AOI22_X1 U10065 ( .A1(n10019), .A2(n10011), .B1(n10009), .B2(n10286), .ZN(
        n9975) );
  AOI22_X1 U10066 ( .A1(n9974), .A2(n10020), .B1(n10010), .B2(n10014), .ZN(
        n9976) );
  AOI22_X1 U10067 ( .A1(n10007), .A2(n9973), .B1(n7764), .B2(DRAM_ADDRESS[13]), 
        .ZN(n9987) );
  XNOR2_X1 U10068 ( .A(\DP_OP_751_130_6421/n1209 ), .B(n9972), .ZN(n9973) );
  AOI21_X1 U10069 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[45] ), .B2(n8337), .A(
        n9971), .ZN(n9988) );
  OAI211_X1 U10070 ( .C1(n9970), .C2(n9969), .A(n9968), .B(n9967), .ZN(n9971)
         );
  AOI211_X1 U10071 ( .C1(n9965), .C2(n9964), .A(n9963), .B(n9962), .ZN(n9969)
         );
  INV_X1 U10072 ( .A(n9961), .ZN(n9962) );
  OAI211_X1 U10073 ( .C1(n9961), .C2(n9960), .A(n9959), .B(n9958), .ZN(n9970)
         );
  INV_X1 U10074 ( .A(n9963), .ZN(n9960) );
  AOI22_X1 U10075 ( .A1(n8299), .A2(n11615), .B1(n165), .B2(n10257), .ZN(n7122) );
  AOI22_X1 U10076 ( .A1(n8299), .A2(n11613), .B1(n172), .B2(n10257), .ZN(n7126) );
  NAND2_X1 U10077 ( .A1(n8299), .A2(IRAM_DATA[19]), .ZN(n11606) );
  OAI21_X1 U10078 ( .B1(n10292), .B2(n7975), .A(n10252), .ZN(n38) );
  NAND2_X1 U10079 ( .A1(n8299), .A2(IRAM_DATA[4]), .ZN(n10252) );
  AOI22_X1 U10080 ( .A1(n8299), .A2(IRAM_DATA[8]), .B1(IR[8]), .B2(n10257), 
        .ZN(n2890) );
  AOI22_X1 U10081 ( .A1(n8299), .A2(IRAM_DATA[13]), .B1(IR[13]), .B2(n10257), 
        .ZN(n2886) );
  AOI22_X1 U10082 ( .A1(n8299), .A2(IRAM_DATA[10]), .B1(IR[10]), .B2(n10257), 
        .ZN(n2889) );
  OAI21_X1 U10083 ( .B1(n8294), .B2(n8094), .A(n10254), .ZN(n35) );
  NAND2_X1 U10084 ( .A1(n8299), .A2(IRAM_DATA[1]), .ZN(n10254) );
  AND2_X1 U10085 ( .A1(\C620/DATA2_14 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[14])
         );
  NAND2_X1 U10086 ( .A1(n8299), .A2(IRAM_DATA[15]), .ZN(n11602) );
  NAND2_X1 U10087 ( .A1(n8299), .A2(IRAM_DATA[16]), .ZN(n11603) );
  NAND2_X1 U10088 ( .A1(n8299), .A2(IRAM_DATA[17]), .ZN(n11604) );
  NAND2_X1 U10089 ( .A1(n8299), .A2(IRAM_DATA[20]), .ZN(n11607) );
  NAND2_X1 U10090 ( .A1(n8299), .A2(IRAM_DATA[12]), .ZN(n11849) );
  NAND2_X1 U10091 ( .A1(n8299), .A2(IRAM_DATA[21]), .ZN(n11608) );
  NAND2_X1 U10092 ( .A1(n8299), .A2(IRAM_DATA[22]), .ZN(n11609) );
  NAND2_X1 U10093 ( .A1(n8299), .A2(IRAM_DATA[11]), .ZN(n11850) );
  NAND2_X1 U10094 ( .A1(n8299), .A2(IRAM_DATA[18]), .ZN(n11605) );
  INV_X1 U10095 ( .A(n9788), .ZN(n9974) );
  NOR2_X1 U10096 ( .A1(n9120), .A2(n9119), .ZN(n9983) );
  OAI22_X1 U10097 ( .A1(n9140), .A2(n9118), .B1(n9139), .B2(n9629), .ZN(n9119)
         );
  INV_X1 U10098 ( .A(n9627), .ZN(n9118) );
  OR2_X1 U10099 ( .A1(n9633), .A2(n9290), .ZN(n9115) );
  AOI22_X1 U10100 ( .A1(n9420), .A2(n11723), .B1(n8325), .B2(n9114), .ZN(n9116) );
  INV_X1 U10101 ( .A(n9389), .ZN(n9114) );
  OAI22_X1 U10102 ( .A1(n9111), .A2(n9683), .B1(n9631), .B2(n9667), .ZN(n9117)
         );
  NOR3_X1 U10103 ( .A1(n9589), .A2(n9634), .A3(n8085), .ZN(n9111) );
  OAI21_X1 U10104 ( .B1(n10292), .B2(n8096), .A(n10251), .ZN(n39) );
  NAND2_X1 U10105 ( .A1(n8299), .A2(IRAM_DATA[5]), .ZN(n10251) );
  OAI21_X1 U10106 ( .B1(n8294), .B2(n8086), .A(n10255), .ZN(n34) );
  NAND2_X1 U10107 ( .A1(n8299), .A2(IRAM_DATA[0]), .ZN(n10255) );
  OAI21_X1 U10108 ( .B1(n8294), .B2(n8098), .A(n10250), .ZN(n41) );
  NAND2_X1 U10109 ( .A1(n8299), .A2(IRAM_DATA[7]), .ZN(n10250) );
  AND2_X1 U10110 ( .A1(\C620/DATA2_15 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[15])
         );
  OAI22_X1 U10111 ( .A1(n7937), .A2(n9343), .B1(n9593), .B2(n9143), .ZN(n9144)
         );
  NAND2_X1 U10112 ( .A1(n8979), .A2(n9607), .ZN(n9143) );
  NOR2_X1 U10113 ( .A1(i_ALU_OP[2]), .A2(n11681), .ZN(n8979) );
  NOR2_X1 U10114 ( .A1(n9633), .A2(n9336), .ZN(n9145) );
  OAI22_X1 U10115 ( .A1(n9140), .A2(n9590), .B1(n9139), .B2(n9138), .ZN(n9146)
         );
  INV_X1 U10116 ( .A(n9591), .ZN(n9138) );
  NAND2_X1 U10117 ( .A1(n9687), .A2(n11731), .ZN(n9139) );
  NOR2_X1 U10118 ( .A1(n9687), .A2(n9691), .ZN(n9140) );
  OAI22_X1 U10119 ( .A1(n9630), .A2(n9592), .B1(n9137), .B2(n9595), .ZN(n9147)
         );
  NAND2_X1 U10120 ( .A1(n9686), .A2(n11718), .ZN(n9137) );
  INV_X1 U10121 ( .A(n9977), .ZN(n9941) );
  NOR2_X1 U10122 ( .A1(n9773), .A2(n9935), .ZN(n9785) );
  NAND2_X1 U10123 ( .A1(n9773), .A2(n9958), .ZN(n9786) );
  INV_X1 U10124 ( .A(n9965), .ZN(n9773) );
  NAND2_X1 U10125 ( .A1(n9770), .A2(n9769), .ZN(n9778) );
  OAI21_X1 U10126 ( .B1(n9961), .B2(n9964), .A(n9768), .ZN(n9777) );
  INV_X1 U10127 ( .A(n9781), .ZN(n9964) );
  AND2_X1 U10128 ( .A1(\C620/DATA2_16 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[16])
         );
  OAI222_X1 U10129 ( .A1(n11735), .A2(n9767), .B1(n11730), .B2(n9766), .C1(
        n11734), .C2(n517), .ZN(n7000) );
  NOR3_X1 U10130 ( .A1(n9765), .A2(n9764), .A3(n9763), .ZN(n9766) );
  OAI22_X1 U10131 ( .A1(n9789), .A2(n9918), .B1(n9881), .B2(n9860), .ZN(n9763)
         );
  OAI22_X1 U10132 ( .A1(n10008), .A2(n9878), .B1(n9790), .B2(n9982), .ZN(n9764) );
  INV_X1 U10133 ( .A(n10014), .ZN(n9790) );
  OAI211_X1 U10134 ( .C1(n8121), .C2(n10017), .A(n9762), .B(n9761), .ZN(n9765)
         );
  AOI22_X1 U10135 ( .A1(n10024), .A2(n9978), .B1(n10022), .B2(n10010), .ZN(
        n9761) );
  AOI22_X1 U10136 ( .A1(n11721), .A2(n10021), .B1(n10013), .B2(n9977), .ZN(
        n9762) );
  NAND4_X1 U10137 ( .A1(n9175), .A2(n9174), .A3(n9173), .A4(n9172), .ZN(n9977)
         );
  NAND2_X1 U10138 ( .A1(n9171), .A2(n9554), .ZN(n9172) );
  OAI21_X1 U10139 ( .B1(n9527), .B2(n9593), .A(n9220), .ZN(n9171) );
  NAND2_X1 U10140 ( .A1(n8325), .A2(n9170), .ZN(n9173) );
  INV_X1 U10141 ( .A(n9564), .ZN(n9170) );
  OAI211_X1 U10142 ( .C1(n11731), .C2(n9559), .A(n9686), .B(n9169), .ZN(n9174)
         );
  OR2_X1 U10143 ( .A1(n9562), .A2(n11733), .ZN(n9169) );
  OAI21_X1 U10144 ( .B1(n9167), .B2(n8085), .A(n9667), .ZN(n9168) );
  AOI211_X1 U10145 ( .C1(\DataPath/ALUhw/i_Q_EXTENDED[48] ), .C2(n8337), .A(
        n9760), .B(n9759), .ZN(n9767) );
  OAI211_X1 U10146 ( .C1(n9999), .C2(n9996), .A(n9758), .B(n9757), .ZN(n9759)
         );
  NAND2_X1 U10147 ( .A1(n9756), .A2(n7774), .ZN(n9757) );
  NOR2_X1 U10148 ( .A1(n9752), .A2(n7774), .ZN(n9760) );
  AOI21_X1 U10149 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9752) );
  OAI211_X1 U10150 ( .C1(n10033), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        n6999) );
  OAI21_X1 U10151 ( .B1(n10029), .B2(n10028), .A(n10280), .ZN(n10030) );
  OAI211_X1 U10152 ( .C1(n8121), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10028) );
  AOI22_X1 U10153 ( .A1(n10024), .A2(n10023), .B1(n10022), .B2(n10021), .ZN(
        n10025) );
  AOI22_X1 U10154 ( .A1(n11721), .A2(n10020), .B1(n10284), .B2(n10019), .ZN(
        n10026) );
  OAI211_X1 U10155 ( .C1(n7777), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        n10029) );
  NAND2_X1 U10156 ( .A1(n10014), .A2(n10013), .ZN(n10015) );
  OAI21_X1 U10157 ( .B1(n9317), .B2(n11733), .A(n9548), .ZN(n9196) );
  INV_X1 U10158 ( .A(n9543), .ZN(n9194) );
  AOI22_X1 U10159 ( .A1(n10012), .A2(n7759), .B1(n10010), .B2(n10009), .ZN(
        n10016) );
  INV_X1 U10160 ( .A(n10008), .ZN(n10012) );
  AOI22_X1 U10161 ( .A1(n10007), .A2(n10006), .B1(n7764), .B2(DRAM_ADDRESS[17]), .ZN(n10031) );
  XNOR2_X1 U10162 ( .A(\DP_OP_751_130_6421/n1005 ), .B(n10005), .ZN(n10006) );
  AOI211_X1 U10163 ( .C1(\DataPath/ALUhw/i_Q_EXTENDED[49] ), .C2(n10004), .A(
        n10003), .B(n10002), .ZN(n10033) );
  OAI22_X1 U10164 ( .A1(n10001), .A2(n10000), .B1(n9999), .B2(n9998), .ZN(
        n10002) );
  XNOR2_X1 U10165 ( .A(n9997), .B(n9996), .ZN(n10000) );
  OAI211_X1 U10166 ( .C1(n9999), .C2(n9995), .A(n9994), .B(n9993), .ZN(n10003)
         );
  NAND2_X1 U10167 ( .A1(n9989), .A2(n9997), .ZN(n9995) );
  INV_X1 U10168 ( .A(n9753), .ZN(n9989) );
  OAI222_X1 U10169 ( .A1(n11735), .A2(n9748), .B1(n11730), .B2(n9747), .C1(
        n11734), .C2(n518), .ZN(n6998) );
  NOR3_X1 U10170 ( .A1(n9746), .A2(n9745), .A3(n9744), .ZN(n9747) );
  OAI22_X1 U10171 ( .A1(n9789), .A2(n9939), .B1(n9881), .B2(n9942), .ZN(n9744)
         );
  INV_X1 U10172 ( .A(n10019), .ZN(n9789) );
  OR4_X1 U10173 ( .A1(n9208), .A2(n9207), .A3(n9206), .A4(n9205), .ZN(n10019)
         );
  OAI21_X1 U10174 ( .B1(n9593), .B2(n9204), .A(n9203), .ZN(n9205) );
  NAND2_X1 U10175 ( .A1(n8325), .A2(n9202), .ZN(n9203) );
  INV_X1 U10176 ( .A(n9498), .ZN(n9202) );
  NAND2_X1 U10177 ( .A1(n9516), .A2(n11731), .ZN(n9204) );
  NOR2_X1 U10178 ( .A1(n9220), .A2(n9495), .ZN(n9206) );
  NOR2_X1 U10179 ( .A1(n9201), .A2(n9589), .ZN(n9207) );
  AOI21_X1 U10180 ( .B1(n11731), .B2(n9500), .A(n9497), .ZN(n9201) );
  AOI21_X1 U10181 ( .B1(n9538), .B2(n9200), .A(n9494), .ZN(n9208) );
  INV_X1 U10182 ( .A(n7942), .ZN(n9197) );
  INV_X1 U10183 ( .A(n9199), .ZN(n9198) );
  OAI22_X1 U10184 ( .A1(n7777), .A2(n10027), .B1(n10008), .B2(n9880), .ZN(
        n9745) );
  OAI211_X1 U10185 ( .C1(n8121), .C2(n9878), .A(n9743), .B(n9742), .ZN(n9746)
         );
  AOI22_X1 U10186 ( .A1(n10024), .A2(n7759), .B1(n10022), .B2(n10020), .ZN(
        n9742) );
  AOI22_X1 U10187 ( .A1(n10286), .A2(n9874), .B1(n11721), .B2(n10284), .ZN(
        n9743) );
  AOI21_X1 U10188 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[50] ), .B2(n10004), .A(
        n9741), .ZN(n9748) );
  OAI211_X1 U10189 ( .C1(n9740), .C2(n10001), .A(n9739), .B(n9738), .ZN(n9741)
         );
  OAI21_X1 U10190 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9733) );
  INV_X1 U10191 ( .A(n9998), .ZN(n9732) );
  INV_X1 U10192 ( .A(n9999), .ZN(n9751) );
  INV_X1 U10193 ( .A(n9754), .ZN(n10001) );
  XNOR2_X1 U10194 ( .A(n9729), .B(n9728), .ZN(n9740) );
  OAI222_X1 U10195 ( .A1(n11735), .A2(n9727), .B1(n11730), .B2(n9726), .C1(
        n11734), .C2(n519), .ZN(n6997) );
  NOR3_X1 U10196 ( .A1(n9725), .A2(n9724), .A3(n9723), .ZN(n9726) );
  OAI22_X1 U10197 ( .A1(n10008), .A2(n9942), .B1(n9881), .B2(n9918), .ZN(n9723) );
  OAI22_X1 U10198 ( .A1(n7777), .A2(n9878), .B1(n9879), .B2(n10017), .ZN(n9724) );
  OAI211_X1 U10199 ( .C1(n8121), .C2(n9860), .A(n9722), .B(n9721), .ZN(n9725)
         );
  AOI22_X1 U10200 ( .A1(n10024), .A2(n10010), .B1(n10022), .B2(n10284), .ZN(
        n9721) );
  AOI22_X1 U10201 ( .A1(n9978), .A2(n9874), .B1(n11721), .B2(n10013), .ZN(
        n9722) );
  OAI211_X1 U10202 ( .C1(n9472), .C2(n9538), .A(n9228), .B(n9227), .ZN(n11721)
         );
  NAND2_X1 U10203 ( .A1(n9226), .A2(n9225), .ZN(n9227) );
  INV_X1 U10204 ( .A(n9596), .ZN(n9226) );
  AOI211_X1 U10205 ( .C1(n9686), .C2(n9224), .A(n9223), .B(n9222), .ZN(n9228)
         );
  OAI22_X1 U10206 ( .A1(n9630), .A2(n9221), .B1(n9220), .B2(n9475), .ZN(n9222)
         );
  INV_X1 U10207 ( .A(n9426), .ZN(n9220) );
  OAI22_X1 U10208 ( .A1(n7937), .A2(n9477), .B1(n11717), .B2(n9593), .ZN(n9223) );
  INV_X1 U10209 ( .A(n9479), .ZN(n9224) );
  AOI21_X1 U10210 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[51] ), .B2(n10004), .A(
        n9720), .ZN(n9727) );
  OAI21_X1 U10211 ( .B1(n9719), .B2(n9999), .A(n9718), .ZN(n9720) );
  AOI21_X1 U10212 ( .B1(n9754), .B2(n9717), .A(n9716), .ZN(n9718) );
  OAI211_X1 U10213 ( .C1(n9715), .C2(n9850), .A(n9714), .B(n9713), .ZN(n9716)
         );
  XNOR2_X1 U10214 ( .A(\DP_OP_751_130_6421/n903 ), .B(n9711), .ZN(n9715) );
  XNOR2_X1 U10215 ( .A(n9710), .B(n9709), .ZN(n9717) );
  AND2_X1 U10216 ( .A1(n9708), .A2(n9958), .ZN(n9754) );
  NAND2_X1 U10217 ( .A1(n9707), .A2(n9958), .ZN(n9999) );
  INV_X1 U10218 ( .A(n9708), .ZN(n9707) );
  XNOR2_X1 U10219 ( .A(n9706), .B(n9709), .ZN(n9719) );
  XNOR2_X1 U10220 ( .A(n9705), .B(n9711), .ZN(n9709) );
  AOI22_X1 U10221 ( .A1(n10267), .A2(i_RD1[9]), .B1(n10266), .B2(
        IRAM_ADDRESS[9]), .ZN(n11669) );
  NOR2_X1 U10222 ( .A1(n8815), .A2(n8814), .ZN(n8810) );
  OAI222_X1 U10223 ( .A1(n11735), .A2(n9704), .B1(n11730), .B2(n9703), .C1(
        n11734), .C2(n520), .ZN(n6996) );
  NOR3_X1 U10224 ( .A1(n9702), .A2(n9701), .A3(n9700), .ZN(n9703) );
  OAI22_X1 U10225 ( .A1(n9879), .A2(n10027), .B1(n9699), .B2(n10017), .ZN(
        n9700) );
  INV_X1 U10226 ( .A(n9875), .ZN(n9699) );
  OAI22_X1 U10227 ( .A1(n7777), .A2(n9860), .B1(n10008), .B2(n9918), .ZN(n9701) );
  OAI211_X1 U10228 ( .C1(n8121), .C2(n9880), .A(n9698), .B(n9697), .ZN(n9702)
         );
  AOI22_X1 U10229 ( .A1(n10024), .A2(n10021), .B1(n10022), .B2(n10013), .ZN(
        n9697) );
  NAND4_X1 U10230 ( .A1(n9696), .A2(n9695), .A3(n9694), .A4(n9693), .ZN(n10022) );
  OAI211_X1 U10231 ( .C1(n9692), .C2(n11731), .A(n9691), .B(n9690), .ZN(n9693)
         );
  NAND2_X1 U10232 ( .A1(n8300), .A2(n11731), .ZN(n9690) );
  NAND2_X1 U10233 ( .A1(n9688), .A2(n9687), .ZN(n9694) );
  AOI22_X1 U10234 ( .A1(n9686), .A2(n9685), .B1(n8325), .B2(n9684), .ZN(n9695)
         );
  AOI22_X1 U10235 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9680), .ZN(n9696)
         );
  INV_X1 U10236 ( .A(n9330), .ZN(n9680) );
  INV_X1 U10237 ( .A(n9670), .ZN(n9681) );
  AOI22_X1 U10238 ( .A1(n9874), .A2(n10023), .B1(n10284), .B2(n10009), .ZN(
        n9698) );
  AOI211_X1 U10239 ( .C1(\DataPath/ALUhw/i_Q_EXTENDED[52] ), .C2(n8337), .A(
        n9664), .B(n9663), .ZN(n9704) );
  OAI211_X1 U10240 ( .C1(n9660), .C2(n9850), .A(n9894), .B(n9659), .ZN(n9661)
         );
  NAND2_X1 U10241 ( .A1(n9992), .A2(n9660), .ZN(n9659) );
  OAI211_X1 U10242 ( .C1(n9660), .C2(n9795), .A(n9658), .B(n9657), .ZN(n9662)
         );
  NAND2_X1 U10243 ( .A1(n9803), .A2(n9660), .ZN(n9657) );
  NAND2_X1 U10244 ( .A1(n9898), .A2(n9656), .ZN(n9658) );
  OAI22_X1 U10245 ( .A1(n9894), .A2(n9656), .B1(n9655), .B2(n9885), .ZN(n9664)
         );
  INV_X1 U10246 ( .A(n9898), .ZN(n9655) );
  OAI21_X1 U10247 ( .B1(n10207), .B2(n11678), .A(n10206), .ZN(n7050) );
  AOI22_X1 U10248 ( .A1(n10267), .A2(i_RD1[6]), .B1(IRAM_ADDRESS[6]), .B2(
        n10266), .ZN(n10206) );
  XNOR2_X1 U10249 ( .A(n7696), .B(n10205), .ZN(n10207) );
  NAND2_X1 U10250 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  INV_X1 U10251 ( .A(n10202), .ZN(n10204) );
  OAI21_X1 U10252 ( .B1(n10193), .B2(n11678), .A(n10192), .ZN(n7046) );
  AOI22_X1 U10253 ( .A1(n10267), .A2(i_RD1[10]), .B1(IRAM_ADDRESS[10]), .B2(
        n10266), .ZN(n10192) );
  NOR2_X1 U10254 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  OAI211_X1 U10255 ( .C1(n9908), .C2(n11730), .A(n9907), .B(n9906), .ZN(n6995)
         );
  AOI22_X1 U10256 ( .A1(n10007), .A2(n9905), .B1(n7764), .B2(DRAM_ADDRESS[21]), 
        .ZN(n9906) );
  XNOR2_X1 U10257 ( .A(\DP_OP_751_130_6421/n801 ), .B(n9904), .ZN(n9905) );
  NAND2_X1 U10258 ( .A1(n9903), .A2(n10279), .ZN(n9907) );
  OAI211_X1 U10259 ( .C1(n9902), .C2(n9901), .A(n9900), .B(n9899), .ZN(n9903)
         );
  AOI211_X1 U10260 ( .C1(n9898), .C2(n9897), .A(n9896), .B(n9895), .ZN(n9899)
         );
  NOR2_X1 U10261 ( .A1(n9894), .A2(n9893), .ZN(n9895) );
  NAND2_X1 U10262 ( .A1(n9888), .A2(n9885), .ZN(n9894) );
  NAND2_X1 U10263 ( .A1(n9892), .A2(n9891), .ZN(n9896) );
  INV_X1 U10264 ( .A(\DP_OP_751_130_6421/n801 ), .ZN(n9890) );
  NAND2_X1 U10265 ( .A1(\DataPath/ALUhw/i_Q_EXTENDED[53] ), .A2(n8337), .ZN(
        n9900) );
  AOI22_X1 U10266 ( .A1(n9888), .A2(n9887), .B1(n9898), .B2(n9886), .ZN(n9901)
         );
  INV_X1 U10267 ( .A(n9885), .ZN(n9887) );
  INV_X1 U10268 ( .A(n9893), .ZN(n9902) );
  NOR3_X1 U10269 ( .A1(n9884), .A2(n9883), .A3(n9882), .ZN(n9908) );
  OAI22_X1 U10270 ( .A1(n10008), .A2(n9982), .B1(n9881), .B2(n9939), .ZN(n9882) );
  INV_X1 U10271 ( .A(n10009), .ZN(n9881) );
  OAI211_X1 U10272 ( .C1(n9679), .C2(n7942), .A(n9677), .B(n9676), .ZN(n10009)
         );
  OAI21_X1 U10273 ( .B1(n9675), .B2(n9674), .A(n9691), .ZN(n9676) );
  NOR2_X1 U10274 ( .A1(n9826), .A2(n11733), .ZN(n9674) );
  AOI21_X1 U10275 ( .B1(n9686), .B2(n9673), .A(n9672), .ZN(n9677) );
  OAI22_X1 U10276 ( .A1(n7937), .A2(n9671), .B1(n9670), .B2(n9669), .ZN(n9672)
         );
  OR2_X1 U10277 ( .A1(n7942), .A2(n9102), .ZN(n9670) );
  INV_X1 U10278 ( .A(n11718), .ZN(n9102) );
  OAI21_X1 U10279 ( .B1(n9668), .B2(n9667), .A(n9666), .ZN(n9673) );
  INV_X1 U10280 ( .A(n9411), .ZN(n9666) );
  INV_X1 U10281 ( .A(n9665), .ZN(n9679) );
  OAI22_X1 U10282 ( .A1(n7777), .A2(n9880), .B1(n9879), .B2(n9878), .ZN(n9883)
         );
  OAI211_X1 U10283 ( .C1(n8121), .C2(n9942), .A(n9877), .B(n9876), .ZN(n9884)
         );
  AOI22_X1 U10284 ( .A1(n10020), .A2(n10024), .B1(n9875), .B2(n9978), .ZN(
        n9876) );
  AOI22_X1 U10285 ( .A1(n9874), .A2(n7759), .B1(n10286), .B2(n9873), .ZN(n9877) );
  OAI222_X1 U10286 ( .A1(n10209), .A2(n7750), .B1(n10210), .B2(\intadd_1/A[3] ), .C1(n11678), .C2(\intadd_1/SUM[3] ), .ZN(n7052) );
  INV_X1 U10287 ( .A(i_RD1[4]), .ZN(n10209) );
  OAI222_X1 U10288 ( .A1(n10208), .A2(n7750), .B1(n10210), .B2(\intadd_1/A[4] ), .C1(n11678), .C2(\intadd_1/SUM[4] ), .ZN(n7051) );
  INV_X1 U10289 ( .A(i_RD1[5]), .ZN(n10208) );
  OAI22_X1 U10290 ( .A1(n9654), .A2(n11735), .B1(n521), .B2(n11734), .ZN(n6994) );
  AOI211_X1 U10291 ( .C1(\DataPath/ALUhw/i_Q_EXTENDED[54] ), .C2(n10004), .A(
        n9653), .B(n9652), .ZN(n9654) );
  OAI211_X1 U10292 ( .C1(n9651), .C2(n9815), .A(n9650), .B(n9649), .ZN(n9652)
         );
  OAI211_X1 U10293 ( .C1(n9645), .C2(n9644), .A(n9898), .B(n9643), .ZN(n9650)
         );
  NOR3_X1 U10294 ( .A1(n9642), .A2(n9641), .A3(n9640), .ZN(n9651) );
  OAI22_X1 U10295 ( .A1(n9879), .A2(n9860), .B1(n9861), .B2(n10017), .ZN(n9640) );
  OAI22_X1 U10296 ( .A1(n7777), .A2(n9942), .B1(n10008), .B2(n9939), .ZN(n9641) );
  OAI22_X1 U10297 ( .A1(n9636), .A2(n9635), .B1(n9634), .B2(n9633), .ZN(n9637)
         );
  NAND2_X1 U10298 ( .A1(n9560), .A2(i_ALU_OP[4]), .ZN(n9633) );
  INV_X1 U10299 ( .A(n9632), .ZN(n9635) );
  AOI21_X1 U10300 ( .B1(n9691), .B2(n9631), .A(n9426), .ZN(n9636) );
  OAI21_X1 U10301 ( .B1(n9630), .B2(n9629), .A(n9628), .ZN(n9638) );
  AOI22_X1 U10302 ( .A1(n9686), .A2(n9627), .B1(n8325), .B2(n9626), .ZN(n9628)
         );
  INV_X1 U10303 ( .A(n9390), .ZN(n9629) );
  OAI211_X1 U10304 ( .C1(n8121), .C2(n9918), .A(n9625), .B(n9624), .ZN(n9642)
         );
  AOI22_X1 U10305 ( .A1(n10284), .A2(n10024), .B1(n9875), .B2(n10023), .ZN(
        n9624) );
  AOI22_X1 U10306 ( .A1(n9874), .A2(n10010), .B1(n9978), .B2(n9873), .ZN(n9625) );
  AOI21_X1 U10307 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9653) );
  INV_X1 U10308 ( .A(n9888), .ZN(n9621) );
  NAND2_X1 U10309 ( .A1(n9620), .A2(n9619), .ZN(n9622) );
  INV_X1 U10310 ( .A(n9644), .ZN(n9619) );
  OAI222_X1 U10311 ( .A1(n10210), .A2(n8133), .B1(n7750), .B2(n8587), .C1(
        n11678), .C2(\intadd_1/SUM[2] ), .ZN(n7053) );
  OAI21_X1 U10312 ( .B1(n8528), .B2(n7750), .A(n10213), .ZN(n7056) );
  NAND2_X1 U10313 ( .A1(n7750), .A2(n10212), .ZN(n10213) );
  OAI222_X1 U10314 ( .A1(n11678), .A2(\intadd_0/SUM[0] ), .B1(n10210), .B2(
        \intadd_0/A[0] ), .C1(n7750), .C2(n8566), .ZN(n7045) );
  OAI222_X1 U10315 ( .A1(n11678), .A2(\intadd_1/SUM[0] ), .B1(n10210), .B2(
        \intadd_1/A[0] ), .C1(n7750), .C2(n11668), .ZN(n7055) );
  OAI222_X1 U10316 ( .A1(n11678), .A2(n10201), .B1(n10210), .B2(n210), .C1(
        n7750), .C2(n8579), .ZN(n7049) );
  XNOR2_X1 U10317 ( .A(n10198), .B(n210), .ZN(n10199) );
  OAI222_X1 U10318 ( .A1(n11678), .A2(\intadd_1/SUM[1] ), .B1(n10210), .B2(
        \intadd_1/A[1] ), .C1(n7750), .C2(n8585), .ZN(n7054) );
  OAI222_X1 U10319 ( .A1(n10210), .A2(n8125), .B1(n7750), .B2(n8543), .C1(
        n11678), .C2(\intadd_0/SUM[4] ), .ZN(n7041) );
  OAI222_X1 U10320 ( .A1(n10210), .A2(n8128), .B1(n7750), .B2(n11671), .C1(
        n11678), .C2(\intadd_0/SUM[1] ), .ZN(n7044) );
  OAI22_X1 U10321 ( .A1(n9618), .A2(n11735), .B1(n522), .B2(n11734), .ZN(n6993) );
  AOI211_X1 U10322 ( .C1(\DataPath/ALUhw/i_Q_EXTENDED[55] ), .C2(n10004), .A(
        n9617), .B(n9616), .ZN(n9618) );
  OAI211_X1 U10323 ( .C1(n9615), .C2(n9815), .A(n9614), .B(n9613), .ZN(n9616)
         );
  AOI211_X1 U10324 ( .C1(n9803), .C2(n9612), .A(n9611), .B(n9610), .ZN(n9613)
         );
  NOR3_X1 U10325 ( .A1(n9797), .A2(n9609), .A3(n9608), .ZN(n9610) );
  NOR3_X1 U10326 ( .A1(n9795), .A2(n9607), .A3(n7782), .ZN(n9611) );
  XNOR2_X1 U10327 ( .A(n7782), .B(n9608), .ZN(n9612) );
  INV_X1 U10328 ( .A(n9604), .ZN(n9605) );
  INV_X1 U10329 ( .A(n9623), .ZN(n9606) );
  NOR3_X1 U10330 ( .A1(n9603), .A2(n9602), .A3(n9601), .ZN(n9615) );
  OAI22_X1 U10331 ( .A1(n9600), .A2(n10017), .B1(n9861), .B2(n10027), .ZN(
        n9601) );
  OAI22_X1 U10332 ( .A1(n7777), .A2(n9918), .B1(n9879), .B2(n9880), .ZN(n9602)
         );
  OAI211_X1 U10333 ( .C1(n8121), .C2(n9982), .A(n9599), .B(n9598), .ZN(n9603)
         );
  AOI22_X1 U10334 ( .A1(n10013), .A2(n10024), .B1(n9875), .B2(n7759), .ZN(
        n9598) );
  NAND2_X1 U10335 ( .A1(n9560), .A2(n11718), .ZN(n9596) );
  INV_X1 U10336 ( .A(n9341), .ZN(n9590) );
  AOI22_X1 U10337 ( .A1(n9874), .A2(n10021), .B1(n10023), .B2(n9873), .ZN(
        n9599) );
  INV_X1 U10338 ( .A(n9859), .ZN(n9874) );
  NOR2_X1 U10339 ( .A1(n9587), .A2(n9586), .ZN(n9617) );
  XNOR2_X1 U10340 ( .A(n9585), .B(n9604), .ZN(n9586) );
  XNOR2_X1 U10341 ( .A(n9584), .B(n9607), .ZN(n9604) );
  NOR2_X1 U10342 ( .A1(n9583), .A2(n11727), .ZN(n9585) );
  INV_X1 U10343 ( .A(n9643), .ZN(n9583) );
  AOI21_X1 U10344 ( .B1(n9888), .B2(n9623), .A(n9898), .ZN(n9587) );
  NOR2_X1 U10345 ( .A1(n9582), .A2(n9935), .ZN(n9898) );
  NAND2_X1 U10346 ( .A1(n9581), .A2(n9644), .ZN(n9623) );
  INV_X1 U10347 ( .A(n9620), .ZN(n9581) );
  NOR2_X1 U10348 ( .A1(n9580), .A2(n9579), .ZN(n9620) );
  NOR2_X1 U10349 ( .A1(n9578), .A2(n9935), .ZN(n9888) );
  INV_X1 U10350 ( .A(n9582), .ZN(n9578) );
  AOI22_X1 U10351 ( .A1(n10267), .A2(i_RD1[18]), .B1(IRAM_ADDRESS[18]), .B2(
        n10266), .ZN(n11674) );
  NAND2_X1 U10352 ( .A1(n10149), .A2(n8830), .ZN(n8828) );
  OAI222_X1 U10353 ( .A1(n10210), .A2(n8127), .B1(n7750), .B2(n8514), .C1(
        n11678), .C2(\intadd_0/SUM[2] ), .ZN(n7043) );
  AOI22_X1 U10354 ( .A1(n10267), .A2(i_RD1[19]), .B1(IRAM_ADDRESS[19]), .B2(
        n10266), .ZN(n11676) );
  XNOR2_X1 U10355 ( .A(n8835), .B(n8834), .ZN(n11677) );
  XNOR2_X1 U10356 ( .A(n10150), .B(IRAM_ADDRESS[19]), .ZN(n8834) );
  AOI21_X1 U10357 ( .B1(n10149), .B2(n10146), .A(n10147), .ZN(n8835) );
  OAI222_X1 U10358 ( .A1(n11735), .A2(n9577), .B1(n11730), .B2(n9576), .C1(
        n11734), .C2(n523), .ZN(n6992) );
  NOR3_X1 U10359 ( .A1(n9575), .A2(n9574), .A3(n9573), .ZN(n9576) );
  OAI211_X1 U10360 ( .C1(n8121), .C2(n9939), .A(n9572), .B(n9571), .ZN(n9573)
         );
  AOI22_X1 U10361 ( .A1(n10010), .A2(n9875), .B1(n9864), .B2(n9978), .ZN(n9571) );
  AOI22_X1 U10362 ( .A1(n9862), .A2(n10286), .B1(n10011), .B2(n9873), .ZN(
        n9572) );
  NAND2_X1 U10363 ( .A1(n9566), .A2(n9565), .ZN(n9567) );
  NAND2_X1 U10364 ( .A1(n9564), .A2(n11733), .ZN(n9565) );
  OAI21_X1 U10365 ( .B1(n9563), .B2(n9593), .A(n9220), .ZN(n9566) );
  INV_X1 U10366 ( .A(n9562), .ZN(n9563) );
  NAND2_X1 U10367 ( .A1(n9561), .A2(n9687), .ZN(n9568) );
  AOI22_X1 U10368 ( .A1(n9560), .A2(n9559), .B1(n8325), .B2(n9558), .ZN(n9569)
         );
  INV_X1 U10369 ( .A(n9557), .ZN(n9558) );
  OAI22_X1 U10370 ( .A1(n8315), .A2(n11684), .B1(n11683), .B2(n9527), .ZN(
        n9559) );
  NAND2_X1 U10371 ( .A1(n9556), .A2(n9555), .ZN(n9570) );
  AND2_X1 U10372 ( .A1(n9686), .A2(n9554), .ZN(n9555) );
  NAND2_X1 U10373 ( .A1(n9305), .A2(n9667), .ZN(n9554) );
  OR2_X1 U10374 ( .A1(n9304), .A2(n9667), .ZN(n9556) );
  OAI22_X1 U10375 ( .A1(n9879), .A2(n9942), .B1(n9861), .B2(n9878), .ZN(n9574)
         );
  OAI22_X1 U10376 ( .A1(n7777), .A2(n9982), .B1(n9859), .B2(n9918), .ZN(n9575)
         );
  AOI21_X1 U10377 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[56] ), .B2(n10004), .A(
        n9536), .ZN(n9577) );
  OAI21_X1 U10378 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9536) );
  AOI21_X1 U10379 ( .B1(n9532), .B2(n9534), .A(n9531), .ZN(n9533) );
  INV_X1 U10380 ( .A(n9850), .ZN(n9803) );
  NAND2_X1 U10381 ( .A1(n9845), .A2(n9843), .ZN(n9534) );
  OAI222_X1 U10382 ( .A1(n10210), .A2(n8126), .B1(n7750), .B2(n8541), .C1(
        n11678), .C2(\intadd_0/SUM[3] ), .ZN(n7042) );
  OAI21_X1 U10383 ( .B1(n7917), .B2(n10188), .A(n8818), .ZN(\intadd_0/n41 ) );
  AND2_X1 U10384 ( .A1(\C620/DATA2_23 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[23])
         );
  OAI222_X1 U10385 ( .A1(n8222), .A2(n11734), .B1(n10032), .B2(n9872), .C1(
        n11730), .C2(n9871), .ZN(n6991) );
  NOR3_X1 U10386 ( .A1(n9870), .A2(n9869), .A3(n9868), .ZN(n9871) );
  OAI211_X1 U10387 ( .C1(n9867), .C2(n9880), .A(n9866), .B(n9865), .ZN(n9868)
         );
  AOI22_X1 U10388 ( .A1(n10021), .A2(n9875), .B1(n9864), .B2(n10023), .ZN(
        n9865) );
  AOI22_X1 U10389 ( .A1(n9863), .A2(n10286), .B1(n9862), .B2(n9978), .ZN(n9866) );
  OAI22_X1 U10390 ( .A1(n9879), .A2(n9918), .B1(n9861), .B2(n9860), .ZN(n9869)
         );
  OAI22_X1 U10391 ( .A1(n7777), .A2(n9939), .B1(n9859), .B2(n9982), .ZN(n9870)
         );
  OAI22_X1 U10392 ( .A1(n9549), .A2(n9548), .B1(n9547), .B2(n10005), .ZN(n9550) );
  AOI21_X1 U10393 ( .B1(n9913), .B2(n11680), .A(n9040), .ZN(n9548) );
  OAI22_X1 U10394 ( .A1(n9546), .A2(n9545), .B1(n7937), .B2(n9544), .ZN(n9551)
         );
  INV_X1 U10395 ( .A(n10283), .ZN(n9544) );
  AOI211_X1 U10396 ( .C1(n9543), .C2(n9667), .A(n9593), .B(n9542), .ZN(n9552)
         );
  NOR2_X1 U10397 ( .A1(n9541), .A2(n11733), .ZN(n9542) );
  OAI22_X1 U10398 ( .A1(n9540), .A2(n9630), .B1(n9539), .B2(n9538), .ZN(n9553)
         );
  INV_X1 U10399 ( .A(n9537), .ZN(n9539) );
  AOI21_X1 U10400 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[57] ), .B2(n8337), .A(
        n9858), .ZN(n9872) );
  OAI21_X1 U10401 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(n9858) );
  AOI21_X1 U10402 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9855) );
  OAI211_X1 U10403 ( .C1(n9851), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9852)
         );
  XNOR2_X1 U10404 ( .A(\DP_OP_751_130_6421/n597 ), .B(n7691), .ZN(n9851) );
  AOI21_X1 U10405 ( .B1(n9843), .B2(n9844), .A(n9842), .ZN(n9856) );
  INV_X1 U10406 ( .A(n9841), .ZN(n9842) );
  INV_X1 U10407 ( .A(n10185), .ZN(n7035) );
  AOI222_X1 U10408 ( .A1(\intadd_2/SUM[0] ), .A2(n8421), .B1(IRAM_ADDRESS[21]), 
        .B2(n10266), .C1(i_RD1[21]), .C2(n10267), .ZN(n10185) );
  OAI22_X1 U10409 ( .A1(n9525), .A2(n11735), .B1(n524), .B2(n11734), .ZN(n6990) );
  AOI211_X1 U10410 ( .C1(\DataPath/ALUhw/i_Q_EXTENDED[58] ), .C2(n10004), .A(
        n9524), .B(n9523), .ZN(n9525) );
  OAI211_X1 U10411 ( .C1(n9522), .C2(n9815), .A(n9521), .B(n9520), .ZN(n9523)
         );
  OAI21_X1 U10412 ( .B1(n9515), .B2(n9514), .A(n9854), .ZN(n9521) );
  INV_X1 U10413 ( .A(n9535), .ZN(n9854) );
  AND3_X1 U10414 ( .A1(n9513), .A2(n9512), .A3(n11729), .ZN(n9514) );
  NOR3_X1 U10415 ( .A1(n9511), .A2(n9510), .A3(n9509), .ZN(n9522) );
  OAI211_X1 U10416 ( .C1(n9867), .C2(n9942), .A(n9508), .B(n9507), .ZN(n9509)
         );
  AOI22_X1 U10417 ( .A1(n10020), .A2(n9875), .B1(n9864), .B2(n7759), .ZN(n9507) );
  AOI22_X1 U10418 ( .A1(n9863), .A2(n9978), .B1(n9828), .B2(n10286), .ZN(n9508) );
  OAI22_X1 U10419 ( .A1(n9859), .A2(n9939), .B1(n9506), .B2(n9878), .ZN(n9510)
         );
  NOR2_X1 U10420 ( .A1(n9505), .A2(n9504), .ZN(n9859) );
  OAI211_X1 U10421 ( .C1(n9538), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9504)
         );
  OAI211_X1 U10422 ( .C1(n11733), .C2(n9500), .A(n9691), .B(n9499), .ZN(n9501)
         );
  NAND2_X1 U10423 ( .A1(n9498), .A2(n9667), .ZN(n9499) );
  AOI22_X1 U10424 ( .A1(n9560), .A2(n9497), .B1(n8325), .B2(n9496), .ZN(n9502)
         );
  INV_X1 U10425 ( .A(n9299), .ZN(n9496) );
  OAI21_X1 U10426 ( .B1(n8309), .B2(n11684), .A(n8964), .ZN(n9497) );
  AOI211_X1 U10427 ( .C1(n9667), .C2(n9495), .A(n9589), .B(n9494), .ZN(n9505)
         );
  NOR2_X1 U10428 ( .A1(n9301), .A2(n9667), .ZN(n9494) );
  OAI22_X1 U10429 ( .A1(n9879), .A2(n9982), .B1(n9861), .B2(n9880), .ZN(n9511)
         );
  NOR2_X1 U10430 ( .A1(n9857), .A2(n9493), .ZN(n9524) );
  XNOR2_X1 U10431 ( .A(n10276), .B(n9492), .ZN(n9493) );
  INV_X1 U10432 ( .A(n9532), .ZN(n9857) );
  AND2_X1 U10433 ( .A1(\C620/DATA2_24 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[24])
         );
  OAI21_X1 U10434 ( .B1(n10182), .B2(n11678), .A(n10181), .ZN(n7031) );
  AOI22_X1 U10435 ( .A1(n10267), .A2(i_RD1[25]), .B1(IRAM_ADDRESS[25]), .B2(
        n10266), .ZN(n10181) );
  XNOR2_X1 U10436 ( .A(\intadd_2/CO ), .B(n10180), .ZN(n10182) );
  INV_X1 U10437 ( .A(n10184), .ZN(n7034) );
  AOI222_X1 U10438 ( .A1(\intadd_2/SUM[1] ), .A2(n8421), .B1(IRAM_ADDRESS[22]), 
        .B2(n10266), .C1(i_RD1[22]), .C2(n10267), .ZN(n10184) );
  INV_X1 U10439 ( .A(n10183), .ZN(n7032) );
  AOI222_X1 U10440 ( .A1(\intadd_2/SUM[3] ), .A2(n8421), .B1(IRAM_ADDRESS[24]), 
        .B2(n10266), .C1(i_RD1[24]), .C2(n10267), .ZN(n10183) );
  OAI21_X1 U10441 ( .B1(n10179), .B2(n11678), .A(n10178), .ZN(n7030) );
  AOI22_X1 U10442 ( .A1(n10267), .A2(i_RD1[26]), .B1(IRAM_ADDRESS[26]), .B2(
        n10266), .ZN(n10178) );
  XNOR2_X1 U10443 ( .A(n10175), .B(IRAM_ADDRESS[26]), .ZN(n10176) );
  AND2_X1 U10444 ( .A1(\C620/DATA2_25 ), .A2(n10822), .ZN(DRAMRF_ADDRESS[25])
         );
  OAI222_X1 U10445 ( .A1(n11735), .A2(n9491), .B1(n11730), .B2(n9490), .C1(
        n11734), .C2(n525), .ZN(n6989) );
  NOR3_X1 U10446 ( .A1(n9489), .A2(n9488), .A3(n9487), .ZN(n9490) );
  OAI211_X1 U10447 ( .C1(n9867), .C2(n9918), .A(n9486), .B(n9485), .ZN(n9487)
         );
  AOI22_X1 U10448 ( .A1(n10284), .A2(n9875), .B1(n9864), .B2(n10010), .ZN(
        n9485) );
  AOI22_X1 U10449 ( .A1(n10023), .A2(n9863), .B1(n9833), .B2(n10286), .ZN(
        n9486) );
  OAI22_X1 U10450 ( .A1(n9484), .A2(n10027), .B1(n9506), .B2(n9860), .ZN(n9488) );
  INV_X1 U10451 ( .A(n10011), .ZN(n9860) );
  OAI22_X1 U10452 ( .A1(n9879), .A2(n9939), .B1(n9861), .B2(n9942), .ZN(n9489)
         );
  INV_X1 U10453 ( .A(n9834), .ZN(n9861) );
  OAI22_X1 U10454 ( .A1(n9549), .A2(n9479), .B1(n9547), .B2(n7693), .ZN(n9480)
         );
  AOI21_X1 U10455 ( .B1(n9085), .B2(n11680), .A(n9006), .ZN(n9479) );
  AOI22_X1 U10456 ( .A1(n9478), .A2(n9220), .B1(n11733), .B2(n9477), .ZN(n9481) );
  NAND2_X1 U10457 ( .A1(n9691), .A2(n9476), .ZN(n9478) );
  OAI22_X1 U10458 ( .A1(n9546), .A2(n9475), .B1(n7937), .B2(n9474), .ZN(n9482)
         );
  INV_X1 U10459 ( .A(n10285), .ZN(n9474) );
  INV_X1 U10460 ( .A(n9473), .ZN(n9546) );
  OAI22_X1 U10461 ( .A1(n9472), .A2(n9630), .B1(n9471), .B2(n9538), .ZN(n9483)
         );
  INV_X1 U10462 ( .A(n9687), .ZN(n9538) );
  INV_X1 U10463 ( .A(n9470), .ZN(n9471) );
  INV_X1 U10464 ( .A(n9683), .ZN(n9630) );
  AOI21_X1 U10465 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[59] ), .B2(n8337), .A(
        n9469), .ZN(n9491) );
  OAI21_X1 U10466 ( .B1(n9535), .B2(n9468), .A(n9467), .ZN(n9469) );
  AOI21_X1 U10467 ( .B1(n9532), .B2(n9466), .A(n9465), .ZN(n9467) );
  OAI211_X1 U10468 ( .C1(n9464), .C2(n9850), .A(n9463), .B(n9462), .ZN(n9465)
         );
  INV_X1 U10469 ( .A(\DP_OP_751_130_6421/n495 ), .ZN(n9461) );
  XNOR2_X1 U10470 ( .A(\DP_OP_751_130_6421/n495 ), .B(n9459), .ZN(n9464) );
  NOR2_X1 U10471 ( .A1(n9458), .A2(n9935), .ZN(n9532) );
  AOI21_X1 U10472 ( .B1(n9512), .B2(n11729), .A(n9513), .ZN(n9515) );
  INV_X1 U10473 ( .A(n9492), .ZN(n9513) );
  INV_X1 U10474 ( .A(n9455), .ZN(n9456) );
  INV_X1 U10475 ( .A(n9466), .ZN(n9457) );
  XNOR2_X1 U10476 ( .A(n9454), .B(n9455), .ZN(n9466) );
  AND2_X1 U10477 ( .A1(n9453), .A2(n9452), .ZN(n9455) );
  AOI21_X1 U10478 ( .B1(n10276), .B2(n9492), .A(n9451), .ZN(n9454) );
  INV_X1 U10479 ( .A(n9450), .ZN(n9451) );
  AND2_X1 U10480 ( .A1(n9450), .A2(n9449), .ZN(n9492) );
  NAND2_X1 U10481 ( .A1(n9458), .A2(n9958), .ZN(n9535) );
  INV_X1 U10482 ( .A(n11728), .ZN(n9458) );
  OAI22_X1 U10483 ( .A1(n9448), .A2(n11735), .B1(n526), .B2(n11734), .ZN(n6988) );
  AOI21_X1 U10484 ( .B1(\DataPath/ALUhw/i_Q_EXTENDED[60] ), .B2(n8337), .A(
        n9447), .ZN(n9448) );
  OAI211_X1 U10485 ( .C1(n9446), .C2(n8300), .A(n9445), .B(n9444), .ZN(n9447)
         );
  AOI21_X1 U10486 ( .B1(n8300), .B2(n9443), .A(n9442), .ZN(n9444) );
  AOI21_X1 U10487 ( .B1(n9822), .B2(n9819), .A(n9825), .ZN(n9442) );
  OAI21_X1 U10488 ( .B1(n9820), .B2(n9441), .A(n9440), .ZN(n9443) );
  INV_X1 U10489 ( .A(n9990), .ZN(n9795) );
  OAI21_X1 U10490 ( .B1(n9438), .B2(n9437), .A(n10287), .ZN(n9445) );
  NAND2_X1 U10491 ( .A1(n9436), .A2(n9435), .ZN(n9437) );
  AOI22_X1 U10492 ( .A1(n9862), .A2(n10010), .B1(n10020), .B2(n9834), .ZN(
        n9435) );
  AOI22_X1 U10493 ( .A1(n9863), .A2(n7759), .B1(n9828), .B2(n10023), .ZN(n9436) );
  OAI211_X1 U10494 ( .C1(n9867), .C2(n9982), .A(n9434), .B(n9433), .ZN(n9438)
         );
  AOI22_X1 U10495 ( .A1(n10013), .A2(n9875), .B1(n9864), .B2(n10021), .ZN(
        n9433) );
  OR2_X1 U10496 ( .A1(n9432), .A2(n9431), .ZN(n9875) );
  NAND2_X1 U10497 ( .A1(n9560), .A2(n9685), .ZN(n9428) );
  NAND2_X1 U10498 ( .A1(n8951), .A2(n8950), .ZN(n9685) );
  NAND2_X1 U10499 ( .A1(n9099), .A2(n11680), .ZN(n8951) );
  NAND2_X1 U10500 ( .A1(n9427), .A2(n9687), .ZN(n9429) );
  NAND2_X1 U10501 ( .A1(n9426), .A2(n9684), .ZN(n9430) );
  INV_X1 U10502 ( .A(n9324), .ZN(n9684) );
  NAND4_X1 U10503 ( .A1(n9425), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(n9432)
         );
  NAND2_X1 U10504 ( .A1(n8325), .A2(n9421), .ZN(n9422) );
  NAND2_X1 U10505 ( .A1(n9420), .A2(n9682), .ZN(n9423) );
  NAND2_X1 U10506 ( .A1(n9473), .A2(n9692), .ZN(n9424) );
  NOR2_X1 U10507 ( .A1(n9589), .A2(n11731), .ZN(n9473) );
  NAND2_X1 U10508 ( .A1(n9683), .A2(n9688), .ZN(n9425) );
  AOI22_X1 U10509 ( .A1(n9833), .A2(n9978), .B1(n10286), .B2(n9832), .ZN(n9434) );
  AOI211_X1 U10510 ( .C1(n9992), .C2(n9439), .A(n9407), .B(n9406), .ZN(n9446)
         );
  NOR2_X1 U10511 ( .A1(n9820), .A2(n9405), .ZN(n9406) );
  NOR2_X1 U10512 ( .A1(n9850), .A2(n9439), .ZN(n9407) );
  OAI21_X1 U10513 ( .B1(n10174), .B2(n11678), .A(n10173), .ZN(n7029) );
  AOI22_X1 U10514 ( .A1(n10267), .A2(i_RD1[27]), .B1(IRAM_ADDRESS[27]), .B2(
        n10266), .ZN(n10173) );
  XNOR2_X1 U10515 ( .A(n10172), .B(n10171), .ZN(n10174) );
  NAND2_X1 U10516 ( .A1(n10170), .A2(n10169), .ZN(n10172) );
  OAI21_X1 U10517 ( .B1(IRAM_ADDRESS[26]), .B2(n10175), .A(n10168), .ZN(n10170) );
  OAI21_X1 U10518 ( .B1(n10167), .B2(n11678), .A(n10166), .ZN(n7028) );
  AOI22_X1 U10519 ( .A1(n10267), .A2(i_RD1[28]), .B1(IRAM_ADDRESS[28]), .B2(
        n10266), .ZN(n10166) );
  XNOR2_X1 U10520 ( .A(n10261), .B(n10165), .ZN(n10167) );
  NAND2_X1 U10521 ( .A1(n10164), .A2(n10163), .ZN(n10165) );
  INV_X1 U10522 ( .A(n10162), .ZN(n10164) );
  OAI21_X1 U10523 ( .B1(n9838), .B2(n9837), .A(n10280), .ZN(n9839) );
  OAI211_X1 U10524 ( .C1(n9867), .C2(n9939), .A(n9836), .B(n9835), .ZN(n9837)
         );
  AOI22_X1 U10525 ( .A1(n9864), .A2(n10020), .B1(n9834), .B2(n10284), .ZN(
        n9835) );
  AOI22_X1 U10526 ( .A1(n9833), .A2(n10023), .B1(n9978), .B2(n9832), .ZN(n9836) );
  INV_X1 U10527 ( .A(n9873), .ZN(n9867) );
  NAND4_X1 U10528 ( .A1(n9419), .A2(n9418), .A3(n9417), .A4(n9416), .ZN(n9873)
         );
  OAI211_X1 U10529 ( .C1(n9667), .C2(n9415), .A(n9691), .B(n9414), .ZN(n9416)
         );
  NAND2_X1 U10530 ( .A1(n9671), .A2(n11733), .ZN(n9414) );
  INV_X1 U10531 ( .A(n9285), .ZN(n9671) );
  NAND2_X1 U10532 ( .A1(n9687), .A2(n9413), .ZN(n9417) );
  INV_X1 U10533 ( .A(n9412), .ZN(n9413) );
  AOI22_X1 U10534 ( .A1(n9560), .A2(n9411), .B1(n8325), .B2(n9410), .ZN(n9418)
         );
  OAI21_X1 U10535 ( .B1(n9665), .B2(n9675), .A(n9686), .ZN(n9419) );
  NOR2_X1 U10536 ( .A1(n9409), .A2(n11731), .ZN(n9675) );
  INV_X1 U10537 ( .A(n9408), .ZN(n9409) );
  OAI211_X1 U10538 ( .C1(n9831), .C2(n10017), .A(n9830), .B(n9829), .ZN(n9838)
         );
  NAND2_X1 U10539 ( .A1(n9862), .A2(n10021), .ZN(n9829) );
  AOI22_X1 U10540 ( .A1(n9863), .A2(n10010), .B1(n9828), .B2(n7759), .ZN(n9830) );
  AOI22_X1 U10541 ( .A1(n10007), .A2(n9827), .B1(n7764), .B2(DRAM_ADDRESS[29]), 
        .ZN(n9840) );
  XNOR2_X1 U10542 ( .A(\DP_OP_751_130_6421/n393 ), .B(n9826), .ZN(n9827) );
  NOR2_X1 U10543 ( .A1(n10032), .A2(n9850), .ZN(n10007) );
  XNOR2_X1 U10544 ( .A(n10160), .B(IRAM_ADDRESS[29]), .ZN(n10161) );
  NAND2_X1 U10545 ( .A1(n10175), .A2(n8178), .ZN(n10163) );
  NOR3_X1 U10546 ( .A1(n9403), .A2(n9402), .A3(n9401), .ZN(n9404) );
  OAI22_X1 U10547 ( .A1(n9506), .A2(n9918), .B1(n9484), .B2(n9880), .ZN(n9401)
         );
  INV_X1 U10548 ( .A(n9828), .ZN(n9484) );
  INV_X1 U10549 ( .A(n9862), .ZN(n9506) );
  OAI211_X1 U10550 ( .C1(n9400), .C2(n9878), .A(n9399), .B(n9398), .ZN(n9402)
         );
  AOI22_X1 U10551 ( .A1(n9864), .A2(n10284), .B1(n9834), .B2(n10013), .ZN(
        n9398) );
  NAND4_X1 U10552 ( .A1(n9397), .A2(n9396), .A3(n9395), .A4(n9394), .ZN(n9834)
         );
  NAND2_X1 U10553 ( .A1(n9393), .A2(n9687), .ZN(n9394) );
  AOI21_X1 U10554 ( .B1(n9426), .B2(n9626), .A(n9392), .ZN(n9395) );
  NOR2_X1 U10555 ( .A1(n7937), .A2(n9391), .ZN(n9392) );
  AOI22_X1 U10556 ( .A1(n9420), .A2(n9390), .B1(n9560), .B2(n9627), .ZN(n9396)
         );
  NAND2_X1 U10557 ( .A1(n9030), .A2(n9029), .ZN(n9627) );
  NAND2_X1 U10558 ( .A1(n9129), .A2(n11680), .ZN(n9030) );
  OAI211_X1 U10559 ( .C1(n9639), .C2(n9667), .A(n9686), .B(n9632), .ZN(n9397)
         );
  NAND2_X1 U10560 ( .A1(n9389), .A2(n9667), .ZN(n9632) );
  AOI22_X1 U10561 ( .A1(n7759), .A2(n9833), .B1(n9863), .B2(n10021), .ZN(n9399) );
  INV_X1 U10562 ( .A(n9832), .ZN(n9400) );
  OAI22_X1 U10563 ( .A1(n9831), .A2(n10027), .B1(n9388), .B2(n10017), .ZN(
        n9403) );
  INV_X1 U10564 ( .A(n9387), .ZN(n9388) );
  OAI211_X1 U10565 ( .C1(n9385), .C2(n9820), .A(n9384), .B(n9383), .ZN(n9386)
         );
  AOI211_X1 U10566 ( .C1(n9382), .C2(n9990), .A(n9381), .B(n9380), .ZN(n9383)
         );
  NOR3_X1 U10567 ( .A1(n9850), .A2(n9382), .A3(n9379), .ZN(n9380) );
  NOR2_X1 U10568 ( .A1(n9797), .A2(n9378), .ZN(n9381) );
  INV_X1 U10569 ( .A(n9379), .ZN(n9378) );
  AND2_X1 U10570 ( .A1(n9377), .A2(n9631), .ZN(n9379) );
  INV_X1 U10571 ( .A(n9992), .ZN(n9797) );
  NOR2_X1 U10572 ( .A1(n9377), .A2(n9631), .ZN(n9382) );
  OAI211_X1 U10573 ( .C1(n9376), .C2(n9375), .A(n9374), .B(n9373), .ZN(n9384)
         );
  INV_X1 U10574 ( .A(n9825), .ZN(n9373) );
  XNOR2_X1 U10575 ( .A(n9372), .B(n9375), .ZN(n9385) );
  OAI21_X1 U10576 ( .B1(n9370), .B2(n9825), .A(n9369), .ZN(n9371) );
  AOI211_X1 U10577 ( .C1(n9368), .C2(n10287), .A(n9367), .B(n9366), .ZN(n9369)
         );
  OAI211_X1 U10578 ( .C1(n9365), .C2(n9850), .A(n9364), .B(n9363), .ZN(n9366)
         );
  NAND2_X1 U10579 ( .A1(n8452), .A2(i_ALU_OP[1]), .ZN(n8956) );
  NOR2_X1 U10580 ( .A1(n8957), .A2(n8174), .ZN(n8943) );
  OR2_X1 U10581 ( .A1(i_ALU_OP[0]), .A2(n11681), .ZN(n8957) );
  AOI21_X1 U10582 ( .B1(i_ALU_OP[3]), .B2(n11722), .A(n8193), .ZN(n8959) );
  NAND2_X1 U10583 ( .A1(n8958), .A2(n8095), .ZN(n8960) );
  XNOR2_X1 U10584 ( .A(n8452), .B(i_ALU_OP[4]), .ZN(n8958) );
  XNOR2_X1 U10585 ( .A(\DP_OP_751_130_6421/n291 ), .B(n9361), .ZN(n9365) );
  NOR2_X1 U10586 ( .A1(n9360), .A2(n9820), .ZN(n9367) );
  OR2_X1 U10587 ( .A1(n9359), .A2(n9935), .ZN(n9820) );
  AOI21_X1 U10588 ( .B1(n9372), .B2(n9375), .A(n9356), .ZN(n9357) );
  OAI22_X1 U10589 ( .A1(n9823), .A2(n9819), .B1(n9355), .B2(n9826), .ZN(n9372)
         );
  NAND2_X1 U10590 ( .A1(n9405), .A2(n9689), .ZN(n9819) );
  INV_X1 U10591 ( .A(n9441), .ZN(n9405) );
  NAND4_X1 U10592 ( .A1(n9354), .A2(n9353), .A3(n9352), .A4(n9351), .ZN(n9368)
         );
  AOI21_X1 U10593 ( .B1(n10011), .B2(n9832), .A(n9350), .ZN(n9351) );
  OAI22_X1 U10594 ( .A1(n9349), .A2(n10017), .B1(n9600), .B2(n9939), .ZN(n9350) );
  NAND2_X1 U10595 ( .A1(n8989), .A2(n8988), .ZN(n9939) );
  NOR2_X1 U10596 ( .A1(n7970), .A2(i_ALU_OP[2]), .ZN(n8988) );
  INV_X1 U10597 ( .A(n7785), .ZN(n8989) );
  INV_X1 U10598 ( .A(n9864), .ZN(n9600) );
  NAND4_X1 U10599 ( .A1(n9348), .A2(n9347), .A3(n9346), .A4(n9345), .ZN(n9864)
         );
  NAND2_X1 U10600 ( .A1(n9344), .A2(n9687), .ZN(n9345) );
  OAI211_X1 U10601 ( .C1(n9597), .C2(n9667), .A(n9686), .B(n9594), .ZN(n9346)
         );
  NAND2_X1 U10602 ( .A1(n9343), .A2(n9667), .ZN(n9594) );
  OAI21_X1 U10603 ( .B1(n9595), .B2(n11725), .A(n9342), .ZN(n9597) );
  NAND2_X1 U10604 ( .A1(n9141), .A2(n8971), .ZN(n9595) );
  NAND2_X1 U10605 ( .A1(i_ALU_OP[2]), .A2(n9608), .ZN(n8971) );
  AOI22_X1 U10606 ( .A1(n9560), .A2(n9341), .B1(n8325), .B2(n9340), .ZN(n9347)
         );
  AOI22_X1 U10607 ( .A1(n9426), .A2(n9588), .B1(n9420), .B2(n9591), .ZN(n9348)
         );
  NOR2_X1 U10608 ( .A1(n9593), .A2(n11733), .ZN(n9420) );
  AOI211_X1 U10609 ( .C1(n9686), .C2(n9344), .A(n9339), .B(n9338), .ZN(n9349)
         );
  OAI22_X1 U10610 ( .A1(n9549), .A2(n9343), .B1(n7937), .B2(n9592), .ZN(n9338)
         );
  NAND2_X1 U10611 ( .A1(n9142), .A2(n9141), .ZN(n9343) );
  OR2_X1 U10612 ( .A1(n9774), .A2(i_ALU_OP[2]), .ZN(n9141) );
  NAND2_X1 U10613 ( .A1(n9157), .A2(i_ALU_OP[2]), .ZN(n9142) );
  AND2_X1 U10614 ( .A1(n9426), .A2(n9340), .ZN(n9339) );
  NAND2_X1 U10615 ( .A1(n11732), .A2(n9337), .ZN(n9340) );
  NAND2_X1 U10616 ( .A1(n9607), .A2(i_ALU_OP[2]), .ZN(n9337) );
  OAI21_X1 U10617 ( .B1(n10299), .B2(n9336), .A(n9342), .ZN(n9344) );
  NAND2_X1 U10618 ( .A1(n9591), .A2(n9335), .ZN(n9342) );
  NAND2_X1 U10619 ( .A1(n8973), .A2(n8972), .ZN(n9591) );
  AOI21_X1 U10620 ( .B1(n9361), .B2(n11682), .A(n11685), .ZN(n8972) );
  NAND2_X1 U10621 ( .A1(n7786), .A2(n11720), .ZN(n8973) );
  INV_X1 U10622 ( .A(n9588), .ZN(n9336) );
  NAND4_X1 U10623 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n9832)
         );
  NAND2_X1 U10624 ( .A1(n9688), .A2(n9691), .ZN(n9331) );
  OAI21_X1 U10625 ( .B1(n11725), .B2(n9330), .A(n9329), .ZN(n9688) );
  NAND2_X1 U10626 ( .A1(n9086), .A2(n8949), .ZN(n9330) );
  NAND2_X1 U10627 ( .A1(n8301), .A2(i_ALU_OP[2]), .ZN(n8949) );
  NAND2_X1 U10628 ( .A1(n9328), .A2(n9682), .ZN(n9332) );
  AOI22_X1 U10629 ( .A1(n9426), .A2(n9421), .B1(n9560), .B2(n9692), .ZN(n9333)
         );
  OR2_X1 U10630 ( .A1(n9782), .A2(i_ALU_OP[2]), .ZN(n9086) );
  OAI21_X1 U10631 ( .B1(n8084), .B2(n8301), .A(n9326), .ZN(n9421) );
  NAND2_X1 U10632 ( .A1(n8084), .A2(n9689), .ZN(n9326) );
  AOI22_X1 U10633 ( .A1(n9325), .A2(n9689), .B1(n9686), .B2(n9427), .ZN(n9334)
         );
  OAI21_X1 U10634 ( .B1(n9782), .B2(n8084), .A(n8946), .ZN(n9324) );
  NAND2_X1 U10635 ( .A1(n8084), .A2(n8301), .ZN(n8946) );
  NAND2_X1 U10636 ( .A1(n9682), .A2(n9335), .ZN(n9329) );
  NAND2_X1 U10637 ( .A1(n9689), .A2(n11682), .ZN(n8950) );
  NAND2_X1 U10638 ( .A1(n9099), .A2(n11720), .ZN(n8947) );
  OAI21_X1 U10639 ( .B1(n9069), .B2(n8084), .A(n7785), .ZN(n8975) );
  AOI22_X1 U10640 ( .A1(n10010), .A2(n9833), .B1(n9863), .B2(n10020), .ZN(
        n9352) );
  OAI211_X1 U10641 ( .C1(n9540), .C2(n9593), .A(n9323), .B(n9322), .ZN(n9863)
         );
  AOI21_X1 U10642 ( .B1(n7691), .B2(n9325), .A(n9321), .ZN(n9322) );
  OAI22_X1 U10643 ( .A1(n9220), .A2(n9320), .B1(n9549), .B2(n9545), .ZN(n9321)
         );
  NAND2_X1 U10644 ( .A1(n9077), .A2(n9076), .ZN(n9545) );
  NAND2_X1 U10645 ( .A1(n8311), .A2(i_ALU_OP[2]), .ZN(n9076) );
  AOI21_X1 U10646 ( .B1(n9991), .B2(n8452), .A(n10283), .ZN(n9320) );
  NOR2_X1 U10647 ( .A1(i_ALU_OP[2]), .A2(n9846), .ZN(n10283) );
  AOI22_X1 U10648 ( .A1(n9328), .A2(n9541), .B1(n9537), .B2(n9686), .ZN(n9323)
         );
  OAI21_X1 U10649 ( .B1(n9543), .B2(n10299), .A(n9319), .ZN(n9537) );
  INV_X1 U10650 ( .A(n9318), .ZN(n9319) );
  AOI21_X1 U10651 ( .B1(i_ALU_OP[2]), .B2(n9932), .A(n9038), .ZN(n9543) );
  NOR2_X1 U10652 ( .A1(n8452), .A2(n10005), .ZN(n9038) );
  INV_X1 U10653 ( .A(n9317), .ZN(n9541) );
  AOI21_X1 U10654 ( .B1(n11720), .B2(n9195), .A(n9318), .ZN(n9540) );
  NOR2_X1 U10655 ( .A1(n9317), .A2(n11726), .ZN(n9318) );
  NOR2_X1 U10656 ( .A1(n9846), .A2(n11683), .ZN(n9040) );
  AND2_X1 U10657 ( .A1(n9077), .A2(n9044), .ZN(n9195) );
  NAND2_X1 U10658 ( .A1(i_ALU_OP[2]), .A2(n10005), .ZN(n9044) );
  NAND2_X1 U10659 ( .A1(n8304), .A2(n8084), .ZN(n9077) );
  OAI211_X1 U10660 ( .C1(n9472), .C2(n9593), .A(n9316), .B(n9315), .ZN(n9833)
         );
  AOI21_X1 U10661 ( .B1(n9328), .B2(n9476), .A(n9314), .ZN(n9315) );
  OAI22_X1 U10662 ( .A1(n9220), .A2(n9313), .B1(n9549), .B2(n9475), .ZN(n9314)
         );
  NAND2_X1 U10663 ( .A1(n9083), .A2(n9082), .ZN(n9475) );
  NAND2_X1 U10664 ( .A1(n8305), .A2(i_ALU_OP[2]), .ZN(n9083) );
  AOI21_X1 U10665 ( .B1(n9711), .B2(n8452), .A(n10285), .ZN(n9313) );
  NOR2_X1 U10666 ( .A1(i_ALU_OP[2]), .A2(n9460), .ZN(n10285) );
  AOI22_X1 U10667 ( .A1(n9325), .A2(n9459), .B1(n9470), .B2(n9686), .ZN(n9316)
         );
  OAI21_X1 U10668 ( .B1(n9477), .B2(n10299), .A(n9312), .ZN(n9470) );
  INV_X1 U10669 ( .A(n9311), .ZN(n9312) );
  AOI21_X1 U10670 ( .B1(i_ALU_OP[2]), .B2(n7799), .A(n9005), .ZN(n9477) );
  NOR2_X1 U10671 ( .A1(i_ALU_OP[2]), .A2(n7693), .ZN(n9005) );
  AOI21_X1 U10672 ( .B1(n11720), .B2(n9225), .A(n9311), .ZN(n9472) );
  NOR2_X1 U10673 ( .A1(n9221), .A2(n11726), .ZN(n9311) );
  INV_X1 U10674 ( .A(n9476), .ZN(n9221) );
  NOR2_X1 U10675 ( .A1(n9460), .A2(n11683), .ZN(n9006) );
  OR2_X1 U10676 ( .A1(n7799), .A2(i_ALU_OP[2]), .ZN(n9082) );
  NAND2_X1 U10677 ( .A1(n8260), .A2(n7974), .ZN(n9054) );
  AOI22_X1 U10678 ( .A1(n10021), .A2(n9828), .B1(n9862), .B2(n10284), .ZN(
        n9353) );
  NAND2_X1 U10679 ( .A1(n9051), .A2(n9050), .ZN(n9052) );
  NAND2_X1 U10680 ( .A1(n7974), .A2(n7860), .ZN(n9051) );
  OR2_X1 U10681 ( .A1(n9064), .A2(n8260), .ZN(n9053) );
  OAI211_X1 U10682 ( .C1(n9310), .C2(n9593), .A(n9309), .B(n9308), .ZN(n9862)
         );
  AOI22_X1 U10683 ( .A1(n9328), .A2(n9562), .B1(n9686), .B2(n9561), .ZN(n9308)
         );
  OAI21_X1 U10684 ( .B1(n9564), .B2(n10299), .A(n9307), .ZN(n9561) );
  OAI21_X1 U10685 ( .B1(n9183), .B2(n8084), .A(n8982), .ZN(n9564) );
  NAND2_X1 U10686 ( .A1(n8084), .A2(n9250), .ZN(n8982) );
  AOI21_X1 U10687 ( .B1(n9526), .B2(n9325), .A(n9306), .ZN(n9309) );
  OAI22_X1 U10688 ( .A1(n9220), .A2(n9557), .B1(n9549), .B2(n9305), .ZN(n9306)
         );
  NAND2_X1 U10689 ( .A1(n8995), .A2(n8994), .ZN(n9305) );
  NAND2_X1 U10690 ( .A1(n8316), .A2(i_ALU_OP[2]), .ZN(n8994) );
  INV_X1 U10691 ( .A(n9527), .ZN(n9526) );
  INV_X1 U10692 ( .A(n9304), .ZN(n9310) );
  OAI21_X1 U10693 ( .B1(n9167), .B2(n11725), .A(n9307), .ZN(n9304) );
  NAND2_X1 U10694 ( .A1(n9562), .A2(n9335), .ZN(n9307) );
  NAND2_X1 U10695 ( .A1(n8992), .A2(n9020), .ZN(n9562) );
  NAND2_X1 U10696 ( .A1(n8991), .A2(n11720), .ZN(n8992) );
  NAND2_X1 U10697 ( .A1(n8995), .A2(n8983), .ZN(n9167) );
  NAND2_X1 U10698 ( .A1(n8452), .A2(n9250), .ZN(n8983) );
  NAND2_X1 U10699 ( .A1(n9161), .A2(n8084), .ZN(n8995) );
  OAI211_X1 U10700 ( .C1(n9503), .C2(n9589), .A(n9303), .B(n9302), .ZN(n9828)
         );
  AOI22_X1 U10701 ( .A1(n9325), .A2(n9516), .B1(n9301), .B2(n9691), .ZN(n9302)
         );
  OAI21_X1 U10702 ( .B1(n11725), .B2(n9199), .A(n9298), .ZN(n9301) );
  NAND2_X1 U10703 ( .A1(n9073), .A2(n8965), .ZN(n9199) );
  NAND2_X1 U10704 ( .A1(n8452), .A2(n8302), .ZN(n8965) );
  AOI21_X1 U10705 ( .B1(n9328), .B2(n9500), .A(n9300), .ZN(n9303) );
  OAI22_X1 U10706 ( .A1(n9220), .A2(n9299), .B1(n9549), .B2(n9495), .ZN(n9300)
         );
  NAND2_X1 U10707 ( .A1(n9074), .A2(n9073), .ZN(n9495) );
  OR2_X1 U10708 ( .A1(n9230), .A2(i_ALU_OP[2]), .ZN(n9073) );
  NAND2_X1 U10709 ( .A1(n8309), .A2(i_ALU_OP[2]), .ZN(n9074) );
  OAI21_X1 U10710 ( .B1(n9230), .B2(n8084), .A(n8963), .ZN(n9498) );
  NAND2_X1 U10711 ( .A1(n8084), .A2(n9246), .ZN(n8963) );
  NAND2_X1 U10712 ( .A1(n9500), .A2(n9335), .ZN(n9298) );
  NAND2_X1 U10713 ( .A1(n9516), .A2(n11682), .ZN(n8964) );
  NAND2_X1 U10714 ( .A1(n9070), .A2(n11720), .ZN(n8962) );
  NAND4_X1 U10715 ( .A1(n9016), .A2(n7970), .A3(n9050), .A4(n9015), .ZN(n9942)
         );
  NAND2_X1 U10716 ( .A1(n7974), .A2(n8084), .ZN(n9015) );
  AOI22_X1 U10717 ( .A1(n9297), .A2(n10023), .B1(n9978), .B2(n9387), .ZN(n9354) );
  OAI211_X1 U10718 ( .C1(n9296), .C2(n9593), .A(n9295), .B(n9294), .ZN(n9387)
         );
  AOI21_X1 U10719 ( .B1(n9328), .B2(n9390), .A(n9293), .ZN(n9294) );
  OAI22_X1 U10720 ( .A1(n9549), .A2(n9389), .B1(n9391), .B2(n9220), .ZN(n9293)
         );
  NAND2_X1 U10721 ( .A1(n9113), .A2(n9112), .ZN(n9389) );
  NAND2_X1 U10722 ( .A1(n7705), .A2(i_ALU_OP[2]), .ZN(n9112) );
  INV_X1 U10723 ( .A(n9560), .ZN(n9549) );
  INV_X1 U10724 ( .A(n9292), .ZN(n9328) );
  AOI22_X1 U10725 ( .A1(n9325), .A2(n9631), .B1(n9686), .B2(n9393), .ZN(n9295)
         );
  INV_X1 U10726 ( .A(n9626), .ZN(n9290) );
  INV_X1 U10727 ( .A(n9289), .ZN(n9325) );
  INV_X1 U10728 ( .A(n9639), .ZN(n9296) );
  OAI21_X1 U10729 ( .B1(n9634), .B2(n11725), .A(n9291), .ZN(n9639) );
  NAND2_X1 U10730 ( .A1(n9390), .A2(n9335), .ZN(n9291) );
  NAND2_X1 U10731 ( .A1(n9631), .A2(n11682), .ZN(n9029) );
  INV_X1 U10732 ( .A(n11685), .ZN(n9020) );
  NAND2_X1 U10733 ( .A1(n9129), .A2(n11720), .ZN(n9021) );
  NAND2_X1 U10734 ( .A1(n9113), .A2(n9022), .ZN(n9634) );
  NAND2_X1 U10735 ( .A1(n8428), .A2(i_ALU_OP[2]), .ZN(n9022) );
  NAND2_X1 U10736 ( .A1(n8303), .A2(n8084), .ZN(n9113) );
  NAND2_X1 U10737 ( .A1(n8967), .A2(n7974), .ZN(n8968) );
  INV_X1 U10738 ( .A(n9050), .ZN(n8967) );
  NAND2_X1 U10739 ( .A1(n9064), .A2(n7860), .ZN(n8969) );
  INV_X1 U10740 ( .A(n9831), .ZN(n9297) );
  AOI211_X1 U10741 ( .C1(n9691), .C2(n9665), .A(n9288), .B(n9287), .ZN(n9831)
         );
  OAI22_X1 U10742 ( .A1(n9289), .A2(n9826), .B1(n9412), .B2(n9589), .ZN(n9287)
         );
  AND2_X1 U10743 ( .A1(n9547), .A2(n9284), .ZN(n9289) );
  OR2_X1 U10744 ( .A1(n7942), .A2(n11725), .ZN(n9284) );
  NAND2_X1 U10745 ( .A1(n8325), .A2(n8452), .ZN(n9547) );
  OAI21_X1 U10746 ( .B1(n9292), .B2(n9668), .A(n9283), .ZN(n9288) );
  AOI22_X1 U10747 ( .A1(n9426), .A2(n9410), .B1(n9560), .B2(n9408), .ZN(n9283)
         );
  NOR2_X1 U10748 ( .A1(n7942), .A2(n11731), .ZN(n9560) );
  OAI21_X1 U10749 ( .B1(i_ALU_OP[2]), .B2(n9826), .A(n9282), .ZN(n9410) );
  NAND2_X1 U10750 ( .A1(n9889), .A2(i_ALU_OP[2]), .ZN(n9282) );
  NOR2_X1 U10751 ( .A1(n9593), .A2(n11731), .ZN(n9426) );
  INV_X1 U10752 ( .A(n9415), .ZN(n9668) );
  AND2_X1 U10753 ( .A1(n9281), .A2(n11726), .ZN(n9292) );
  NAND2_X1 U10754 ( .A1(n8325), .A2(n8084), .ZN(n9281) );
  OAI21_X1 U10755 ( .B1(n9669), .B2(n11725), .A(n9286), .ZN(n9665) );
  NAND2_X1 U10756 ( .A1(n9415), .A2(n9335), .ZN(n9286) );
  INV_X1 U10757 ( .A(n11726), .ZN(n9335) );
  INV_X1 U10758 ( .A(n11722), .ZN(n10299) );
  NAND2_X1 U10759 ( .A1(n8977), .A2(n8976), .ZN(n9415) );
  AOI21_X1 U10760 ( .B1(n7775), .B2(n11682), .A(n11685), .ZN(n8976) );
  NAND2_X1 U10761 ( .A1(n7792), .A2(n11720), .ZN(n8977) );
  NAND2_X1 U10762 ( .A1(n9105), .A2(n8978), .ZN(n9669) );
  NAND2_X1 U10763 ( .A1(n8452), .A2(n9904), .ZN(n8978) );
  NAND2_X1 U10764 ( .A1(n9972), .A2(n8084), .ZN(n9105) );
  NAND2_X1 U10765 ( .A1(n7688), .A2(n7690), .ZN(n9593) );
  NAND2_X1 U10766 ( .A1(n9359), .A2(n9958), .ZN(n9825) );
  NOR2_X1 U10767 ( .A1(i_ALU_OP[0]), .A2(i_ALU_OP[1]), .ZN(n9958) );
  NAND2_X1 U10768 ( .A1(n9280), .A2(n9459), .ZN(n9452) );
  INV_X1 U10769 ( .A(n9279), .ZN(n9280) );
  NAND2_X1 U10770 ( .A1(n9279), .A2(n9460), .ZN(n9453) );
  XNOR2_X1 U10771 ( .A(\DP_OP_751_130_6421/n495 ), .B(n8452), .ZN(n9279) );
  NAND2_X1 U10772 ( .A1(n9278), .A2(n7634), .ZN(n9449) );
  INV_X1 U10773 ( .A(n9276), .ZN(n9278) );
  AND2_X1 U10774 ( .A1(n9841), .A2(n9512), .ZN(n10276) );
  OR2_X1 U10775 ( .A1(n9844), .A2(n9843), .ZN(n9841) );
  NAND2_X1 U10776 ( .A1(n9269), .A2(n9527), .ZN(n9843) );
  NAND2_X1 U10777 ( .A1(n9512), .A2(n9268), .ZN(n9844) );
  NAND2_X1 U10778 ( .A1(n9267), .A2(n9846), .ZN(n9512) );
  OAI21_X1 U10779 ( .B1(n9266), .B2(n9608), .A(n9265), .ZN(n11728) );
  OAI22_X1 U10780 ( .A1(n9264), .A2(n11727), .B1(n9607), .B2(n9584), .ZN(n9265) );
  AOI21_X1 U10781 ( .B1(n9582), .B2(n9580), .A(n9643), .ZN(n9264) );
  NAND2_X1 U10782 ( .A1(n9645), .A2(n9644), .ZN(n9643) );
  XNOR2_X1 U10783 ( .A(n11724), .B(n11723), .ZN(n9644) );
  XNOR2_X1 U10784 ( .A(n9646), .B(n8452), .ZN(n11724) );
  NOR2_X1 U10785 ( .A1(n9897), .A2(n9579), .ZN(n9645) );
  INV_X1 U10786 ( .A(n9263), .ZN(n9579) );
  NOR2_X1 U10787 ( .A1(n9893), .A2(n9886), .ZN(n9897) );
  NAND2_X1 U10788 ( .A1(n9656), .A2(n8301), .ZN(n9886) );
  NAND2_X1 U10789 ( .A1(n9263), .A2(n9262), .ZN(n9893) );
  NAND2_X1 U10790 ( .A1(n9261), .A2(n9904), .ZN(n9263) );
  AND2_X1 U10791 ( .A1(n9262), .A2(n9885), .ZN(n9580) );
  NAND2_X1 U10792 ( .A1(n9260), .A2(n9327), .ZN(n9885) );
  INV_X1 U10793 ( .A(n9656), .ZN(n9260) );
  XNOR2_X1 U10794 ( .A(n9660), .B(i_ALU_OP[2]), .ZN(n9656) );
  NAND2_X1 U10795 ( .A1(n9259), .A2(n9889), .ZN(n9262) );
  INV_X1 U10796 ( .A(n9261), .ZN(n9259) );
  XNOR2_X1 U10797 ( .A(\DP_OP_751_130_6421/n801 ), .B(i_ALU_OP[2]), .ZN(n9261)
         );
  AOI21_X1 U10798 ( .B1(n9258), .B2(n9257), .A(n9256), .ZN(n9582) );
  NOR2_X1 U10799 ( .A1(n9705), .A2(n7693), .ZN(n9256) );
  AND2_X1 U10800 ( .A1(n9706), .A2(n9255), .ZN(n9257) );
  NAND2_X1 U10801 ( .A1(n9705), .A2(n7693), .ZN(n9255) );
  XNOR2_X1 U10802 ( .A(\DP_OP_751_130_6421/n903 ), .B(i_ALU_OP[2]), .ZN(n9705)
         );
  NAND2_X1 U10803 ( .A1(n9734), .A2(n9254), .ZN(n9706) );
  INV_X1 U10804 ( .A(n9253), .ZN(n9254) );
  NAND2_X1 U10805 ( .A1(n9252), .A2(n9998), .ZN(n9734) );
  NAND2_X1 U10806 ( .A1(n9251), .A2(n9753), .ZN(n9998) );
  AND2_X1 U10807 ( .A1(n9750), .A2(n9250), .ZN(n9753) );
  INV_X1 U10808 ( .A(n9249), .ZN(n9750) );
  INV_X1 U10809 ( .A(n9997), .ZN(n9251) );
  NOR2_X1 U10810 ( .A1(n9730), .A2(n9731), .ZN(n9252) );
  AND2_X1 U10811 ( .A1(n9248), .A2(n10005), .ZN(n9731) );
  INV_X1 U10812 ( .A(n9728), .ZN(n9730) );
  NAND2_X1 U10813 ( .A1(n9708), .A2(n9710), .ZN(n9258) );
  AOI21_X1 U10814 ( .B1(n9729), .B2(n9728), .A(n9253), .ZN(n9710) );
  AND2_X1 U10815 ( .A1(n9247), .A2(n7749), .ZN(n9253) );
  XNOR2_X1 U10816 ( .A(n9247), .B(n8302), .ZN(n9728) );
  XNOR2_X1 U10817 ( .A(n9735), .B(n8084), .ZN(n9247) );
  OAI22_X1 U10818 ( .A1(n9997), .A2(n9996), .B1(n9248), .B2(n10005), .ZN(n9729) );
  NAND2_X1 U10819 ( .A1(n9249), .A2(n7774), .ZN(n9996) );
  XNOR2_X1 U10820 ( .A(n9755), .B(n8084), .ZN(n9249) );
  XNOR2_X1 U10821 ( .A(n9248), .B(n10005), .ZN(n9997) );
  XNOR2_X1 U10822 ( .A(\DP_OP_751_130_6421/n1005 ), .B(i_ALU_OP[2]), .ZN(n9248) );
  AOI21_X1 U10823 ( .B1(n9245), .B2(n9244), .A(n9243), .ZN(n9708) );
  NOR2_X1 U10824 ( .A1(n9772), .A2(n9775), .ZN(n9243) );
  AND2_X1 U10825 ( .A1(n9769), .A2(n9242), .ZN(n9244) );
  NAND2_X1 U10826 ( .A1(n9772), .A2(n9775), .ZN(n9242) );
  XNOR2_X1 U10827 ( .A(\DP_OP_751_130_6421/n1107 ), .B(i_ALU_OP[2]), .ZN(n9772) );
  NAND2_X1 U10828 ( .A1(n9241), .A2(n8303), .ZN(n9769) );
  INV_X1 U10829 ( .A(n9240), .ZN(n9241) );
  NAND2_X1 U10830 ( .A1(n9959), .A2(n9771), .ZN(n9245) );
  AND2_X1 U10831 ( .A1(n9776), .A2(n9770), .ZN(n9771) );
  NAND2_X1 U10832 ( .A1(n9240), .A2(n9779), .ZN(n9770) );
  INV_X1 U10833 ( .A(n8303), .ZN(n9779) );
  XNOR2_X1 U10834 ( .A(n9780), .B(n8084), .ZN(n9240) );
  OAI21_X1 U10835 ( .B1(n9961), .B2(n9963), .A(n9768), .ZN(n9776) );
  NAND2_X1 U10836 ( .A1(n9965), .A2(n9238), .ZN(n9959) );
  NOR2_X1 U10837 ( .A1(n9961), .A2(n9781), .ZN(n9238) );
  AND2_X1 U10838 ( .A1(n9239), .A2(n9783), .ZN(n9781) );
  XNOR2_X1 U10839 ( .A(n9784), .B(i_ALU_OP[2]), .ZN(n9239) );
  NAND2_X1 U10840 ( .A1(n9237), .A2(n9972), .ZN(n9768) );
  XNOR2_X1 U10841 ( .A(\DP_OP_751_130_6421/n1209 ), .B(i_ALU_OP[2]), .ZN(n9237) );
  NAND2_X1 U10842 ( .A1(n9236), .A2(n9235), .ZN(n9965) );
  NAND2_X1 U10843 ( .A1(n9793), .A2(n7799), .ZN(n9235) );
  OAI21_X1 U10844 ( .B1(n9793), .B2(n7799), .A(n9792), .ZN(n9236) );
  XNOR2_X1 U10845 ( .A(\DP_OP_751_130_6421/n1311 ), .B(n8084), .ZN(n9792) );
  AOI21_X1 U10846 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9793) );
  NOR2_X1 U10847 ( .A1(n9231), .A2(n9230), .ZN(n9232) );
  NAND2_X1 U10848 ( .A1(n9231), .A2(n9230), .ZN(n9233) );
  XNOR2_X1 U10849 ( .A(n9191), .B(n8084), .ZN(n9231) );
  NAND2_X1 U10850 ( .A1(n9163), .A2(n9183), .ZN(n9927) );
  INV_X1 U10851 ( .A(n9161), .ZN(n9183) );
  INV_X1 U10852 ( .A(n9162), .ZN(n9163) );
  INV_X1 U10853 ( .A(n9951), .ZN(n9932) );
  XNOR2_X1 U10854 ( .A(\DP_OP_751_130_6421/n1413 ), .B(n8084), .ZN(n9929) );
  AND2_X1 U10855 ( .A1(n9162), .A2(n9161), .ZN(n9926) );
  XNOR2_X1 U10856 ( .A(n9182), .B(i_ALU_OP[2]), .ZN(n9162) );
  NAND2_X1 U10857 ( .A1(n9160), .A2(n9159), .ZN(n9928) );
  NAND2_X1 U10858 ( .A1(n9158), .A2(n9157), .ZN(n9159) );
  OAI22_X1 U10859 ( .A1(n9156), .A2(n9155), .B1(n9157), .B2(n9158), .ZN(n9160)
         );
  XNOR2_X1 U10860 ( .A(\DP_OP_751_130_6421/n1515 ), .B(n8452), .ZN(n9158) );
  AOI21_X1 U10861 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9156) );
  NAND2_X1 U10862 ( .A1(n10277), .A2(n9148), .ZN(n9152) );
  NAND2_X1 U10863 ( .A1(n9124), .A2(n9129), .ZN(n9148) );
  XNOR2_X1 U10864 ( .A(n9130), .B(n8452), .ZN(n9124) );
  AND2_X1 U10865 ( .A1(n9123), .A2(n9127), .ZN(n10277) );
  NAND2_X1 U10866 ( .A1(n9122), .A2(n7792), .ZN(n9127) );
  INV_X1 U10867 ( .A(n9126), .ZN(n9122) );
  NAND2_X1 U10868 ( .A1(n9100), .A2(n9811), .ZN(n9123) );
  AND2_X1 U10869 ( .A1(n9805), .A2(n9099), .ZN(n9811) );
  XNOR2_X1 U10870 ( .A(n9126), .B(n7792), .ZN(n9100) );
  XNOR2_X1 U10871 ( .A(n8057), .B(n8452), .ZN(n9126) );
  NAND2_X1 U10872 ( .A1(n9801), .A2(n9806), .ZN(n9809) );
  INV_X1 U10873 ( .A(n9805), .ZN(n9801) );
  XNOR2_X1 U10874 ( .A(n7685), .B(n8084), .ZN(n9805) );
  AOI21_X1 U10875 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9154) );
  AND2_X1 U10876 ( .A1(n9094), .A2(n9093), .ZN(n9096) );
  NAND2_X1 U10877 ( .A1(n9068), .A2(n9070), .ZN(n9093) );
  INV_X1 U10878 ( .A(n8308), .ZN(n9070) );
  NAND2_X1 U10879 ( .A1(n9080), .A2(n9085), .ZN(n9094) );
  INV_X1 U10880 ( .A(n8305), .ZN(n9085) );
  XNOR2_X1 U10881 ( .A(n7690), .B(n8084), .ZN(n9080) );
  NAND2_X1 U10882 ( .A1(n9066), .A2(n8311), .ZN(n9090) );
  INV_X1 U10883 ( .A(n9065), .ZN(n9066) );
  NAND2_X1 U10884 ( .A1(n9067), .A2(n8308), .ZN(n9091) );
  INV_X1 U10885 ( .A(n9068), .ZN(n9067) );
  NAND2_X1 U10886 ( .A1(n9050), .A2(n8966), .ZN(n9068) );
  NAND2_X1 U10887 ( .A1(n7860), .A2(n8084), .ZN(n8966) );
  OR2_X1 U10888 ( .A1(n7860), .A2(n8084), .ZN(n9050) );
  OR2_X1 U10889 ( .A1(n7970), .A2(n8084), .ZN(n9088) );
  NAND2_X1 U10890 ( .A1(n9065), .A2(n9913), .ZN(n9089) );
  INV_X1 U10891 ( .A(n8311), .ZN(n9913) );
  NOR2_X1 U10892 ( .A1(n7974), .A2(i_ALU_OP[2]), .ZN(n9064) );
  INV_X1 U10893 ( .A(n9584), .ZN(n9266) );
  XNOR2_X1 U10894 ( .A(n7782), .B(n8084), .ZN(n9584) );
  NAND2_X1 U10895 ( .A1(n9845), .A2(n9268), .ZN(n11729) );
  NAND2_X1 U10896 ( .A1(n9229), .A2(n7691), .ZN(n9268) );
  INV_X1 U10897 ( .A(n9267), .ZN(n9229) );
  XNOR2_X1 U10898 ( .A(\DP_OP_751_130_6421/n597 ), .B(i_ALU_OP[2]), .ZN(n9267)
         );
  OR2_X1 U10899 ( .A1(n9269), .A2(n9527), .ZN(n9845) );
  XNOR2_X1 U10900 ( .A(n9528), .B(i_ALU_OP[2]), .ZN(n9269) );
  NAND2_X1 U10901 ( .A1(n9276), .A2(n9516), .ZN(n9450) );
  XNOR2_X1 U10902 ( .A(n9517), .B(n8084), .ZN(n9276) );
  XNOR2_X1 U10903 ( .A(n9275), .B(n9358), .ZN(n9370) );
  XNOR2_X1 U10904 ( .A(n9274), .B(n9362), .ZN(n9358) );
  INV_X1 U10905 ( .A(\DP_OP_751_130_6421/n291 ), .ZN(n9362) );
  OAI21_X1 U10906 ( .B1(n9361), .B2(n8084), .A(n11732), .ZN(n9274) );
  NAND2_X1 U10907 ( .A1(n8084), .A2(n9361), .ZN(n11732) );
  NAND2_X1 U10908 ( .A1(n9374), .A2(n9273), .ZN(n9275) );
  INV_X1 U10909 ( .A(n9356), .ZN(n9273) );
  AND2_X1 U10910 ( .A1(n9272), .A2(n9631), .ZN(n9356) );
  INV_X1 U10911 ( .A(n9271), .ZN(n9272) );
  NAND2_X1 U10912 ( .A1(n9376), .A2(n9375), .ZN(n9374) );
  XNOR2_X1 U10913 ( .A(n9271), .B(n9631), .ZN(n9375) );
  XNOR2_X1 U10914 ( .A(n9377), .B(n8452), .ZN(n9271) );
  AOI21_X1 U10915 ( .B1(n9355), .B2(n9826), .A(n9821), .ZN(n9376) );
  NOR2_X1 U10916 ( .A1(n9823), .A2(n9822), .ZN(n9821) );
  NAND2_X1 U10917 ( .A1(n9441), .A2(n8300), .ZN(n9822) );
  XNOR2_X1 U10918 ( .A(n9439), .B(i_ALU_OP[2]), .ZN(n9441) );
  XNOR2_X1 U10919 ( .A(n9355), .B(n9826), .ZN(n9823) );
  XNOR2_X1 U10920 ( .A(\DP_OP_751_130_6421/n393 ), .B(i_ALU_OP[2]), .ZN(n9355)
         );
  NOR2_X1 U10921 ( .A1(n7758), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][18] ) );
  OAI22_X1 U10922 ( .A1(n8901), .A2(n8315), .B1(n8314), .B2(n8902), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][17] ) );
  OAI22_X1 U10923 ( .A1(n8895), .A2(n8311), .B1(n8309), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][16] ) );
  NOR2_X1 U10924 ( .A1(n7763), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][16] ) );
  AND2_X1 U10925 ( .A1(n8991), .A2(n7970), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][0] ) );
  INV_X1 U10926 ( .A(n9910), .ZN(n8991) );
  NOR2_X1 U10927 ( .A1(n8321), .A2(n8316), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][2] ) );
  OAI22_X1 U10928 ( .A1(n7637), .A2(n8316), .B1(n8322), .B2(n8311), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][3] ) );
  OAI22_X1 U10929 ( .A1(n7733), .A2(n9910), .B1(n8311), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][5] ) );
  OAI22_X1 U10930 ( .A1(n7741), .A2(n8305), .B1(n8260), .B2(n9806), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][4] ) );
  NOR2_X1 U10931 ( .A1(n8331), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][6] ) );
  OAI22_X1 U10932 ( .A1(n8872), .A2(n8315), .B1(n8312), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][7] ) );
  OAI22_X1 U10933 ( .A1(n7734), .A2(n8311), .B1(n8309), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][6] ) );
  OAI22_X1 U10934 ( .A1(n7741), .A2(n9806), .B1(n8260), .B2(n9125), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][5] ) );
  OAI22_X1 U10935 ( .A1(n8334), .A2(n8315), .B1(n8312), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][9] ) );
  OAI22_X1 U10936 ( .A1(n7743), .A2(n8311), .B1(n8308), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][8] ) );
  OAI22_X1 U10937 ( .A1(n8327), .A2(n8310), .B1(n8306), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][7] ) );
  OAI22_X1 U10938 ( .A1(n7740), .A2(n9125), .B1(n8260), .B2(n7705), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][6] ) );
  OAI22_X1 U10939 ( .A1(n7637), .A2(n8305), .B1(n8321), .B2(n9806), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][6] ) );
  NOR2_X1 U10940 ( .A1(n8884), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][10] ) );
  OAI22_X1 U10941 ( .A1(n7742), .A2(n9910), .B1(n8311), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][11] ) );
  OAI22_X1 U10942 ( .A1(n8878), .A2(n8314), .B1(n8308), .B2(n8879), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][10] ) );
  OAI22_X1 U10943 ( .A1(n7743), .A2(n8309), .B1(n8305), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][9] ) );
  OAI22_X1 U10944 ( .A1(n7733), .A2(n8305), .B1(n9806), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][8] ) );
  OAI22_X1 U10945 ( .A1(n7741), .A2(n7705), .B1(n8260), .B2(n9157), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][7] ) );
  OAI22_X1 U10946 ( .A1(n8317), .A2(n9806), .B1(n8324), .B2(n9125), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][7] ) );
  NOR2_X1 U10947 ( .A1(n7760), .A2(n9910), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][12] ) );
  OAI22_X1 U10948 ( .A1(n8891), .A2(n9910), .B1(n8311), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][13] ) );
  OAI22_X1 U10949 ( .A1(n7742), .A2(n8311), .B1(n8308), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][12] ) );
  OAI22_X1 U10950 ( .A1(n8878), .A2(n8309), .B1(n8305), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][11] ) );
  OAI22_X1 U10951 ( .A1(n8872), .A2(n8305), .B1(n9806), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][10] ) );
  OAI22_X1 U10952 ( .A1(n8327), .A2(n9806), .B1(n9125), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][9] ) );
  OAI22_X1 U10953 ( .A1(n7741), .A2(n9157), .B1(n9161), .B2(n8260), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][8] ) );
  OAI22_X1 U10954 ( .A1(n8318), .A2(n9125), .B1(n8324), .B2(n7705), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][8] ) );
  NOR2_X1 U10955 ( .A1(n7765), .A2(n8316), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][14] ) );
  OAI22_X1 U10956 ( .A1(n8891), .A2(n8308), .B1(n8307), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][15] ) );
  OAI22_X1 U10957 ( .A1(n8895), .A2(n8316), .B1(n8311), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][15] ) );
  OAI22_X1 U10958 ( .A1(n7742), .A2(n8306), .B1(n9806), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][14] ) );
  OAI22_X1 U10959 ( .A1(n8891), .A2(n8313), .B1(n8309), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][14] ) );
  OAI22_X1 U10960 ( .A1(n8333), .A2(n9806), .B1(n9125), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][13] ) );
  OAI22_X1 U10961 ( .A1(n7742), .A2(n8308), .B1(n8307), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][13] ) );
  OAI22_X1 U10962 ( .A1(n7743), .A2(n9125), .B1(n7705), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][12] ) );
  OAI22_X1 U10963 ( .A1(n8333), .A2(n8305), .B1(n9806), .B2(n8879), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][12] ) );
  OAI22_X1 U10964 ( .A1(n7734), .A2(n7705), .B1(n9157), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][11] ) );
  OAI22_X1 U10965 ( .A1(n8872), .A2(n9806), .B1(n9125), .B2(n8331), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][11] ) );
  OAI22_X1 U10966 ( .A1(n7740), .A2(n9951), .B1(n8260), .B2(n8941), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][10] ) );
  OAI22_X1 U10967 ( .A1(n9157), .A2(n8319), .B1(n8324), .B2(n9161), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][10] ) );
  OAI22_X1 U10968 ( .A1(n8327), .A2(n9125), .B1(n7705), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][10] ) );
  OAI22_X1 U10969 ( .A1(n7740), .A2(n9161), .B1(n8261), .B2(n9951), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][9] ) );
  OAI22_X1 U10970 ( .A1(n8319), .A2(n7705), .B1(n8324), .B2(n9157), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][9] ) );
  OAI22_X1 U10971 ( .A1(n8908), .A2(n9910), .B1(n8311), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][19] ) );
  OAI22_X1 U10972 ( .A1(n8901), .A2(n8311), .B1(n8308), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][18] ) );
  OAI22_X1 U10973 ( .A1(n8895), .A2(n8310), .B1(n8306), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][17] ) );
  OAI22_X1 U10974 ( .A1(n8891), .A2(n8305), .B1(n9806), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][16] ) );
  OAI22_X1 U10975 ( .A1(n7742), .A2(n9806), .B1(n9125), .B2(n8335), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][15] ) );
  OAI22_X1 U10976 ( .A1(n8334), .A2(n9125), .B1(n7705), .B2(n8879), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][14] ) );
  OAI22_X1 U10977 ( .A1(n7743), .A2(n7705), .B1(n9157), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][13] ) );
  OAI22_X1 U10978 ( .A1(n8326), .A2(n9157), .B1(n9161), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][12] ) );
  OAI22_X1 U10979 ( .A1(n7740), .A2(n8941), .B1(n8260), .B2(n9796), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][11] ) );
  OAI22_X1 U10980 ( .A1(n8319), .A2(n9161), .B1(n8323), .B2(n9951), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][11] ) );
  NOR2_X1 U10981 ( .A1(n8336), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][20] ) );
  OAI22_X1 U10982 ( .A1(n8915), .A2(n8315), .B1(n8314), .B2(n8336), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][21] ) );
  OAI22_X1 U10983 ( .A1(n8908), .A2(n8314), .B1(n8308), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][20] ) );
  OAI22_X1 U10984 ( .A1(n8901), .A2(n8309), .B1(n8306), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][19] ) );
  OAI22_X1 U10985 ( .A1(n8895), .A2(n8307), .B1(n9806), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][18] ) );
  OAI22_X1 U10986 ( .A1(n8891), .A2(n9806), .B1(n9125), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][17] ) );
  OAI22_X1 U10987 ( .A1(n7742), .A2(n9125), .B1(n7705), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][16] ) );
  OAI22_X1 U10988 ( .A1(n8333), .A2(n7705), .B1(n9157), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][15] ) );
  OAI22_X1 U10989 ( .A1(n7743), .A2(n9157), .B1(n9161), .B2(n8331), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][14] ) );
  OAI22_X1 U10990 ( .A1(n8326), .A2(n9161), .B1(n9951), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][13] ) );
  OAI22_X1 U10991 ( .A1(n7740), .A2(n9796), .B1(n8260), .B2(n9783), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][12] ) );
  OAI22_X1 U10992 ( .A1(n8318), .A2(n9951), .B1(n8324), .B2(n8941), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][12] ) );
  NOR2_X1 U10993 ( .A1(n8923), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][22] ) );
  OAI22_X1 U10994 ( .A1(n8922), .A2(n8316), .B1(n8311), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][23] ) );
  BUF_X1 U10995 ( .A(n9910), .Z(n8316) );
  OAI22_X1 U10996 ( .A1(n8915), .A2(n8314), .B1(n8308), .B2(n8916), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][22] ) );
  OAI22_X1 U10997 ( .A1(n8908), .A2(n8308), .B1(n8305), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][21] ) );
  OAI22_X1 U10998 ( .A1(n8901), .A2(n8305), .B1(n9806), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][20] ) );
  OAI22_X1 U10999 ( .A1(n8895), .A2(n9806), .B1(n9125), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][19] ) );
  OAI22_X1 U11000 ( .A1(n8891), .A2(n9125), .B1(n7705), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][18] ) );
  OAI22_X1 U11001 ( .A1(n7742), .A2(n7705), .B1(n9157), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][17] ) );
  OAI22_X1 U11002 ( .A1(n8333), .A2(n9157), .B1(n9161), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][16] ) );
  OAI22_X1 U11003 ( .A1(n7743), .A2(n9161), .B1(n8304), .B2(n8331), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][15] ) );
  OAI22_X1 U11004 ( .A1(n8326), .A2(n9951), .B1(n8941), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][14] ) );
  OAI22_X1 U11005 ( .A1(n7740), .A2(n9783), .B1(n8260), .B2(n9972), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][13] ) );
  NOR2_X1 U11006 ( .A1(n8927), .A2(n9910), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][24] ) );
  OAI22_X1 U11007 ( .A1(n8926), .A2(n8315), .B1(n8313), .B2(n8927), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][25] ) );
  OAI22_X1 U11008 ( .A1(n8922), .A2(n8312), .B1(n8310), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][24] ) );
  BUF_X1 U11009 ( .A(n8311), .Z(n8312) );
  OAI22_X1 U11010 ( .A1(n8915), .A2(n8308), .B1(n8305), .B2(n8336), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][23] ) );
  OAI22_X1 U11011 ( .A1(n8908), .A2(n8306), .B1(n9806), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][22] ) );
  OAI22_X1 U11012 ( .A1(n8901), .A2(n9806), .B1(n9125), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][21] ) );
  OAI22_X1 U11013 ( .A1(n8895), .A2(n9125), .B1(n7705), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][20] ) );
  OAI22_X1 U11014 ( .A1(n8891), .A2(n7705), .B1(n9157), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][19] ) );
  OAI22_X1 U11015 ( .A1(n7742), .A2(n9157), .B1(n9161), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][18] ) );
  OAI22_X1 U11016 ( .A1(n8333), .A2(n9161), .B1(n8304), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][17] ) );
  OAI22_X1 U11017 ( .A1(n7743), .A2(n9951), .B1(n8941), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][16] ) );
  OAI22_X1 U11018 ( .A1(n8326), .A2(n8941), .B1(n9796), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][15] ) );
  NOR2_X1 U11019 ( .A1(n8931), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[13][26] ) );
  OAI22_X1 U11020 ( .A1(n8930), .A2(n8315), .B1(n8313), .B2(n8931), .ZN(
        \DataPath/ALUhw/MULT/mux_out[13][27] ) );
  BUF_X1 U11021 ( .A(n8311), .Z(n8313) );
  OAI22_X1 U11022 ( .A1(n8926), .A2(n8311), .B1(n8308), .B2(n8927), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][26] ) );
  OAI22_X1 U11023 ( .A1(n8922), .A2(n8308), .B1(n8306), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][25] ) );
  BUF_X1 U11024 ( .A(n8305), .Z(n8306) );
  OAI22_X1 U11025 ( .A1(n8915), .A2(n8307), .B1(n9806), .B2(n8336), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][24] ) );
  OAI22_X1 U11026 ( .A1(n8908), .A2(n9806), .B1(n9125), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][23] ) );
  OAI22_X1 U11027 ( .A1(n8901), .A2(n9125), .B1(n7705), .B2(n8902), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][22] ) );
  OAI22_X1 U11028 ( .A1(n8895), .A2(n7705), .B1(n9157), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][21] ) );
  OAI22_X1 U11029 ( .A1(n8891), .A2(n9157), .B1(n9161), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][20] ) );
  OAI22_X1 U11030 ( .A1(n7742), .A2(n9161), .B1(n8304), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][19] ) );
  OAI22_X1 U11031 ( .A1(n8333), .A2(n9951), .B1(n8941), .B2(n8879), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][18] ) );
  OAI22_X1 U11032 ( .A1(n7743), .A2(n8941), .B1(n9796), .B2(n8331), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][17] ) );
  OAI22_X1 U11033 ( .A1(n7733), .A2(n9796), .B1(n9783), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][16] ) );
  OAI22_X1 U11034 ( .A1(n7740), .A2(n8303), .B1(n8261), .B2(n9775), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][15] ) );
  OAI22_X1 U11035 ( .A1(n8317), .A2(n9783), .B1(n8321), .B2(n9972), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][15] ) );
  NOR2_X1 U11036 ( .A1(n8938), .A2(n8316), .ZN(
        \DataPath/ALUhw/MULT/mux_out[14][28] ) );
  OAI22_X1 U11037 ( .A1(n8937), .A2(n8315), .B1(n8314), .B2(n8938), .ZN(
        \DataPath/ALUhw/MULT/mux_out[14][29] ) );
  OAI22_X1 U11038 ( .A1(n8930), .A2(n8314), .B1(n8309), .B2(n8931), .ZN(
        \DataPath/ALUhw/MULT/mux_out[13][28] ) );
  BUF_X1 U11039 ( .A(n8311), .Z(n8314) );
  OAI22_X1 U11040 ( .A1(n8926), .A2(n8310), .B1(n8307), .B2(n8927), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][27] ) );
  BUF_X1 U11041 ( .A(n8308), .Z(n8310) );
  OAI22_X1 U11042 ( .A1(n8922), .A2(n8305), .B1(n9806), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][26] ) );
  OAI22_X1 U11043 ( .A1(n8915), .A2(n9806), .B1(n9125), .B2(n8336), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][25] ) );
  OAI22_X1 U11044 ( .A1(n8908), .A2(n9125), .B1(n7705), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][24] ) );
  OAI22_X1 U11045 ( .A1(n8901), .A2(n7705), .B1(n9157), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][23] ) );
  OAI22_X1 U11046 ( .A1(n8895), .A2(n9157), .B1(n9161), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][22] ) );
  OAI22_X1 U11047 ( .A1(n8891), .A2(n9161), .B1(n9951), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][21] ) );
  OAI22_X1 U11048 ( .A1(n7742), .A2(n9951), .B1(n8941), .B2(n8884), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][20] ) );
  OAI22_X1 U11049 ( .A1(n8334), .A2(n8941), .B1(n9796), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][19] ) );
  OAI22_X1 U11050 ( .A1(n7743), .A2(n9796), .B1(n9783), .B2(n8331), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][18] ) );
  OAI22_X1 U11051 ( .A1(n8327), .A2(n9783), .B1(n9972), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][17] ) );
  OAI22_X1 U11052 ( .A1(n7740), .A2(n9775), .B1(n8260), .B2(n9250), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][16] ) );
  OAI22_X1 U11053 ( .A1(n8319), .A2(n9972), .B1(n8321), .B2(n8303), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][16] ) );
  NOR2_X1 U11054 ( .A1(n8942), .A2(n8315), .ZN(
        \DataPath/ALUhw/MULT/mux_out[15][30] ) );
  OAI22_X1 U11055 ( .A1(n7740), .A2(n9026), .B1(n8260), .B2(n9592), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][31] ) );
  OAI22_X1 U11056 ( .A1(n8319), .A2(n8300), .B1(n8321), .B2(n9826), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][31] ) );
  OAI22_X1 U11057 ( .A1(n8327), .A2(n9277), .B1(n9460), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][31] ) );
  OAI22_X1 U11058 ( .A1(n8332), .A2(n9527), .B1(n8331), .B2(n9846), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][31] ) );
  OAI22_X1 U11059 ( .A1(n8333), .A2(n8428), .B1(n9608), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][31] ) );
  OAI22_X1 U11060 ( .A1(n7742), .A2(n8301), .B1(n9904), .B2(n8884), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][31] ) );
  OAI22_X1 U11061 ( .A1(n8891), .A2(n9246), .B1(n7693), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][31] ) );
  OAI22_X1 U11062 ( .A1(n8895), .A2(n9250), .B1(n10005), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][31] ) );
  OAI22_X1 U11063 ( .A1(n8901), .A2(n8303), .B1(n9775), .B2(n8902), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][31] ) );
  OAI22_X1 U11064 ( .A1(n8908), .A2(n9783), .B1(n9972), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][31] ) );
  OAI22_X1 U11065 ( .A1(n8915), .A2(n8941), .B1(n9796), .B2(n8916), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][31] ) );
  OAI22_X1 U11066 ( .A1(n8922), .A2(n9161), .B1(n8304), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][31] ) );
  OAI22_X1 U11067 ( .A1(n8926), .A2(n7705), .B1(n9157), .B2(n8927), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][31] ) );
  OAI22_X1 U11068 ( .A1(n8930), .A2(n9806), .B1(n9125), .B2(n8931), .ZN(
        \DataPath/ALUhw/MULT/mux_out[13][31] ) );
  OAI22_X1 U11069 ( .A1(n8937), .A2(n8308), .B1(n8305), .B2(n8938), .ZN(
        \DataPath/ALUhw/MULT/mux_out[14][31] ) );
  XNOR2_X1 U11070 ( .A(\DP_OP_751_130_6421/n393 ), .B(n9377), .ZN(n8942) );
  NAND2_X1 U11071 ( .A1(\DataPath/i_PIPLIN_A[0] ), .A2(n7692), .ZN(n8856) );
  NAND2_X1 U11072 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[0] ), .ZN(n8857) );
  OAI21_X1 U11073 ( .B1(n8190), .B2(n7907), .A(n8940), .ZN(n9377) );
  OAI22_X1 U11074 ( .A1(n8318), .A2(n9460), .B1(n8322), .B2(n8300), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][30] ) );
  OAI22_X1 U11075 ( .A1(n8327), .A2(n9846), .B1(n9277), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][30] ) );
  OAI22_X1 U11076 ( .A1(n8872), .A2(n9608), .B1(n7746), .B2(n9527), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][30] ) );
  OAI22_X1 U11077 ( .A1(n8334), .A2(n9904), .B1(n8428), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][30] ) );
  OAI22_X1 U11078 ( .A1(n7742), .A2(n7693), .B1(n8301), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][30] ) );
  OAI22_X1 U11079 ( .A1(n8891), .A2(n10005), .B1(n9246), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][30] ) );
  OAI22_X1 U11080 ( .A1(n8895), .A2(n9775), .B1(n9250), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][30] ) );
  OAI22_X1 U11081 ( .A1(n8901), .A2(n9972), .B1(n8303), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][30] ) );
  OAI22_X1 U11082 ( .A1(n8908), .A2(n9796), .B1(n9783), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][30] ) );
  OAI22_X1 U11083 ( .A1(n8915), .A2(n8304), .B1(n8941), .B2(n8916), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][30] ) );
  OAI22_X1 U11084 ( .A1(n8922), .A2(n9157), .B1(n9161), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][30] ) );
  OAI22_X1 U11085 ( .A1(n8926), .A2(n9125), .B1(n7705), .B2(n8927), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][30] ) );
  OAI22_X1 U11086 ( .A1(n8930), .A2(n8305), .B1(n9806), .B2(n8931), .ZN(
        \DataPath/ALUhw/MULT/mux_out[13][30] ) );
  OAI22_X1 U11087 ( .A1(n8937), .A2(n8311), .B1(n8309), .B2(n8938), .ZN(
        \DataPath/ALUhw/MULT/mux_out[14][30] ) );
  NAND2_X1 U11088 ( .A1(\DataPath/i_PIPLIN_A[1] ), .A2(n7692), .ZN(n8854) );
  NAND2_X1 U11089 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[1] ), .ZN(n8855) );
  OAI21_X1 U11090 ( .B1(n8936), .B2(\DP_OP_751_130_6421/n495 ), .A(n8935), 
        .ZN(n8937) );
  OAI21_X1 U11091 ( .B1(n9824), .B2(\DP_OP_751_130_6421/n495 ), .A(n8934), 
        .ZN(n8935) );
  NAND2_X1 U11092 ( .A1(n9824), .A2(n9439), .ZN(n8934) );
  INV_X1 U11093 ( .A(n9439), .ZN(n8936) );
  OAI21_X1 U11094 ( .B1(n8188), .B2(n7907), .A(n8933), .ZN(n9439) );
  OAI22_X1 U11095 ( .A1(n9277), .A2(n7637), .B1(n7656), .B2(n9460), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][29] ) );
  OAI22_X1 U11096 ( .A1(n8868), .A2(n9527), .B1(n9846), .B2(n8329), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][29] ) );
  OAI22_X1 U11097 ( .A1(n8872), .A2(n8428), .B1(n7746), .B2(n9608), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][29] ) );
  OAI22_X1 U11098 ( .A1(n8333), .A2(n8301), .B1(n9904), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][29] ) );
  OAI22_X1 U11099 ( .A1(n7742), .A2(n8302), .B1(n7693), .B2(n8335), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][29] ) );
  OAI22_X1 U11100 ( .A1(n8891), .A2(n9250), .B1(n10005), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][29] ) );
  OAI22_X1 U11101 ( .A1(n8895), .A2(n8303), .B1(n9775), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][29] ) );
  OAI22_X1 U11102 ( .A1(n8901), .A2(n9783), .B1(n9972), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][29] ) );
  OAI22_X1 U11103 ( .A1(n8908), .A2(n8941), .B1(n9796), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][29] ) );
  OAI22_X1 U11104 ( .A1(n8915), .A2(n9161), .B1(n9951), .B2(n8916), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][29] ) );
  OAI22_X1 U11105 ( .A1(n8922), .A2(n7705), .B1(n9157), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][29] ) );
  OAI22_X1 U11106 ( .A1(n8926), .A2(n9806), .B1(n9125), .B2(n8927), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][29] ) );
  OAI22_X1 U11107 ( .A1(n8930), .A2(n8308), .B1(n8305), .B2(n8931), .ZN(
        \DataPath/ALUhw/MULT/mux_out[13][29] ) );
  NAND2_X1 U11108 ( .A1(\DataPath/i_PIPLIN_A[2] ), .A2(n7692), .ZN(n8852) );
  NAND2_X1 U11109 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[2] ), .ZN(n8853) );
  NAND2_X1 U11110 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[27] ), .ZN(n8928)
         );
  OAI21_X1 U11111 ( .B1(n8186), .B2(n7907), .A(n8929), .ZN(n9517) );
  OAI22_X1 U11112 ( .A1(n9608), .A2(n8868), .B1(n9527), .B2(n8329), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][28] ) );
  OAI22_X1 U11113 ( .A1(n8872), .A2(n9904), .B1(n7746), .B2(n8428), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][28] ) );
  OAI22_X1 U11114 ( .A1(n8333), .A2(n7693), .B1(n8301), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][28] ) );
  OAI22_X1 U11115 ( .A1(n7742), .A2(n10005), .B1(n8302), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][28] ) );
  OAI22_X1 U11116 ( .A1(n8891), .A2(n9775), .B1(n9250), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][28] ) );
  OAI22_X1 U11117 ( .A1(n8895), .A2(n9972), .B1(n8303), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][28] ) );
  OAI22_X1 U11118 ( .A1(n8901), .A2(n9796), .B1(n9783), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][28] ) );
  OAI22_X1 U11119 ( .A1(n8908), .A2(n8304), .B1(n8941), .B2(n8909), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][28] ) );
  OAI22_X1 U11120 ( .A1(n8915), .A2(n9157), .B1(n9161), .B2(n8336), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][28] ) );
  OAI22_X1 U11121 ( .A1(n8922), .A2(n9125), .B1(n7705), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][28] ) );
  OAI22_X1 U11122 ( .A1(n8926), .A2(n8307), .B1(n9806), .B2(n8927), .ZN(
        \DataPath/ALUhw/MULT/mux_out[12][28] ) );
  NAND2_X1 U11123 ( .A1(\DataPath/i_PIPLIN_A[3] ), .A2(n465), .ZN(n8850) );
  NAND2_X1 U11124 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[3] ), .ZN(n8851) );
  NAND2_X1 U11125 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[25] ), .ZN(n8924)
         );
  OAI21_X1 U11126 ( .B1(n8157), .B2(n7907), .A(n8925), .ZN(n9528) );
  NAND2_X1 U11127 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[24] ), .ZN(n8925)
         );
  OAI22_X1 U11128 ( .A1(n7733), .A2(n8428), .B1(n9608), .B2(n7687), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][27] ) );
  OAI22_X1 U11129 ( .A1(n8872), .A2(n8301), .B1(n7746), .B2(n9904), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][27] ) );
  OAI22_X1 U11130 ( .A1(n8333), .A2(n8302), .B1(n7693), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][27] ) );
  OAI22_X1 U11131 ( .A1(n7742), .A2(n9250), .B1(n10005), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][27] ) );
  OAI22_X1 U11132 ( .A1(n8891), .A2(n8303), .B1(n9775), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][27] ) );
  OAI22_X1 U11133 ( .A1(n8895), .A2(n9783), .B1(n9972), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][27] ) );
  OAI22_X1 U11134 ( .A1(n8901), .A2(n8941), .B1(n9796), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][27] ) );
  OAI22_X1 U11135 ( .A1(n8908), .A2(n9161), .B1(n8304), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][27] ) );
  OAI22_X1 U11136 ( .A1(n8915), .A2(n7705), .B1(n9157), .B2(n8336), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][27] ) );
  OAI22_X1 U11137 ( .A1(n8922), .A2(n9806), .B1(n9125), .B2(n8923), .ZN(
        \DataPath/ALUhw/MULT/mux_out[11][27] ) );
  OAI21_X1 U11138 ( .B1(n8921), .B2(\DP_OP_751_130_6421/n801 ), .A(n8920), 
        .ZN(n8922) );
  OAI21_X1 U11139 ( .B1(n9609), .B2(\DP_OP_751_130_6421/n801 ), .A(n8919), 
        .ZN(n8920) );
  NAND2_X1 U11140 ( .A1(n9609), .A2(n9646), .ZN(n8919) );
  NAND2_X1 U11141 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[23] ), .ZN(n8917)
         );
  INV_X1 U11142 ( .A(n9646), .ZN(n8921) );
  OAI21_X1 U11143 ( .B1(n8155), .B2(n7907), .A(n8918), .ZN(n9646) );
  NAND2_X1 U11144 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[22] ), .ZN(n8918)
         );
  OAI22_X1 U11145 ( .A1(n8858), .A2(n9846), .B1(n8974), .B2(n9277), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][26] ) );
  OAI22_X1 U11146 ( .A1(n7637), .A2(n9608), .B1(n7689), .B2(n9527), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][26] ) );
  OAI22_X1 U11147 ( .A1(n7734), .A2(n9904), .B1(n8428), .B2(n7687), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][26] ) );
  OAI22_X1 U11148 ( .A1(n8872), .A2(n7693), .B1(n7746), .B2(n8301), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][26] ) );
  OAI22_X1 U11149 ( .A1(n8333), .A2(n10005), .B1(n8302), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][26] ) );
  OAI22_X1 U11150 ( .A1(n7742), .A2(n9775), .B1(n9250), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][26] ) );
  OAI22_X1 U11151 ( .A1(n8891), .A2(n9972), .B1(n8303), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][26] ) );
  OAI22_X1 U11152 ( .A1(n8895), .A2(n9796), .B1(n9783), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][26] ) );
  OAI22_X1 U11153 ( .A1(n8901), .A2(n8304), .B1(n8941), .B2(n8902), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][26] ) );
  OAI22_X1 U11154 ( .A1(n8908), .A2(n9157), .B1(n9161), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][26] ) );
  OAI22_X1 U11155 ( .A1(n8915), .A2(n9125), .B1(n7705), .B2(n8336), .ZN(
        \DataPath/ALUhw/MULT/mux_out[10][26] ) );
  NAND2_X1 U11156 ( .A1(n8849), .A2(n8848), .ZN(n9121) );
  NAND2_X1 U11157 ( .A1(\DataPath/i_PIPLIN_A[5] ), .A2(n7732), .ZN(n8848) );
  NAND2_X1 U11158 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[5] ), .ZN(n8849) );
  OAI21_X1 U11159 ( .B1(n9712), .B2(n9660), .A(n8914), .ZN(n8915) );
  OAI21_X1 U11160 ( .B1(n9712), .B2(\DP_OP_751_130_6421/n801 ), .A(n8913), 
        .ZN(n8914) );
  NAND2_X1 U11161 ( .A1(n8912), .A2(\DP_OP_751_130_6421/n801 ), .ZN(n8913) );
  INV_X1 U11162 ( .A(n9660), .ZN(n8912) );
  NAND2_X1 U11163 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[21] ), .ZN(n8910)
         );
  OAI21_X1 U11164 ( .B1(n8153), .B2(n7907), .A(n8911), .ZN(n9660) );
  NAND2_X1 U11165 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[20] ), .ZN(n8911)
         );
  INV_X1 U11166 ( .A(\DP_OP_751_130_6421/n903 ), .ZN(n9712) );
  OAI22_X1 U11167 ( .A1(n7741), .A2(n9527), .B1(n8261), .B2(n9846), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][25] ) );
  OAI22_X1 U11168 ( .A1(n8317), .A2(n8428), .B1(n7689), .B2(n9608), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][25] ) );
  OAI22_X1 U11169 ( .A1(n8326), .A2(n8301), .B1(n9904), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][25] ) );
  OAI22_X1 U11170 ( .A1(n8332), .A2(n8302), .B1(n8331), .B2(n7693), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][25] ) );
  OAI22_X1 U11171 ( .A1(n8334), .A2(n9250), .B1(n10005), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][25] ) );
  OAI22_X1 U11172 ( .A1(n7742), .A2(n8303), .B1(n9775), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][25] ) );
  OAI22_X1 U11173 ( .A1(n8891), .A2(n9783), .B1(n9972), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][25] ) );
  OAI22_X1 U11174 ( .A1(n8895), .A2(n8941), .B1(n9796), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][25] ) );
  OAI22_X1 U11175 ( .A1(n8901), .A2(n9161), .B1(n8304), .B2(n7763), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][25] ) );
  OAI22_X1 U11176 ( .A1(n8908), .A2(n7705), .B1(n9157), .B2(n7758), .ZN(
        \DataPath/ALUhw/MULT/mux_out[9][25] ) );
  XNOR2_X1 U11177 ( .A(\DP_OP_751_130_6421/n1005 ), .B(n9735), .ZN(n8909) );
  NAND2_X1 U11178 ( .A1(\DataPath/i_PIPLIN_A[6] ), .A2(n7692), .ZN(n8846) );
  NAND2_X1 U11179 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[6] ), .ZN(n8847) );
  OAI21_X1 U11180 ( .B1(n8449), .B2(\DP_OP_751_130_6421/n903 ), .A(n8906), 
        .ZN(n8907) );
  NAND2_X1 U11181 ( .A1(n8905), .A2(\DP_OP_751_130_6421/n903 ), .ZN(n8906) );
  INV_X1 U11182 ( .A(n9735), .ZN(n8905) );
  NAND2_X1 U11183 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[19] ), .ZN(n8903)
         );
  OAI21_X1 U11184 ( .B1(n8152), .B2(n7940), .A(n8904), .ZN(n9735) );
  NAND2_X1 U11185 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[18] ), .ZN(n8904)
         );
  OAI22_X1 U11186 ( .A1(n7741), .A2(n9608), .B1(n8261), .B2(n9527), .ZN(
        \DataPath/ALUhw/MULT/mux_out[0][24] ) );
  OAI22_X1 U11187 ( .A1(n8319), .A2(n9904), .B1(n7656), .B2(n8428), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][24] ) );
  OAI22_X1 U11188 ( .A1(n8326), .A2(n7693), .B1(n8301), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][24] ) );
  OAI22_X1 U11189 ( .A1(n8332), .A2(n10005), .B1(n8331), .B2(n8302), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][24] ) );
  OAI22_X1 U11190 ( .A1(n8334), .A2(n9775), .B1(n9250), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][24] ) );
  BUF_X1 U11191 ( .A(n8878), .Z(n8334) );
  OAI22_X1 U11192 ( .A1(n7742), .A2(n9972), .B1(n8303), .B2(n7744), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][24] ) );
  OAI22_X1 U11193 ( .A1(n8891), .A2(n9796), .B1(n9783), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][24] ) );
  OAI22_X1 U11194 ( .A1(n8895), .A2(n8304), .B1(n8941), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][24] ) );
  OAI22_X1 U11195 ( .A1(n8901), .A2(n9157), .B1(n9161), .B2(n8902), .ZN(
        \DataPath/ALUhw/MULT/mux_out[8][24] ) );
  XNOR2_X1 U11196 ( .A(\DP_OP_751_130_6421/n1107 ), .B(n9755), .ZN(n8902) );
  OAI21_X1 U11197 ( .B1(n7767), .B2(\DP_OP_751_130_6421/n1005 ), .A(n8899), 
        .ZN(n8900) );
  NAND2_X1 U11198 ( .A1(n8898), .A2(\DP_OP_751_130_6421/n1005 ), .ZN(n8899) );
  INV_X1 U11199 ( .A(n9755), .ZN(n8898) );
  OAI21_X1 U11200 ( .B1(n8150), .B2(n7940), .A(n8897), .ZN(n9755) );
  NAND2_X1 U11201 ( .A1(n7940), .A2(\DataPath/i_PIPLIN_IN2[16] ), .ZN(n8897)
         );
  OAI22_X1 U11202 ( .A1(n8319), .A2(n8301), .B1(n8322), .B2(n9904), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][23] ) );
  OAI22_X1 U11203 ( .A1(n7734), .A2(n8302), .B1(n7693), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][23] ) );
  OAI22_X1 U11204 ( .A1(n8332), .A2(n9250), .B1(n8331), .B2(n10005), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][23] ) );
  OAI22_X1 U11205 ( .A1(n8333), .A2(n8303), .B1(n9775), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][23] ) );
  OAI22_X1 U11206 ( .A1(n7742), .A2(n9783), .B1(n9972), .B2(n8335), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][23] ) );
  OAI22_X1 U11207 ( .A1(n8891), .A2(n8941), .B1(n9796), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][23] ) );
  OAI22_X1 U11208 ( .A1(n8895), .A2(n9161), .B1(n8304), .B2(n7765), .ZN(
        \DataPath/ALUhw/MULT/mux_out[7][23] ) );
  NAND2_X1 U11209 ( .A1(\DataPath/i_PIPLIN_A[8] ), .A2(n7732), .ZN(n8844) );
  NAND2_X1 U11210 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[8] ), .ZN(n8845) );
  OAI21_X1 U11211 ( .B1(n7767), .B2(n9780), .A(n8893), .ZN(n8894) );
  NAND2_X1 U11212 ( .A1(n7767), .A2(\DP_OP_751_130_6421/n1209 ), .ZN(n8893) );
  OAI22_X1 U11213 ( .A1(n7693), .A2(n8318), .B1(n8324), .B2(n8301), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][22] ) );
  OAI22_X1 U11214 ( .A1(n7734), .A2(n10005), .B1(n8302), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][22] ) );
  OAI22_X1 U11215 ( .A1(n7743), .A2(n9775), .B1(n8331), .B2(n9250), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][22] ) );
  OAI22_X1 U11216 ( .A1(n8333), .A2(n9972), .B1(n8303), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][22] ) );
  OAI22_X1 U11217 ( .A1(n7742), .A2(n9796), .B1(n9783), .B2(n8335), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][22] ) );
  OAI22_X1 U11218 ( .A1(n8891), .A2(n9951), .B1(n8941), .B2(n7760), .ZN(
        \DataPath/ALUhw/MULT/mux_out[6][22] ) );
  OAI21_X1 U11219 ( .B1(n8890), .B2(\DP_OP_751_130_6421/n1209 ), .A(n8888), 
        .ZN(n8889) );
  NAND2_X1 U11220 ( .A1(n7771), .A2(\DP_OP_751_130_6421/n1209 ), .ZN(n8888) );
  NAND2_X1 U11221 ( .A1(n7940), .A2(\DataPath/i_PIPLIN_IN2[13] ), .ZN(n8885)
         );
  NAND2_X1 U11222 ( .A1(n8455), .A2(\DataPath/i_PIPLIN_B[13] ), .ZN(n8886) );
  INV_X1 U11223 ( .A(n9784), .ZN(n8890) );
  OAI21_X1 U11224 ( .B1(n8147), .B2(n7940), .A(n8887), .ZN(n9784) );
  NAND2_X1 U11225 ( .A1(n7940), .A2(\DataPath/i_PIPLIN_IN2[12] ), .ZN(n8887)
         );
  OAI22_X1 U11226 ( .A1(n8319), .A2(n8302), .B1(n7693), .B2(n8323), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][21] ) );
  OAI22_X1 U11227 ( .A1(n7734), .A2(n9250), .B1(n10005), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][21] ) );
  OAI22_X1 U11228 ( .A1(n7743), .A2(n8303), .B1(n9775), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][21] ) );
  OAI22_X1 U11229 ( .A1(n8333), .A2(n9783), .B1(n9972), .B2(n8879), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][21] ) );
  OAI22_X1 U11230 ( .A1(n7742), .A2(n8941), .B1(n9796), .B2(n8335), .ZN(
        \DataPath/ALUhw/MULT/mux_out[5][21] ) );
  NAND2_X1 U11231 ( .A1(\DataPath/i_PIPLIN_A[10] ), .A2(n7731), .ZN(n8843) );
  OAI21_X1 U11232 ( .B1(n9191), .B2(\DP_OP_751_130_6421/n1311 ), .A(n8882), 
        .ZN(n8883) );
  AOI21_X1 U11233 ( .B1(n8447), .B2(n9191), .A(n8881), .ZN(n8882) );
  NOR2_X1 U11234 ( .A1(n8447), .A2(n7771), .ZN(n8881) );
  OAI21_X1 U11235 ( .B1(n8146), .B2(n7940), .A(n8880), .ZN(n9191) );
  NAND2_X1 U11236 ( .A1(n7940), .A2(\DataPath/i_PIPLIN_IN2[10] ), .ZN(n8880)
         );
  OAI22_X1 U11237 ( .A1(n8318), .A2(n10005), .B1(n7689), .B2(n9246), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][20] ) );
  OAI22_X1 U11238 ( .A1(n8327), .A2(n9775), .B1(n9250), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][20] ) );
  OAI22_X1 U11239 ( .A1(n8332), .A2(n9972), .B1(n8303), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][20] ) );
  OAI22_X1 U11240 ( .A1(n8333), .A2(n9796), .B1(n9783), .B2(n7745), .ZN(
        \DataPath/ALUhw/MULT/mux_out[4][20] ) );
  OAI21_X1 U11241 ( .B1(n8160), .B2(n7732), .A(n8842), .ZN(n9794) );
  NAND2_X1 U11242 ( .A1(\DataPath/i_PIPLIN_A[11] ), .A2(n7732), .ZN(n8842) );
  OAI21_X1 U11243 ( .B1(n8877), .B2(\DP_OP_751_130_6421/n1515 ), .A(n8876), 
        .ZN(n8878) );
  OAI21_X1 U11244 ( .B1(n8447), .B2(\DP_OP_751_130_6421/n1515 ), .A(n8875), 
        .ZN(n8876) );
  NAND2_X1 U11245 ( .A1(n8447), .A2(n9182), .ZN(n8875) );
  OAI21_X1 U11246 ( .B1(n8144), .B2(n8454), .A(n8874), .ZN(n406) );
  NAND2_X1 U11247 ( .A1(n8454), .A2(\DataPath/i_PIPLIN_IN2[9] ), .ZN(n8874) );
  INV_X1 U11248 ( .A(n9182), .ZN(n8877) );
  OAI22_X1 U11249 ( .A1(n7686), .A2(n9250), .B1(n8323), .B2(n10005), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][19] ) );
  OAI22_X1 U11250 ( .A1(n8327), .A2(n8303), .B1(n9775), .B2(n8330), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][19] ) );
  OAI22_X1 U11251 ( .A1(n7743), .A2(n9783), .B1(n9972), .B2(n7746), .ZN(
        \DataPath/ALUhw/MULT/mux_out[3][19] ) );
  XNOR2_X1 U11252 ( .A(n8445), .B(n9130), .ZN(n8873) );
  NAND2_X1 U11253 ( .A1(\DataPath/i_PIPLIN_A[12] ), .A2(n7731), .ZN(n8841) );
  OAI21_X1 U11254 ( .B1(n8140), .B2(n8454), .A(n8871), .ZN(n9130) );
  NAND2_X1 U11255 ( .A1(n8454), .A2(n497), .ZN(n8871) );
  NAND2_X1 U11256 ( .A1(n8453), .A2(\DataPath/i_PIPLIN_IN2[7] ), .ZN(n8870) );
  OAI22_X1 U11257 ( .A1(n8317), .A2(n9775), .B1(n8323), .B2(n9250), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][18] ) );
  OAI22_X1 U11258 ( .A1(n9972), .A2(n8326), .B1(n8303), .B2(n8328), .ZN(
        \DataPath/ALUhw/MULT/mux_out[2][18] ) );
  NAND2_X1 U11259 ( .A1(n7738), .A2(\DataPath/i_PIPLIN_IN2[5] ), .ZN(n8865) );
  NAND2_X1 U11260 ( .A1(n7630), .A2(n9802), .ZN(n9678) );
  NAND2_X1 U11261 ( .A1(n8867), .A2(n8866), .ZN(n9802) );
  NAND2_X1 U11262 ( .A1(n7738), .A2(\DataPath/i_PIPLIN_IN2[4] ), .ZN(n8866) );
  NAND2_X1 U11263 ( .A1(n7739), .A2(\DataPath/i_PIPLIN_B[4] ), .ZN(n8867) );
  AND2_X1 U11264 ( .A1(n7731), .A2(\DataPath/i_PIPLIN_A[17] ), .ZN(n9991) );
  NAND2_X1 U11265 ( .A1(n8837), .A2(n8836), .ZN(n9062) );
  NAND2_X1 U11266 ( .A1(n7739), .A2(\DataPath/i_PIPLIN_B[0] ), .ZN(n8837) );
  OAI22_X1 U11267 ( .A1(n8318), .A2(n8303), .B1(n8324), .B2(n9775), .ZN(
        \DataPath/ALUhw/MULT/mux_out[1][17] ) );
  OAI21_X1 U11268 ( .B1(n8158), .B2(n7732), .A(n8838), .ZN(n9774) );
  NAND2_X1 U11269 ( .A1(\DataPath/i_PIPLIN_A[15] ), .A2(n7692), .ZN(n8838) );
  NAND2_X1 U11270 ( .A1(\DataPath/i_PIPLIN_A[14] ), .A2(n7731), .ZN(n8839) );
  NAND2_X1 U11271 ( .A1(n8443), .A2(\DataPath/i_PIPLIN_IN1[14] ), .ZN(n8840)
         );
  NAND2_X1 U11272 ( .A1(n8087), .A2(\DataPath/i_PIPLIN_B[3] ), .ZN(n8860) );
  OAI21_X1 U11273 ( .B1(n10269), .B2(n11678), .A(n10268), .ZN(n7025) );
  AOI22_X1 U11274 ( .A1(n10267), .A2(i_RD1[31]), .B1(IRAM_ADDRESS[31]), .B2(
        n10266), .ZN(n10268) );
  INV_X1 U11275 ( .A(n10140), .ZN(n8485) );
  NOR2_X1 U11276 ( .A1(n10260), .A2(n10263), .ZN(n10262) );
  NAND2_X1 U11277 ( .A1(n10162), .A2(IRAM_ADDRESS[29]), .ZN(n10260) );
  NOR2_X1 U11278 ( .A1(n10175), .A2(n8178), .ZN(n10162) );
  NAND2_X1 U11279 ( .A1(n10175), .A2(IRAM_ADDRESS[26]), .ZN(n10169) );
  OAI22_X1 U11280 ( .A1(n10156), .A2(n10175), .B1(IRAM_ADDRESS[27]), .B2(
        n10168), .ZN(n10159) );
  INV_X1 U11281 ( .A(n10177), .ZN(n10168) );
  OR2_X1 U11282 ( .A1(n10153), .A2(n173), .ZN(n10154) );
  OR2_X1 U11283 ( .A1(\intadd_2/B[3] ), .A2(IRAM_ADDRESS[24]), .ZN(n8120) );
  OAI21_X1 U11284 ( .B1(n174), .B2(n10153), .A(n10155), .ZN(\intadd_2/B[3] )
         );
  OAI21_X1 U11285 ( .B1(n175), .B2(n10153), .A(n10155), .ZN(\intadd_2/B[2] )
         );
  OR2_X1 U11286 ( .A1(\intadd_2/B[1] ), .A2(IRAM_ADDRESS[22]), .ZN(n8092) );
  OAI21_X1 U11287 ( .B1(n176), .B2(n10153), .A(n10155), .ZN(\intadd_2/B[1] )
         );
  OR2_X1 U11288 ( .A1(\intadd_2/B[0] ), .A2(IRAM_ADDRESS[21]), .ZN(n8123) );
  OAI21_X1 U11289 ( .B1(n177), .B2(n10153), .A(n10155), .ZN(\intadd_2/B[0] )
         );
  OAI21_X1 U11290 ( .B1(n178), .B2(n10153), .A(n10155), .ZN(n10186) );
  NAND2_X1 U11291 ( .A1(n10150), .A2(n8180), .ZN(n10151) );
  AOI21_X1 U11292 ( .B1(n8833), .B2(n8184), .A(n8832), .ZN(n10150) );
  INV_X1 U11293 ( .A(n10155), .ZN(n8832) );
  INV_X1 U11294 ( .A(n10153), .ZN(n8833) );
  AND2_X1 U11295 ( .A1(n8830), .A2(n8829), .ZN(n10146) );
  OAI22_X1 U11296 ( .A1(n8827), .A2(n11673), .B1(IRAM_ADDRESS[17]), .B2(n11672), .ZN(n8830) );
  INV_X1 U11297 ( .A(n8823), .ZN(n8827) );
  INV_X1 U11298 ( .A(n8831), .ZN(n10147) );
  NAND2_X1 U11299 ( .A1(n8831), .A2(n8829), .ZN(n10148) );
  NAND2_X1 U11300 ( .A1(n8826), .A2(IRAM_ADDRESS[18]), .ZN(n8829) );
  OR2_X1 U11301 ( .A1(n8826), .A2(IRAM_ADDRESS[18]), .ZN(n8831) );
  XNOR2_X1 U11302 ( .A(n11672), .B(n8181), .ZN(n8824) );
  OR2_X1 U11303 ( .A1(n8253), .A2(n10187), .ZN(n8251) );
  OAI21_X1 U11304 ( .B1(IRAM_ADDRESS[16]), .B2(n8822), .A(n8823), .ZN(n10187)
         );
  NAND2_X1 U11305 ( .A1(n8822), .A2(IRAM_ADDRESS[16]), .ZN(n8823) );
  INV_X1 U11306 ( .A(n7636), .ZN(n8820) );
  NOR2_X1 U11307 ( .A1(n10191), .A2(n8254), .ZN(n8252) );
  AND2_X1 U11308 ( .A1(n8817), .A2(IRAM_ADDRESS[10]), .ZN(n10188) );
  INV_X1 U11309 ( .A(n10189), .ZN(n8818) );
  NOR2_X1 U11310 ( .A1(n8817), .A2(IRAM_ADDRESS[10]), .ZN(n10189) );
  OR2_X1 U11311 ( .A1(\intadd_0/B[4] ), .A2(n8125), .ZN(n8093) );
  OR2_X1 U11312 ( .A1(\intadd_0/B[1] ), .A2(n8128), .ZN(n8091) );
  OR2_X1 U11313 ( .A1(\intadd_0/B[0] ), .A2(\intadd_0/A[0] ), .ZN(n8122) );
  NOR2_X1 U11314 ( .A1(n8804), .A2(IRAM_ADDRESS[9]), .ZN(n8815) );
  INV_X1 U11315 ( .A(n8805), .ZN(n8804) );
  NOR2_X1 U11316 ( .A1(n10194), .A2(n8169), .ZN(n10196) );
  NOR2_X1 U11317 ( .A1(n8805), .A2(n208), .ZN(n8814) );
  NAND2_X1 U11318 ( .A1(n10194), .A2(n8169), .ZN(n10195) );
  AOI21_X1 U11319 ( .B1(\intadd_1/CO ), .B2(n10203), .A(n10202), .ZN(n10200)
         );
  NOR2_X1 U11320 ( .A1(n8806), .A2(IRAM_ADDRESS[6]), .ZN(n10202) );
  NAND2_X1 U11321 ( .A1(n8806), .A2(IRAM_ADDRESS[6]), .ZN(n10203) );
  OAI21_X1 U11322 ( .B1(\intadd_1/n19 ), .B2(n8118), .A(\intadd_1/n8 ), .ZN(
        \intadd_1/CO ) );
  OAI21_X1 U11323 ( .B1(\intadd_1/n29 ), .B2(\intadd_1/n31 ), .A(
        \intadd_1/n30 ), .ZN(\intadd_1/n28 ) );
  NAND2_X1 U11324 ( .A1(n10211), .A2(IRAM_ADDRESS[0]), .ZN(\intadd_1/CI ) );
  INV_X1 U11325 ( .A(n10198), .ZN(n8808) );
  NAND2_X1 U11326 ( .A1(n10295), .A2(n8482), .ZN(n8483) );
  NAND2_X1 U11327 ( .A1(n8491), .A2(n8479), .ZN(n8481) );
  NAND2_X1 U11328 ( .A1(n7990), .A2(n8115), .ZN(n8479) );
  AOI21_X1 U11329 ( .B1(n8798), .B2(n8797), .A(n8796), .ZN(n8799) );
  AOI21_X1 U11330 ( .B1(n8795), .B2(n8794), .A(n8793), .ZN(n8796) );
  AOI21_X1 U11331 ( .B1(n10105), .B2(n10138), .A(n8792), .ZN(n8797) );
  NAND2_X1 U11332 ( .A1(n10223), .A2(n8130), .ZN(n8792) );
  NOR2_X1 U11333 ( .A1(n8794), .A2(n8279), .ZN(n10223) );
  INV_X1 U11334 ( .A(n7954), .ZN(n8794) );
  NAND2_X1 U11335 ( .A1(n10093), .A2(n10139), .ZN(n8798) );
  INV_X1 U11336 ( .A(n10105), .ZN(n10093) );
  NOR2_X1 U11337 ( .A1(n8789), .A2(n10065), .ZN(n10231) );
  INV_X1 U11338 ( .A(n8788), .ZN(n8789) );
  NOR2_X1 U11339 ( .A1(n10105), .A2(n10232), .ZN(n8790) );
  INV_X1 U11340 ( .A(n8784), .ZN(n8229) );
  AND2_X1 U11341 ( .A1(n7751), .A2(n8785), .ZN(n8225) );
  OAI21_X1 U11342 ( .B1(n8717), .B2(n8716), .A(n8784), .ZN(n8785) );
  NAND2_X1 U11343 ( .A1(n8717), .A2(n8715), .ZN(n8784) );
  AOI21_X1 U11344 ( .B1(n10246), .B2(n8714), .A(\CU_I/CW_ID[UNSIGNED_ID] ), 
        .ZN(n8715) );
  NOR2_X1 U11345 ( .A1(n11621), .A2(n7975), .ZN(n8714) );
  OAI21_X1 U11346 ( .B1(IR[1]), .B2(IR[2]), .A(n11623), .ZN(n11621) );
  INV_X1 U11347 ( .A(n10098), .ZN(n10246) );
  NAND2_X1 U11348 ( .A1(n8713), .A2(i_RD1[30]), .ZN(n8716) );
  INV_X1 U11349 ( .A(n8712), .ZN(n8713) );
  OAI21_X1 U11350 ( .B1(n8231), .B2(n8783), .A(n8782), .ZN(n8230) );
  AOI21_X1 U11351 ( .B1(n8233), .B2(n8697), .A(n8778), .ZN(n8231) );
  NAND2_X1 U11352 ( .A1(n8773), .A2(i_RD1[27]), .ZN(n8774) );
  INV_X1 U11353 ( .A(n8772), .ZN(n8773) );
  INV_X1 U11354 ( .A(n8771), .ZN(n8777) );
  INV_X1 U11355 ( .A(n8233), .ZN(n8232) );
  AND2_X1 U11356 ( .A1(n8119), .A2(n8234), .ZN(n8233) );
  NAND2_X1 U11357 ( .A1(n8769), .A2(n8770), .ZN(n8234) );
  NAND2_X1 U11358 ( .A1(n8765), .A2(n8764), .ZN(n8766) );
  OAI211_X1 U11359 ( .C1(n8763), .C2(n8762), .A(n8761), .B(n8760), .ZN(n8768)
         );
  NAND2_X1 U11360 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  NAND2_X1 U11361 ( .A1(n8757), .A2(n8756), .ZN(n8759) );
  NAND4_X1 U11362 ( .A1(n8755), .A2(n8754), .A3(n8753), .A4(n8758), .ZN(n8761)
         );
  NAND2_X1 U11363 ( .A1(n8752), .A2(n8751), .ZN(n8755) );
  OR2_X1 U11364 ( .A1(n8750), .A2(n8749), .ZN(n8762) );
  AOI21_X1 U11365 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n8763) );
  OR2_X1 U11366 ( .A1(n8745), .A2(n8744), .ZN(n8746) );
  INV_X1 U11367 ( .A(n8726), .ZN(n8727) );
  NAND2_X1 U11368 ( .A1(n8711), .A2(n10138), .ZN(n8786) );
  XNOR2_X1 U11369 ( .A(n8726), .B(i_RD1[5]), .ZN(n8728) );
  NAND2_X1 U11370 ( .A1(n8707), .A2(n8706), .ZN(n8726) );
  NAND2_X1 U11371 ( .A1(i_SEL_CMPB), .A2(i_RD2[5]), .ZN(n8706) );
  NAND2_X1 U11372 ( .A1(n10090), .A2(n8456), .ZN(n8707) );
  AOI21_X1 U11373 ( .B1(n8295), .B2(IRAM_ADDRESS[5]), .A(n8703), .ZN(n8704) );
  XNOR2_X1 U11374 ( .A(n8712), .B(i_RD1[30]), .ZN(n8780) );
  NAND2_X1 U11375 ( .A1(n8702), .A2(n8701), .ZN(n8712) );
  NAND2_X1 U11376 ( .A1(i_SEL_CMPB), .A2(i_RD2[30]), .ZN(n8701) );
  NAND2_X1 U11377 ( .A1(n10073), .A2(n8456), .ZN(n8702) );
  NAND2_X1 U11378 ( .A1(n8700), .A2(n8699), .ZN(n10073) );
  AOI21_X1 U11379 ( .B1(n8296), .B2(IRAM_ADDRESS[30]), .A(n8698), .ZN(n8699)
         );
  NAND2_X1 U11380 ( .A1(n8695), .A2(n8694), .ZN(n8745) );
  NAND2_X1 U11381 ( .A1(n8693), .A2(i_RD1[16]), .ZN(n8694) );
  INV_X1 U11382 ( .A(n8775), .ZN(n8696) );
  AND2_X1 U11383 ( .A1(n8692), .A2(n8691), .ZN(n8775) );
  NAND2_X1 U11384 ( .A1(n8690), .A2(i_RD1[28]), .ZN(n8691) );
  NAND2_X1 U11385 ( .A1(n8688), .A2(n8687), .ZN(n8689) );
  INV_X1 U11386 ( .A(i_RD1[31]), .ZN(n8687) );
  AOI22_X1 U11387 ( .A1(n8297), .A2(IRAM_ADDRESS[31]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[31] ), .ZN(n8684) );
  AND2_X1 U11388 ( .A1(n8683), .A2(n8682), .ZN(n8769) );
  NAND2_X1 U11389 ( .A1(n8681), .A2(n8680), .ZN(n8682) );
  AOI21_X1 U11390 ( .B1(n7856), .B2(i_RD2[24]), .A(n8679), .ZN(n8680) );
  INV_X1 U11391 ( .A(i_RD1[24]), .ZN(n8679) );
  NAND2_X1 U11392 ( .A1(n10079), .A2(n8456), .ZN(n8681) );
  NAND2_X1 U11393 ( .A1(n8676), .A2(i_RD1[26]), .ZN(n8776) );
  INV_X1 U11394 ( .A(n8675), .ZN(n8676) );
  OAI211_X1 U11395 ( .C1(n7856), .C2(n10079), .A(n8683), .B(n8674), .ZN(n8677)
         );
  AOI21_X1 U11396 ( .B1(i_SEL_CMPB), .B2(n8673), .A(i_RD1[24]), .ZN(n8674) );
  INV_X1 U11397 ( .A(i_RD2[24]), .ZN(n8673) );
  NAND2_X1 U11398 ( .A1(n8672), .A2(i_RD1[25]), .ZN(n8683) );
  NAND2_X1 U11399 ( .A1(n8700), .A2(n8671), .ZN(n10079) );
  AOI22_X1 U11400 ( .A1(n8297), .A2(IRAM_ADDRESS[24]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[24] ), .ZN(n8671) );
  XNOR2_X1 U11401 ( .A(n8772), .B(i_RD1[27]), .ZN(n8771) );
  NAND2_X1 U11402 ( .A1(n8670), .A2(n8669), .ZN(n8772) );
  NAND2_X1 U11403 ( .A1(n7856), .A2(i_RD2[27]), .ZN(n8669) );
  NAND2_X1 U11404 ( .A1(n10076), .A2(n8456), .ZN(n8670) );
  NAND2_X1 U11405 ( .A1(n8700), .A2(n8668), .ZN(n10076) );
  AOI21_X1 U11406 ( .B1(n8295), .B2(IRAM_ADDRESS[27]), .A(n8667), .ZN(n8668)
         );
  AOI22_X1 U11407 ( .A1(n8675), .A2(n8666), .B1(n8665), .B2(n8664), .ZN(n8678)
         );
  INV_X1 U11408 ( .A(i_RD1[25]), .ZN(n8664) );
  INV_X1 U11409 ( .A(n8672), .ZN(n8665) );
  OAI21_X1 U11410 ( .B1(n10078), .B2(n7856), .A(n8663), .ZN(n8672) );
  NAND2_X1 U11411 ( .A1(i_SEL_CMPB), .A2(n8662), .ZN(n8663) );
  INV_X1 U11412 ( .A(i_RD2[25]), .ZN(n8662) );
  NAND2_X1 U11413 ( .A1(n8700), .A2(n8661), .ZN(n10078) );
  AOI21_X1 U11414 ( .B1(n8297), .B2(IRAM_ADDRESS[25]), .A(n8660), .ZN(n8661)
         );
  INV_X1 U11415 ( .A(i_RD1[26]), .ZN(n8666) );
  NAND2_X1 U11416 ( .A1(n8700), .A2(n8659), .ZN(n10077) );
  AOI22_X1 U11417 ( .A1(n8297), .A2(IRAM_ADDRESS[26]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[26] ), .ZN(n8659) );
  NOR2_X1 U11418 ( .A1(n8658), .A2(n8750), .ZN(n8709) );
  NAND4_X1 U11419 ( .A1(n8657), .A2(n8656), .A3(n8752), .A4(n8655), .ZN(n8750)
         );
  INV_X1 U11420 ( .A(i_RD1[16]), .ZN(n8653) );
  INV_X1 U11421 ( .A(n8693), .ZN(n8654) );
  OAI21_X1 U11422 ( .B1(n10086), .B2(i_SEL_CMPB), .A(n8652), .ZN(n8693) );
  NAND2_X1 U11423 ( .A1(n7856), .A2(n8651), .ZN(n8652) );
  INV_X1 U11424 ( .A(i_RD2[16]), .ZN(n8651) );
  NAND2_X1 U11425 ( .A1(n8700), .A2(n8650), .ZN(n10086) );
  AOI22_X1 U11426 ( .A1(n8295), .A2(IRAM_ADDRESS[16]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[16] ), .ZN(n8650) );
  NAND2_X1 U11427 ( .A1(n8649), .A2(i_RD1[17]), .ZN(n8695) );
  NAND2_X1 U11428 ( .A1(n8648), .A2(i_RD1[18]), .ZN(n8752) );
  INV_X1 U11429 ( .A(n8647), .ZN(n8648) );
  AOI22_X1 U11430 ( .A1(n8647), .A2(n8646), .B1(n8645), .B2(n8644), .ZN(n8656)
         );
  INV_X1 U11431 ( .A(i_RD1[17]), .ZN(n8644) );
  INV_X1 U11432 ( .A(n8649), .ZN(n8645) );
  OAI21_X1 U11433 ( .B1(n10085), .B2(n7856), .A(n8643), .ZN(n8649) );
  NAND2_X1 U11434 ( .A1(n7856), .A2(n8642), .ZN(n8643) );
  INV_X1 U11435 ( .A(i_RD2[17]), .ZN(n8642) );
  NAND2_X1 U11436 ( .A1(n8700), .A2(n8641), .ZN(n10085) );
  AOI21_X1 U11437 ( .B1(n8296), .B2(IRAM_ADDRESS[17]), .A(n8640), .ZN(n8641)
         );
  INV_X1 U11438 ( .A(i_RD1[18]), .ZN(n8646) );
  NAND2_X1 U11439 ( .A1(n8700), .A2(n8639), .ZN(n10084) );
  AOI22_X1 U11440 ( .A1(n8297), .A2(IRAM_ADDRESS[18]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[18] ), .ZN(n8639) );
  BUF_X1 U11441 ( .A(n8295), .Z(n8297) );
  AND2_X1 U11442 ( .A1(n8754), .A2(n8751), .ZN(n8657) );
  NAND2_X1 U11443 ( .A1(n8638), .A2(i_RD1[19]), .ZN(n8751) );
  OR2_X1 U11444 ( .A1(n8638), .A2(i_RD1[19]), .ZN(n8754) );
  OAI21_X1 U11445 ( .B1(n10083), .B2(i_SEL_CMPB), .A(n8637), .ZN(n8638) );
  NAND2_X1 U11446 ( .A1(i_SEL_CMPB), .A2(n8636), .ZN(n8637) );
  INV_X1 U11447 ( .A(i_RD2[19]), .ZN(n8636) );
  NAND2_X1 U11448 ( .A1(n8700), .A2(n8635), .ZN(n10083) );
  AOI21_X1 U11449 ( .B1(n8296), .B2(IRAM_ADDRESS[19]), .A(n8634), .ZN(n8635)
         );
  NAND4_X1 U11450 ( .A1(n8633), .A2(n8163), .A3(n8632), .A4(n8765), .ZN(n8658)
         );
  NAND2_X1 U11451 ( .A1(n8631), .A2(i_RD1[22]), .ZN(n8765) );
  NOR2_X1 U11452 ( .A1(n8630), .A2(n8629), .ZN(n8632) );
  INV_X1 U11453 ( .A(n8764), .ZN(n8629) );
  NAND2_X1 U11454 ( .A1(n8628), .A2(n8627), .ZN(n8764) );
  AOI21_X1 U11455 ( .B1(n7856), .B2(i_RD2[23]), .A(n8626), .ZN(n8627) );
  NAND2_X1 U11456 ( .A1(n10080), .A2(n8456), .ZN(n8628) );
  INV_X1 U11457 ( .A(n8723), .ZN(n8630) );
  NAND2_X1 U11458 ( .A1(n8625), .A2(i_RD1[4]), .ZN(n8723) );
  AND4_X1 U11459 ( .A1(n8767), .A2(n8757), .A3(n8756), .A4(n8624), .ZN(n8163)
         );
  INV_X1 U11460 ( .A(n8731), .ZN(n8624) );
  NOR2_X1 U11461 ( .A1(n8623), .A2(i_RD1[6]), .ZN(n8731) );
  NAND2_X1 U11462 ( .A1(n8622), .A2(i_RD1[21]), .ZN(n8756) );
  NAND2_X1 U11463 ( .A1(n8621), .A2(i_RD1[20]), .ZN(n8757) );
  OR2_X1 U11464 ( .A1(n8631), .A2(i_RD1[22]), .ZN(n8767) );
  OAI21_X1 U11465 ( .B1(n10081), .B2(n7856), .A(n8620), .ZN(n8631) );
  NAND2_X1 U11466 ( .A1(n7856), .A2(n8619), .ZN(n8620) );
  INV_X1 U11467 ( .A(i_RD2[22]), .ZN(n8619) );
  NAND2_X1 U11468 ( .A1(n8700), .A2(n8618), .ZN(n10081) );
  AOI22_X1 U11469 ( .A1(n8295), .A2(IRAM_ADDRESS[22]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[22] ), .ZN(n8618) );
  INV_X1 U11470 ( .A(n8749), .ZN(n8633) );
  NAND2_X1 U11471 ( .A1(n8758), .A2(n8753), .ZN(n8749) );
  OR2_X1 U11472 ( .A1(n8621), .A2(i_RD1[20]), .ZN(n8753) );
  OAI21_X1 U11473 ( .B1(n10134), .B2(i_SEL_CMPB), .A(n8617), .ZN(n8621) );
  NAND2_X1 U11474 ( .A1(i_SEL_CMPB), .A2(n8616), .ZN(n8617) );
  INV_X1 U11475 ( .A(i_RD2[20]), .ZN(n8616) );
  NAND2_X1 U11476 ( .A1(n8700), .A2(n8615), .ZN(n10134) );
  AOI22_X1 U11477 ( .A1(n8296), .A2(IRAM_ADDRESS[20]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[20] ), .ZN(n8615) );
  OR2_X1 U11478 ( .A1(n8622), .A2(i_RD1[21]), .ZN(n8758) );
  OAI21_X1 U11479 ( .B1(n10082), .B2(n7856), .A(n8614), .ZN(n8622) );
  NAND2_X1 U11480 ( .A1(n7856), .A2(n8613), .ZN(n8614) );
  INV_X1 U11481 ( .A(i_RD2[21]), .ZN(n8613) );
  NAND2_X1 U11482 ( .A1(n8700), .A2(n8612), .ZN(n10082) );
  AOI21_X1 U11483 ( .B1(n8296), .B2(IRAM_ADDRESS[21]), .A(n8611), .ZN(n8612)
         );
  NOR2_X1 U11484 ( .A1(n8610), .A2(n8609), .ZN(n8710) );
  OR2_X1 U11485 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  INV_X1 U11486 ( .A(n7646), .ZN(n8606) );
  OAI21_X1 U11487 ( .B1(n8605), .B2(i_RD1[1]), .A(n8604), .ZN(n8718) );
  OAI21_X1 U11488 ( .B1(n10113), .B2(i_SEL_CMPB), .A(n8603), .ZN(n8604) );
  AOI21_X1 U11489 ( .B1(i_SEL_CMPB), .B2(n8602), .A(i_RD1[0]), .ZN(n8603) );
  INV_X1 U11490 ( .A(i_RD2[0]), .ZN(n8602) );
  AOI22_X1 U11491 ( .A1(n8605), .A2(i_RD1[1]), .B1(n8601), .B2(i_RD1[2]), .ZN(
        n8719) );
  AND2_X1 U11492 ( .A1(i_SEL_CMPB), .A2(i_RD2[1]), .ZN(n8600) );
  NAND2_X1 U11493 ( .A1(n8295), .A2(IRAM_ADDRESS[1]), .ZN(n8598) );
  AOI22_X1 U11494 ( .A1(i_RD1[6]), .A2(n8623), .B1(n8597), .B2(i_RD1[7]), .ZN(
        n8730) );
  OAI21_X1 U11495 ( .B1(n10120), .B2(n7856), .A(n8596), .ZN(n8623) );
  NAND2_X1 U11496 ( .A1(i_SEL_CMPB), .A2(n11629), .ZN(n8596) );
  INV_X1 U11497 ( .A(i_RD2[6]), .ZN(n11629) );
  NAND2_X1 U11498 ( .A1(n8297), .A2(IRAM_ADDRESS[6]), .ZN(n8594) );
  NAND2_X1 U11499 ( .A1(n10245), .A2(\DECODEhw/i_tickcounter[6] ), .ZN(n8595)
         );
  AOI22_X1 U11500 ( .A1(n7638), .A2(i_RD1[9]), .B1(n8592), .B2(i_RD1[10]), 
        .ZN(n8736) );
  INV_X1 U11501 ( .A(n8744), .ZN(n8591) );
  AND2_X1 U11502 ( .A1(n8590), .A2(i_RD1[15]), .ZN(n8744) );
  NAND2_X1 U11503 ( .A1(n8589), .A2(i_RD1[12]), .ZN(n8739) );
  AOI22_X1 U11504 ( .A1(n8588), .A2(n8587), .B1(n8586), .B2(n8585), .ZN(n8721)
         );
  INV_X1 U11505 ( .A(n7718), .ZN(n8586) );
  AND2_X1 U11506 ( .A1(n7856), .A2(i_RD2[2]), .ZN(n8584) );
  NAND2_X1 U11507 ( .A1(n10245), .A2(\DECODEhw/i_tickcounter[2] ), .ZN(n8582)
         );
  NAND2_X1 U11508 ( .A1(n8295), .A2(IRAM_ADDRESS[2]), .ZN(n8583) );
  NAND2_X1 U11509 ( .A1(n8580), .A2(n8579), .ZN(n8734) );
  INV_X1 U11510 ( .A(n8597), .ZN(n8580) );
  AOI21_X1 U11511 ( .B1(n10089), .B2(n8456), .A(n8578), .ZN(n8597) );
  AND2_X1 U11512 ( .A1(i_SEL_CMPB), .A2(i_RD2[7]), .ZN(n8578) );
  NAND2_X1 U11513 ( .A1(n8296), .A2(IRAM_ADDRESS[7]), .ZN(n8576) );
  INV_X1 U11514 ( .A(n8720), .ZN(n8581) );
  AND2_X1 U11515 ( .A1(n8575), .A2(i_RD1[3]), .ZN(n8720) );
  INV_X1 U11516 ( .A(n8588), .ZN(n8575) );
  AOI21_X1 U11517 ( .B1(n8295), .B2(IRAM_ADDRESS[3]), .A(n8573), .ZN(n8574) );
  NAND2_X1 U11518 ( .A1(n8571), .A2(i_RD1[11]), .ZN(n8738) );
  INV_X1 U11519 ( .A(n8570), .ZN(n8571) );
  NAND4_X1 U11520 ( .A1(n8781), .A2(n8569), .A3(n8568), .A4(n8567), .ZN(n8610)
         );
  NOR2_X1 U11521 ( .A1(n7639), .A2(n7752), .ZN(n8567) );
  AOI22_X1 U11522 ( .A1(n8570), .A2(n8566), .B1(n8565), .B2(n8564), .ZN(n8741)
         );
  INV_X1 U11523 ( .A(i_RD1[10]), .ZN(n8564) );
  INV_X1 U11524 ( .A(n8592), .ZN(n8565) );
  AOI21_X1 U11525 ( .B1(n10124), .B2(n8456), .A(n8563), .ZN(n8592) );
  AND2_X1 U11526 ( .A1(n7856), .A2(i_RD2[10]), .ZN(n8563) );
  NAND2_X1 U11527 ( .A1(n10245), .A2(\DECODEhw/i_tickcounter[10] ), .ZN(n8561)
         );
  NAND2_X1 U11528 ( .A1(n8298), .A2(IRAM_ADDRESS[10]), .ZN(n8562) );
  AOI21_X1 U11529 ( .B1(n8298), .B2(IRAM_ADDRESS[11]), .A(n8559), .ZN(n8560)
         );
  OAI21_X1 U11530 ( .B1(n8572), .B2(i_RD1[8]), .A(n8558), .ZN(n8737) );
  NAND2_X1 U11531 ( .A1(n8557), .A2(n8556), .ZN(n8558) );
  INV_X1 U11532 ( .A(i_RD1[9]), .ZN(n8556) );
  INV_X1 U11533 ( .A(n8593), .ZN(n8557) );
  AOI21_X1 U11534 ( .B1(n10088), .B2(n8456), .A(n8555), .ZN(n8593) );
  AND2_X1 U11535 ( .A1(i_SEL_CMPB), .A2(i_RD2[9]), .ZN(n8555) );
  NAND2_X1 U11536 ( .A1(n8298), .A2(IRAM_ADDRESS[9]), .ZN(n8553) );
  OAI21_X1 U11537 ( .B1(n10122), .B2(i_SEL_CMPB), .A(n8552), .ZN(n8572) );
  NAND2_X1 U11538 ( .A1(n7856), .A2(n8551), .ZN(n8552) );
  INV_X1 U11539 ( .A(i_RD2[8]), .ZN(n8551) );
  NAND2_X1 U11540 ( .A1(n8297), .A2(IRAM_ADDRESS[8]), .ZN(n8549) );
  NAND2_X1 U11541 ( .A1(n10245), .A2(\DECODEhw/i_tickcounter[8] ), .ZN(n8550)
         );
  NOR2_X1 U11542 ( .A1(n8548), .A2(n8547), .ZN(n8568) );
  INV_X1 U11543 ( .A(n8742), .ZN(n8547) );
  AOI22_X1 U11544 ( .A1(i_RD1[13]), .A2(n8546), .B1(n8545), .B2(i_RD1[14]), 
        .ZN(n8742) );
  INV_X1 U11545 ( .A(n8747), .ZN(n8548) );
  AOI22_X1 U11546 ( .A1(n8544), .A2(n8543), .B1(n8542), .B2(n8541), .ZN(n8747)
         );
  INV_X1 U11547 ( .A(n8545), .ZN(n8542) );
  AOI21_X1 U11548 ( .B1(n10130), .B2(n8456), .A(n8540), .ZN(n8545) );
  AND2_X1 U11549 ( .A1(n7856), .A2(i_RD2[14]), .ZN(n8540) );
  NAND2_X1 U11550 ( .A1(n10245), .A2(\DECODEhw/i_tickcounter[14] ), .ZN(n8538)
         );
  NAND2_X1 U11551 ( .A1(n8296), .A2(IRAM_ADDRESS[14]), .ZN(n8539) );
  INV_X1 U11552 ( .A(n8590), .ZN(n8544) );
  OAI21_X1 U11553 ( .B1(n10132), .B2(n7856), .A(n8537), .ZN(n8590) );
  NAND2_X1 U11554 ( .A1(i_SEL_CMPB), .A2(n8536), .ZN(n8537) );
  INV_X1 U11555 ( .A(i_RD2[15]), .ZN(n8536) );
  NAND2_X1 U11556 ( .A1(n8295), .A2(IRAM_ADDRESS[15]), .ZN(n8535) );
  NOR2_X1 U11557 ( .A1(n8743), .A2(n8533), .ZN(n8569) );
  NAND2_X1 U11558 ( .A1(n8530), .A2(n8529), .ZN(n8531) );
  AOI21_X1 U11559 ( .B1(n7856), .B2(i_RD2[0]), .A(n8528), .ZN(n8529) );
  NAND2_X1 U11560 ( .A1(n10113), .A2(n8456), .ZN(n8530) );
  AOI21_X1 U11561 ( .B1(n8295), .B2(IRAM_ADDRESS[0]), .A(n8526), .ZN(n8527) );
  BUF_X1 U11562 ( .A(n8295), .Z(n8298) );
  NOR2_X1 U11563 ( .A1(n8625), .A2(i_RD1[4]), .ZN(n8724) );
  OAI22_X1 U11564 ( .A1(n10117), .A2(n8525), .B1(i_RD2[4]), .B2(n8456), .ZN(
        n8625) );
  OR2_X1 U11565 ( .A1(n10291), .A2(i_SEL_CMPB), .ZN(n8525) );
  INV_X1 U11566 ( .A(n8521), .ZN(n8522) );
  NAND2_X1 U11567 ( .A1(n8298), .A2(IRAM_ADDRESS[4]), .ZN(n8524) );
  INV_X1 U11568 ( .A(n8770), .ZN(n8532) );
  AOI21_X1 U11569 ( .B1(n8520), .B2(n8456), .A(n8519), .ZN(n8770) );
  OAI21_X1 U11570 ( .B1(i_RD2[23]), .B2(n8456), .A(n8626), .ZN(n8519) );
  INV_X1 U11571 ( .A(i_RD1[23]), .ZN(n8626) );
  INV_X1 U11572 ( .A(n10080), .ZN(n8520) );
  NAND2_X1 U11573 ( .A1(n8700), .A2(n8518), .ZN(n10080) );
  AOI21_X1 U11574 ( .B1(n8295), .B2(IRAM_ADDRESS[23]), .A(n8517), .ZN(n8518)
         );
  OAI21_X1 U11575 ( .B1(n8589), .B2(i_RD1[12]), .A(n8516), .ZN(n8743) );
  NAND2_X1 U11576 ( .A1(n8515), .A2(n8514), .ZN(n8516) );
  INV_X1 U11577 ( .A(n8546), .ZN(n8515) );
  AOI21_X1 U11578 ( .B1(n10128), .B2(n8456), .A(n8513), .ZN(n8546) );
  AND2_X1 U11579 ( .A1(i_SEL_CMPB), .A2(i_RD2[13]), .ZN(n8513) );
  NAND2_X1 U11580 ( .A1(n8295), .A2(IRAM_ADDRESS[13]), .ZN(n8511) );
  OAI21_X1 U11581 ( .B1(n10126), .B2(i_SEL_CMPB), .A(n8510), .ZN(n8589) );
  NAND2_X1 U11582 ( .A1(i_SEL_CMPB), .A2(n8509), .ZN(n8510) );
  INV_X1 U11583 ( .A(i_RD2[12]), .ZN(n8509) );
  NAND2_X1 U11584 ( .A1(n8298), .A2(IRAM_ADDRESS[12]), .ZN(n8507) );
  NAND2_X1 U11585 ( .A1(n10245), .A2(\DECODEhw/i_tickcounter[12] ), .ZN(n8508)
         );
  NAND2_X1 U11586 ( .A1(n8506), .A2(n8692), .ZN(n8781) );
  NAND2_X1 U11587 ( .A1(n8505), .A2(i_RD1[29]), .ZN(n8692) );
  OAI22_X1 U11588 ( .A1(i_RD1[29]), .A2(n8505), .B1(n8690), .B2(i_RD1[28]), 
        .ZN(n8506) );
  OAI21_X1 U11589 ( .B1(n10075), .B2(n7856), .A(n8504), .ZN(n8690) );
  NAND2_X1 U11590 ( .A1(n7856), .A2(n8503), .ZN(n8504) );
  INV_X1 U11591 ( .A(i_RD2[28]), .ZN(n8503) );
  NAND2_X1 U11592 ( .A1(n8700), .A2(n8502), .ZN(n10075) );
  AOI21_X1 U11593 ( .B1(n8295), .B2(IRAM_ADDRESS[28]), .A(n8501), .ZN(n8502)
         );
  OAI21_X1 U11594 ( .B1(n10074), .B2(i_SEL_CMPB), .A(n8500), .ZN(n8505) );
  NAND2_X1 U11595 ( .A1(i_SEL_CMPB), .A2(n8499), .ZN(n8500) );
  INV_X1 U11596 ( .A(i_RD2[29]), .ZN(n8499) );
  NAND2_X1 U11597 ( .A1(n8700), .A2(n8498), .ZN(n10074) );
  AOI22_X1 U11598 ( .A1(n8297), .A2(IRAM_ADDRESS[29]), .B1(n10245), .B2(
        \DECODEhw/i_tickcounter[29] ), .ZN(n8498) );
  NAND2_X1 U11599 ( .A1(n10221), .A2(n7954), .ZN(n8496) );
  INV_X1 U11600 ( .A(n10232), .ZN(n10221) );
  NOR2_X1 U11601 ( .A1(n183), .A2(\CU_I/CW_ID[UNSIGNED_ID] ), .ZN(n8494) );
  NAND2_X1 U11602 ( .A1(n10098), .A2(n10271), .ZN(n8521) );
  NOR2_X1 U11603 ( .A1(n10232), .A2(n10065), .ZN(n8493) );
  NAND2_X1 U11604 ( .A1(n10235), .A2(n10226), .ZN(n10098) );
  NOR2_X1 U11605 ( .A1(n10139), .A2(n8492), .ZN(n10235) );
  NAND2_X1 U11606 ( .A1(n10219), .A2(n8130), .ZN(n10220) );
  NOR2_X1 U11607 ( .A1(n10067), .A2(n8279), .ZN(n10219) );
  INV_X1 U11608 ( .A(n8492), .ZN(n8489) );
  NAND2_X1 U11609 ( .A1(n10224), .A2(n8115), .ZN(n8491) );
  NAND2_X1 U11610 ( .A1(n8244), .A2(n10232), .ZN(n8787) );
  NOR2_X1 U11611 ( .A1(n8129), .A2(n471), .ZN(n10293) );
  XNOR2_X1 U11612 ( .A(\DP_OP_751_130_6421/n1311 ), .B(n9784), .ZN(n8892) );
  XNOR2_X1 U11613 ( .A(n9182), .B(\DP_OP_751_130_6421/n1515 ), .ZN(n8879) );
  XNOR2_X1 U11614 ( .A(\DP_OP_751_130_6421/n597 ), .B(n9517), .ZN(n8931) );
  XNOR2_X1 U11615 ( .A(\DP_OP_751_130_6421/n1209 ), .B(n9780), .ZN(n8896) );
  XNOR2_X1 U11616 ( .A(\DP_OP_751_130_6421/n1413 ), .B(n9191), .ZN(n8884) );
  NAND2_X1 U11617 ( .A1(n8049), .A2(n9678), .ZN(n8869) );
  OR2_X1 U11618 ( .A1(n8232), .A2(n8783), .ZN(n8088) );
  NAND2_X1 U11619 ( .A1(n8084), .A2(n11716), .ZN(n11733) );
  INV_X1 U11620 ( .A(n9062), .ZN(n8974) );
  OAI211_X1 U11621 ( .C1(n8777), .C2(n8776), .A(n8775), .B(n8774), .ZN(n8778)
         );
  NAND2_X1 U11622 ( .A1(\DataPath/i_PIPLIN_A[18] ), .A2(n7692), .ZN(n9246) );
  NOR2_X1 U11623 ( .A1(n10359), .A2(n10354), .ZN(n8114) );
  NAND2_X1 U11624 ( .A1(\DataPath/i_PIPLIN_A[27] ), .A2(n7692), .ZN(n9460) );
  NAND2_X1 U11625 ( .A1(\DataPath/i_PIPLIN_A[25] ), .A2(n8442), .ZN(n9846) );
  INV_X1 U11626 ( .A(i_RD1[14]), .ZN(n8541) );
  INV_X1 U11627 ( .A(i_RD1[2]), .ZN(n8585) );
  OR2_X1 U11628 ( .A1(\intadd_1/n16 ), .A2(\intadd_1/n11 ), .ZN(n8118) );
  OR2_X1 U11629 ( .A1(\intadd_0/n25 ), .A2(\intadd_0/n22 ), .ZN(n8124) );
  XNOR2_X1 U11630 ( .A(n7782), .B(n9528), .ZN(n8927) );
  AND3_X1 U11631 ( .A1(n165), .A2(n8287), .A3(n172), .ZN(n8135) );
  AND4_X1 U11632 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(n8161)
         );
  NAND2_X1 U11633 ( .A1(n8686), .A2(i_RD1[31]), .ZN(n8782) );
  AND2_X1 U11634 ( .A1(\intadd_2/n15 ), .A2(n8120), .ZN(n8164) );
  INV_X1 U11635 ( .A(n8769), .ZN(n8697) );
  AND4_X1 U11636 ( .A1(n8738), .A2(n8733), .A3(n8581), .A4(n8734), .ZN(n8165)
         );
  INV_X1 U11637 ( .A(n9361), .ZN(n9592) );
  XNOR2_X1 U11638 ( .A(\DP_OP_751_130_6421/n495 ), .B(n9439), .ZN(n8938) );
  AND2_X1 U11639 ( .A1(n10822), .A2(n8462), .ZN(n8171) );
  NOR2_X1 U11640 ( .A1(n9053), .A2(n8975), .ZN(n10011) );
  OR2_X1 U11641 ( .A1(i_ALU_OP[0]), .A2(n8174), .ZN(n8193) );
  INV_X1 U11642 ( .A(i_RD1[11]), .ZN(n8566) );
  INV_X1 U11643 ( .A(i_RD1[7]), .ZN(n8579) );
  INV_X1 U11644 ( .A(i_RD1[13]), .ZN(n8514) );
  INV_X1 U11645 ( .A(i_RD1[15]), .ZN(n8543) );
  INV_X1 U11646 ( .A(i_RD1[3]), .ZN(n8587) );
  INV_X1 U11647 ( .A(i_RD1[0]), .ZN(n8528) );
  OAI21_X1 U11648 ( .B1(n7716), .B2(n8088), .A(n8225), .ZN(n8228) );
  NAND2_X1 U11649 ( .A1(n8228), .A2(n8226), .ZN(n10106) );
  AOI21_X1 U11650 ( .B1(n8088), .B2(n7751), .A(n8229), .ZN(n8227) );
  OAI21_X1 U11651 ( .B1(n8173), .B2(\DataPath/RF/c_swin[1] ), .A(n8237), .ZN(
        n8236) );
  NAND2_X1 U11652 ( .A1(\DataPath/RF/c_swin[2] ), .A2(n8273), .ZN(n8237) );
  OAI21_X1 U11653 ( .B1(n590), .B2(\DataPath/RF/c_swin[0] ), .A(n8249), .ZN(
        n8248) );
  NAND2_X1 U11654 ( .A1(\DataPath/RF/c_win[0] ), .A2(n836), .ZN(n8249) );
  NOR2_X1 U11655 ( .A1(n8252), .A2(n8251), .ZN(n8825) );
  OAI22_X1 U11656 ( .A1(n11830), .A2(n11624), .B1(n11828), .B2(n8455), .ZN(
        n7081) );
  INV_X1 U11657 ( .A(n10304), .ZN(n8270) );
  OAI21_X1 U11658 ( .B1(n7630), .B2(n7635), .A(n8862), .ZN(n8863) );
  NAND2_X1 U11659 ( .A1(n7727), .A2(n7635), .ZN(n9016) );
  OR2_X1 U11660 ( .A1(n2872), .A2(\CU_I/i_FILL_delay ), .ZN(n8480) );
  AOI21_X1 U11661 ( .B1(n8053), .B2(n8481), .A(n8480), .ZN(n8482) );
  XNOR2_X1 U11662 ( .A(n7917), .B(n10190), .ZN(n10193) );
  NAND2_X1 U11663 ( .A1(\intadd_1/n36 ), .A2(\intadd_1/n30 ), .ZN(
        \intadd_1/n5 ) );
  OAI22_X1 U11664 ( .A1(n10099), .A2(n173), .B1(n183), .B2(n10098), .ZN(n10094) );
  OAI22_X1 U11665 ( .A1(n10099), .A2(n174), .B1(n184), .B2(n10098), .ZN(n10096) );
  OAI22_X1 U11666 ( .A1(n10099), .A2(n175), .B1(n10098), .B2(n8136), .ZN(
        n10100) );
  NAND2_X1 U11667 ( .A1(n10105), .A2(n10059), .ZN(n8711) );
  NOR2_X1 U11668 ( .A1(n10099), .A2(n584), .ZN(n8698) );
  NOR2_X1 U11669 ( .A1(n10099), .A2(n582), .ZN(n8667) );
  OR2_X1 U11670 ( .A1(n10099), .A2(n570), .ZN(n8534) );
  NOR2_X1 U11671 ( .A1(n10099), .A2(n578), .ZN(n8517) );
  NOR2_X1 U11672 ( .A1(n10099), .A2(n580), .ZN(n8660) );
  NOR2_X1 U11673 ( .A1(n10099), .A2(n576), .ZN(n8611) );
  NOR2_X1 U11674 ( .A1(n10099), .A2(n583), .ZN(n8501) );
  OR2_X1 U11675 ( .A1(n10099), .A2(n568), .ZN(n8512) );
  NOR2_X1 U11676 ( .A1(n10099), .A2(n574), .ZN(n8634) );
  NOR2_X1 U11677 ( .A1(n10099), .A2(n572), .ZN(n8640) );
  NOR2_X1 U11678 ( .A1(n10099), .A2(n566), .ZN(n8559) );
  OR2_X1 U11679 ( .A1(n10099), .A2(n564), .ZN(n8554) );
  OR2_X1 U11680 ( .A1(n10099), .A2(n562), .ZN(n8577) );
  OAI211_X1 U11681 ( .C1(n10099), .C2(n8166), .A(n8524), .B(n8523), .ZN(n10117) );
  NOR2_X1 U11682 ( .A1(n10099), .A2(n560), .ZN(n8703) );
  OR2_X1 U11683 ( .A1(n10099), .A2(n556), .ZN(n8599) );
  NOR2_X1 U11684 ( .A1(n10099), .A2(n555), .ZN(n8526) );
  NOR2_X1 U11685 ( .A1(n10099), .A2(n558), .ZN(n8573) );
  INV_X1 U11686 ( .A(n10059), .ZN(n10139) );
  OR2_X1 U11687 ( .A1(\DataPath/RF/c_win[0] ), .A2(n8117), .ZN(n8283) );
  OR2_X1 U11688 ( .A1(n8273), .A2(\DataPath/RF/c_swin[0] ), .ZN(n8284) );
  NAND3_X1 U11689 ( .A1(n10306), .A2(n8284), .A3(n8283), .ZN(n10307) );
  AOI22_X1 U11690 ( .A1(n10258), .A2(IRAM_DATA[27]), .B1(n7969), .B2(n10257), 
        .ZN(n10259) );
  AOI21_X1 U11691 ( .B1(n7969), .B2(n8130), .A(n166), .ZN(n8471) );
  OR2_X1 U11692 ( .A1(n7969), .A2(n172), .ZN(n10138) );
  NAND2_X1 U11693 ( .A1(n7969), .A2(n8279), .ZN(n10066) );
  OR2_X1 U11694 ( .A1(n7969), .A2(n8280), .ZN(n10140) );
  AND2_X1 U11695 ( .A1(\DataPath/RF/c_win[1] ), .A2(n835), .ZN(n8289) );
  NOR3_X1 U11696 ( .A1(n10305), .A2(n8289), .A3(n8288), .ZN(n10306) );
  INV_X1 U11697 ( .A(n11647), .ZN(n10309) );
  NAND2_X1 U11698 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[31] ), .ZN(n8939)
         );
  NAND2_X1 U11699 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[30] ), .ZN(n8940)
         );
  NAND2_X1 U11700 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[28] ), .ZN(n8933)
         );
  NAND2_X1 U11701 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[29] ), .ZN(n8932)
         );
  NAND2_X1 U11702 ( .A1(n7907), .A2(\DataPath/i_PIPLIN_IN2[26] ), .ZN(n8929)
         );
  NAND2_X1 U11703 ( .A1(i_S2), .A2(\DataPath/i_PIPLIN_IN2[0] ), .ZN(n8836) );
  NAND2_X1 U11704 ( .A1(i_S2), .A2(\DataPath/i_PIPLIN_IN2[2] ), .ZN(n8861) );
  NAND2_X1 U11705 ( .A1(i_S2), .A2(\DataPath/i_PIPLIN_IN2[3] ), .ZN(n8859) );
  AOI22_X1 U11706 ( .A1(n7647), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[1] ), .ZN(n2398) );
  XNOR2_X1 U11707 ( .A(n10177), .B(n10176), .ZN(n10179) );
  OAI21_X1 U11708 ( .B1(n7894), .B2(n10196), .A(n10195), .ZN(n8809) );
  NOR3_X1 U11709 ( .A1(n10177), .A2(n8103), .A3(n8185), .ZN(n10156) );
  NOR2_X1 U11710 ( .A1(n8816), .A2(n8815), .ZN(n10191) );
  NOR2_X1 U11711 ( .A1(\intadd_1/n22 ), .A2(\intadd_1/n25 ), .ZN(
        \intadd_1/n20 ) );
  OAI21_X1 U11712 ( .B1(\intadd_1/n22 ), .B2(\intadd_1/n26 ), .A(
        \intadd_1/n23 ), .ZN(\intadd_1/n21 ) );
  NAND2_X1 U11713 ( .A1(\intadd_1/B[2] ), .A2(n8133), .ZN(\intadd_1/n23 ) );
  NOR2_X1 U11714 ( .A1(\intadd_1/B[2] ), .A2(n8133), .ZN(\intadd_1/n22 ) );
  OAI21_X1 U11715 ( .B1(n8725), .B2(n8724), .A(n8723), .ZN(n8729) );
  AOI21_X1 U11716 ( .B1(n10092), .B2(n8456), .A(n8600), .ZN(n8605) );
  AND2_X1 U11717 ( .A1(n8129), .A2(n471), .ZN(n8292) );
  AOI21_X1 U11718 ( .B1(n8270), .B2(n7698), .A(n11846), .ZN(n11637) );
  NOR2_X1 U11719 ( .A1(n10295), .A2(n11840), .ZN(n10294) );
  INV_X1 U11720 ( .A(n10216), .ZN(n10234) );
  OAI22_X1 U11721 ( .A1(n10236), .A2(n10216), .B1(n10067), .B2(n10065), .ZN(
        n10035) );
  AND2_X1 U11722 ( .A1(n7969), .A2(n8287), .ZN(n10225) );
  AOI21_X1 U11723 ( .B1(n8287), .B2(n8090), .A(n7969), .ZN(n10222) );
  OAI21_X1 U11724 ( .B1(n8473), .B2(n10059), .A(n7720), .ZN(n8474) );
  AOI22_X1 U11725 ( .A1(n10258), .A2(n11614), .B1(n8287), .B2(n10257), .ZN(
        n7124) );
  AND2_X1 U11726 ( .A1(n7954), .A2(n7720), .ZN(n10060) );
  NOR2_X1 U11727 ( .A1(n7720), .A2(n8135), .ZN(n8486) );
  NAND2_X1 U11728 ( .A1(n8485), .A2(n8287), .ZN(n8487) );
  INV_X1 U11729 ( .A(n7720), .ZN(n8795) );
  OAI21_X1 U11730 ( .B1(n8287), .B2(n8280), .A(n7969), .ZN(n8793) );
  NAND2_X1 U11731 ( .A1(n8496), .A2(n8287), .ZN(n8497) );
  AOI22_X1 U11732 ( .A1(n10091), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_IN2[2] ), .ZN(n2396) );
  XNOR2_X1 U11733 ( .A(n7697), .B(n10199), .ZN(n10201) );
  OAI211_X1 U11734 ( .C1(n10162), .C2(n8050), .A(n10158), .B(n10210), .ZN(
        n10160) );
  NAND2_X1 U11735 ( .A1(n10159), .A2(n10169), .ZN(n10261) );
  NOR2_X1 U11736 ( .A1(\intadd_1/B[0] ), .A2(\intadd_1/A[0] ), .ZN(
        \intadd_1/n29 ) );
  NAND2_X1 U11737 ( .A1(\intadd_1/B[0] ), .A2(\intadd_1/A[0] ), .ZN(
        \intadd_1/n30 ) );
  NAND4_X1 U11738 ( .A1(n8736), .A2(n8730), .A3(n7717), .A4(n8606), .ZN(n8607)
         );
  NAND2_X1 U11739 ( .A1(n8719), .A2(n8718), .ZN(n8722) );
  AOI21_X1 U11740 ( .B1(n10091), .B2(n8456), .A(n8584), .ZN(n8601) );
  XNOR2_X1 U11741 ( .A(\intadd_0/n41 ), .B(\intadd_0/n5 ), .ZN(
        \intadd_0/SUM[0] ) );
  AOI22_X1 U11742 ( .A1(n10264), .A2(n10263), .B1(n10262), .B2(n10261), .ZN(
        n10265) );
  XNOR2_X1 U11743 ( .A(\intadd_2/n33 ), .B(\intadd_2/n4 ), .ZN(
        \intadd_2/SUM[0] ) );
  AOI21_X1 U11744 ( .B1(\intadd_0/n41 ), .B2(n8122), .A(\intadd_0/n38 ), .ZN(
        \intadd_0/n36 ) );
  AOI21_X1 U11745 ( .B1(\intadd_0/n41 ), .B2(\intadd_0/n16 ), .A(
        \intadd_0/n17 ), .ZN(\intadd_0/n15 ) );
  AOI21_X1 U11746 ( .B1(\intadd_2/n33 ), .B2(n8123), .A(\intadd_2/n30 ), .ZN(
        \intadd_2/n28 ) );
  AOI21_X1 U11747 ( .B1(\intadd_2/n33 ), .B2(\intadd_2/n15 ), .A(
        \intadd_2/n16 ), .ZN(\intadd_2/n14 ) );
  AOI21_X1 U11748 ( .B1(\intadd_0/n41 ), .B2(\intadd_0/n28 ), .A(
        \intadd_0/n29 ), .ZN(\intadd_0/n27 ) );
  NOR2_X1 U11749 ( .A1(n7737), .A2(n8137), .ZN(n8817) );
  OR2_X1 U11750 ( .A1(n7737), .A2(n8101), .ZN(n8805) );
  OR2_X1 U11751 ( .A1(n7736), .A2(n8139), .ZN(n10194) );
  NOR2_X1 U11752 ( .A1(n7737), .A2(n8098), .ZN(n10198) );
  NAND2_X1 U11753 ( .A1(n8813), .A2(IR[13]), .ZN(\intadd_0/B[2] ) );
  NAND2_X1 U11754 ( .A1(n8813), .A2(n8134), .ZN(\intadd_0/B[3] ) );
  NAND2_X1 U11755 ( .A1(n8813), .A2(n8099), .ZN(\intadd_0/B[0] ) );
  NAND2_X1 U11756 ( .A1(n8813), .A2(n8100), .ZN(\intadd_0/B[1] ) );
  NOR2_X1 U11757 ( .A1(n7737), .A2(n8107), .ZN(n8806) );
  NOR2_X1 U11758 ( .A1(n7735), .A2(IR[2]), .ZN(\intadd_1/B[1] ) );
  NAND4_X1 U11759 ( .A1(n8165), .A2(n8721), .A3(n8739), .A4(n8591), .ZN(n8608)
         );
  OAI21_X1 U11760 ( .B1(n8732), .B2(n8731), .A(n8730), .ZN(n8735) );
  OAI211_X1 U11761 ( .C1(n8705), .C2(n183), .A(n8535), .B(n8534), .ZN(n10132)
         );
  OAI211_X1 U11762 ( .C1(n8705), .C2(n184), .A(n8539), .B(n8538), .ZN(n10130)
         );
  OAI211_X1 U11763 ( .C1(n8705), .C2(n8136), .A(n8512), .B(n8511), .ZN(n10128)
         );
  OAI211_X1 U11764 ( .C1(n8705), .C2(n185), .A(n8508), .B(n8507), .ZN(n10126)
         );
  OAI211_X1 U11765 ( .C1(n8705), .C2(n8137), .A(n8562), .B(n8561), .ZN(n10124)
         );
  OAI21_X1 U11766 ( .B1(n8705), .B2(n186), .A(n8560), .ZN(n10087) );
  OAI211_X1 U11767 ( .C1(n8705), .C2(n8139), .A(n8550), .B(n8549), .ZN(n10122)
         );
  AOI21_X1 U11768 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(n8725) );
  OAI211_X1 U11769 ( .C1(n8705), .C2(n8101), .A(n8554), .B(n8553), .ZN(n10088)
         );
  OAI211_X1 U11770 ( .C1(n8705), .C2(n8098), .A(n8577), .B(n8576), .ZN(n10089)
         );
  OAI211_X1 U11771 ( .C1(n8705), .C2(n8107), .A(n8595), .B(n8594), .ZN(n10120)
         );
  OAI21_X1 U11772 ( .B1(n8705), .B2(n8096), .A(n8704), .ZN(n10090) );
  OAI21_X1 U11773 ( .B1(n7721), .B2(n8097), .A(n8574), .ZN(n10115) );
  OAI21_X1 U11774 ( .B1(n7721), .B2(n8086), .A(n8527), .ZN(n10113) );
  OAI211_X1 U11775 ( .C1(n7721), .C2(n8094), .A(n8599), .B(n8598), .ZN(n10092)
         );
  OAI211_X1 U11776 ( .C1(n7721), .C2(n8196), .A(n8583), .B(n8582), .ZN(n10091)
         );
  NAND2_X1 U11777 ( .A1(n165), .A2(n167), .ZN(n8492) );
  NAND2_X1 U11778 ( .A1(n8279), .A2(n167), .ZN(n10065) );
  INV_X1 U11779 ( .A(n9689), .ZN(n8300) );
  INV_X1 U11780 ( .A(n8320), .ZN(n8322) );
  INV_X1 U11781 ( .A(n8320), .ZN(n8323) );
  INV_X1 U11782 ( .A(n7768), .ZN(n8324) );
  INV_X1 U11783 ( .A(n7937), .ZN(n8325) );
  INV_X1 U11784 ( .A(\intadd_1/n16 ), .ZN(\intadd_1/n33 ) );
  INV_X1 U11785 ( .A(n7719), .ZN(\intadd_1/n15 ) );
  INV_X1 U11786 ( .A(\intadd_1/n19 ), .ZN(\intadd_1/n18 ) );
  INV_X1 U11787 ( .A(\intadd_1/n28 ), .ZN(\intadd_1/n27 ) );
  INV_X1 U11788 ( .A(\intadd_1/CI ), .ZN(\intadd_1/n31 ) );
  INV_X1 U11789 ( .A(\intadd_1/n11 ), .ZN(\intadd_1/n32 ) );
  INV_X1 U11790 ( .A(\intadd_1/n22 ), .ZN(\intadd_1/n34 ) );
  INV_X1 U11791 ( .A(n7939), .ZN(\intadd_1/n35 ) );
  INV_X1 U11792 ( .A(\intadd_1/n29 ), .ZN(\intadd_1/n36 ) );
  INV_X1 U11793 ( .A(\intadd_1/n10 ), .ZN(\intadd_1/n8 ) );
  INV_X1 U11794 ( .A(\intadd_0/n21 ), .ZN(\intadd_0/n19 ) );
  INV_X1 U11795 ( .A(\intadd_0/n30 ), .ZN(\intadd_0/n28 ) );
  INV_X1 U11796 ( .A(\intadd_0/n31 ), .ZN(\intadd_0/n29 ) );
  INV_X1 U11797 ( .A(\intadd_0/n35 ), .ZN(\intadd_0/n33 ) );
  INV_X1 U11798 ( .A(\intadd_0/n40 ), .ZN(\intadd_0/n38 ) );
  INV_X1 U11799 ( .A(\intadd_0/n22 ), .ZN(\intadd_0/n44 ) );
  INV_X1 U11800 ( .A(\intadd_0/n25 ), .ZN(\intadd_0/n45 ) );
  INV_X1 U11801 ( .A(\intadd_2/n13 ), .ZN(\intadd_2/n11 ) );
  INV_X1 U11802 ( .A(\intadd_2/n27 ), .ZN(\intadd_2/n25 ) );
  INV_X1 U11803 ( .A(\intadd_2/n32 ), .ZN(\intadd_2/n30 ) );
  MUX2_X1 U11804 ( .A(n8487), .B(n8486), .S(n8115), .Z(n8488) );
  NAND3_X1 U11805 ( .A1(n10226), .A2(IR[27]), .A3(n8489), .ZN(n8490) );
  NAND3_X1 U11806 ( .A1(n10272), .A2(n8522), .A3(IR[4]), .ZN(n8523) );
  NAND3_X1 U11807 ( .A1(n8532), .A2(n7640), .A3(n8531), .ZN(n8533) );
  MUX2_X1 U11808 ( .A(n10087), .B(i_RD2[11]), .S(n7856), .Z(n8570) );
  MUX2_X1 U11809 ( .A(n10115), .B(i_RD2[3]), .S(i_SEL_CMPB), .Z(n8588) );
  MUX2_X1 U11810 ( .A(i_RD2[18]), .B(n10084), .S(n8456), .Z(n8647) );
  NAND3_X1 U11811 ( .A1(n8695), .A2(n8654), .A3(n8653), .ZN(n8655) );
  MUX2_X1 U11812 ( .A(i_RD2[26]), .B(n10077), .S(n8456), .Z(n8675) );
  NAND3_X1 U11813 ( .A1(n8781), .A2(n8780), .A3(n8779), .ZN(n8783) );
  MUX2_X1 U11814 ( .A(n8787), .B(n8786), .S(n10106), .Z(n8791) );
  XOR2_X1 U11815 ( .A(n8810), .B(n8809), .Z(n11670) );
  XOR2_X1 U11816 ( .A(n10148), .B(n8828), .Z(n11675) );
  MUX2_X1 U11817 ( .A(n7709), .B(n8116), .S(n9071), .Z(n8862) );
  NAND3_X1 U11818 ( .A1(n8947), .A2(n9020), .A3(n8950), .ZN(n9682) );
  NAND3_X1 U11819 ( .A1(n8962), .A2(n9020), .A3(n8964), .ZN(n9500) );
  MUX2_X1 U11820 ( .A(n7634), .B(n9246), .S(n8452), .Z(n9299) );
  MUX2_X1 U11821 ( .A(n9607), .B(n9774), .S(i_ALU_OP[2]), .Z(n9588) );
  MUX2_X1 U11822 ( .A(n9527), .B(n9250), .S(n8452), .Z(n9557) );
  NAND3_X1 U11823 ( .A1(n9168), .A2(n9686), .A3(n8990), .ZN(n9001) );
  NAND3_X1 U11824 ( .A1(n9169), .A2(n8993), .A3(n9197), .ZN(n9000) );
  NAND3_X1 U11825 ( .A1(n9197), .A2(i_ALU_OP[2]), .A3(i_ALU_OP[4]), .ZN(n9010)
         );
  MUX2_X1 U11826 ( .A(n9779), .B(n11723), .S(n8084), .Z(n9626) );
  NAND3_X1 U11827 ( .A1(n9021), .A2(n9020), .A3(n9029), .ZN(n9390) );
  MUX2_X1 U11828 ( .A(n9026), .B(n8428), .S(n8452), .Z(n9391) );
  NAND3_X1 U11829 ( .A1(n9089), .A2(n9088), .A3(n7766), .ZN(n9092) );
  NAND3_X1 U11830 ( .A1(n9092), .A2(n9091), .A3(n9090), .ZN(n9097) );
  NAND3_X1 U11831 ( .A1(n9117), .A2(n9116), .A3(n9115), .ZN(n9120) );
  XOR2_X1 U11832 ( .A(n11713), .B(n9150), .Z(n9136) );
  MUX2_X1 U11833 ( .A(n9850), .B(n9797), .S(n9129), .Z(n9132) );
  MUX2_X1 U11834 ( .A(n9850), .B(n9795), .S(n7705), .Z(n9131) );
  MUX2_X1 U11835 ( .A(n9132), .B(n9131), .S(n9130), .Z(n9133) );
  NAND3_X1 U11836 ( .A1(n9556), .A2(n9197), .A3(n9168), .ZN(n9175) );
  MUX2_X1 U11837 ( .A(n9795), .B(n9850), .S(n9182), .Z(n9185) );
  MUX2_X1 U11838 ( .A(n9850), .B(n9797), .S(n9182), .Z(n9184) );
  MUX2_X1 U11839 ( .A(n9185), .B(n9184), .S(n9183), .Z(n9186) );
  MUX2_X1 U11840 ( .A(n9795), .B(n9850), .S(n9191), .Z(n9193) );
  MUX2_X1 U11841 ( .A(n9850), .B(n9797), .S(n9191), .Z(n9192) );
  MUX2_X1 U11842 ( .A(n9193), .B(n9192), .S(n9230), .Z(n9217) );
  NAND3_X1 U11843 ( .A1(n9198), .A2(n9197), .A3(i_ALU_OP[4]), .ZN(n9200) );
  XOR2_X1 U11844 ( .A(n9358), .B(n9357), .Z(n9360) );
  NAND3_X1 U11845 ( .A1(n9992), .A2(n9361), .A3(\DP_OP_751_130_6421/n291 ), 
        .ZN(n9364) );
  NAND3_X1 U11846 ( .A1(n9362), .A2(n9990), .A3(n9592), .ZN(n9363) );
  NAND3_X1 U11847 ( .A1(n9430), .A2(n9429), .A3(n9428), .ZN(n9431) );
  MUX2_X1 U11848 ( .A(n9795), .B(n9850), .S(n9439), .Z(n9440) );
  MUX2_X1 U11849 ( .A(n9457), .B(n9456), .S(n9515), .Z(n9468) );
  NAND3_X1 U11850 ( .A1(n9992), .A2(n9459), .A3(\DP_OP_751_130_6421/n495 ), 
        .ZN(n9463) );
  NAND3_X1 U11851 ( .A1(n9461), .A2(n9990), .A3(n9460), .ZN(n9462) );
  MUX2_X1 U11852 ( .A(n9795), .B(n9850), .S(n9516), .Z(n9519) );
  MUX2_X1 U11853 ( .A(n9850), .B(n9797), .S(n9516), .Z(n9518) );
  MUX2_X1 U11854 ( .A(n9519), .B(n9518), .S(n9517), .Z(n9520) );
  MUX2_X1 U11855 ( .A(n9990), .B(n9803), .S(n9526), .Z(n9530) );
  MUX2_X1 U11856 ( .A(n9992), .B(n9803), .S(n9527), .Z(n9529) );
  MUX2_X1 U11857 ( .A(n9530), .B(n9529), .S(n9528), .Z(n9531) );
  NAND3_X1 U11858 ( .A1(n9888), .A2(n9606), .A3(n9605), .ZN(n9614) );
  MUX2_X1 U11859 ( .A(n9795), .B(n9850), .S(n11723), .Z(n9648) );
  MUX2_X1 U11860 ( .A(n9850), .B(n9797), .S(n11723), .Z(n9647) );
  MUX2_X1 U11861 ( .A(n9648), .B(n9647), .S(n9646), .Z(n9649) );
  MUX2_X1 U11862 ( .A(n9662), .B(n9661), .S(n9327), .Z(n9663) );
  NAND3_X1 U11863 ( .A1(n9992), .A2(n9711), .A3(\DP_OP_751_130_6421/n903 ), 
        .ZN(n9714) );
  NAND3_X1 U11864 ( .A1(n9712), .A2(n9990), .A3(n7693), .ZN(n9713) );
  NAND3_X1 U11865 ( .A1(n9751), .A2(n9734), .A3(n9733), .ZN(n9739) );
  MUX2_X1 U11866 ( .A(n9795), .B(n9850), .S(n7749), .Z(n9737) );
  MUX2_X1 U11867 ( .A(n9850), .B(n9797), .S(n7749), .Z(n9736) );
  MUX2_X1 U11868 ( .A(n9737), .B(n9736), .S(n9735), .Z(n9738) );
  MUX2_X1 U11869 ( .A(n9990), .B(n9803), .S(n9755), .Z(n9749) );
  NAND3_X1 U11870 ( .A1(n9754), .A2(n9996), .A3(n9989), .ZN(n9758) );
  MUX2_X1 U11871 ( .A(n9803), .B(n9992), .S(n9755), .Z(n9756) );
  MUX2_X1 U11872 ( .A(n9992), .B(n9803), .S(n7688), .Z(n9800) );
  MUX2_X1 U11873 ( .A(n9990), .B(n9803), .S(n7685), .Z(n9804) );
  MUX2_X1 U11874 ( .A(n9808), .B(n9807), .S(n9806), .Z(n9814) );
  XOR2_X1 U11875 ( .A(n9845), .B(n9844), .Z(n9853) );
  NAND3_X1 U11876 ( .A1(n9992), .A2(n7691), .A3(\DP_OP_751_130_6421/n597 ), 
        .ZN(n9849) );
  NAND3_X1 U11877 ( .A1(n9847), .A2(n9990), .A3(n9846), .ZN(n9848) );
  NAND3_X1 U11878 ( .A1(n9992), .A2(n9889), .A3(\DP_OP_751_130_6421/n801 ), 
        .ZN(n9892) );
  NAND3_X1 U11879 ( .A1(n9890), .A2(n9990), .A3(n9904), .ZN(n9891) );
  NAND3_X1 U11880 ( .A1(n8447), .A2(n9990), .A3(n9951), .ZN(n9934) );
  NAND3_X1 U11881 ( .A1(n9992), .A2(n9932), .A3(\DP_OP_751_130_6421/n1413 ), 
        .ZN(n9933) );
  NAND3_X1 U11882 ( .A1(n9950), .A2(n9949), .A3(n9948), .ZN(n9955) );
  XOR2_X1 U11883 ( .A(\DP_OP_751_130_6421/n1413 ), .B(n8304), .Z(n9952) );
  NAND3_X1 U11884 ( .A1(n9992), .A2(n9966), .A3(\DP_OP_751_130_6421/n1209 ), 
        .ZN(n9968) );
  NAND3_X1 U11885 ( .A1(n8448), .A2(n9990), .A3(n9972), .ZN(n9967) );
  NAND3_X1 U11886 ( .A1(n8449), .A2(n9990), .A3(n10005), .ZN(n9994) );
  NAND3_X1 U11887 ( .A1(n9992), .A2(n9991), .A3(\DP_OP_751_130_6421/n1005 ), 
        .ZN(n9993) );
  NAND3_X1 U11888 ( .A1(n10300), .A2(n10069), .A3(n10068), .ZN(n10070) );
  NAND3_X1 U11889 ( .A1(n10106), .A2(n7753), .A3(n10105), .ZN(n10107) );
  XOR2_X1 U11890 ( .A(IRAM_ADDRESS[25]), .B(n10175), .Z(n10180) );
  XOR2_X1 U11891 ( .A(IRAM_ADDRESS[27]), .B(n10175), .Z(n10171) );
  XOR2_X1 U11892 ( .A(IRAM_ADDRESS[0]), .B(n10211), .Z(n10212) );
  NAND3_X1 U11893 ( .A1(n7954), .A2(n8287), .A3(n10236), .ZN(n10214) );
  NAND3_X1 U11894 ( .A1(n10230), .A2(n10271), .A3(n10229), .ZN(
        \CU_I/CW[RF_RD2_EN] ) );
  NAND3_X1 U11895 ( .A1(n10297), .A2(n10238), .A3(n10237), .ZN(
        \CU_I/CW[RF_RD1_EN] ) );
  OAI211_X1 U11897 ( .C1(n166), .C2(n8287), .A(IR[31]), .B(n165), .ZN(n10301)
         );
  NAND3_X1 U11898 ( .A1(n166), .A2(n165), .A3(IR[31]), .ZN(n10302) );
  NOR2_X1 U11899 ( .A1(n10297), .A2(n10302), .ZN(\CU_I/CW[WB_MUX_SEL] ) );
  NOR2_X1 U11900 ( .A1(n7969), .A2(n10302), .ZN(n10303) );
  NOR2_X1 U11901 ( .A1(n10296), .A2(n11667), .ZN(\CU_I/CW_IF[WB_EN] ) );
  AND2_X1 U11902 ( .A1(n10300), .A2(\CU_I/CW_MEM[WB_EN] ), .ZN(\CU_I/N301 ) );
  AND2_X1 U11903 ( .A1(n10300), .A2(\CU_I/CW_MEM[WB_MUX_SEL] ), .ZN(
        \CU_I/N302 ) );
  OAI22_X1 U11904 ( .A1(\DataPath/RF/c_win[3] ), .A2(n8272), .B1(n835), .B2(
        \DataPath/RF/c_win[1] ), .ZN(n10305) );
  NOR2_X1 U11905 ( .A1(RST), .A2(n8054), .ZN(\CU_I/N314 ) );
  NOR2_X1 U11906 ( .A1(n10295), .A2(RST), .ZN(\CU_I/N315 ) );
  NAND2_X1 U11907 ( .A1(n10308), .A2(DRAMRF_READY), .ZN(n10821) );
  XOR2_X1 U11908 ( .A(\DataPath/RF/PUSH_ADDRGEN/curr_state[0] ), .B(n849), .Z(
        n11646) );
  INV_X1 U11909 ( .A(n10815), .ZN(n10818) );
  AOI22_X1 U11910 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[2] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[3] ), .B2(n10314), .ZN(n10329)
         );
  AOI22_X1 U11911 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[1] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[2] ), .B2(n10314), .ZN(n10330)
         );
  NAND2_X1 U11912 ( .A1(n10329), .A2(n10330), .ZN(n10311) );
  AOI22_X1 U11913 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[0] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[1] ), .B2(n10314), .ZN(n10350)
         );
  AOI22_X1 U11914 ( .A1(n10309), .A2(n11646), .B1(
        \DataPath/RF/PUSH_ADDRGEN/curr_addr[0] ), .B2(n10314), .ZN(n10347) );
  NAND2_X1 U11915 ( .A1(n10350), .A2(n10347), .ZN(n10317) );
  NOR2_X1 U11916 ( .A1(n10311), .A2(n10317), .ZN(n10335) );
  AOI22_X1 U11917 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[6] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[7] ), .B2(n10314), .ZN(n10318)
         );
  AOI22_X1 U11918 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[5] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[6] ), .B2(n10314), .ZN(n10325)
         );
  NAND2_X1 U11919 ( .A1(n10318), .A2(n10325), .ZN(n10316) );
  INV_X1 U11920 ( .A(n10316), .ZN(n10310) );
  AOI22_X1 U11921 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[4] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[5] ), .B2(n10314), .ZN(n10328)
         );
  AOI22_X1 U11922 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[3] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[4] ), .B2(n10314), .ZN(n10327)
         );
  AND2_X1 U11923 ( .A1(n10328), .A2(n10327), .ZN(n10315) );
  NAND2_X1 U11924 ( .A1(n10310), .A2(n10315), .ZN(n10336) );
  OAI21_X1 U11925 ( .B1(n10821), .B2(n8104), .A(n8224), .ZN(n10820) );
  NAND2_X1 U11926 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[13] ), 
        .ZN(n10819) );
  INV_X1 U11927 ( .A(n10819), .ZN(n10312) );
  AOI21_X1 U11928 ( .B1(n10314), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[14] ), 
        .A(n10312), .ZN(n10322) );
  INV_X1 U11929 ( .A(n10322), .ZN(n10313) );
  NOR2_X1 U11930 ( .A1(n10820), .A2(n10313), .ZN(n10331) );
  AOI22_X1 U11931 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[9] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[10] ), .B2(n10314), .ZN(n10319) );
  AOI22_X1 U11932 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[10] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[11] ), .B2(n10314), .ZN(n10324) );
  NAND2_X1 U11933 ( .A1(n10319), .A2(n10324), .ZN(n10333) );
  AOI22_X1 U11934 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[12] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[13] ), .B2(n10314), .ZN(n10320) );
  AOI22_X1 U11935 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[11] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[12] ), .B2(n10314), .ZN(n10321) );
  NAND2_X1 U11936 ( .A1(n10320), .A2(n10321), .ZN(n10334) );
  AOI22_X1 U11937 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[8] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[9] ), .B2(n10314), .ZN(n10323)
         );
  AOI22_X1 U11938 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[7] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[8] ), .B2(n10314), .ZN(n10326)
         );
  NAND2_X1 U11939 ( .A1(n10323), .A2(n10326), .ZN(n10332) );
  NAND2_X1 U11940 ( .A1(n10353), .A2(n10349), .ZN(n10341) );
  NOR2_X1 U11941 ( .A1(n10333), .A2(n10332), .ZN(n10338) );
  INV_X1 U11942 ( .A(n10338), .ZN(n10339) );
  NAND2_X1 U11943 ( .A1(n10337), .A2(n10357), .ZN(n10354) );
  NOR2_X1 U11944 ( .A1(n10354), .A2(n10341), .ZN(n10671) );
  AOI22_X1 U11945 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[192] ), 
        .B1(n8108), .B2(\DataPath/RF/bus_sel_savedwin_data[64] ), .ZN(n10346)
         );
  NOR2_X1 U11946 ( .A1(n10337), .A2(n10336), .ZN(n10340) );
  NAND2_X1 U11947 ( .A1(n10338), .A2(n10340), .ZN(n10358) );
  NOR2_X1 U11948 ( .A1(n10358), .A2(n10341), .ZN(n10670) );
  NAND2_X1 U11949 ( .A1(n10340), .A2(n10339), .ZN(n10355) );
  NOR2_X1 U11950 ( .A1(n10341), .A2(n10355), .ZN(n10673) );
  AOI22_X1 U11951 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[448] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[320] ), .ZN(n10345) );
  INV_X1 U11952 ( .A(n10353), .ZN(n10351) );
  NOR2_X1 U11953 ( .A1(n10355), .A2(n10342), .ZN(n10667) );
  NOR2_X1 U11954 ( .A1(n10358), .A2(n10342), .ZN(n10672) );
  AOI22_X1 U11955 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[352] ), 
        .B1(n8343), .B2(\DataPath/RF/bus_sel_savedwin_data[480] ), .ZN(n10344)
         );
  NOR2_X1 U11956 ( .A1(n10354), .A2(n10342), .ZN(n10668) );
  AOI22_X1 U11957 ( .A1(n8345), .A2(\DataPath/RF/bus_sel_savedwin_data[96] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[224] ), .ZN(n10343)
         );
  NAND4_X1 U11958 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10365) );
  INV_X1 U11959 ( .A(n10347), .ZN(n10348) );
  AOI21_X1 U11960 ( .B1(n10350), .B2(n10349), .A(n10348), .ZN(n10352) );
  NAND2_X1 U11961 ( .A1(n10352), .A2(n10351), .ZN(n10359) );
  NOR2_X1 U11962 ( .A1(n10359), .A2(n10357), .ZN(n10679) );
  AOI22_X1 U11963 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[32] ), 
        .B1(n8351), .B2(\DataPath/RF/bus_sel_savedwin_data[160] ), .ZN(n10363)
         );
  NOR2_X1 U11964 ( .A1(n10354), .A2(n10356), .ZN(n10678) );
  NOR2_X1 U11965 ( .A1(n10356), .A2(n10358), .ZN(n10684) );
  AOI22_X1 U11966 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[0] ), 
        .B1(n8111), .B2(\DataPath/RF/bus_sel_savedwin_data[384] ), .ZN(n10362)
         );
  NOR2_X1 U11967 ( .A1(n10356), .A2(n10355), .ZN(n10683) );
  NOR2_X1 U11968 ( .A1(n10359), .A2(n10355), .ZN(n10681) );
  AOI22_X1 U11969 ( .A1(n8353), .A2(\DataPath/RF/bus_sel_savedwin_data[256] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[288] ), .ZN(n10361)
         );
  NOR2_X1 U11970 ( .A1(n10357), .A2(n10356), .ZN(n10680) );
  NOR2_X1 U11971 ( .A1(n10359), .A2(n10358), .ZN(n10682) );
  AOI22_X1 U11972 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[128] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[416] ), .ZN(n10360)
         );
  NAND4_X1 U11973 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10364) );
  OR2_X1 U11974 ( .A1(n10365), .A2(n10364), .ZN(DRAMRF_DATA_OUT[0]) );
  AOI22_X1 U11975 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[362] ), 
        .B1(n8343), .B2(\DataPath/RF/bus_sel_savedwin_data[490] ), .ZN(n10369)
         );
  AOI22_X1 U11976 ( .A1(n8345), .A2(\DataPath/RF/bus_sel_savedwin_data[106] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[234] ), .ZN(n10368)
         );
  AOI22_X1 U11977 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[74] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[330] ), .ZN(n10367) );
  AOI22_X1 U11978 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[202] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[458] ), .ZN(n10366)
         );
  NAND4_X1 U11979 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10375) );
  AOI22_X1 U11980 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[42] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[10] ), .ZN(n10373)
         );
  AOI22_X1 U11981 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[394] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[266] ), .ZN(n10372)
         );
  AOI22_X1 U11982 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[170] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[426] ), .ZN(n10371)
         );
  AOI22_X1 U11983 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[138] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[298] ), .ZN(n10370)
         );
  NAND4_X1 U11984 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10374) );
  OR2_X1 U11985 ( .A1(n10375), .A2(n10374), .ZN(DRAMRF_DATA_OUT[10]) );
  AOI22_X1 U11986 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[203] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[459] ), .ZN(n10379)
         );
  AOI22_X1 U11987 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[75] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[331] ), .ZN(n10378) );
  AOI22_X1 U11988 ( .A1(n8345), .A2(\DataPath/RF/bus_sel_savedwin_data[107] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[235] ), .ZN(n10377)
         );
  AOI22_X1 U11989 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[363] ), 
        .B1(n8343), .B2(\DataPath/RF/bus_sel_savedwin_data[491] ), .ZN(n10376)
         );
  NAND4_X1 U11990 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10385) );
  AOI22_X1 U11991 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[395] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[299] ), .ZN(n10383)
         );
  AOI22_X1 U11992 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[171] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[427] ), .ZN(n10382)
         );
  AOI22_X1 U11993 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[139] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[267] ), .ZN(n10381)
         );
  AOI22_X1 U11994 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[43] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[11] ), .ZN(n10380)
         );
  NAND4_X1 U11995 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10384) );
  OR2_X1 U11996 ( .A1(n10385), .A2(n10384), .ZN(DRAMRF_DATA_OUT[11]) );
  AOI22_X1 U11997 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[204] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[236] ), .ZN(n10389)
         );
  AOI22_X1 U11998 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[332] ), 
        .B1(n8343), .B2(\DataPath/RF/bus_sel_savedwin_data[492] ), .ZN(n10388)
         );
  AOI22_X1 U11999 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[460] ), 
        .B1(n8109), .B2(\DataPath/RF/bus_sel_savedwin_data[364] ), .ZN(n10387)
         );
  AOI22_X1 U12000 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[76] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[108] ), .ZN(n10386)
         );
  NAND4_X1 U12001 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10395) );
  AOI22_X1 U12002 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[140] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[300] ), .ZN(n10393)
         );
  AOI22_X1 U12003 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[12] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[428] ), .ZN(n10392)
         );
  AOI22_X1 U12004 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[44] ), 
        .B1(n10679), .B2(\DataPath/RF/bus_sel_savedwin_data[172] ), .ZN(n10391) );
  AOI22_X1 U12005 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[396] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[268] ), .ZN(n10390) );
  NAND4_X1 U12006 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10394) );
  OR2_X1 U12007 ( .A1(n10395), .A2(n10394), .ZN(DRAMRF_DATA_OUT[12]) );
  AOI22_X1 U12008 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[461] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[333] ), .ZN(n10399) );
  AOI22_X1 U12009 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[493] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[109] ), .ZN(n10398)
         );
  AOI22_X1 U12010 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[365] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[237] ), .ZN(n10397)
         );
  AOI22_X1 U12011 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[205] ), 
        .B1(n8108), .B2(\DataPath/RF/bus_sel_savedwin_data[77] ), .ZN(n10396)
         );
  NAND4_X1 U12012 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10405) );
  AOI22_X1 U12013 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[173] ), 
        .B1(n10680), .B2(\DataPath/RF/bus_sel_savedwin_data[141] ), .ZN(n10403) );
  AOI22_X1 U12014 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[13] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[429] ), .ZN(n10402)
         );
  AOI22_X1 U12015 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[45] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[301] ), .ZN(n10401)
         );
  AOI22_X1 U12016 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[397] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[269] ), .ZN(n10400) );
  NAND4_X1 U12017 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10404) );
  OR2_X1 U12018 ( .A1(n10405), .A2(n10404), .ZN(DRAMRF_DATA_OUT[13]) );
  AOI22_X1 U12019 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[494] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[110] ), .ZN(n10409)
         );
  AOI22_X1 U12020 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[206] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[238] ), .ZN(n10408)
         );
  AOI22_X1 U12021 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[462] ), 
        .B1(n8110), .B2(\DataPath/RF/bus_sel_savedwin_data[334] ), .ZN(n10407)
         );
  AOI22_X1 U12022 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[78] ), 
        .B1(n8109), .B2(\DataPath/RF/bus_sel_savedwin_data[366] ), .ZN(n10406)
         );
  NAND4_X1 U12023 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10415) );
  AOI22_X1 U12024 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[14] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[302] ), .ZN(n10413)
         );
  AOI22_X1 U12025 ( .A1(n8357), .A2(\DataPath/RF/bus_sel_savedwin_data[142] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[270] ), .ZN(n10412) );
  AOI22_X1 U12026 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[46] ), 
        .B1(n10679), .B2(\DataPath/RF/bus_sel_savedwin_data[174] ), .ZN(n10411) );
  AOI22_X1 U12027 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[398] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[430] ), .ZN(n10410)
         );
  NAND4_X1 U12028 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10414) );
  OR2_X1 U12029 ( .A1(n10415), .A2(n10414), .ZN(DRAMRF_DATA_OUT[14]) );
  AOI22_X1 U12030 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[79] ), 
        .B1(n8110), .B2(\DataPath/RF/bus_sel_savedwin_data[335] ), .ZN(n10419)
         );
  AOI22_X1 U12031 ( .A1(n8345), .A2(\DataPath/RF/bus_sel_savedwin_data[111] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[239] ), .ZN(n10418)
         );
  AOI22_X1 U12032 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[463] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[367] ), .ZN(n10417)
         );
  AOI22_X1 U12033 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[207] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[495] ), .ZN(n10416)
         );
  NAND4_X1 U12034 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10425) );
  AOI22_X1 U12035 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[15] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[303] ), .ZN(n10423)
         );
  AOI22_X1 U12036 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[47] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[431] ), .ZN(n10422) );
  AOI22_X1 U12037 ( .A1(n8111), .A2(\DataPath/RF/bus_sel_savedwin_data[399] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[271] ), .ZN(n10421) );
  AOI22_X1 U12038 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[175] ), 
        .B1(n8356), .B2(\DataPath/RF/bus_sel_savedwin_data[143] ), .ZN(n10420)
         );
  NAND4_X1 U12039 ( .A1(n10423), .A2(n10422), .A3(n10421), .A4(n10420), .ZN(
        n10424) );
  OR2_X1 U12040 ( .A1(n10425), .A2(n10424), .ZN(DRAMRF_DATA_OUT[15]) );
  AOI22_X1 U12041 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[496] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[112] ), .ZN(n10429)
         );
  AOI22_X1 U12042 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[464] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[368] ), .ZN(n10428)
         );
  AOI22_X1 U12043 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[208] ), 
        .B1(n10671), .B2(\DataPath/RF/bus_sel_savedwin_data[80] ), .ZN(n10427)
         );
  AOI22_X1 U12044 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[336] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[240] ), .ZN(n10426)
         );
  NAND4_X1 U12045 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10435) );
  AOI22_X1 U12046 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[48] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[144] ), .ZN(n10433)
         );
  AOI22_X1 U12047 ( .A1(n8111), .A2(\DataPath/RF/bus_sel_savedwin_data[400] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[272] ), .ZN(n10432)
         );
  AOI22_X1 U12048 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[176] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[432] ), .ZN(n10431) );
  AOI22_X1 U12049 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[16] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[304] ), .ZN(n10430)
         );
  NAND4_X1 U12050 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10434) );
  OR2_X1 U12051 ( .A1(n10435), .A2(n10434), .ZN(DRAMRF_DATA_OUT[16]) );
  AOI22_X1 U12052 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[209] ), 
        .B1(n10671), .B2(\DataPath/RF/bus_sel_savedwin_data[81] ), .ZN(n10439)
         );
  AOI22_X1 U12053 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[369] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[241] ), .ZN(n10438) );
  AOI22_X1 U12054 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[337] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[113] ), .ZN(n10437) );
  AOI22_X1 U12055 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[465] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[497] ), .ZN(n10436)
         );
  NAND4_X1 U12056 ( .A1(n10439), .A2(n10438), .A3(n10437), .A4(n10436), .ZN(
        n10445) );
  AOI22_X1 U12057 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[17] ), 
        .B1(n8111), .B2(\DataPath/RF/bus_sel_savedwin_data[401] ), .ZN(n10443)
         );
  AOI22_X1 U12058 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[49] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[273] ), .ZN(n10442)
         );
  AOI22_X1 U12059 ( .A1(n8357), .A2(\DataPath/RF/bus_sel_savedwin_data[145] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[433] ), .ZN(n10441)
         );
  AOI22_X1 U12060 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[177] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[305] ), .ZN(n10440) );
  NAND4_X1 U12061 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10444) );
  OR2_X1 U12062 ( .A1(n10445), .A2(n10444), .ZN(DRAMRF_DATA_OUT[17]) );
  AOI22_X1 U12063 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[338] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[370] ), .ZN(n10449)
         );
  AOI22_X1 U12064 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[498] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[114] ), .ZN(n10448) );
  AOI22_X1 U12065 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[466] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[242] ), .ZN(n10447) );
  AOI22_X1 U12066 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[210] ), 
        .B1(n10671), .B2(\DataPath/RF/bus_sel_savedwin_data[82] ), .ZN(n10446)
         );
  NAND4_X1 U12067 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10455) );
  AOI22_X1 U12068 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[178] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[274] ), .ZN(n10453)
         );
  AOI22_X1 U12069 ( .A1(n8357), .A2(\DataPath/RF/bus_sel_savedwin_data[146] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[434] ), .ZN(n10452)
         );
  AOI22_X1 U12070 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[50] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[18] ), .ZN(n10451)
         );
  AOI22_X1 U12071 ( .A1(n8111), .A2(\DataPath/RF/bus_sel_savedwin_data[402] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[306] ), .ZN(n10450) );
  NAND4_X1 U12072 ( .A1(n10453), .A2(n10452), .A3(n10451), .A4(n10450), .ZN(
        n10454) );
  OR2_X1 U12073 ( .A1(n10455), .A2(n10454), .ZN(DRAMRF_DATA_OUT[18]) );
  AOI22_X1 U12074 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[211] ), 
        .B1(n10667), .B2(\DataPath/RF/bus_sel_savedwin_data[371] ), .ZN(n10459) );
  AOI22_X1 U12075 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[467] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[243] ), .ZN(n10458)
         );
  AOI22_X1 U12076 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[83] ), 
        .B1(n8110), .B2(\DataPath/RF/bus_sel_savedwin_data[339] ), .ZN(n10457)
         );
  AOI22_X1 U12077 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[499] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[115] ), .ZN(n10456) );
  NAND4_X1 U12078 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10465) );
  AOI22_X1 U12079 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[147] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[435] ), .ZN(n10463)
         );
  AOI22_X1 U12080 ( .A1(n8111), .A2(\DataPath/RF/bus_sel_savedwin_data[403] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[275] ), .ZN(n10462)
         );
  AOI22_X1 U12081 ( .A1(n10679), .A2(\DataPath/RF/bus_sel_savedwin_data[179] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[307] ), .ZN(n10461)
         );
  AOI22_X1 U12082 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[51] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[19] ), .ZN(n10460)
         );
  NAND4_X1 U12083 ( .A1(n10463), .A2(n10462), .A3(n10461), .A4(n10460), .ZN(
        n10464) );
  OR2_X1 U12084 ( .A1(n10465), .A2(n10464), .ZN(DRAMRF_DATA_OUT[19]) );
  AOI22_X1 U12085 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[193] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[449] ), .ZN(n10469)
         );
  AOI22_X1 U12086 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[353] ), 
        .B1(n10672), .B2(\DataPath/RF/bus_sel_savedwin_data[481] ), .ZN(n10468) );
  AOI22_X1 U12087 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[65] ), 
        .B1(n8110), .B2(\DataPath/RF/bus_sel_savedwin_data[321] ), .ZN(n10467)
         );
  AOI22_X1 U12088 ( .A1(n8346), .A2(\DataPath/RF/bus_sel_savedwin_data[97] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[225] ), .ZN(n10466)
         );
  NAND4_X1 U12089 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10475) );
  AOI22_X1 U12090 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[1] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[289] ), .ZN(n10473)
         );
  AOI22_X1 U12091 ( .A1(n8358), .A2(\DataPath/RF/bus_sel_savedwin_data[417] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[257] ), .ZN(n10472)
         );
  AOI22_X1 U12092 ( .A1(n10679), .A2(\DataPath/RF/bus_sel_savedwin_data[161] ), 
        .B1(n8111), .B2(\DataPath/RF/bus_sel_savedwin_data[385] ), .ZN(n10471)
         );
  AOI22_X1 U12093 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[33] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[129] ), .ZN(n10470)
         );
  NAND4_X1 U12094 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10474) );
  OR2_X1 U12095 ( .A1(n10475), .A2(n10474), .ZN(DRAMRF_DATA_OUT[1]) );
  AOI22_X1 U12096 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[212] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[340] ), .ZN(n10479)
         );
  AOI22_X1 U12097 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[468] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[244] ), .ZN(n10478)
         );
  AOI22_X1 U12098 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[84] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[116] ), .ZN(n10477) );
  AOI22_X1 U12099 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[372] ), 
        .B1(n10672), .B2(\DataPath/RF/bus_sel_savedwin_data[500] ), .ZN(n10476) );
  NAND4_X1 U12100 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10485) );
  AOI22_X1 U12101 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[148] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[308] ), .ZN(n10483)
         );
  AOI22_X1 U12102 ( .A1(n10679), .A2(\DataPath/RF/bus_sel_savedwin_data[180] ), 
        .B1(n8111), .B2(\DataPath/RF/bus_sel_savedwin_data[404] ), .ZN(n10482)
         );
  AOI22_X1 U12103 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[52] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[436] ), .ZN(n10481)
         );
  AOI22_X1 U12104 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[20] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[276] ), .ZN(n10480)
         );
  NAND4_X1 U12105 ( .A1(n10483), .A2(n10482), .A3(n10481), .A4(n10480), .ZN(
        n10484) );
  OR2_X1 U12106 ( .A1(n10485), .A2(n10484), .ZN(DRAMRF_DATA_OUT[20]) );
  AOI22_X1 U12107 ( .A1(n10671), .A2(\DataPath/RF/bus_sel_savedwin_data[85] ), 
        .B1(n8109), .B2(\DataPath/RF/bus_sel_savedwin_data[373] ), .ZN(n10489)
         );
  AOI22_X1 U12108 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[501] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[245] ), .ZN(n10488) );
  AOI22_X1 U12109 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[213] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[341] ), .ZN(n10487)
         );
  AOI22_X1 U12110 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[469] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[117] ), .ZN(n10486)
         );
  NAND4_X1 U12111 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10495) );
  AOI22_X1 U12112 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[181] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[437] ), .ZN(n10493)
         );
  AOI22_X1 U12113 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[405] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[277] ), .ZN(n10492)
         );
  AOI22_X1 U12114 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[21] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[309] ), .ZN(n10491) );
  AOI22_X1 U12115 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[53] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[149] ), .ZN(n10490)
         );
  NAND4_X1 U12116 ( .A1(n10493), .A2(n10492), .A3(n10491), .A4(n10490), .ZN(
        n10494) );
  OR2_X1 U12117 ( .A1(n10495), .A2(n10494), .ZN(DRAMRF_DATA_OUT[21]) );
  AOI22_X1 U12118 ( .A1(n10671), .A2(\DataPath/RF/bus_sel_savedwin_data[86] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[470] ), .ZN(n10499)
         );
  AOI22_X1 U12119 ( .A1(n8344), .A2(\DataPath/RF/bus_sel_savedwin_data[502] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[246] ), .ZN(n10498)
         );
  AOI22_X1 U12120 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[342] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[118] ), .ZN(n10497)
         );
  AOI22_X1 U12121 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[214] ), 
        .B1(n8109), .B2(\DataPath/RF/bus_sel_savedwin_data[374] ), .ZN(n10496)
         );
  NAND4_X1 U12122 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10505) );
  AOI22_X1 U12123 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[54] ), 
        .B1(n10679), .B2(\DataPath/RF/bus_sel_savedwin_data[182] ), .ZN(n10503) );
  AOI22_X1 U12124 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[150] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[278] ), .ZN(n10502)
         );
  AOI22_X1 U12125 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[406] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[310] ), .ZN(n10501)
         );
  AOI22_X1 U12126 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[22] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[438] ), .ZN(n10500)
         );
  NAND4_X1 U12127 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  OR2_X1 U12128 ( .A1(n10505), .A2(n10504), .ZN(DRAMRF_DATA_OUT[22]) );
  AOI22_X1 U12129 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[215] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[247] ), .ZN(n10509)
         );
  AOI22_X1 U12130 ( .A1(n10671), .A2(\DataPath/RF/bus_sel_savedwin_data[87] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[503] ), .ZN(n10508)
         );
  AOI22_X1 U12131 ( .A1(n8342), .A2(\DataPath/RF/bus_sel_savedwin_data[375] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[119] ), .ZN(n10507)
         );
  AOI22_X1 U12132 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[471] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[343] ), .ZN(n10506)
         );
  NAND4_X1 U12133 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10515) );
  AOI22_X1 U12134 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[183] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[23] ), .ZN(n10513)
         );
  AOI22_X1 U12135 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[55] ), 
        .B1(n10684), .B2(\DataPath/RF/bus_sel_savedwin_data[407] ), .ZN(n10512) );
  AOI22_X1 U12136 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[151] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[439] ), .ZN(n10511) );
  AOI22_X1 U12137 ( .A1(n8353), .A2(\DataPath/RF/bus_sel_savedwin_data[279] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[311] ), .ZN(n10510)
         );
  NAND4_X1 U12138 ( .A1(n10513), .A2(n10512), .A3(n10511), .A4(n10510), .ZN(
        n10514) );
  OR2_X1 U12139 ( .A1(n10515), .A2(n10514), .ZN(DRAMRF_DATA_OUT[23]) );
  AOI22_X1 U12140 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[472] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[504] ), .ZN(n10519)
         );
  AOI22_X1 U12141 ( .A1(n10671), .A2(\DataPath/RF/bus_sel_savedwin_data[88] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[248] ), .ZN(n10518)
         );
  AOI22_X1 U12142 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[216] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[120] ), .ZN(n10517)
         );
  AOI22_X1 U12143 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[344] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[376] ), .ZN(n10516)
         );
  NAND4_X1 U12144 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n10525) );
  AOI22_X1 U12145 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[152] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[440] ), .ZN(n10523) );
  AOI22_X1 U12146 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[184] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[280] ), .ZN(n10522)
         );
  AOI22_X1 U12147 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[24] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[312] ), .ZN(n10521)
         );
  AOI22_X1 U12148 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[56] ), 
        .B1(n10684), .B2(\DataPath/RF/bus_sel_savedwin_data[408] ), .ZN(n10520) );
  NAND4_X1 U12149 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10524) );
  OR2_X1 U12150 ( .A1(n10525), .A2(n10524), .ZN(DRAMRF_DATA_OUT[24]) );
  AOI22_X1 U12151 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[217] ), 
        .B1(n10671), .B2(\DataPath/RF/bus_sel_savedwin_data[89] ), .ZN(n10529)
         );
  AOI22_X1 U12152 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[473] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[345] ), .ZN(n10528)
         );
  AOI22_X1 U12153 ( .A1(n8342), .A2(\DataPath/RF/bus_sel_savedwin_data[377] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[505] ), .ZN(n10527)
         );
  AOI22_X1 U12154 ( .A1(n8346), .A2(\DataPath/RF/bus_sel_savedwin_data[121] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[249] ), .ZN(n10526) );
  NAND4_X1 U12155 ( .A1(n10529), .A2(n10528), .A3(n10527), .A4(n10526), .ZN(
        n10535) );
  AOI22_X1 U12156 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[25] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[153] ), .ZN(n10533)
         );
  AOI22_X1 U12157 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[185] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[313] ), .ZN(n10532) );
  AOI22_X1 U12158 ( .A1(n8111), .A2(\DataPath/RF/bus_sel_savedwin_data[409] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[441] ), .ZN(n10531) );
  AOI22_X1 U12159 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[57] ), 
        .B1(n8353), .B2(\DataPath/RF/bus_sel_savedwin_data[281] ), .ZN(n10530)
         );
  NAND4_X1 U12160 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10534) );
  OR2_X1 U12161 ( .A1(n10535), .A2(n10534), .ZN(DRAMRF_DATA_OUT[25]) );
  AOI22_X1 U12162 ( .A1(n8344), .A2(\DataPath/RF/bus_sel_savedwin_data[506] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[250] ), .ZN(n10539) );
  AOI22_X1 U12163 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[218] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[378] ), .ZN(n10538)
         );
  AOI22_X1 U12164 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[474] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[346] ), .ZN(n10537)
         );
  AOI22_X1 U12165 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[90] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[122] ), .ZN(n10536) );
  NAND4_X1 U12166 ( .A1(n10539), .A2(n10538), .A3(n10537), .A4(n10536), .ZN(
        n10545) );
  AOI22_X1 U12167 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[58] ), 
        .B1(n10678), .B2(\DataPath/RF/bus_sel_savedwin_data[26] ), .ZN(n10543)
         );
  AOI22_X1 U12168 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[186] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[314] ), .ZN(n10542) );
  AOI22_X1 U12169 ( .A1(n8357), .A2(\DataPath/RF/bus_sel_savedwin_data[154] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[442] ), .ZN(n10541)
         );
  AOI22_X1 U12170 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[410] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[282] ), .ZN(n10540)
         );
  NAND4_X1 U12171 ( .A1(n10543), .A2(n10542), .A3(n10541), .A4(n10540), .ZN(
        n10544) );
  OR2_X1 U12172 ( .A1(n10545), .A2(n10544), .ZN(DRAMRF_DATA_OUT[26]) );
  AOI22_X1 U12173 ( .A1(n8344), .A2(\DataPath/RF/bus_sel_savedwin_data[507] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[251] ), .ZN(n10549)
         );
  AOI22_X1 U12174 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[91] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[347] ), .ZN(n10548)
         );
  AOI22_X1 U12175 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[219] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[379] ), .ZN(n10547)
         );
  AOI22_X1 U12176 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[475] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[123] ), .ZN(n10546) );
  NAND4_X1 U12177 ( .A1(n10549), .A2(n10548), .A3(n10547), .A4(n10546), .ZN(
        n10555) );
  AOI22_X1 U12178 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[27] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[315] ), .ZN(n10553)
         );
  AOI22_X1 U12179 ( .A1(n10684), .A2(\DataPath/RF/bus_sel_savedwin_data[411] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[283] ), .ZN(n10552)
         );
  AOI22_X1 U12180 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[187] ), 
        .B1(n10680), .B2(\DataPath/RF/bus_sel_savedwin_data[155] ), .ZN(n10551) );
  AOI22_X1 U12181 ( .A1(n8348), .A2(\DataPath/RF/bus_sel_savedwin_data[59] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[443] ), .ZN(n10550)
         );
  NAND4_X1 U12182 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n10550), .ZN(
        n10554) );
  OR2_X1 U12183 ( .A1(n10555), .A2(n10554), .ZN(DRAMRF_DATA_OUT[27]) );
  AOI22_X1 U12184 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[348] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[380] ), .ZN(n10559)
         );
  AOI22_X1 U12185 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[476] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[124] ), .ZN(n10558)
         );
  AOI22_X1 U12186 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[220] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[508] ), .ZN(n10557)
         );
  AOI22_X1 U12187 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[92] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[252] ), .ZN(n10556)
         );
  NAND4_X1 U12188 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10565) );
  AOI22_X1 U12189 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[188] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[284] ), .ZN(n10563)
         );
  AOI22_X1 U12190 ( .A1(n10680), .A2(\DataPath/RF/bus_sel_savedwin_data[156] ), 
        .B1(n8358), .B2(\DataPath/RF/bus_sel_savedwin_data[444] ), .ZN(n10562)
         );
  AOI22_X1 U12191 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[28] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[316] ), .ZN(n10561)
         );
  AOI22_X1 U12192 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[60] ), 
        .B1(n10684), .B2(\DataPath/RF/bus_sel_savedwin_data[412] ), .ZN(n10560) );
  NAND4_X1 U12193 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10564) );
  OR2_X1 U12194 ( .A1(n10565), .A2(n10564), .ZN(DRAMRF_DATA_OUT[28]) );
  AOI22_X1 U12195 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[221] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[349] ), .ZN(n10569)
         );
  AOI22_X1 U12196 ( .A1(n8344), .A2(\DataPath/RF/bus_sel_savedwin_data[509] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[125] ), .ZN(n10568)
         );
  AOI22_X1 U12197 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[93] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[253] ), .ZN(n10567)
         );
  AOI22_X1 U12198 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[477] ), 
        .B1(n8342), .B2(\DataPath/RF/bus_sel_savedwin_data[381] ), .ZN(n10566)
         );
  NAND4_X1 U12199 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10575) );
  AOI22_X1 U12200 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[61] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[317] ), .ZN(n10573)
         );
  AOI22_X1 U12201 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[189] ), 
        .B1(n10684), .B2(\DataPath/RF/bus_sel_savedwin_data[413] ), .ZN(n10572) );
  AOI22_X1 U12202 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[29] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[445] ), .ZN(n10571)
         );
  AOI22_X1 U12203 ( .A1(n10680), .A2(\DataPath/RF/bus_sel_savedwin_data[157] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[285] ), .ZN(n10570)
         );
  NAND4_X1 U12204 ( .A1(n10573), .A2(n10572), .A3(n10571), .A4(n10570), .ZN(
        n10574) );
  OR2_X1 U12205 ( .A1(n10575), .A2(n10574), .ZN(DRAMRF_DATA_OUT[29]) );
  AOI22_X1 U12206 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[450] ), 
        .B1(n8112), .B2(\DataPath/RF/bus_sel_savedwin_data[322] ), .ZN(n10579)
         );
  AOI22_X1 U12207 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[66] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[482] ), .ZN(n10578)
         );
  AOI22_X1 U12208 ( .A1(n10667), .A2(\DataPath/RF/bus_sel_savedwin_data[354] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[226] ), .ZN(n10577) );
  AOI22_X1 U12209 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[194] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[98] ), .ZN(n10576)
         );
  NAND4_X1 U12210 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10585) );
  AOI22_X1 U12211 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[2] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[258] ), .ZN(n10583)
         );
  AOI22_X1 U12212 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[34] ), 
        .B1(n10679), .B2(\DataPath/RF/bus_sel_savedwin_data[162] ), .ZN(n10582) );
  AOI22_X1 U12213 ( .A1(n10684), .A2(\DataPath/RF/bus_sel_savedwin_data[386] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[418] ), .ZN(n10581)
         );
  AOI22_X1 U12214 ( .A1(n10680), .A2(\DataPath/RF/bus_sel_savedwin_data[130] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[290] ), .ZN(n10580) );
  NAND4_X1 U12215 ( .A1(n10583), .A2(n10582), .A3(n10581), .A4(n10580), .ZN(
        n10584) );
  OR2_X1 U12216 ( .A1(n10585), .A2(n10584), .ZN(DRAMRF_DATA_OUT[2]) );
  AOI22_X1 U12217 ( .A1(n10667), .A2(\DataPath/RF/bus_sel_savedwin_data[382] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[254] ), .ZN(n10589)
         );
  AOI22_X1 U12218 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[94] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[350] ), .ZN(n10588) );
  AOI22_X1 U12219 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[222] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[478] ), .ZN(n10587)
         );
  AOI22_X1 U12220 ( .A1(n10672), .A2(\DataPath/RF/bus_sel_savedwin_data[510] ), 
        .B1(n8345), .B2(\DataPath/RF/bus_sel_savedwin_data[126] ), .ZN(n10586)
         );
  NAND4_X1 U12221 ( .A1(n10589), .A2(n10588), .A3(n10587), .A4(n10586), .ZN(
        n10595) );
  AOI22_X1 U12222 ( .A1(n10684), .A2(\DataPath/RF/bus_sel_savedwin_data[414] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[446] ), .ZN(n10593)
         );
  AOI22_X1 U12223 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[62] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[286] ), .ZN(n10592)
         );
  AOI22_X1 U12224 ( .A1(n10680), .A2(\DataPath/RF/bus_sel_savedwin_data[158] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[318] ), .ZN(n10591)
         );
  AOI22_X1 U12225 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[190] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[30] ), .ZN(n10590)
         );
  NAND4_X1 U12226 ( .A1(n10593), .A2(n10592), .A3(n10591), .A4(n10590), .ZN(
        n10594) );
  OR2_X1 U12227 ( .A1(n10595), .A2(n10594), .ZN(DRAMRF_DATA_OUT[30]) );
  AOI22_X1 U12228 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[95] ), 
        .B1(n10667), .B2(\DataPath/RF/bus_sel_savedwin_data[383] ), .ZN(n10599) );
  AOI22_X1 U12229 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[479] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[255] ), .ZN(n10598)
         );
  AOI22_X1 U12230 ( .A1(n8110), .A2(\DataPath/RF/bus_sel_savedwin_data[351] ), 
        .B1(n8344), .B2(\DataPath/RF/bus_sel_savedwin_data[511] ), .ZN(n10597)
         );
  AOI22_X1 U12231 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[223] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[127] ), .ZN(n10596)
         );
  NAND4_X1 U12232 ( .A1(n10599), .A2(n10598), .A3(n10597), .A4(n10596), .ZN(
        n10605) );
  AOI22_X1 U12233 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[31] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[287] ), .ZN(n10603)
         );
  AOI22_X1 U12234 ( .A1(n10684), .A2(\DataPath/RF/bus_sel_savedwin_data[415] ), 
        .B1(n8113), .B2(\DataPath/RF/bus_sel_savedwin_data[447] ), .ZN(n10602)
         );
  AOI22_X1 U12235 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[191] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[319] ), .ZN(n10601)
         );
  AOI22_X1 U12236 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[63] ), 
        .B1(n10680), .B2(\DataPath/RF/bus_sel_savedwin_data[159] ), .ZN(n10600) );
  NAND4_X1 U12237 ( .A1(n10603), .A2(n10602), .A3(n10601), .A4(n10600), .ZN(
        n10604) );
  OR2_X1 U12238 ( .A1(n10605), .A2(n10604), .ZN(DRAMRF_DATA_OUT[31]) );
  AOI22_X1 U12239 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[195] ), 
        .B1(n10667), .B2(\DataPath/RF/bus_sel_savedwin_data[355] ), .ZN(n10609) );
  AOI22_X1 U12240 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[67] ), 
        .B1(n10672), .B2(\DataPath/RF/bus_sel_savedwin_data[483] ), .ZN(n10608) );
  AOI22_X1 U12241 ( .A1(n8112), .A2(\DataPath/RF/bus_sel_savedwin_data[323] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[99] ), .ZN(n10607)
         );
  AOI22_X1 U12242 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[451] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[227] ), .ZN(n10606)
         );
  NAND4_X1 U12243 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10615) );
  AOI22_X1 U12244 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[35] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[3] ), .ZN(n10613)
         );
  AOI22_X1 U12245 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[131] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[291] ), .ZN(n10612)
         );
  AOI22_X1 U12246 ( .A1(n8350), .A2(\DataPath/RF/bus_sel_savedwin_data[163] ), 
        .B1(n8111), .B2(\DataPath/RF/bus_sel_savedwin_data[387] ), .ZN(n10611)
         );
  AOI22_X1 U12247 ( .A1(n8358), .A2(\DataPath/RF/bus_sel_savedwin_data[419] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[259] ), .ZN(n10610)
         );
  NAND4_X1 U12248 ( .A1(n10613), .A2(n10612), .A3(n10611), .A4(n10610), .ZN(
        n10614) );
  OR2_X1 U12249 ( .A1(n10615), .A2(n10614), .ZN(DRAMRF_DATA_OUT[3]) );
  AOI22_X1 U12250 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[196] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[324] ), .ZN(n10619) );
  AOI22_X1 U12251 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[68] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[452] ), .ZN(n10618)
         );
  AOI22_X1 U12252 ( .A1(n10672), .A2(\DataPath/RF/bus_sel_savedwin_data[484] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[100] ), .ZN(n10617)
         );
  AOI22_X1 U12253 ( .A1(n10667), .A2(\DataPath/RF/bus_sel_savedwin_data[356] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[228] ), .ZN(n10616) );
  NAND4_X1 U12254 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10625) );
  AOI22_X1 U12255 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[36] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[132] ), .ZN(n10623)
         );
  AOI22_X1 U12256 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[388] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[292] ), .ZN(n10622) );
  AOI22_X1 U12257 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[164] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[420] ), .ZN(n10621) );
  AOI22_X1 U12258 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[4] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[260] ), .ZN(n10620)
         );
  NAND4_X1 U12259 ( .A1(n10623), .A2(n10622), .A3(n10621), .A4(n10620), .ZN(
        n10624) );
  OR2_X1 U12260 ( .A1(n10625), .A2(n10624), .ZN(DRAMRF_DATA_OUT[4]) );
  AOI22_X1 U12261 ( .A1(n8340), .A2(\DataPath/RF/bus_sel_savedwin_data[69] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[101] ), .ZN(n10629)
         );
  AOI22_X1 U12262 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[197] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[453] ), .ZN(n10628)
         );
  AOI22_X1 U12263 ( .A1(n8112), .A2(\DataPath/RF/bus_sel_savedwin_data[325] ), 
        .B1(n10672), .B2(\DataPath/RF/bus_sel_savedwin_data[485] ), .ZN(n10627) );
  AOI22_X1 U12264 ( .A1(n8109), .A2(\DataPath/RF/bus_sel_savedwin_data[357] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[229] ), .ZN(n10626) );
  NAND4_X1 U12265 ( .A1(n10629), .A2(n10628), .A3(n10627), .A4(n10626), .ZN(
        n10635) );
  AOI22_X1 U12266 ( .A1(n8349), .A2(\DataPath/RF/bus_sel_savedwin_data[37] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[293] ), .ZN(n10633) );
  AOI22_X1 U12267 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[389] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[133] ), .ZN(n10632)
         );
  AOI22_X1 U12268 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[5] ), 
        .B1(n8354), .B2(\DataPath/RF/bus_sel_savedwin_data[261] ), .ZN(n10631)
         );
  AOI22_X1 U12269 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[165] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[421] ), .ZN(n10630) );
  NAND4_X1 U12270 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10634) );
  OR2_X1 U12271 ( .A1(n10635), .A2(n10634), .ZN(DRAMRF_DATA_OUT[5]) );
  AOI22_X1 U12272 ( .A1(n8341), .A2(\DataPath/RF/bus_sel_savedwin_data[454] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[326] ), .ZN(n10639) );
  AOI22_X1 U12273 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[486] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[230] ), .ZN(n10638)
         );
  AOI22_X1 U12274 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[70] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[102] ), .ZN(n10637)
         );
  AOI22_X1 U12275 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[198] ), 
        .B1(n10667), .B2(\DataPath/RF/bus_sel_savedwin_data[358] ), .ZN(n10636) );
  NAND4_X1 U12276 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10645) );
  AOI22_X1 U12277 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[166] ), 
        .B1(n8352), .B2(\DataPath/RF/bus_sel_savedwin_data[6] ), .ZN(n10643)
         );
  AOI22_X1 U12278 ( .A1(n8356), .A2(\DataPath/RF/bus_sel_savedwin_data[134] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[294] ), .ZN(n10642)
         );
  AOI22_X1 U12279 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[38] ), 
        .B1(n10682), .B2(\DataPath/RF/bus_sel_savedwin_data[422] ), .ZN(n10641) );
  AOI22_X1 U12280 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[390] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[262] ), .ZN(n10640) );
  NAND4_X1 U12281 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10644) );
  OR2_X1 U12282 ( .A1(n10645), .A2(n10644), .ZN(DRAMRF_DATA_OUT[6]) );
  AOI22_X1 U12283 ( .A1(n8343), .A2(\DataPath/RF/bus_sel_savedwin_data[487] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[231] ), .ZN(n10649) );
  AOI22_X1 U12284 ( .A1(n10670), .A2(\DataPath/RF/bus_sel_savedwin_data[455] ), 
        .B1(n10667), .B2(\DataPath/RF/bus_sel_savedwin_data[359] ), .ZN(n10648) );
  AOI22_X1 U12285 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[71] ), 
        .B1(n8346), .B2(\DataPath/RF/bus_sel_savedwin_data[103] ), .ZN(n10647)
         );
  AOI22_X1 U12286 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[199] ), 
        .B1(n10673), .B2(\DataPath/RF/bus_sel_savedwin_data[327] ), .ZN(n10646) );
  NAND4_X1 U12287 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10655) );
  AOI22_X1 U12288 ( .A1(n8352), .A2(\DataPath/RF/bus_sel_savedwin_data[7] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[135] ), .ZN(n10653)
         );
  AOI22_X1 U12289 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[167] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[295] ), .ZN(n10652) );
  AOI22_X1 U12290 ( .A1(n8358), .A2(\DataPath/RF/bus_sel_savedwin_data[423] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[263] ), .ZN(n10651) );
  AOI22_X1 U12291 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[39] ), 
        .B1(n8111), .B2(\DataPath/RF/bus_sel_savedwin_data[391] ), .ZN(n10650)
         );
  NAND4_X1 U12292 ( .A1(n10653), .A2(n10652), .A3(n10651), .A4(n10650), .ZN(
        n10654) );
  OR2_X1 U12293 ( .A1(n10655), .A2(n10654), .ZN(DRAMRF_DATA_OUT[7]) );
  AOI22_X1 U12294 ( .A1(n8342), .A2(\DataPath/RF/bus_sel_savedwin_data[360] ), 
        .B1(n8347), .B2(\DataPath/RF/bus_sel_savedwin_data[232] ), .ZN(n10659)
         );
  AOI22_X1 U12295 ( .A1(n8112), .A2(\DataPath/RF/bus_sel_savedwin_data[328] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[104] ), .ZN(n10658) );
  AOI22_X1 U12296 ( .A1(n8339), .A2(\DataPath/RF/bus_sel_savedwin_data[200] ), 
        .B1(n10672), .B2(\DataPath/RF/bus_sel_savedwin_data[488] ), .ZN(n10657) );
  AOI22_X1 U12297 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[72] ), 
        .B1(n10670), .B2(\DataPath/RF/bus_sel_savedwin_data[456] ), .ZN(n10656) );
  NAND4_X1 U12298 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10665) );
  AOI22_X1 U12299 ( .A1(n10678), .A2(\DataPath/RF/bus_sel_savedwin_data[8] ), 
        .B1(n8357), .B2(\DataPath/RF/bus_sel_savedwin_data[136] ), .ZN(n10663)
         );
  AOI22_X1 U12300 ( .A1(n8358), .A2(\DataPath/RF/bus_sel_savedwin_data[424] ), 
        .B1(n8355), .B2(\DataPath/RF/bus_sel_savedwin_data[296] ), .ZN(n10662)
         );
  AOI22_X1 U12301 ( .A1(n8351), .A2(\DataPath/RF/bus_sel_savedwin_data[168] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[264] ), .ZN(n10661) );
  AOI22_X1 U12302 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[40] ), 
        .B1(n8111), .B2(\DataPath/RF/bus_sel_savedwin_data[392] ), .ZN(n10660)
         );
  NAND4_X1 U12303 ( .A1(n10663), .A2(n10662), .A3(n10661), .A4(n10660), .ZN(
        n10664) );
  OR2_X1 U12304 ( .A1(n10665), .A2(n10664), .ZN(DRAMRF_DATA_OUT[8]) );
  AOI22_X1 U12305 ( .A1(n8342), .A2(\DataPath/RF/bus_sel_savedwin_data[361] ), 
        .B1(n10666), .B2(\DataPath/RF/bus_sel_savedwin_data[233] ), .ZN(n10677) );
  AOI22_X1 U12306 ( .A1(n10669), .A2(\DataPath/RF/bus_sel_savedwin_data[201] ), 
        .B1(n10668), .B2(\DataPath/RF/bus_sel_savedwin_data[105] ), .ZN(n10676) );
  AOI22_X1 U12307 ( .A1(n8108), .A2(\DataPath/RF/bus_sel_savedwin_data[73] ), 
        .B1(n8341), .B2(\DataPath/RF/bus_sel_savedwin_data[457] ), .ZN(n10675)
         );
  AOI22_X1 U12308 ( .A1(n8112), .A2(\DataPath/RF/bus_sel_savedwin_data[329] ), 
        .B1(n10672), .B2(\DataPath/RF/bus_sel_savedwin_data[489] ), .ZN(n10674) );
  NAND4_X1 U12309 ( .A1(n10677), .A2(n10676), .A3(n10675), .A4(n10674), .ZN(
        n10690) );
  AOI22_X1 U12310 ( .A1(n10679), .A2(\DataPath/RF/bus_sel_savedwin_data[169] ), 
        .B1(n10678), .B2(\DataPath/RF/bus_sel_savedwin_data[9] ), .ZN(n10688)
         );
  AOI22_X1 U12311 ( .A1(n8114), .A2(\DataPath/RF/bus_sel_savedwin_data[41] ), 
        .B1(n10680), .B2(\DataPath/RF/bus_sel_savedwin_data[137] ), .ZN(n10687) );
  AOI22_X1 U12312 ( .A1(n8113), .A2(\DataPath/RF/bus_sel_savedwin_data[425] ), 
        .B1(n10681), .B2(\DataPath/RF/bus_sel_savedwin_data[297] ), .ZN(n10686) );
  AOI22_X1 U12313 ( .A1(n8089), .A2(\DataPath/RF/bus_sel_savedwin_data[393] ), 
        .B1(n10683), .B2(\DataPath/RF/bus_sel_savedwin_data[265] ), .ZN(n10685) );
  NAND4_X1 U12314 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10689) );
  OR2_X1 U12315 ( .A1(n10690), .A2(n10689), .ZN(DRAMRF_DATA_OUT[9]) );
  NOR2_X1 U12316 ( .A1(n11662), .A2(n8172), .ZN(n11650) );
  INV_X1 U12317 ( .A(n11650), .ZN(n11649) );
  NAND2_X1 U12318 ( .A1(n11841), .A2(n11649), .ZN(n11845) );
  INV_X1 U12319 ( .A(n11845), .ZN(DRAMRF_READNOTWRITE) );
  NOR2_X1 U12320 ( .A1(n507), .A2(n381), .ZN(DRAM_ADDRESS[0]) );
  AOI21_X1 U12321 ( .B1(n381), .B2(n380), .A(n508), .ZN(DRAM_ADDRESS[1]) );
  AOI221_X1 U12322 ( .B1(n381), .B2(n8168), .C1(n381), .C2(n380), .A(n11616), 
        .ZN(n10693) );
  NOR4_X1 U12323 ( .A1(n507), .A2(n11616), .A3(n8168), .A4(n10703), .ZN(n10691) );
  AOI22_X1 U12324 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[16]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[16] ), .B2(n11616), .ZN(n10735) );
  NAND2_X1 U12325 ( .A1(n507), .A2(n10693), .ZN(n10694) );
  MUX2_X1 U12326 ( .A(DRAM_DATA_IN[8]), .B(\DataPath/i_REG_ME_DATA_DATAMEM[8] ), .S(n11616), .Z(n10758) );
  AOI22_X1 U12327 ( .A1(n10736), .A2(n10758), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[0] ), .B2(n11616), .ZN(n10696) );
  NAND2_X1 U12328 ( .A1(n10800), .A2(n8168), .ZN(n10692) );
  MUX2_X1 U12329 ( .A(DRAM_DATA_IN[24]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[24] ), .S(n11616), .Z(n10789) );
  AOI22_X1 U12330 ( .A1(n10738), .A2(DRAM_DATA_IN[0]), .B1(n10737), .B2(n10789), .ZN(n10695) );
  OAI211_X1 U12331 ( .C1(n10741), .C2(n10735), .A(n10696), .B(n10695), .ZN(
        DRAM_DATA_OUT[0]) );
  AOI22_X1 U12332 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[23]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[23] ), .B2(n11616), .ZN(n10757) );
  MUX2_X1 U12333 ( .A(DRAM_DATA_IN[15]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[15] ), .S(n11616), .Z(n10730) );
  AOI22_X1 U12334 ( .A1(n10736), .A2(n10730), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[7] ), .B2(n11616), .ZN(n10698) );
  MUX2_X1 U12335 ( .A(DRAM_DATA_IN[31]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[31] ), .S(n11616), .Z(n10782) );
  AOI22_X1 U12336 ( .A1(n10738), .A2(DRAM_DATA_IN[7]), .B1(n10737), .B2(n10782), .ZN(n10697) );
  OAI211_X1 U12337 ( .C1(n10757), .C2(n10741), .A(n10698), .B(n10697), .ZN(
        DRAM_DATA_OUT[7]) );
  AOI22_X1 U12338 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[18]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[18] ), .B2(n11616), .ZN(n10745) );
  MUX2_X1 U12339 ( .A(DRAM_DATA_IN[26]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[26] ), .S(n11616), .Z(n10764) );
  AOI22_X1 U12340 ( .A1(n10737), .A2(n10764), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[2] ), .B2(n11616), .ZN(n10700) );
  MUX2_X1 U12341 ( .A(DRAM_DATA_IN[10]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[10] ), .S(n11616), .Z(n10701) );
  AOI22_X1 U12342 ( .A1(n10738), .A2(DRAM_DATA_IN[2]), .B1(n10736), .B2(n10701), .ZN(n10699) );
  OAI211_X1 U12343 ( .C1(n10741), .C2(n10745), .A(n10700), .B(n10699), .ZN(
        DRAM_DATA_OUT[2]) );
  NAND2_X1 U12344 ( .A1(n10795), .A2(n10701), .ZN(n10766) );
  INV_X1 U12345 ( .A(n10766), .ZN(n10702) );
  AOI21_X1 U12346 ( .B1(n10797), .B2(n10764), .A(n10702), .ZN(n10705) );
  NAND2_X1 U12347 ( .A1(n10790), .A2(DRAM_DATA_OUT[2]), .ZN(n10704) );
  NAND3_X1 U12348 ( .A1(n10800), .A2(n217), .A3(DRAM_DATA_OUT[7]), .ZN(n10755)
         );
  OAI211_X1 U12349 ( .C1(n10800), .C2(n10705), .A(n10704), .B(n10791), .ZN(
        DRAM_DATA_OUT[10]) );
  AOI22_X1 U12350 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[19]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[19] ), .B2(n11616), .ZN(n10747) );
  MUX2_X1 U12351 ( .A(DRAM_DATA_IN[11]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[11] ), .S(n11616), .Z(n10708) );
  AOI22_X1 U12352 ( .A1(n10736), .A2(n10708), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[3] ), .B2(n11616), .ZN(n10707) );
  MUX2_X1 U12353 ( .A(DRAM_DATA_IN[27]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[27] ), .S(n11616), .Z(n10767) );
  AOI22_X1 U12354 ( .A1(n10738), .A2(DRAM_DATA_IN[3]), .B1(n10737), .B2(n10767), .ZN(n10706) );
  OAI211_X1 U12355 ( .C1(n10741), .C2(n10747), .A(n10707), .B(n10706), .ZN(
        DRAM_DATA_OUT[3]) );
  NAND2_X1 U12356 ( .A1(n10795), .A2(n10708), .ZN(n10769) );
  INV_X1 U12357 ( .A(n10769), .ZN(n10709) );
  AOI21_X1 U12358 ( .B1(n10797), .B2(n10767), .A(n10709), .ZN(n10711) );
  NAND2_X1 U12359 ( .A1(n10790), .A2(DRAM_DATA_OUT[3]), .ZN(n10710) );
  OAI211_X1 U12360 ( .C1(n10800), .C2(n10711), .A(n10710), .B(n10791), .ZN(
        DRAM_DATA_OUT[11]) );
  AOI22_X1 U12361 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[20]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[20] ), .B2(n11616), .ZN(n10749) );
  AOI22_X1 U12362 ( .A1(DRAM_DATA_IN[4]), .A2(n10738), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[4] ), .B2(n11616), .ZN(n10713) );
  MUX2_X1 U12363 ( .A(DRAM_DATA_IN[28]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[28] ), .S(n11616), .Z(n10770) );
  MUX2_X1 U12364 ( .A(DRAM_DATA_IN[12]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[12] ), .S(n11616), .Z(n10714) );
  AOI22_X1 U12365 ( .A1(n10737), .A2(n10770), .B1(n10736), .B2(n10714), .ZN(
        n10712) );
  OAI211_X1 U12366 ( .C1(n10741), .C2(n10749), .A(n10713), .B(n10712), .ZN(
        DRAM_DATA_OUT[4]) );
  NAND2_X1 U12367 ( .A1(n10795), .A2(n10714), .ZN(n10772) );
  INV_X1 U12368 ( .A(n10772), .ZN(n10715) );
  AOI21_X1 U12369 ( .B1(n10797), .B2(n10770), .A(n10715), .ZN(n10717) );
  NAND2_X1 U12370 ( .A1(n10790), .A2(DRAM_DATA_OUT[4]), .ZN(n10716) );
  OAI211_X1 U12371 ( .C1(n10800), .C2(n10717), .A(n10716), .B(n10791), .ZN(
        DRAM_DATA_OUT[12]) );
  AOI22_X1 U12372 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[21]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[21] ), .B2(n11616), .ZN(n10751) );
  AOI22_X1 U12373 ( .A1(DRAM_DATA_IN[5]), .A2(n10738), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[5] ), .B2(n11616), .ZN(n10719) );
  MUX2_X1 U12374 ( .A(DRAM_DATA_IN[29]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[29] ), .S(n11616), .Z(n10773) );
  MUX2_X1 U12375 ( .A(DRAM_DATA_IN[13]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[13] ), .S(n11616), .Z(n10720) );
  AOI22_X1 U12376 ( .A1(n10737), .A2(n10773), .B1(n10736), .B2(n10720), .ZN(
        n10718) );
  OAI211_X1 U12377 ( .C1(n10741), .C2(n10751), .A(n10719), .B(n10718), .ZN(
        DRAM_DATA_OUT[5]) );
  NAND2_X1 U12378 ( .A1(n10795), .A2(n10720), .ZN(n10775) );
  INV_X1 U12379 ( .A(n10775), .ZN(n10721) );
  AOI21_X1 U12380 ( .B1(n10797), .B2(n10773), .A(n10721), .ZN(n10723) );
  NAND2_X1 U12381 ( .A1(n10790), .A2(DRAM_DATA_OUT[5]), .ZN(n10722) );
  OAI211_X1 U12382 ( .C1(n10800), .C2(n10723), .A(n10722), .B(n10791), .ZN(
        DRAM_DATA_OUT[13]) );
  AOI22_X1 U12383 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[22]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[22] ), .B2(n11616), .ZN(n10753) );
  MUX2_X1 U12384 ( .A(DRAM_DATA_IN[14]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[14] ), .S(n11616), .Z(n10726) );
  AOI22_X1 U12385 ( .A1(n10736), .A2(n10726), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[6] ), .B2(n11616), .ZN(n10725) );
  MUX2_X1 U12386 ( .A(DRAM_DATA_IN[30]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[30] ), .S(n11616), .Z(n10776) );
  AOI22_X1 U12387 ( .A1(n10738), .A2(DRAM_DATA_IN[6]), .B1(n10737), .B2(n10776), .ZN(n10724) );
  OAI211_X1 U12388 ( .C1(n10741), .C2(n10753), .A(n10725), .B(n10724), .ZN(
        DRAM_DATA_OUT[6]) );
  NAND2_X1 U12389 ( .A1(n10795), .A2(n10726), .ZN(n10781) );
  INV_X1 U12390 ( .A(n10781), .ZN(n10727) );
  AOI21_X1 U12391 ( .B1(n10797), .B2(n10776), .A(n10727), .ZN(n10729) );
  NAND2_X1 U12392 ( .A1(n10790), .A2(DRAM_DATA_OUT[6]), .ZN(n10728) );
  OAI211_X1 U12393 ( .C1(n10800), .C2(n10729), .A(n10728), .B(n10791), .ZN(
        DRAM_DATA_OUT[14]) );
  AOI22_X1 U12394 ( .A1(n10795), .A2(n10730), .B1(n10782), .B2(n10797), .ZN(
        n10733) );
  OAI211_X1 U12395 ( .C1(n217), .C2(n11616), .A(n10800), .B(DRAM_DATA_OUT[7]), 
        .ZN(n10784) );
  OAI21_X1 U12396 ( .B1(n10800), .B2(n10733), .A(n10784), .ZN(
        DRAM_DATA_OUT[15]) );
  INV_X1 U12397 ( .A(n10790), .ZN(n10731) );
  NAND3_X1 U12398 ( .A1(n11616), .A2(DATA_SIZE[0]), .A3(n381), .ZN(n10780) );
  AOI21_X1 U12399 ( .B1(n381), .B2(n380), .A(n11616), .ZN(n10732) );
  NOR2_X1 U12400 ( .A1(n11616), .A2(n10783), .ZN(n10761) );
  NAND2_X1 U12401 ( .A1(n10754), .A2(DRAM_DATA_OUT[0]), .ZN(n10734) );
  OAI211_X1 U12402 ( .C1(n10735), .C2(n10785), .A(n10779), .B(n10734), .ZN(
        DRAM_DATA_OUT[16]) );
  AOI22_X1 U12403 ( .A1(i_DATAMEM_RM), .A2(DRAM_DATA_IN[17]), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[17] ), .B2(n11616), .ZN(n10743) );
  MUX2_X1 U12404 ( .A(DRAM_DATA_IN[9]), .B(\DataPath/i_REG_ME_DATA_DATAMEM[9] ), .S(n11616), .Z(n10794) );
  AOI22_X1 U12405 ( .A1(n10736), .A2(n10794), .B1(
        \DataPath/i_REG_ME_DATA_DATAMEM[1] ), .B2(n11616), .ZN(n10740) );
  MUX2_X1 U12406 ( .A(DRAM_DATA_IN[25]), .B(
        \DataPath/i_REG_ME_DATA_DATAMEM[25] ), .S(n11616), .Z(n10796) );
  AOI22_X1 U12407 ( .A1(n10738), .A2(DRAM_DATA_IN[1]), .B1(n10737), .B2(n10796), .ZN(n10739) );
  OAI211_X1 U12408 ( .C1(n10741), .C2(n10743), .A(n10740), .B(n10739), .ZN(
        DRAM_DATA_OUT[1]) );
  NAND2_X1 U12409 ( .A1(DRAM_DATA_OUT[1]), .A2(n10754), .ZN(n10742) );
  OAI211_X1 U12410 ( .C1(n10743), .C2(n10785), .A(n10779), .B(n10742), .ZN(
        DRAM_DATA_OUT[17]) );
  NAND2_X1 U12411 ( .A1(n10754), .A2(DRAM_DATA_OUT[2]), .ZN(n10744) );
  OAI211_X1 U12412 ( .C1(n10745), .C2(n10785), .A(n10779), .B(n10744), .ZN(
        DRAM_DATA_OUT[18]) );
  NAND2_X1 U12413 ( .A1(n10754), .A2(DRAM_DATA_OUT[3]), .ZN(n10746) );
  OAI211_X1 U12414 ( .C1(n10747), .C2(n10785), .A(n10779), .B(n10746), .ZN(
        DRAM_DATA_OUT[19]) );
  NAND2_X1 U12415 ( .A1(n10754), .A2(DRAM_DATA_OUT[4]), .ZN(n10748) );
  OAI211_X1 U12416 ( .C1(n10749), .C2(n10785), .A(n10779), .B(n10748), .ZN(
        DRAM_DATA_OUT[20]) );
  NAND2_X1 U12417 ( .A1(n10754), .A2(DRAM_DATA_OUT[5]), .ZN(n10750) );
  OAI211_X1 U12418 ( .C1(n10751), .C2(n10785), .A(n10779), .B(n10750), .ZN(
        DRAM_DATA_OUT[21]) );
  NAND2_X1 U12419 ( .A1(n10754), .A2(DRAM_DATA_OUT[6]), .ZN(n10752) );
  OAI211_X1 U12420 ( .C1(n10753), .C2(n10785), .A(n10779), .B(n10752), .ZN(
        DRAM_DATA_OUT[22]) );
  AOI21_X1 U12421 ( .B1(DRAM_DATA_OUT[7]), .B2(n10754), .A(n10761), .ZN(n10756) );
  OAI211_X1 U12422 ( .C1(n10757), .C2(n10785), .A(n10756), .B(n10755), .ZN(
        DRAM_DATA_OUT[23]) );
  NAND2_X1 U12423 ( .A1(n10795), .A2(n10758), .ZN(n10787) );
  AOI22_X1 U12424 ( .A1(n10790), .A2(DRAM_DATA_OUT[0]), .B1(n10777), .B2(
        n10789), .ZN(n10759) );
  OAI211_X1 U12425 ( .C1(n10787), .C2(n10780), .A(n10779), .B(n10759), .ZN(
        DRAM_DATA_OUT[24]) );
  NAND2_X1 U12426 ( .A1(n10795), .A2(n10794), .ZN(n10763) );
  AOI21_X1 U12427 ( .B1(n10790), .B2(DRAM_DATA_OUT[1]), .A(n10760), .ZN(n10798) );
  AOI21_X1 U12428 ( .B1(n10777), .B2(n10796), .A(n10761), .ZN(n10762) );
  OAI211_X1 U12429 ( .C1(n10780), .C2(n10763), .A(n10798), .B(n10762), .ZN(
        DRAM_DATA_OUT[25]) );
  AOI22_X1 U12430 ( .A1(n10790), .A2(DRAM_DATA_OUT[2]), .B1(n10777), .B2(
        n10764), .ZN(n10765) );
  OAI211_X1 U12431 ( .C1(n10766), .C2(n10780), .A(n10779), .B(n10765), .ZN(
        DRAM_DATA_OUT[26]) );
  AOI22_X1 U12432 ( .A1(n10790), .A2(DRAM_DATA_OUT[3]), .B1(n10777), .B2(
        n10767), .ZN(n10768) );
  OAI211_X1 U12433 ( .C1(n10769), .C2(n10780), .A(n10779), .B(n10768), .ZN(
        DRAM_DATA_OUT[27]) );
  AOI22_X1 U12434 ( .A1(n10790), .A2(DRAM_DATA_OUT[4]), .B1(n10777), .B2(
        n10770), .ZN(n10771) );
  OAI211_X1 U12435 ( .C1(n10772), .C2(n10780), .A(n10779), .B(n10771), .ZN(
        DRAM_DATA_OUT[28]) );
  AOI22_X1 U12436 ( .A1(n10790), .A2(DRAM_DATA_OUT[5]), .B1(n10777), .B2(
        n10773), .ZN(n10774) );
  OAI211_X1 U12437 ( .C1(n10775), .C2(n10780), .A(n10779), .B(n10774), .ZN(
        DRAM_DATA_OUT[29]) );
  AOI22_X1 U12438 ( .A1(n10790), .A2(DRAM_DATA_OUT[6]), .B1(n10777), .B2(
        n10776), .ZN(n10778) );
  OAI211_X1 U12439 ( .C1(n10781), .C2(n10780), .A(n10779), .B(n10778), .ZN(
        DRAM_DATA_OUT[30]) );
  INV_X1 U12440 ( .A(n10782), .ZN(n10786) );
  OAI211_X1 U12441 ( .C1(n10786), .C2(n10785), .A(n10784), .B(n10783), .ZN(
        DRAM_DATA_OUT[31]) );
  INV_X1 U12442 ( .A(n10787), .ZN(n10788) );
  AOI21_X1 U12443 ( .B1(n10797), .B2(n10789), .A(n10788), .ZN(n10793) );
  NAND2_X1 U12444 ( .A1(n10790), .A2(DRAM_DATA_OUT[0]), .ZN(n10792) );
  OAI211_X1 U12445 ( .C1(n10800), .C2(n10793), .A(n10792), .B(n10791), .ZN(
        DRAM_DATA_OUT[8]) );
  AOI22_X1 U12446 ( .A1(n10797), .A2(n10796), .B1(n10795), .B2(n10794), .ZN(
        n10799) );
  OAI21_X1 U12447 ( .B1(n10800), .B2(n10799), .A(n10798), .ZN(DRAM_DATA_OUT[9]) );
  OAI211_X1 U12448 ( .C1(n10915), .C2(n8212), .A(n8457), .B(n11661), .ZN(
        \DataPath/RF/POP_ADDRGEN/N46 ) );
  AOI22_X1 U12449 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[0] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[1] ), .ZN(n10919)
         );
  NOR2_X1 U12450 ( .A1(RST), .A2(n10919), .ZN(\DataPath/RF/POP_ADDRGEN/N47 )
         );
  AOI22_X1 U12451 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[1] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[2] ), .ZN(n10924)
         );
  NOR2_X1 U12452 ( .A1(RST), .A2(n10924), .ZN(\DataPath/RF/POP_ADDRGEN/N48 )
         );
  AOI22_X1 U12453 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[2] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[3] ), .ZN(n10928)
         );
  NOR2_X1 U12454 ( .A1(RST), .A2(n10928), .ZN(\DataPath/RF/POP_ADDRGEN/N49 )
         );
  AOI22_X1 U12455 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[3] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[4] ), .ZN(n10933)
         );
  NOR2_X1 U12456 ( .A1(RST), .A2(n10933), .ZN(\DataPath/RF/POP_ADDRGEN/N50 )
         );
  AOI22_X1 U12457 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[4] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[5] ), .ZN(n10827)
         );
  NOR2_X1 U12458 ( .A1(RST), .A2(n10827), .ZN(\DataPath/RF/POP_ADDRGEN/N51 )
         );
  AOI22_X1 U12459 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[5] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[6] ), .ZN(n10842)
         );
  NOR2_X1 U12460 ( .A1(RST), .A2(n10842), .ZN(\DataPath/RF/POP_ADDRGEN/N52 )
         );
  AOI22_X1 U12461 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[6] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[7] ), .ZN(n10865)
         );
  NOR2_X1 U12462 ( .A1(RST), .A2(n10865), .ZN(\DataPath/RF/POP_ADDRGEN/N53 )
         );
  AOI22_X1 U12463 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[7] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[8] ), .ZN(n10869)
         );
  NOR2_X1 U12464 ( .A1(RST), .A2(n10869), .ZN(\DataPath/RF/POP_ADDRGEN/N54 )
         );
  AOI22_X1 U12465 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[8] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[9] ), .ZN(n10875)
         );
  NOR2_X1 U12466 ( .A1(RST), .A2(n10875), .ZN(\DataPath/RF/POP_ADDRGEN/N55 )
         );
  AOI22_X1 U12467 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[9] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[10] ), .ZN(n10881)
         );
  NOR2_X1 U12468 ( .A1(RST), .A2(n10881), .ZN(\DataPath/RF/POP_ADDRGEN/N56 )
         );
  AOI22_X1 U12469 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[10] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[11] ), .ZN(n10887)
         );
  NOR2_X1 U12470 ( .A1(RST), .A2(n10887), .ZN(\DataPath/RF/POP_ADDRGEN/N57 )
         );
  AOI22_X1 U12471 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[11] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[12] ), .ZN(n10892)
         );
  NOR2_X1 U12472 ( .A1(RST), .A2(n10892), .ZN(\DataPath/RF/POP_ADDRGEN/N58 )
         );
  AOI22_X1 U12473 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[12] ), 
        .B1(n10802), .B2(\DataPath/RF/POP_ADDRGEN/curr_addr[13] ), .ZN(n10898)
         );
  NOR2_X1 U12474 ( .A1(RST), .A2(n10898), .ZN(\DataPath/RF/POP_ADDRGEN/N59 )
         );
  AOI22_X1 U12475 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[13] ), 
        .B1(\DataPath/RF/POP_ADDRGEN/curr_addr[14] ), .B2(n10802), .ZN(n10903)
         );
  NOR2_X1 U12476 ( .A1(RST), .A2(n10903), .ZN(\DataPath/RF/POP_ADDRGEN/N60 )
         );
  NAND2_X1 U12477 ( .A1(n10915), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[14] ), 
        .ZN(n10908) );
  AOI221_X1 U12478 ( .B1(n11665), .B2(n10908), .C1(n8172), .C2(n10908), .A(RST), .ZN(\DataPath/RF/POP_ADDRGEN/N61 ) );
  NOR2_X1 U12479 ( .A1(RST), .A2(n11646), .ZN(n11848) );
  OAI21_X1 U12480 ( .B1(n8338), .B2(n8210), .A(n11848), .ZN(
        \DataPath/RF/PUSH_ADDRGEN/N46 ) );
  AOI22_X1 U12481 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[0] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[1] ), .ZN(n10803)
         );
  NOR2_X1 U12482 ( .A1(RST), .A2(n10803), .ZN(\DataPath/RF/PUSH_ADDRGEN/N47 )
         );
  AOI22_X1 U12483 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[1] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[2] ), .ZN(n10804)
         );
  NOR2_X1 U12484 ( .A1(RST), .A2(n10804), .ZN(\DataPath/RF/PUSH_ADDRGEN/N48 )
         );
  AOI22_X1 U12485 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[2] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[3] ), .ZN(n10805)
         );
  NOR2_X1 U12486 ( .A1(RST), .A2(n10805), .ZN(\DataPath/RF/PUSH_ADDRGEN/N49 )
         );
  AOI22_X1 U12487 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[3] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[4] ), .ZN(n10806)
         );
  NOR2_X1 U12488 ( .A1(RST), .A2(n10806), .ZN(\DataPath/RF/PUSH_ADDRGEN/N50 )
         );
  AOI22_X1 U12489 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[4] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[5] ), .ZN(n10807)
         );
  NOR2_X1 U12490 ( .A1(RST), .A2(n10807), .ZN(\DataPath/RF/PUSH_ADDRGEN/N51 )
         );
  AOI22_X1 U12491 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[5] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[6] ), .ZN(n10808)
         );
  NOR2_X1 U12492 ( .A1(RST), .A2(n10808), .ZN(\DataPath/RF/PUSH_ADDRGEN/N52 )
         );
  AOI22_X1 U12493 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[6] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[7] ), .ZN(n10809)
         );
  NOR2_X1 U12494 ( .A1(RST), .A2(n10809), .ZN(\DataPath/RF/PUSH_ADDRGEN/N53 )
         );
  AOI22_X1 U12495 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[7] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[8] ), .ZN(n10810)
         );
  NOR2_X1 U12496 ( .A1(RST), .A2(n10810), .ZN(\DataPath/RF/PUSH_ADDRGEN/N54 )
         );
  AOI22_X1 U12497 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[8] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[9] ), .ZN(n10811)
         );
  NOR2_X1 U12498 ( .A1(RST), .A2(n10811), .ZN(\DataPath/RF/PUSH_ADDRGEN/N55 )
         );
  AOI22_X1 U12499 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[9] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[10] ), .ZN(n10812) );
  NOR2_X1 U12500 ( .A1(RST), .A2(n10812), .ZN(\DataPath/RF/PUSH_ADDRGEN/N56 )
         );
  AOI22_X1 U12501 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[10] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[11] ), .ZN(n10813) );
  NOR2_X1 U12502 ( .A1(RST), .A2(n10813), .ZN(\DataPath/RF/PUSH_ADDRGEN/N57 )
         );
  AOI22_X1 U12503 ( .A1(n8338), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[11] ), 
        .B1(n10815), .B2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[12] ), .ZN(n10814) );
  NOR2_X1 U12504 ( .A1(RST), .A2(n10814), .ZN(\DataPath/RF/PUSH_ADDRGEN/N58 )
         );
  AOI22_X1 U12505 ( .A1(n10816), .A2(\DataPath/RF/PUSH_ADDRGEN/curr_addr[12] ), 
        .B1(\DataPath/RF/PUSH_ADDRGEN/curr_addr[13] ), .B2(n10815), .ZN(n10817) );
  NOR2_X1 U12506 ( .A1(RST), .A2(n10817), .ZN(\DataPath/RF/PUSH_ADDRGEN/N59 )
         );
  AOI221_X1 U12507 ( .B1(n8104), .B2(n10819), .C1(n10818), .C2(n10819), .A(RST), .ZN(\DataPath/RF/PUSH_ADDRGEN/N60 ) );
  AND2_X1 U12508 ( .A1(n11848), .A2(n10820), .ZN(
        \DataPath/RF/PUSH_ADDRGEN/N61 ) );
  AOI22_X1 U12509 ( .A1(n10294), .A2(n8129), .B1(\DP_OP_1091J1_126_6973/n72 ), 
        .B2(n11649), .ZN(n10825) );
  NOR2_X1 U12510 ( .A1(n8054), .A2(\DP_OP_1091J1_126_6973/n72 ), .ZN(n10823)
         );
  AOI22_X1 U12511 ( .A1(n10823), .A2(n10822), .B1(n10293), .B2(n9270), .ZN(
        n10824) );
  AOI21_X1 U12512 ( .B1(n10825), .B2(n10824), .A(RST), .ZN(
        \DataPath/WRF_CUhw/N145 ) );
  MUX2_X1 U12513 ( .A(DRAMRF_DATA_IN[18]), .B(
        \DataPath/WRF_CUhw/curr_data[18] ), .S(n11840), .Z(n11538) );
  MUX2_X1 U12514 ( .A(\DataPath/i_REG_MEM_ALUOUT[18] ), .B(
        \DataPath/i_REG_LDSTR_OUT[18] ), .S(i_S3), .Z(n10826) );
  OAI22_X1 U12515 ( .A1(n8437), .A2(n11290), .B1(n11497), .B2(n8183), .ZN(
        n11787) );
  NAND2_X1 U12516 ( .A1(n10932), .A2(n11472), .ZN(n11322) );
  INV_X1 U12517 ( .A(n10827), .ZN(n10828) );
  AOI22_X1 U12518 ( .A1(n11746), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2386] ), .ZN(n6127) );
  MUX2_X1 U12519 ( .A(DRAMRF_DATA_IN[19]), .B(
        \DataPath/WRF_CUhw/curr_data[19] ), .S(n11840), .Z(n11539) );
  MUX2_X1 U12520 ( .A(\DataPath/i_REG_MEM_ALUOUT[19] ), .B(
        \DataPath/i_REG_LDSTR_OUT[19] ), .S(i_S3), .Z(n10829) );
  OAI22_X1 U12521 ( .A1(n8437), .A2(n11291), .B1(n11498), .B2(n8183), .ZN(
        n11788) );
  AOI22_X1 U12522 ( .A1(n11747), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2387] ), .ZN(n6126) );
  MUX2_X1 U12523 ( .A(DRAMRF_DATA_IN[20]), .B(
        \DataPath/WRF_CUhw/curr_data[20] ), .S(n11840), .Z(n11540) );
  MUX2_X1 U12524 ( .A(\DataPath/i_REG_MEM_ALUOUT[20] ), .B(
        \DataPath/i_REG_LDSTR_OUT[20] ), .S(i_S3), .Z(n10830) );
  OAI22_X1 U12525 ( .A1(n8436), .A2(n11292), .B1(n11499), .B2(n8183), .ZN(
        n11789) );
  AOI22_X1 U12526 ( .A1(n11748), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2388] ), .ZN(n6125) );
  MUX2_X1 U12527 ( .A(DRAMRF_DATA_IN[21]), .B(
        \DataPath/WRF_CUhw/curr_data[21] ), .S(n11840), .Z(n11541) );
  MUX2_X1 U12528 ( .A(\DataPath/i_REG_MEM_ALUOUT[21] ), .B(
        \DataPath/i_REG_LDSTR_OUT[21] ), .S(i_S3), .Z(n10831) );
  OAI22_X1 U12529 ( .A1(n8436), .A2(n11293), .B1(n11500), .B2(n8183), .ZN(
        n11790) );
  AOI22_X1 U12530 ( .A1(n11749), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2389] ), .ZN(n6124) );
  MUX2_X1 U12531 ( .A(DRAMRF_DATA_IN[22]), .B(
        \DataPath/WRF_CUhw/curr_data[22] ), .S(n11840), .Z(n11542) );
  MUX2_X1 U12532 ( .A(\DataPath/i_REG_MEM_ALUOUT[22] ), .B(
        \DataPath/i_REG_LDSTR_OUT[22] ), .S(i_S3), .Z(n10832) );
  OAI22_X1 U12533 ( .A1(n8436), .A2(n11294), .B1(n11501), .B2(n8183), .ZN(
        n11765) );
  AOI22_X1 U12534 ( .A1(n11791), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2390] ), .ZN(n6123) );
  MUX2_X1 U12535 ( .A(DRAMRF_DATA_IN[23]), .B(
        \DataPath/WRF_CUhw/curr_data[23] ), .S(n11840), .Z(n11543) );
  MUX2_X1 U12536 ( .A(\DataPath/i_REG_MEM_ALUOUT[23] ), .B(
        \DataPath/i_REG_LDSTR_OUT[23] ), .S(n8451), .Z(n10833) );
  OAI22_X1 U12537 ( .A1(n8436), .A2(n11295), .B1(n11502), .B2(n8183), .ZN(
        n11792) );
  AOI22_X1 U12538 ( .A1(n11750), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2391] ), .ZN(n6122) );
  MUX2_X1 U12539 ( .A(DRAMRF_DATA_IN[24]), .B(
        \DataPath/WRF_CUhw/curr_data[24] ), .S(n11840), .Z(n11544) );
  MUX2_X1 U12540 ( .A(\DataPath/i_REG_MEM_ALUOUT[24] ), .B(
        \DataPath/i_REG_LDSTR_OUT[24] ), .S(i_S3), .Z(n10834) );
  OAI22_X1 U12541 ( .A1(n8436), .A2(n11296), .B1(n11503), .B2(n8183), .ZN(
        n11766) );
  AOI22_X1 U12542 ( .A1(n11793), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2392] ), .ZN(n6121) );
  MUX2_X1 U12543 ( .A(DRAMRF_DATA_IN[25]), .B(
        \DataPath/WRF_CUhw/curr_data[25] ), .S(n11840), .Z(n11545) );
  MUX2_X1 U12544 ( .A(\DataPath/i_REG_MEM_ALUOUT[25] ), .B(
        \DataPath/i_REG_LDSTR_OUT[25] ), .S(i_S3), .Z(n10835) );
  OAI22_X1 U12545 ( .A1(n8437), .A2(n11297), .B1(n11504), .B2(n8183), .ZN(
        n11767) );
  AOI22_X1 U12546 ( .A1(n11794), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2393] ), .ZN(n6120) );
  MUX2_X1 U12547 ( .A(DRAMRF_DATA_IN[26]), .B(
        \DataPath/WRF_CUhw/curr_data[26] ), .S(n11840), .Z(n11546) );
  MUX2_X1 U12548 ( .A(\DataPath/i_REG_MEM_ALUOUT[26] ), .B(
        \DataPath/i_REG_LDSTR_OUT[26] ), .S(i_S3), .Z(n10836) );
  OAI22_X1 U12549 ( .A1(n8436), .A2(n11298), .B1(n11505), .B2(n8183), .ZN(
        n11795) );
  AOI22_X1 U12550 ( .A1(n11751), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2394] ), .ZN(n6119) );
  MUX2_X1 U12551 ( .A(DRAMRF_DATA_IN[27]), .B(
        \DataPath/WRF_CUhw/curr_data[27] ), .S(n11840), .Z(n11547) );
  MUX2_X1 U12552 ( .A(\DataPath/i_REG_MEM_ALUOUT[27] ), .B(
        \DataPath/i_REG_LDSTR_OUT[27] ), .S(i_S3), .Z(n10837) );
  OAI22_X1 U12553 ( .A1(n8437), .A2(n11299), .B1(n11506), .B2(n8183), .ZN(
        n11768) );
  AOI22_X1 U12554 ( .A1(n11796), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2395] ), .ZN(n6118) );
  MUX2_X1 U12555 ( .A(DRAMRF_DATA_IN[28]), .B(
        \DataPath/WRF_CUhw/curr_data[28] ), .S(n11840), .Z(n11548) );
  MUX2_X1 U12556 ( .A(\DataPath/i_REG_MEM_ALUOUT[28] ), .B(
        \DataPath/i_REG_LDSTR_OUT[28] ), .S(i_S3), .Z(n10838) );
  OAI22_X1 U12557 ( .A1(n8437), .A2(n11300), .B1(n11507), .B2(n8183), .ZN(
        n11797) );
  AOI22_X1 U12558 ( .A1(n11752), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2396] ), .ZN(n6117) );
  MUX2_X1 U12559 ( .A(DRAMRF_DATA_IN[29]), .B(
        \DataPath/WRF_CUhw/curr_data[29] ), .S(n11840), .Z(n11549) );
  MUX2_X1 U12560 ( .A(\DataPath/i_REG_MEM_ALUOUT[29] ), .B(
        \DataPath/i_REG_LDSTR_OUT[29] ), .S(n8451), .Z(n10839) );
  OAI22_X1 U12561 ( .A1(n8436), .A2(n11301), .B1(n11508), .B2(n8183), .ZN(
        n11798) );
  AOI22_X1 U12562 ( .A1(n11753), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2397] ), .ZN(n6116) );
  MUX2_X1 U12563 ( .A(DRAMRF_DATA_IN[30]), .B(
        \DataPath/WRF_CUhw/curr_data[30] ), .S(n11840), .Z(n11550) );
  MUX2_X1 U12564 ( .A(\DataPath/i_REG_MEM_ALUOUT[30] ), .B(
        \DataPath/i_REG_LDSTR_OUT[30] ), .S(n8451), .Z(n10840) );
  OAI22_X1 U12565 ( .A1(n8437), .A2(n11302), .B1(n11509), .B2(n8183), .ZN(
        n11799) );
  AOI22_X1 U12566 ( .A1(n11754), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2398] ), .ZN(n6115) );
  MUX2_X1 U12567 ( .A(DRAMRF_DATA_IN[31]), .B(
        \DataPath/WRF_CUhw/curr_data[31] ), .S(n11840), .Z(n11551) );
  MUX2_X1 U12568 ( .A(\DataPath/i_REG_MEM_ALUOUT[31] ), .B(
        \DataPath/i_REG_LDSTR_OUT[31] ), .S(n8451), .Z(n10841) );
  OAI22_X1 U12569 ( .A1(n8437), .A2(n11304), .B1(n11512), .B2(n8183), .ZN(
        n11769) );
  AOI22_X1 U12570 ( .A1(n11803), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2399] ), .ZN(n6114) );
  NAND2_X1 U12571 ( .A1(n10932), .A2(n11477), .ZN(n11327) );
  INV_X1 U12572 ( .A(n10842), .ZN(n10843) );
  MUX2_X1 U12573 ( .A(DRAMRF_DATA_IN[0]), .B(\DataPath/WRF_CUhw/curr_data[0] ), 
        .S(n11840), .Z(n11520) );
  MUX2_X1 U12574 ( .A(\DataPath/i_REG_MEM_ALUOUT[0] ), .B(
        \DataPath/i_REG_LDSTR_OUT[0] ), .S(n8451), .Z(n10844) );
  OAI22_X1 U12575 ( .A1(n8437), .A2(n11272), .B1(n11479), .B2(n8183), .ZN(
        n11774) );
  AOI22_X1 U12576 ( .A1(\DataPath/RF/bus_reg_dataout[2336] ), .A2(n8359), .B1(
        n10862), .B2(n11774), .ZN(n6111) );
  MUX2_X1 U12577 ( .A(DRAMRF_DATA_IN[1]), .B(\DataPath/WRF_CUhw/curr_data[1] ), 
        .S(n11840), .Z(n11521) );
  MUX2_X1 U12578 ( .A(\DataPath/i_REG_MEM_ALUOUT[1] ), .B(
        \DataPath/i_REG_LDSTR_OUT[1] ), .S(n8451), .Z(n10845) );
  OAI22_X1 U12579 ( .A1(n8437), .A2(n11273), .B1(n11480), .B2(n8183), .ZN(
        n11775) );
  AOI22_X1 U12580 ( .A1(\DataPath/RF/bus_reg_dataout[2337] ), .A2(n8359), .B1(
        n10862), .B2(n11775), .ZN(n6110) );
  MUX2_X1 U12581 ( .A(DRAMRF_DATA_IN[2]), .B(\DataPath/WRF_CUhw/curr_data[2] ), 
        .S(n11840), .Z(n11522) );
  MUX2_X1 U12582 ( .A(\DataPath/i_REG_MEM_ALUOUT[2] ), .B(
        \DataPath/i_REG_LDSTR_OUT[2] ), .S(n8451), .Z(n10846) );
  OAI22_X1 U12583 ( .A1(n8437), .A2(n11274), .B1(n11481), .B2(n8183), .ZN(
        n11776) );
  AOI22_X1 U12584 ( .A1(\DataPath/RF/bus_reg_dataout[2338] ), .A2(n8359), .B1(
        n10862), .B2(n11776), .ZN(n6109) );
  MUX2_X1 U12585 ( .A(DRAMRF_DATA_IN[3]), .B(\DataPath/WRF_CUhw/curr_data[3] ), 
        .S(n11840), .Z(n11523) );
  MUX2_X1 U12586 ( .A(\DataPath/i_REG_MEM_ALUOUT[3] ), .B(
        \DataPath/i_REG_LDSTR_OUT[3] ), .S(n8451), .Z(n10847) );
  OAI22_X1 U12587 ( .A1(n8437), .A2(n11275), .B1(n11482), .B2(n8183), .ZN(
        n11777) );
  AOI22_X1 U12588 ( .A1(\DataPath/RF/bus_reg_dataout[2339] ), .A2(n10863), 
        .B1(n10862), .B2(n11777), .ZN(n6108) );
  MUX2_X1 U12589 ( .A(DRAMRF_DATA_IN[4]), .B(\DataPath/WRF_CUhw/curr_data[4] ), 
        .S(n11840), .Z(n11524) );
  MUX2_X1 U12590 ( .A(\DataPath/i_REG_MEM_ALUOUT[4] ), .B(
        \DataPath/i_REG_LDSTR_OUT[4] ), .S(n8451), .Z(n10848) );
  OAI22_X1 U12591 ( .A1(n8437), .A2(n11276), .B1(n11483), .B2(n8183), .ZN(
        n11778) );
  AOI22_X1 U12592 ( .A1(\DataPath/RF/bus_reg_dataout[2340] ), .A2(n10863), 
        .B1(n10862), .B2(n11778), .ZN(n6107) );
  MUX2_X1 U12593 ( .A(DRAMRF_DATA_IN[5]), .B(\DataPath/WRF_CUhw/curr_data[5] ), 
        .S(n11840), .Z(n11525) );
  MUX2_X1 U12594 ( .A(\DataPath/i_REG_MEM_ALUOUT[5] ), .B(
        \DataPath/i_REG_LDSTR_OUT[5] ), .S(n8451), .Z(n10849) );
  OAI22_X1 U12595 ( .A1(n8437), .A2(n11277), .B1(n11484), .B2(n8183), .ZN(
        n11779) );
  AOI22_X1 U12596 ( .A1(\DataPath/RF/bus_reg_dataout[2341] ), .A2(n8359), .B1(
        n10862), .B2(n11779), .ZN(n6106) );
  MUX2_X1 U12597 ( .A(DRAMRF_DATA_IN[6]), .B(\DataPath/WRF_CUhw/curr_data[6] ), 
        .S(n11840), .Z(n11526) );
  MUX2_X1 U12598 ( .A(\DataPath/i_REG_MEM_ALUOUT[6] ), .B(
        \DataPath/i_REG_LDSTR_OUT[6] ), .S(n8451), .Z(n10850) );
  OAI22_X1 U12599 ( .A1(n8437), .A2(n11278), .B1(n11485), .B2(n8183), .ZN(
        n11780) );
  AOI22_X1 U12600 ( .A1(\DataPath/RF/bus_reg_dataout[2342] ), .A2(n8359), .B1(
        n10862), .B2(n11780), .ZN(n6105) );
  MUX2_X1 U12601 ( .A(DRAMRF_DATA_IN[7]), .B(\DataPath/WRF_CUhw/curr_data[7] ), 
        .S(n11840), .Z(n11527) );
  MUX2_X1 U12602 ( .A(\DataPath/i_REG_MEM_ALUOUT[7] ), .B(
        \DataPath/i_REG_LDSTR_OUT[7] ), .S(n8451), .Z(n10851) );
  OAI22_X1 U12603 ( .A1(n8436), .A2(n11279), .B1(n11486), .B2(n8183), .ZN(
        n11781) );
  AOI22_X1 U12604 ( .A1(\DataPath/RF/bus_reg_dataout[2343] ), .A2(n8359), .B1(
        n10862), .B2(n11781), .ZN(n6104) );
  MUX2_X1 U12605 ( .A(DRAMRF_DATA_IN[8]), .B(\DataPath/WRF_CUhw/curr_data[8] ), 
        .S(n11840), .Z(n11528) );
  MUX2_X1 U12606 ( .A(\DataPath/i_REG_MEM_ALUOUT[8] ), .B(
        \DataPath/i_REG_LDSTR_OUT[8] ), .S(i_S3), .Z(n10852) );
  OAI22_X1 U12607 ( .A1(n8436), .A2(n11280), .B1(n11487), .B2(n8183), .ZN(
        n11782) );
  AOI22_X1 U12608 ( .A1(\DataPath/RF/bus_reg_dataout[2344] ), .A2(n10863), 
        .B1(n10862), .B2(n11782), .ZN(n6103) );
  MUX2_X1 U12609 ( .A(DRAMRF_DATA_IN[9]), .B(\DataPath/WRF_CUhw/curr_data[9] ), 
        .S(n11840), .Z(n11529) );
  MUX2_X1 U12610 ( .A(\DataPath/i_REG_MEM_ALUOUT[9] ), .B(
        \DataPath/i_REG_LDSTR_OUT[9] ), .S(i_S3), .Z(n10853) );
  OAI22_X1 U12611 ( .A1(n8436), .A2(n11281), .B1(n11488), .B2(n8183), .ZN(
        n11760) );
  AOI22_X1 U12612 ( .A1(\DataPath/RF/bus_reg_dataout[2345] ), .A2(n8359), .B1(
        n10862), .B2(n11760), .ZN(n6102) );
  MUX2_X1 U12613 ( .A(DRAMRF_DATA_IN[10]), .B(
        \DataPath/WRF_CUhw/curr_data[10] ), .S(n11840), .Z(n11530) );
  MUX2_X1 U12614 ( .A(\DataPath/i_REG_MEM_ALUOUT[10] ), .B(
        \DataPath/i_REG_LDSTR_OUT[10] ), .S(i_S3), .Z(n10854) );
  OAI22_X1 U12615 ( .A1(n8436), .A2(n11282), .B1(n11489), .B2(n8183), .ZN(
        n11783) );
  AOI22_X1 U12616 ( .A1(\DataPath/RF/bus_reg_dataout[2346] ), .A2(n8359), .B1(
        n10862), .B2(n11783), .ZN(n6101) );
  MUX2_X1 U12617 ( .A(DRAMRF_DATA_IN[11]), .B(
        \DataPath/WRF_CUhw/curr_data[11] ), .S(n11840), .Z(n11531) );
  MUX2_X1 U12618 ( .A(\DataPath/i_REG_MEM_ALUOUT[11] ), .B(
        \DataPath/i_REG_LDSTR_OUT[11] ), .S(i_S3), .Z(n10855) );
  OAI22_X1 U12619 ( .A1(n8436), .A2(n11283), .B1(n11490), .B2(n8183), .ZN(
        n11784) );
  AOI22_X1 U12620 ( .A1(\DataPath/RF/bus_reg_dataout[2347] ), .A2(n8359), .B1(
        n10862), .B2(n11784), .ZN(n6100) );
  MUX2_X1 U12621 ( .A(DRAMRF_DATA_IN[12]), .B(
        \DataPath/WRF_CUhw/curr_data[12] ), .S(n11840), .Z(n11532) );
  MUX2_X1 U12622 ( .A(\DataPath/i_REG_MEM_ALUOUT[12] ), .B(
        \DataPath/i_REG_LDSTR_OUT[12] ), .S(i_S3), .Z(n10856) );
  OAI22_X1 U12623 ( .A1(n8436), .A2(n11284), .B1(n11491), .B2(n8183), .ZN(
        n11761) );
  AOI22_X1 U12624 ( .A1(\DataPath/RF/bus_reg_dataout[2348] ), .A2(n10863), 
        .B1(n10862), .B2(n11761), .ZN(n6099) );
  MUX2_X1 U12625 ( .A(DRAMRF_DATA_IN[13]), .B(
        \DataPath/WRF_CUhw/curr_data[13] ), .S(n11840), .Z(n11533) );
  MUX2_X1 U12626 ( .A(\DataPath/i_REG_MEM_ALUOUT[13] ), .B(
        \DataPath/i_REG_LDSTR_OUT[13] ), .S(i_S3), .Z(n10857) );
  OAI22_X1 U12627 ( .A1(n8436), .A2(n11285), .B1(n11492), .B2(n8183), .ZN(
        n11785) );
  AOI22_X1 U12628 ( .A1(\DataPath/RF/bus_reg_dataout[2349] ), .A2(n10863), 
        .B1(n10862), .B2(n11785), .ZN(n6098) );
  MUX2_X1 U12629 ( .A(DRAMRF_DATA_IN[14]), .B(
        \DataPath/WRF_CUhw/curr_data[14] ), .S(n11840), .Z(n11534) );
  MUX2_X1 U12630 ( .A(\DataPath/i_REG_MEM_ALUOUT[14] ), .B(
        \DataPath/i_REG_LDSTR_OUT[14] ), .S(i_S3), .Z(n10858) );
  OAI22_X1 U12631 ( .A1(n8436), .A2(n11286), .B1(n11493), .B2(n8183), .ZN(
        n11786) );
  AOI22_X1 U12632 ( .A1(\DataPath/RF/bus_reg_dataout[2350] ), .A2(n10863), 
        .B1(n10862), .B2(n11786), .ZN(n6097) );
  MUX2_X1 U12633 ( .A(DRAMRF_DATA_IN[15]), .B(
        \DataPath/WRF_CUhw/curr_data[15] ), .S(n11840), .Z(n11535) );
  MUX2_X1 U12634 ( .A(\DataPath/i_REG_MEM_ALUOUT[15] ), .B(
        \DataPath/i_REG_LDSTR_OUT[15] ), .S(i_S3), .Z(n10859) );
  OAI22_X1 U12635 ( .A1(n8436), .A2(n11287), .B1(n11494), .B2(n8183), .ZN(
        n11762) );
  AOI22_X1 U12636 ( .A1(\DataPath/RF/bus_reg_dataout[2351] ), .A2(n8359), .B1(
        n10862), .B2(n11762), .ZN(n6096) );
  MUX2_X1 U12637 ( .A(DRAMRF_DATA_IN[16]), .B(
        \DataPath/WRF_CUhw/curr_data[16] ), .S(n11840), .Z(n11536) );
  MUX2_X1 U12638 ( .A(\DataPath/i_REG_MEM_ALUOUT[16] ), .B(
        \DataPath/i_REG_LDSTR_OUT[16] ), .S(i_S3), .Z(n10860) );
  OAI22_X1 U12639 ( .A1(n8436), .A2(n11288), .B1(n11495), .B2(n8183), .ZN(
        n11763) );
  AOI22_X1 U12640 ( .A1(\DataPath/RF/bus_reg_dataout[2352] ), .A2(n8359), .B1(
        n10862), .B2(n11763), .ZN(n6095) );
  MUX2_X1 U12641 ( .A(DRAMRF_DATA_IN[17]), .B(
        \DataPath/WRF_CUhw/curr_data[17] ), .S(n11840), .Z(n11537) );
  MUX2_X1 U12642 ( .A(\DataPath/i_REG_MEM_ALUOUT[17] ), .B(
        \DataPath/i_REG_LDSTR_OUT[17] ), .S(i_S3), .Z(n10861) );
  OAI22_X1 U12643 ( .A1(n8436), .A2(n11289), .B1(n11496), .B2(n8183), .ZN(
        n11764) );
  AOI22_X1 U12644 ( .A1(\DataPath/RF/bus_reg_dataout[2353] ), .A2(n10863), 
        .B1(n10862), .B2(n11764), .ZN(n6094) );
  AOI22_X1 U12645 ( .A1(\DataPath/RF/bus_reg_dataout[2354] ), .A2(n8359), .B1(
        n10862), .B2(n11787), .ZN(n6093) );
  AOI22_X1 U12646 ( .A1(n11747), .A2(n10864), .B1(n10863), .B2(
        \DataPath/RF/bus_reg_dataout[2355] ), .ZN(n6092) );
  AOI22_X1 U12647 ( .A1(\DataPath/RF/bus_reg_dataout[2356] ), .A2(n8359), .B1(
        n10862), .B2(n11789), .ZN(n6091) );
  AOI22_X1 U12648 ( .A1(\DataPath/RF/bus_reg_dataout[2357] ), .A2(n8359), .B1(
        n10862), .B2(n11790), .ZN(n6090) );
  AOI22_X1 U12649 ( .A1(\DataPath/RF/bus_reg_dataout[2358] ), .A2(n8359), .B1(
        n10862), .B2(n11765), .ZN(n6089) );
  AOI22_X1 U12650 ( .A1(\DataPath/RF/bus_reg_dataout[2359] ), .A2(n8359), .B1(
        n10862), .B2(n11792), .ZN(n6088) );
  AOI22_X1 U12651 ( .A1(n11793), .A2(n10864), .B1(n8359), .B2(
        \DataPath/RF/bus_reg_dataout[2360] ), .ZN(n6087) );
  AOI22_X1 U12652 ( .A1(n11794), .A2(n10864), .B1(n8359), .B2(
        \DataPath/RF/bus_reg_dataout[2361] ), .ZN(n6086) );
  AOI22_X1 U12653 ( .A1(\DataPath/RF/bus_reg_dataout[2362] ), .A2(n10863), 
        .B1(n10862), .B2(n11795), .ZN(n6085) );
  AOI22_X1 U12654 ( .A1(\DataPath/RF/bus_reg_dataout[2363] ), .A2(n8359), .B1(
        n10862), .B2(n11768), .ZN(n6084) );
  AOI22_X1 U12655 ( .A1(n11752), .A2(n10864), .B1(n8359), .B2(
        \DataPath/RF/bus_reg_dataout[2364] ), .ZN(n6083) );
  AOI22_X1 U12656 ( .A1(\DataPath/RF/bus_reg_dataout[2365] ), .A2(n8359), .B1(
        n10862), .B2(n11798), .ZN(n6082) );
  AOI22_X1 U12657 ( .A1(\DataPath/RF/bus_reg_dataout[2366] ), .A2(n8359), .B1(
        n10862), .B2(n11799), .ZN(n6081) );
  AOI22_X1 U12658 ( .A1(n11803), .A2(n10864), .B1(n10863), .B2(
        \DataPath/RF/bus_reg_dataout[2367] ), .ZN(n6078) );
  NAND2_X1 U12659 ( .A1(n10932), .A2(n10911), .ZN(n11333) );
  INV_X1 U12660 ( .A(n10865), .ZN(n10866) );
  AOI22_X1 U12661 ( .A1(n11804), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2304] ), .ZN(n6075) );
  AOI22_X1 U12662 ( .A1(n11805), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2305] ), .ZN(n6074) );
  AOI22_X1 U12663 ( .A1(n11806), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2306] ), .ZN(n6073) );
  AOI22_X1 U12664 ( .A1(n11807), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2307] ), .ZN(n6072) );
  AOI22_X1 U12665 ( .A1(n11808), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2308] ), .ZN(n6071) );
  AOI22_X1 U12666 ( .A1(n11809), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2309] ), .ZN(n6070) );
  AOI22_X1 U12667 ( .A1(n11810), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2310] ), .ZN(n6069) );
  AOI22_X1 U12668 ( .A1(n11811), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2311] ), .ZN(n6068) );
  AOI22_X1 U12669 ( .A1(n11812), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2312] ), .ZN(n6067) );
  AOI22_X1 U12670 ( .A1(n11813), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2313] ), .ZN(n6066) );
  AOI22_X1 U12671 ( .A1(n11814), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2314] ), .ZN(n6065) );
  AOI22_X1 U12672 ( .A1(n11815), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2315] ), .ZN(n6064) );
  AOI22_X1 U12673 ( .A1(n11816), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2316] ), .ZN(n6063) );
  AOI22_X1 U12674 ( .A1(n11817), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2317] ), .ZN(n6062) );
  AOI22_X1 U12675 ( .A1(n11818), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2318] ), .ZN(n6061) );
  AOI22_X1 U12676 ( .A1(n11819), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2319] ), .ZN(n6060) );
  AOI22_X1 U12677 ( .A1(n11820), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2320] ), .ZN(n6059) );
  AOI22_X1 U12678 ( .A1(n11823), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2321] ), .ZN(n6058) );
  AOI22_X1 U12679 ( .A1(n11746), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2322] ), .ZN(n6057) );
  AOI22_X1 U12680 ( .A1(n11747), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2323] ), .ZN(n6056) );
  AOI22_X1 U12681 ( .A1(n11748), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2324] ), .ZN(n6055) );
  AOI22_X1 U12682 ( .A1(n11749), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2325] ), .ZN(n6054) );
  AOI22_X1 U12683 ( .A1(n11791), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2326] ), .ZN(n6053) );
  AOI22_X1 U12684 ( .A1(n11750), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2327] ), .ZN(n6052) );
  AOI22_X1 U12685 ( .A1(n11793), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2328] ), .ZN(n6051) );
  AOI22_X1 U12686 ( .A1(n11794), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2329] ), .ZN(n6050) );
  AOI22_X1 U12687 ( .A1(n11751), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2330] ), .ZN(n6049) );
  AOI22_X1 U12688 ( .A1(n11796), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2331] ), .ZN(n6048) );
  AOI22_X1 U12689 ( .A1(n11752), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2332] ), .ZN(n6047) );
  AOI22_X1 U12690 ( .A1(n11753), .A2(n10868), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2333] ), .ZN(n6046) );
  AOI22_X1 U12691 ( .A1(n11754), .A2(n8360), .B1(n8361), .B2(
        \DataPath/RF/bus_reg_dataout[2334] ), .ZN(n6045) );
  AOI22_X1 U12692 ( .A1(n11803), .A2(n8360), .B1(n10867), .B2(
        \DataPath/RF/bus_reg_dataout[2335] ), .ZN(n6042) );
  NAND2_X1 U12693 ( .A1(n11452), .A2(n10909), .ZN(n11339) );
  NAND2_X1 U12694 ( .A1(n11452), .A2(n10910), .ZN(n11338) );
  OAI22_X1 U12695 ( .A1(n8293), .A2(n11339), .B1(n8450), .B2(n11338), .ZN(
        n10871) );
  AOI22_X1 U12696 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2272] ), 
        .B1(n11804), .B2(n10872), .ZN(n6038) );
  AOI22_X1 U12697 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2273] ), 
        .B1(n11805), .B2(n10872), .ZN(n6037) );
  AOI22_X1 U12698 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2274] ), 
        .B1(n11806), .B2(n10872), .ZN(n6036) );
  AOI22_X1 U12699 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2275] ), 
        .B1(n11807), .B2(n10872), .ZN(n6035) );
  AOI22_X1 U12700 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2276] ), 
        .B1(n11808), .B2(n10872), .ZN(n6034) );
  AOI22_X1 U12701 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2277] ), 
        .B1(n11809), .B2(n10872), .ZN(n6033) );
  AOI22_X1 U12702 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2278] ), 
        .B1(n11810), .B2(n10872), .ZN(n6032) );
  NOR2_X1 U12703 ( .A1(RST), .A2(n10874), .ZN(n10873) );
  AOI22_X1 U12704 ( .A1(\DataPath/RF/bus_reg_dataout[2279] ), .A2(n10874), 
        .B1(n10873), .B2(n11781), .ZN(n6031) );
  AOI22_X1 U12705 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2280] ), 
        .B1(n11812), .B2(n10872), .ZN(n6030) );
  AOI22_X1 U12706 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2281] ), 
        .B1(n11813), .B2(n10872), .ZN(n6029) );
  AOI22_X1 U12707 ( .A1(\DataPath/RF/bus_reg_dataout[2282] ), .A2(n10874), 
        .B1(n10873), .B2(n11783), .ZN(n6028) );
  AOI22_X1 U12708 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2283] ), 
        .B1(n11815), .B2(n10872), .ZN(n6027) );
  AOI22_X1 U12709 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2284] ), 
        .B1(n11816), .B2(n10872), .ZN(n6026) );
  AOI22_X1 U12710 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2285] ), 
        .B1(n11817), .B2(n10872), .ZN(n6025) );
  AOI22_X1 U12711 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2286] ), 
        .B1(n11818), .B2(n10872), .ZN(n6024) );
  AOI22_X1 U12712 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2287] ), 
        .B1(n11819), .B2(n10872), .ZN(n6023) );
  AOI22_X1 U12713 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2288] ), 
        .B1(n11820), .B2(n10872), .ZN(n6022) );
  AOI22_X1 U12714 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2289] ), 
        .B1(n11823), .B2(n10872), .ZN(n6021) );
  AOI22_X1 U12715 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2290] ), 
        .B1(n11746), .B2(n10872), .ZN(n6020) );
  AOI22_X1 U12716 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2291] ), 
        .B1(n11747), .B2(n10872), .ZN(n6019) );
  AOI22_X1 U12717 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2292] ), 
        .B1(n11748), .B2(n10872), .ZN(n6018) );
  AOI22_X1 U12718 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2293] ), 
        .B1(n11749), .B2(n10872), .ZN(n6017) );
  AOI22_X1 U12719 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2294] ), 
        .B1(n11791), .B2(n10872), .ZN(n6016) );
  AOI22_X1 U12720 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2295] ), 
        .B1(n11750), .B2(n10872), .ZN(n6015) );
  AOI22_X1 U12721 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2296] ), 
        .B1(n11793), .B2(n10872), .ZN(n6014) );
  AOI22_X1 U12722 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2297] ), 
        .B1(n11794), .B2(n10872), .ZN(n6013) );
  AOI22_X1 U12723 ( .A1(\DataPath/RF/bus_reg_dataout[2298] ), .A2(n10874), 
        .B1(n10873), .B2(n11795), .ZN(n6012) );
  AOI22_X1 U12724 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2299] ), 
        .B1(n11796), .B2(n10872), .ZN(n6011) );
  AOI22_X1 U12725 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2300] ), 
        .B1(n11752), .B2(n10872), .ZN(n6010) );
  AOI22_X1 U12726 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2301] ), 
        .B1(n11753), .B2(n10872), .ZN(n6009) );
  AOI22_X1 U12727 ( .A1(n10874), .A2(\DataPath/RF/bus_reg_dataout[2302] ), 
        .B1(n11754), .B2(n10872), .ZN(n6008) );
  AOI22_X1 U12728 ( .A1(\DataPath/RF/bus_reg_dataout[2303] ), .A2(n10874), 
        .B1(n10873), .B2(n11769), .ZN(n6005) );
  NAND2_X1 U12729 ( .A1(n10910), .A2(n11456), .ZN(n11194) );
  NAND2_X1 U12730 ( .A1(n10909), .A2(n11456), .ZN(n11346) );
  INV_X1 U12731 ( .A(n10875), .ZN(n10876) );
  OAI22_X1 U12732 ( .A1(n8293), .A2(n11346), .B1(n11345), .B2(n8436), .ZN(
        n10877) );
  AOI22_X1 U12733 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2240] ), 
        .B1(n11804), .B2(n10879), .ZN(n6002) );
  AOI22_X1 U12734 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2241] ), 
        .B1(n11805), .B2(n10879), .ZN(n6001) );
  AOI22_X1 U12735 ( .A1(\DataPath/RF/bus_reg_dataout[2242] ), .A2(n10880), 
        .B1(n10878), .B2(n11776), .ZN(n6000) );
  AOI22_X1 U12736 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2243] ), 
        .B1(n11807), .B2(n10879), .ZN(n5999) );
  AOI22_X1 U12737 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2244] ), 
        .B1(n11808), .B2(n10879), .ZN(n5998) );
  AOI22_X1 U12738 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2245] ), 
        .B1(n11809), .B2(n10879), .ZN(n5997) );
  AOI22_X1 U12739 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2246] ), 
        .B1(n11810), .B2(n10879), .ZN(n5996) );
  AOI22_X1 U12740 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2247] ), 
        .B1(n11811), .B2(n10879), .ZN(n5995) );
  AOI22_X1 U12741 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2248] ), 
        .B1(n11812), .B2(n10879), .ZN(n5994) );
  AOI22_X1 U12742 ( .A1(\DataPath/RF/bus_reg_dataout[2249] ), .A2(n10880), 
        .B1(n10878), .B2(n11760), .ZN(n5993) );
  AOI22_X1 U12743 ( .A1(\DataPath/RF/bus_reg_dataout[2250] ), .A2(n10880), 
        .B1(n10878), .B2(n11783), .ZN(n5992) );
  AOI22_X1 U12744 ( .A1(\DataPath/RF/bus_reg_dataout[2251] ), .A2(n10880), 
        .B1(n10878), .B2(n11784), .ZN(n5991) );
  AOI22_X1 U12745 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2252] ), 
        .B1(n11816), .B2(n10879), .ZN(n5990) );
  AOI22_X1 U12746 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2253] ), 
        .B1(n11817), .B2(n10879), .ZN(n5989) );
  AOI22_X1 U12747 ( .A1(\DataPath/RF/bus_reg_dataout[2254] ), .A2(n10880), 
        .B1(n10878), .B2(n11786), .ZN(n5988) );
  AOI22_X1 U12748 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2255] ), 
        .B1(n11819), .B2(n10879), .ZN(n5987) );
  AOI22_X1 U12749 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2256] ), 
        .B1(n11820), .B2(n10879), .ZN(n5986) );
  AOI22_X1 U12750 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2257] ), 
        .B1(n11823), .B2(n10879), .ZN(n5985) );
  AOI22_X1 U12751 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2258] ), 
        .B1(n11746), .B2(n10879), .ZN(n5984) );
  AOI22_X1 U12752 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2259] ), 
        .B1(n11747), .B2(n10879), .ZN(n5983) );
  AOI22_X1 U12753 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2260] ), 
        .B1(n11748), .B2(n10879), .ZN(n5982) );
  AOI22_X1 U12754 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2261] ), 
        .B1(n11749), .B2(n10879), .ZN(n5981) );
  AOI22_X1 U12755 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2262] ), 
        .B1(n11791), .B2(n10879), .ZN(n5980) );
  AOI22_X1 U12756 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2263] ), 
        .B1(n11750), .B2(n10879), .ZN(n5979) );
  AOI22_X1 U12757 ( .A1(\DataPath/RF/bus_reg_dataout[2264] ), .A2(n10880), 
        .B1(n10878), .B2(n11766), .ZN(n5978) );
  AOI22_X1 U12758 ( .A1(\DataPath/RF/bus_reg_dataout[2265] ), .A2(n10880), 
        .B1(n10878), .B2(n11767), .ZN(n5977) );
  AOI22_X1 U12759 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2266] ), 
        .B1(n11751), .B2(n10879), .ZN(n5976) );
  AOI22_X1 U12760 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2267] ), 
        .B1(n11796), .B2(n10879), .ZN(n5975) );
  AOI22_X1 U12761 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2268] ), 
        .B1(n11752), .B2(n10879), .ZN(n5974) );
  AOI22_X1 U12762 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2269] ), 
        .B1(n11753), .B2(n10879), .ZN(n5973) );
  AOI22_X1 U12763 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2270] ), 
        .B1(n11754), .B2(n10879), .ZN(n5972) );
  AOI22_X1 U12764 ( .A1(n10880), .A2(\DataPath/RF/bus_reg_dataout[2271] ), 
        .B1(n11803), .B2(n10879), .ZN(n5969) );
  NAND2_X1 U12765 ( .A1(n10910), .A2(n11460), .ZN(n11070) );
  NAND2_X1 U12766 ( .A1(n10909), .A2(n11460), .ZN(n11353) );
  INV_X1 U12767 ( .A(n10881), .ZN(n10882) );
  AOI22_X1 U12768 ( .A1(n10295), .A2(\DataPath/RF/POP_ADDRGEN/curr_addr[10] ), 
        .B1(n10882), .B2(n10934), .ZN(n11352) );
  OAI22_X1 U12769 ( .A1(n8293), .A2(n11353), .B1(n11352), .B2(n8436), .ZN(
        n10883) );
  AOI22_X1 U12770 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2208] ), 
        .B1(n11804), .B2(n10885), .ZN(n5966) );
  AOI22_X1 U12771 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2209] ), 
        .B1(n11805), .B2(n10885), .ZN(n5965) );
  AOI22_X1 U12772 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2210] ), 
        .B1(n11806), .B2(n10885), .ZN(n5964) );
  AOI22_X1 U12773 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2211] ), 
        .B1(n11807), .B2(n10885), .ZN(n5963) );
  AOI22_X1 U12774 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2212] ), 
        .B1(n11808), .B2(n10885), .ZN(n5962) );
  AOI22_X1 U12775 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2213] ), 
        .B1(n11809), .B2(n10885), .ZN(n5961) );
  AOI22_X1 U12776 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2214] ), 
        .B1(n11810), .B2(n10885), .ZN(n5960) );
  NOR2_X1 U12777 ( .A1(RST), .A2(n10886), .ZN(n10884) );
  AOI22_X1 U12778 ( .A1(\DataPath/RF/bus_reg_dataout[2215] ), .A2(n10886), 
        .B1(n10884), .B2(n11781), .ZN(n5959) );
  AOI22_X1 U12779 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2216] ), 
        .B1(n11812), .B2(n10885), .ZN(n5958) );
  AOI22_X1 U12780 ( .A1(\DataPath/RF/bus_reg_dataout[2217] ), .A2(n10886), 
        .B1(n10884), .B2(n11760), .ZN(n5957) );
  AOI22_X1 U12781 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2218] ), 
        .B1(n11814), .B2(n10885), .ZN(n5956) );
  AOI22_X1 U12782 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2219] ), 
        .B1(n11815), .B2(n10885), .ZN(n5955) );
  AOI22_X1 U12783 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2220] ), 
        .B1(n11816), .B2(n10885), .ZN(n5954) );
  AOI22_X1 U12784 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2221] ), 
        .B1(n11817), .B2(n10885), .ZN(n5953) );
  AOI22_X1 U12785 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2222] ), 
        .B1(n11818), .B2(n10885), .ZN(n5952) );
  AOI22_X1 U12786 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2223] ), 
        .B1(n11819), .B2(n10885), .ZN(n5951) );
  AOI22_X1 U12787 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2224] ), 
        .B1(n11820), .B2(n10885), .ZN(n5950) );
  AOI22_X1 U12788 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2225] ), 
        .B1(n11823), .B2(n10885), .ZN(n5949) );
  AOI22_X1 U12789 ( .A1(\DataPath/RF/bus_reg_dataout[2226] ), .A2(n10886), 
        .B1(n10884), .B2(n11787), .ZN(n5948) );
  AOI22_X1 U12790 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2227] ), 
        .B1(n11747), .B2(n10885), .ZN(n5947) );
  AOI22_X1 U12791 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2228] ), 
        .B1(n11748), .B2(n10885), .ZN(n5946) );
  AOI22_X1 U12792 ( .A1(\DataPath/RF/bus_reg_dataout[2229] ), .A2(n10886), 
        .B1(n10884), .B2(n11790), .ZN(n5945) );
  AOI22_X1 U12793 ( .A1(\DataPath/RF/bus_reg_dataout[2230] ), .A2(n10886), 
        .B1(n10884), .B2(n11765), .ZN(n5944) );
  AOI22_X1 U12794 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2231] ), 
        .B1(n11750), .B2(n10885), .ZN(n5943) );
  AOI22_X1 U12795 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2232] ), 
        .B1(n11793), .B2(n10885), .ZN(n5942) );
  AOI22_X1 U12796 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2233] ), 
        .B1(n11794), .B2(n10885), .ZN(n5941) );
  AOI22_X1 U12797 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2234] ), 
        .B1(n11751), .B2(n10885), .ZN(n5940) );
  AOI22_X1 U12798 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2235] ), 
        .B1(n11796), .B2(n10885), .ZN(n5939) );
  AOI22_X1 U12799 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2236] ), 
        .B1(n11752), .B2(n10885), .ZN(n5938) );
  AOI22_X1 U12800 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2237] ), 
        .B1(n11753), .B2(n10885), .ZN(n5937) );
  AOI22_X1 U12801 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2238] ), 
        .B1(n11754), .B2(n10885), .ZN(n5936) );
  AOI22_X1 U12802 ( .A1(n10886), .A2(\DataPath/RF/bus_reg_dataout[2239] ), 
        .B1(n11803), .B2(n10885), .ZN(n5933) );
  NAND2_X1 U12803 ( .A1(n10910), .A2(n11464), .ZN(n11359) );
  NAND2_X1 U12804 ( .A1(n10909), .A2(n11464), .ZN(n11360) );
  INV_X1 U12805 ( .A(n10887), .ZN(n10888) );
  OAI22_X1 U12806 ( .A1(n8293), .A2(n11360), .B1(n11361), .B2(n8437), .ZN(
        n10889) );
  AOI22_X1 U12807 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2176] ), 
        .B1(n11804), .B2(n10890), .ZN(n5930) );
  AOI22_X1 U12808 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2177] ), 
        .B1(n11805), .B2(n10890), .ZN(n5929) );
  AOI22_X1 U12809 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2178] ), 
        .B1(n11806), .B2(n10890), .ZN(n5928) );
  AOI22_X1 U12810 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2179] ), 
        .B1(n11807), .B2(n10890), .ZN(n5927) );
  AOI22_X1 U12811 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2180] ), 
        .B1(n11808), .B2(n10890), .ZN(n5926) );
  AOI22_X1 U12812 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2181] ), 
        .B1(n11809), .B2(n10890), .ZN(n5925) );
  AOI22_X1 U12813 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2182] ), 
        .B1(n11810), .B2(n10890), .ZN(n5924) );
  AOI22_X1 U12814 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2183] ), 
        .B1(n11811), .B2(n10890), .ZN(n5923) );
  AOI22_X1 U12815 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2184] ), 
        .B1(n11812), .B2(n10890), .ZN(n5922) );
  AOI22_X1 U12816 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2185] ), 
        .B1(n11813), .B2(n10890), .ZN(n5921) );
  AOI22_X1 U12817 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2186] ), 
        .B1(n11814), .B2(n10890), .ZN(n5920) );
  AOI22_X1 U12818 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2187] ), 
        .B1(n11815), .B2(n10890), .ZN(n5919) );
  AOI22_X1 U12819 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2188] ), 
        .B1(n11816), .B2(n10890), .ZN(n5918) );
  AOI22_X1 U12820 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2189] ), 
        .B1(n11817), .B2(n10890), .ZN(n5917) );
  AOI22_X1 U12821 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2190] ), 
        .B1(n11818), .B2(n10890), .ZN(n5916) );
  AOI22_X1 U12822 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2191] ), 
        .B1(n11819), .B2(n10890), .ZN(n5915) );
  AOI22_X1 U12823 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2192] ), 
        .B1(n11820), .B2(n10890), .ZN(n5914) );
  AOI22_X1 U12824 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2193] ), 
        .B1(n11823), .B2(n10890), .ZN(n5913) );
  AOI22_X1 U12825 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2194] ), 
        .B1(n11746), .B2(n10890), .ZN(n5912) );
  AOI22_X1 U12826 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2195] ), 
        .B1(n11747), .B2(n10890), .ZN(n5911) );
  AOI22_X1 U12827 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2196] ), 
        .B1(n11748), .B2(n10890), .ZN(n5910) );
  AOI22_X1 U12828 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2197] ), 
        .B1(n11749), .B2(n10890), .ZN(n5909) );
  AOI22_X1 U12829 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2198] ), 
        .B1(n11791), .B2(n10890), .ZN(n5908) );
  AOI22_X1 U12830 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2199] ), 
        .B1(n11750), .B2(n10890), .ZN(n5907) );
  AOI22_X1 U12831 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2200] ), 
        .B1(n11793), .B2(n10890), .ZN(n5906) );
  AOI22_X1 U12832 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2201] ), 
        .B1(n11794), .B2(n10890), .ZN(n5905) );
  AOI22_X1 U12833 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2202] ), 
        .B1(n11751), .B2(n10890), .ZN(n5904) );
  AOI22_X1 U12834 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2203] ), 
        .B1(n11796), .B2(n10890), .ZN(n5903) );
  AOI22_X1 U12835 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2204] ), 
        .B1(n11752), .B2(n10890), .ZN(n5902) );
  AOI22_X1 U12836 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2205] ), 
        .B1(n11753), .B2(n10890), .ZN(n5901) );
  AOI22_X1 U12837 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2206] ), 
        .B1(n11754), .B2(n10890), .ZN(n5900) );
  AOI22_X1 U12838 ( .A1(n10891), .A2(\DataPath/RF/bus_reg_dataout[2207] ), 
        .B1(n11803), .B2(n10890), .ZN(n5897) );
  NAND2_X1 U12839 ( .A1(n10909), .A2(n11468), .ZN(n11367) );
  INV_X1 U12840 ( .A(n10892), .ZN(n10893) );
  OAI22_X1 U12841 ( .A1(n8293), .A2(n11367), .B1(n11366), .B2(n8437), .ZN(
        n10894) );
  AOI22_X1 U12842 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2144] ), 
        .B1(n11804), .B2(n10896), .ZN(n5894) );
  AOI22_X1 U12843 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2145] ), 
        .B1(n11805), .B2(n10896), .ZN(n5893) );
  AOI22_X1 U12844 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2146] ), 
        .B1(n11806), .B2(n10896), .ZN(n5892) );
  AOI22_X1 U12845 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2147] ), 
        .B1(n11807), .B2(n10896), .ZN(n5891) );
  AOI22_X1 U12846 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2148] ), 
        .B1(n11808), .B2(n10896), .ZN(n5890) );
  AOI22_X1 U12847 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2149] ), 
        .B1(n11809), .B2(n10896), .ZN(n5889) );
  AOI22_X1 U12848 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2150] ), 
        .B1(n11810), .B2(n10896), .ZN(n5888) );
  NOR2_X1 U12849 ( .A1(RST), .A2(n10897), .ZN(n10895) );
  AOI22_X1 U12850 ( .A1(\DataPath/RF/bus_reg_dataout[2151] ), .A2(n10897), 
        .B1(n10895), .B2(n11781), .ZN(n5887) );
  AOI22_X1 U12851 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2152] ), 
        .B1(n11812), .B2(n10896), .ZN(n5886) );
  AOI22_X1 U12852 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2153] ), 
        .B1(n11813), .B2(n10896), .ZN(n5885) );
  AOI22_X1 U12853 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2154] ), 
        .B1(n11814), .B2(n10896), .ZN(n5884) );
  AOI22_X1 U12854 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2155] ), 
        .B1(n11815), .B2(n10896), .ZN(n5883) );
  AOI22_X1 U12855 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2156] ), 
        .B1(n11816), .B2(n10896), .ZN(n5882) );
  AOI22_X1 U12856 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2157] ), 
        .B1(n11817), .B2(n10896), .ZN(n5881) );
  AOI22_X1 U12857 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2158] ), 
        .B1(n11818), .B2(n10896), .ZN(n5880) );
  AOI22_X1 U12858 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2159] ), 
        .B1(n11819), .B2(n10896), .ZN(n5879) );
  AOI22_X1 U12859 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2160] ), 
        .B1(n11820), .B2(n10896), .ZN(n5878) );
  AOI22_X1 U12860 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2161] ), 
        .B1(n11823), .B2(n10896), .ZN(n5877) );
  AOI22_X1 U12861 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2162] ), 
        .B1(n11746), .B2(n10896), .ZN(n5876) );
  AOI22_X1 U12862 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2163] ), 
        .B1(n11747), .B2(n10896), .ZN(n5875) );
  AOI22_X1 U12863 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2164] ), 
        .B1(n11748), .B2(n10896), .ZN(n5874) );
  AOI22_X1 U12864 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2165] ), 
        .B1(n11749), .B2(n10896), .ZN(n5873) );
  AOI22_X1 U12865 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2166] ), 
        .B1(n11791), .B2(n10896), .ZN(n5872) );
  AOI22_X1 U12866 ( .A1(\DataPath/RF/bus_reg_dataout[2167] ), .A2(n10897), 
        .B1(n10895), .B2(n11792), .ZN(n5871) );
  AOI22_X1 U12867 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2168] ), 
        .B1(n11793), .B2(n10896), .ZN(n5870) );
  AOI22_X1 U12868 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2169] ), 
        .B1(n11794), .B2(n10896), .ZN(n5869) );
  AOI22_X1 U12869 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2170] ), 
        .B1(n11751), .B2(n10896), .ZN(n5868) );
  AOI22_X1 U12870 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2171] ), 
        .B1(n11796), .B2(n10896), .ZN(n5867) );
  AOI22_X1 U12871 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2172] ), 
        .B1(n11752), .B2(n10896), .ZN(n5866) );
  AOI22_X1 U12872 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2173] ), 
        .B1(n11753), .B2(n10896), .ZN(n5865) );
  AOI22_X1 U12873 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2174] ), 
        .B1(n11754), .B2(n10896), .ZN(n5864) );
  AOI22_X1 U12874 ( .A1(n10897), .A2(\DataPath/RF/bus_reg_dataout[2175] ), 
        .B1(n11803), .B2(n10896), .ZN(n5861) );
  NAND2_X1 U12875 ( .A1(n10909), .A2(n11472), .ZN(n11375) );
  NAND2_X1 U12876 ( .A1(n10910), .A2(n11472), .ZN(n11374) );
  OAI22_X1 U12877 ( .A1(n8293), .A2(n11375), .B1(n8173), .B2(n11374), .ZN(
        n10899) );
  AOI22_X1 U12878 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2112] ), 
        .B1(n11804), .B2(n10901), .ZN(n5858) );
  AOI22_X1 U12879 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2113] ), 
        .B1(n11805), .B2(n10901), .ZN(n5857) );
  AOI22_X1 U12880 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2114] ), 
        .B1(n11806), .B2(n10901), .ZN(n5856) );
  AOI22_X1 U12881 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2115] ), 
        .B1(n11807), .B2(n10901), .ZN(n5855) );
  AOI22_X1 U12882 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2116] ), 
        .B1(n11808), .B2(n10901), .ZN(n5854) );
  AOI22_X1 U12883 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2117] ), 
        .B1(n11809), .B2(n10901), .ZN(n5853) );
  NOR2_X1 U12884 ( .A1(RST), .A2(n10902), .ZN(n10900) );
  AOI22_X1 U12885 ( .A1(\DataPath/RF/bus_reg_dataout[2118] ), .A2(n10902), 
        .B1(n10900), .B2(n11780), .ZN(n5852) );
  AOI22_X1 U12886 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2119] ), 
        .B1(n11811), .B2(n10901), .ZN(n5851) );
  AOI22_X1 U12887 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2120] ), 
        .B1(n11812), .B2(n10901), .ZN(n5850) );
  AOI22_X1 U12888 ( .A1(\DataPath/RF/bus_reg_dataout[2121] ), .A2(n10902), 
        .B1(n10900), .B2(n11760), .ZN(n5849) );
  AOI22_X1 U12889 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2122] ), 
        .B1(n11814), .B2(n10901), .ZN(n5848) );
  AOI22_X1 U12890 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2123] ), 
        .B1(n11815), .B2(n10901), .ZN(n5847) );
  AOI22_X1 U12891 ( .A1(\DataPath/RF/bus_reg_dataout[2124] ), .A2(n10902), 
        .B1(n10900), .B2(n11761), .ZN(n5846) );
  AOI22_X1 U12892 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2125] ), 
        .B1(n11817), .B2(n10901), .ZN(n5845) );
  AOI22_X1 U12893 ( .A1(\DataPath/RF/bus_reg_dataout[2126] ), .A2(n10902), 
        .B1(n10900), .B2(n11786), .ZN(n5844) );
  AOI22_X1 U12894 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2127] ), 
        .B1(n11819), .B2(n10901), .ZN(n5843) );
  AOI22_X1 U12895 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2128] ), 
        .B1(n11820), .B2(n10901), .ZN(n5842) );
  AOI22_X1 U12896 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2129] ), 
        .B1(n11823), .B2(n10901), .ZN(n5841) );
  AOI22_X1 U12897 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2130] ), 
        .B1(n11746), .B2(n10901), .ZN(n5840) );
  AOI22_X1 U12898 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2131] ), 
        .B1(n11747), .B2(n10901), .ZN(n5839) );
  AOI22_X1 U12899 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2132] ), 
        .B1(n11748), .B2(n10901), .ZN(n5838) );
  AOI22_X1 U12900 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2133] ), 
        .B1(n11749), .B2(n10901), .ZN(n5837) );
  AOI22_X1 U12901 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2134] ), 
        .B1(n11791), .B2(n10901), .ZN(n5836) );
  AOI22_X1 U12902 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2135] ), 
        .B1(n11750), .B2(n10901), .ZN(n5835) );
  AOI22_X1 U12903 ( .A1(\DataPath/RF/bus_reg_dataout[2136] ), .A2(n10902), 
        .B1(n10900), .B2(n11766), .ZN(n5834) );
  AOI22_X1 U12904 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2137] ), 
        .B1(n11794), .B2(n10901), .ZN(n5833) );
  AOI22_X1 U12905 ( .A1(\DataPath/RF/bus_reg_dataout[2138] ), .A2(n10902), 
        .B1(n10900), .B2(n11795), .ZN(n5832) );
  AOI22_X1 U12906 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2139] ), 
        .B1(n11796), .B2(n10901), .ZN(n5831) );
  AOI22_X1 U12907 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2140] ), 
        .B1(n11752), .B2(n10901), .ZN(n5830) );
  AOI22_X1 U12908 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2141] ), 
        .B1(n11753), .B2(n10901), .ZN(n5829) );
  AOI22_X1 U12909 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2142] ), 
        .B1(n11754), .B2(n10901), .ZN(n5828) );
  AOI22_X1 U12910 ( .A1(n10902), .A2(\DataPath/RF/bus_reg_dataout[2143] ), 
        .B1(n11803), .B2(n10901), .ZN(n5825) );
  INV_X1 U12911 ( .A(n10903), .ZN(n10904) );
  NAND2_X1 U12912 ( .A1(n10909), .A2(n11477), .ZN(n11407) );
  NAND2_X1 U12913 ( .A1(n10910), .A2(n11477), .ZN(n11406) );
  OAI22_X1 U12914 ( .A1(n8293), .A2(n11407), .B1(n8450), .B2(n11406), .ZN(
        n10905) );
  AOI22_X1 U12915 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2080] ), 
        .B1(n11804), .B2(n10906), .ZN(n5822) );
  AOI22_X1 U12916 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2081] ), 
        .B1(n11805), .B2(n10906), .ZN(n5821) );
  AOI22_X1 U12917 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2082] ), 
        .B1(n11806), .B2(n10906), .ZN(n5820) );
  AOI22_X1 U12918 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2083] ), 
        .B1(n11807), .B2(n10906), .ZN(n5819) );
  AOI22_X1 U12919 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2084] ), 
        .B1(n11808), .B2(n10906), .ZN(n5818) );
  AOI22_X1 U12920 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2085] ), 
        .B1(n11809), .B2(n10906), .ZN(n5817) );
  AOI22_X1 U12921 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2086] ), 
        .B1(n11810), .B2(n10906), .ZN(n5816) );
  AOI22_X1 U12922 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2087] ), 
        .B1(n11811), .B2(n10906), .ZN(n5815) );
  AOI22_X1 U12923 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2088] ), 
        .B1(n11812), .B2(n10906), .ZN(n5814) );
  AOI22_X1 U12924 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2089] ), 
        .B1(n11813), .B2(n10906), .ZN(n5813) );
  AOI22_X1 U12925 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2090] ), 
        .B1(n11814), .B2(n10906), .ZN(n5812) );
  AOI22_X1 U12926 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2091] ), 
        .B1(n11815), .B2(n10906), .ZN(n5811) );
  AOI22_X1 U12927 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2092] ), 
        .B1(n11816), .B2(n10906), .ZN(n5810) );
  AOI22_X1 U12928 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2093] ), 
        .B1(n11817), .B2(n10906), .ZN(n5809) );
  AOI22_X1 U12929 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2094] ), 
        .B1(n11818), .B2(n10906), .ZN(n5808) );
  AOI22_X1 U12930 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2095] ), 
        .B1(n11819), .B2(n10906), .ZN(n5807) );
  AOI22_X1 U12931 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2096] ), 
        .B1(n11820), .B2(n10906), .ZN(n5806) );
  AOI22_X1 U12932 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2097] ), 
        .B1(n11823), .B2(n10906), .ZN(n5805) );
  AOI22_X1 U12933 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2098] ), 
        .B1(n11746), .B2(n10906), .ZN(n5804) );
  AOI22_X1 U12934 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2099] ), 
        .B1(n11747), .B2(n10906), .ZN(n5803) );
  AOI22_X1 U12935 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2100] ), 
        .B1(n11748), .B2(n10906), .ZN(n5802) );
  AOI22_X1 U12936 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2101] ), 
        .B1(n11749), .B2(n10906), .ZN(n5801) );
  AOI22_X1 U12937 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2102] ), 
        .B1(n11791), .B2(n10906), .ZN(n5800) );
  AOI22_X1 U12938 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2103] ), 
        .B1(n11750), .B2(n10906), .ZN(n5799) );
  AOI22_X1 U12939 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2104] ), 
        .B1(n11793), .B2(n10906), .ZN(n5798) );
  AOI22_X1 U12940 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2105] ), 
        .B1(n11794), .B2(n10906), .ZN(n5797) );
  AOI22_X1 U12941 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2106] ), 
        .B1(n11751), .B2(n10906), .ZN(n5796) );
  AOI22_X1 U12942 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2107] ), 
        .B1(n11796), .B2(n10906), .ZN(n5795) );
  AOI22_X1 U12943 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2108] ), 
        .B1(n11752), .B2(n10906), .ZN(n5794) );
  AOI22_X1 U12944 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2109] ), 
        .B1(n11753), .B2(n10906), .ZN(n5793) );
  AOI22_X1 U12945 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2110] ), 
        .B1(n11754), .B2(n10906), .ZN(n5792) );
  AOI22_X1 U12946 ( .A1(n10907), .A2(\DataPath/RF/bus_reg_dataout[2111] ), 
        .B1(n11803), .B2(n10906), .ZN(n5789) );
  NAND2_X1 U12947 ( .A1(n10911), .A2(n10909), .ZN(n11416) );
  NAND2_X1 U12948 ( .A1(n10911), .A2(n10910), .ZN(n11414) );
  OAI22_X1 U12949 ( .A1(n8293), .A2(n11416), .B1(n8450), .B2(n11414), .ZN(
        n10912) );
  AOI22_X1 U12950 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2048] ), 
        .B1(n11804), .B2(n10913), .ZN(n5783) );
  AOI22_X1 U12951 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2049] ), 
        .B1(n11805), .B2(n10913), .ZN(n5782) );
  AOI22_X1 U12952 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2050] ), 
        .B1(n11806), .B2(n10913), .ZN(n5781) );
  AOI22_X1 U12953 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2051] ), 
        .B1(n11807), .B2(n10913), .ZN(n5780) );
  AOI22_X1 U12954 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2052] ), 
        .B1(n11808), .B2(n10913), .ZN(n5779) );
  AOI22_X1 U12955 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2053] ), 
        .B1(n11809), .B2(n10913), .ZN(n5778) );
  AOI22_X1 U12956 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2054] ), 
        .B1(n11810), .B2(n10913), .ZN(n5777) );
  AOI22_X1 U12957 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2055] ), 
        .B1(n11811), .B2(n10913), .ZN(n5776) );
  AOI22_X1 U12958 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2056] ), 
        .B1(n11812), .B2(n10913), .ZN(n5775) );
  AOI22_X1 U12959 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2057] ), 
        .B1(n11813), .B2(n10913), .ZN(n5774) );
  AOI22_X1 U12960 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2058] ), 
        .B1(n11814), .B2(n10913), .ZN(n5773) );
  AOI22_X1 U12961 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2059] ), 
        .B1(n11815), .B2(n10913), .ZN(n5772) );
  AOI22_X1 U12962 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2060] ), 
        .B1(n11816), .B2(n10913), .ZN(n5771) );
  AOI22_X1 U12963 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2061] ), 
        .B1(n11817), .B2(n10913), .ZN(n5770) );
  AOI22_X1 U12964 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2062] ), 
        .B1(n11818), .B2(n10913), .ZN(n5769) );
  AOI22_X1 U12965 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2063] ), 
        .B1(n11819), .B2(n10913), .ZN(n5768) );
  AOI22_X1 U12966 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2064] ), 
        .B1(n11820), .B2(n10913), .ZN(n5767) );
  AOI22_X1 U12967 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2065] ), 
        .B1(n11823), .B2(n10913), .ZN(n5766) );
  AOI22_X1 U12968 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2066] ), 
        .B1(n11746), .B2(n10913), .ZN(n5765) );
  AOI22_X1 U12969 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2067] ), 
        .B1(n11747), .B2(n10913), .ZN(n5764) );
  AOI22_X1 U12970 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2068] ), 
        .B1(n11748), .B2(n10913), .ZN(n5763) );
  AOI22_X1 U12971 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2069] ), 
        .B1(n11749), .B2(n10913), .ZN(n5762) );
  AOI22_X1 U12972 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2070] ), 
        .B1(n11791), .B2(n10913), .ZN(n5761) );
  AOI22_X1 U12973 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2071] ), 
        .B1(n11750), .B2(n10913), .ZN(n5760) );
  AOI22_X1 U12974 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2072] ), 
        .B1(n11793), .B2(n10913), .ZN(n5759) );
  AOI22_X1 U12975 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2073] ), 
        .B1(n11794), .B2(n10913), .ZN(n5758) );
  AOI22_X1 U12976 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2074] ), 
        .B1(n11751), .B2(n10913), .ZN(n5757) );
  AOI22_X1 U12977 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2075] ), 
        .B1(n11796), .B2(n10913), .ZN(n5756) );
  AOI22_X1 U12978 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2076] ), 
        .B1(n11752), .B2(n10913), .ZN(n5755) );
  AOI22_X1 U12979 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2077] ), 
        .B1(n11753), .B2(n10913), .ZN(n5754) );
  AOI22_X1 U12980 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2078] ), 
        .B1(n11754), .B2(n10913), .ZN(n5753) );
  AOI22_X1 U12981 ( .A1(n10914), .A2(\DataPath/RF/bus_reg_dataout[2079] ), 
        .B1(n11803), .B2(n10913), .ZN(n5750) );
  OAI22_X1 U12982 ( .A1(n10999), .A2(n11272), .B1(n11479), .B2(n11003), .ZN(
        n10956) );
  NAND2_X1 U12983 ( .A1(n10932), .A2(n11452), .ZN(n11737) );
  INV_X1 U12984 ( .A(n10915), .ZN(n11660) );
  OAI22_X1 U12985 ( .A1(n11004), .A2(n10918), .B1(
        \DataPath/RF/bus_reg_dataout[2016] ), .B2(n8362), .ZN(n5746) );
  OAI22_X1 U12986 ( .A1(n10999), .A2(n11273), .B1(n11480), .B2(n11003), .ZN(
        n10980) );
  OAI22_X1 U12987 ( .A1(n10918), .A2(n11005), .B1(
        \DataPath/RF/bus_reg_dataout[2017] ), .B2(n10917), .ZN(n5745) );
  OAI22_X1 U12988 ( .A1(n10999), .A2(n11274), .B1(n11481), .B2(n11003), .ZN(
        n10981) );
  OAI22_X1 U12989 ( .A1(n10918), .A2(n11006), .B1(
        \DataPath/RF/bus_reg_dataout[2018] ), .B2(n8362), .ZN(n5744) );
  OAI22_X1 U12990 ( .A1(n10999), .A2(n11275), .B1(n11482), .B2(n11003), .ZN(
        n10957) );
  OAI22_X1 U12991 ( .A1(n8363), .A2(n11007), .B1(
        \DataPath/RF/bus_reg_dataout[2019] ), .B2(n8362), .ZN(n5743) );
  OAI22_X1 U12992 ( .A1(n10999), .A2(n11276), .B1(n11483), .B2(n11003), .ZN(
        n10958) );
  AOI22_X1 U12993 ( .A1(\DataPath/RF/bus_reg_dataout[2020] ), .A2(n8363), .B1(
        n11008), .B2(n8362), .ZN(n5742) );
  OAI22_X1 U12994 ( .A1(n10999), .A2(n11277), .B1(n11484), .B2(n11003), .ZN(
        n10959) );
  OAI22_X1 U12995 ( .A1(n8363), .A2(n11009), .B1(
        \DataPath/RF/bus_reg_dataout[2021] ), .B2(n8362), .ZN(n5741) );
  OAI22_X1 U12996 ( .A1(n10999), .A2(n11278), .B1(n11485), .B2(n11003), .ZN(
        n10989) );
  OAI22_X1 U12997 ( .A1(n8363), .A2(n11010), .B1(
        \DataPath/RF/bus_reg_dataout[2022] ), .B2(n10917), .ZN(n5740) );
  OAI22_X1 U12998 ( .A1(n10999), .A2(n11279), .B1(n11486), .B2(n11003), .ZN(
        n10960) );
  OAI22_X1 U12999 ( .A1(n8363), .A2(n11011), .B1(
        \DataPath/RF/bus_reg_dataout[2023] ), .B2(n10917), .ZN(n5739) );
  OAI22_X1 U13000 ( .A1(n10999), .A2(n11280), .B1(n11487), .B2(n11003), .ZN(
        n10961) );
  OAI22_X1 U13001 ( .A1(n8363), .A2(n11012), .B1(
        \DataPath/RF/bus_reg_dataout[2024] ), .B2(n8362), .ZN(n5738) );
  OAI22_X1 U13002 ( .A1(n10999), .A2(n11281), .B1(n11488), .B2(n11003), .ZN(
        n10982) );
  OAI22_X1 U13003 ( .A1(n8363), .A2(n11013), .B1(
        \DataPath/RF/bus_reg_dataout[2025] ), .B2(n8362), .ZN(n5737) );
  OAI22_X1 U13004 ( .A1(n10999), .A2(n11282), .B1(n11489), .B2(n11003), .ZN(
        n10962) );
  OAI22_X1 U13005 ( .A1(n10918), .A2(n11014), .B1(
        \DataPath/RF/bus_reg_dataout[2026] ), .B2(n8362), .ZN(n5736) );
  OAI22_X1 U13006 ( .A1(n10999), .A2(n11283), .B1(n11490), .B2(n11003), .ZN(
        n10963) );
  OAI22_X1 U13007 ( .A1(n10918), .A2(n11015), .B1(
        \DataPath/RF/bus_reg_dataout[2027] ), .B2(n10917), .ZN(n5735) );
  OAI22_X1 U13008 ( .A1(n10999), .A2(n11284), .B1(n11491), .B2(n11003), .ZN(
        n10964) );
  AOI22_X1 U13009 ( .A1(\DataPath/RF/bus_reg_dataout[2028] ), .A2(n8363), .B1(
        n11016), .B2(n8362), .ZN(n5734) );
  OAI22_X1 U13010 ( .A1(n10999), .A2(n11285), .B1(n11492), .B2(n11003), .ZN(
        n10965) );
  OAI22_X1 U13011 ( .A1(n10918), .A2(n11017), .B1(
        \DataPath/RF/bus_reg_dataout[2029] ), .B2(n8362), .ZN(n5733) );
  OAI22_X1 U13012 ( .A1(n10999), .A2(n11286), .B1(n11493), .B2(n11003), .ZN(
        n10990) );
  OAI22_X1 U13013 ( .A1(n8363), .A2(n11018), .B1(
        \DataPath/RF/bus_reg_dataout[2030] ), .B2(n8362), .ZN(n5732) );
  OAI22_X1 U13014 ( .A1(n10999), .A2(n11287), .B1(n11494), .B2(n11003), .ZN(
        n10991) );
  OAI22_X1 U13015 ( .A1(n8363), .A2(n11019), .B1(
        \DataPath/RF/bus_reg_dataout[2031] ), .B2(n8362), .ZN(n5731) );
  OAI22_X1 U13016 ( .A1(n10999), .A2(n11288), .B1(n11495), .B2(n11003), .ZN(
        n10966) );
  OAI22_X1 U13017 ( .A1(n8363), .A2(n11020), .B1(
        \DataPath/RF/bus_reg_dataout[2032] ), .B2(n10917), .ZN(n5730) );
  OAI22_X1 U13018 ( .A1(n10999), .A2(n11289), .B1(n11496), .B2(n11003), .ZN(
        n10967) );
  OAI22_X1 U13019 ( .A1(n8363), .A2(n11021), .B1(
        \DataPath/RF/bus_reg_dataout[2033] ), .B2(n10917), .ZN(n5729) );
  OAI22_X1 U13020 ( .A1(n10999), .A2(n11290), .B1(n11497), .B2(n11003), .ZN(
        n10968) );
  AOI22_X1 U13021 ( .A1(\DataPath/RF/bus_reg_dataout[2034] ), .A2(n8363), .B1(
        n11022), .B2(n8362), .ZN(n5728) );
  OAI22_X1 U13022 ( .A1(n10999), .A2(n11291), .B1(n11498), .B2(n11003), .ZN(
        n10983) );
  OAI22_X1 U13023 ( .A1(n8363), .A2(n11023), .B1(
        \DataPath/RF/bus_reg_dataout[2035] ), .B2(n8362), .ZN(n5727) );
  OAI22_X1 U13024 ( .A1(n10999), .A2(n11292), .B1(n11499), .B2(n11003), .ZN(
        n10969) );
  OAI22_X1 U13025 ( .A1(n8363), .A2(n11024), .B1(
        \DataPath/RF/bus_reg_dataout[2036] ), .B2(n8362), .ZN(n5726) );
  OAI22_X1 U13026 ( .A1(n10999), .A2(n11293), .B1(n11500), .B2(n11003), .ZN(
        n10970) );
  OAI22_X1 U13027 ( .A1(n10918), .A2(n11025), .B1(
        \DataPath/RF/bus_reg_dataout[2037] ), .B2(n8362), .ZN(n5725) );
  OAI22_X1 U13028 ( .A1(n10999), .A2(n11294), .B1(n11501), .B2(n11003), .ZN(
        n10984) );
  OAI22_X1 U13029 ( .A1(n10918), .A2(n11026), .B1(
        \DataPath/RF/bus_reg_dataout[2038] ), .B2(n10917), .ZN(n5724) );
  OAI22_X1 U13030 ( .A1(n10999), .A2(n11295), .B1(n11502), .B2(n11003), .ZN(
        n10971) );
  OAI22_X1 U13031 ( .A1(n10918), .A2(n11027), .B1(
        \DataPath/RF/bus_reg_dataout[2039] ), .B2(n8362), .ZN(n5723) );
  OAI22_X1 U13032 ( .A1(n10999), .A2(n11296), .B1(n11503), .B2(n11003), .ZN(
        n10972) );
  OAI22_X1 U13033 ( .A1(n8363), .A2(n11028), .B1(
        \DataPath/RF/bus_reg_dataout[2040] ), .B2(n8362), .ZN(n5722) );
  OAI22_X1 U13034 ( .A1(n10999), .A2(n11297), .B1(n11504), .B2(n11003), .ZN(
        n10985) );
  OAI22_X1 U13035 ( .A1(n8363), .A2(n11029), .B1(
        \DataPath/RF/bus_reg_dataout[2041] ), .B2(n8362), .ZN(n5721) );
  OAI22_X1 U13036 ( .A1(n10999), .A2(n11298), .B1(n11505), .B2(n11003), .ZN(
        n10992) );
  OAI22_X1 U13037 ( .A1(n8363), .A2(n11030), .B1(
        \DataPath/RF/bus_reg_dataout[2042] ), .B2(n10917), .ZN(n5720) );
  OAI22_X1 U13038 ( .A1(n10999), .A2(n11299), .B1(n11506), .B2(n11003), .ZN(
        n10974) );
  OAI22_X1 U13039 ( .A1(n8363), .A2(n11031), .B1(
        \DataPath/RF/bus_reg_dataout[2043] ), .B2(n10917), .ZN(n5719) );
  OAI22_X1 U13040 ( .A1(n10999), .A2(n11300), .B1(n11507), .B2(n11003), .ZN(
        n10993) );
  OAI22_X1 U13041 ( .A1(n8363), .A2(n11032), .B1(
        \DataPath/RF/bus_reg_dataout[2044] ), .B2(n8362), .ZN(n5718) );
  OAI22_X1 U13042 ( .A1(n10999), .A2(n11301), .B1(n11508), .B2(n11003), .ZN(
        n10975) );
  OAI22_X1 U13043 ( .A1(n8363), .A2(n11033), .B1(
        \DataPath/RF/bus_reg_dataout[2045] ), .B2(n8362), .ZN(n5717) );
  OAI22_X1 U13044 ( .A1(n10999), .A2(n11302), .B1(n11509), .B2(n11003), .ZN(
        n10976) );
  OAI22_X1 U13045 ( .A1(n8363), .A2(n11034), .B1(
        \DataPath/RF/bus_reg_dataout[2046] ), .B2(n8362), .ZN(n5716) );
  OAI22_X1 U13046 ( .A1(n10999), .A2(n11304), .B1(n11512), .B2(n11003), .ZN(
        n10995) );
  OAI22_X1 U13047 ( .A1(n10918), .A2(n11036), .B1(
        \DataPath/RF/bus_reg_dataout[2047] ), .B2(n8362), .ZN(n5713) );
  NAND2_X1 U13048 ( .A1(n10932), .A2(n11456), .ZN(n11741) );
  INV_X1 U13049 ( .A(n10919), .ZN(n10920) );
  AOI22_X1 U13050 ( .A1(\DataPath/RF/bus_reg_dataout[1984] ), .A2(n8364), .B1(
        n10922), .B2(n10956), .ZN(n5709) );
  AOI22_X1 U13051 ( .A1(\DataPath/RF/bus_reg_dataout[1985] ), .A2(n8364), .B1(
        n10922), .B2(n10980), .ZN(n5708) );
  AOI22_X1 U13052 ( .A1(\DataPath/RF/bus_reg_dataout[1986] ), .A2(n8364), .B1(
        n10922), .B2(n10981), .ZN(n5707) );
  AOI22_X1 U13053 ( .A1(\DataPath/RF/bus_reg_dataout[1987] ), .A2(n10923), 
        .B1(n10922), .B2(n10957), .ZN(n5706) );
  AOI22_X1 U13054 ( .A1(\DataPath/RF/bus_reg_dataout[1988] ), .A2(n10923), 
        .B1(n10922), .B2(n10958), .ZN(n5705) );
  AOI22_X1 U13055 ( .A1(\DataPath/RF/bus_reg_dataout[1989] ), .A2(n8364), .B1(
        n10922), .B2(n10959), .ZN(n5704) );
  AOI22_X1 U13056 ( .A1(\DataPath/RF/bus_reg_dataout[1990] ), .A2(n8364), .B1(
        n10922), .B2(n10989), .ZN(n5703) );
  AOI22_X1 U13057 ( .A1(\DataPath/RF/bus_reg_dataout[1991] ), .A2(n8364), .B1(
        n10922), .B2(n10960), .ZN(n5702) );
  AOI22_X1 U13058 ( .A1(\DataPath/RF/bus_reg_dataout[1992] ), .A2(n10923), 
        .B1(n10922), .B2(n10961), .ZN(n5701) );
  AOI22_X1 U13059 ( .A1(\DataPath/RF/bus_reg_dataout[1993] ), .A2(n8364), .B1(
        n10922), .B2(n10982), .ZN(n5700) );
  AOI22_X1 U13060 ( .A1(\DataPath/RF/bus_reg_dataout[1994] ), .A2(n8364), .B1(
        n10922), .B2(n10962), .ZN(n5699) );
  AOI22_X1 U13061 ( .A1(\DataPath/RF/bus_reg_dataout[1995] ), .A2(n8364), .B1(
        n10922), .B2(n10963), .ZN(n5698) );
  AOI22_X1 U13062 ( .A1(n11016), .A2(n10921), .B1(n8364), .B2(
        \DataPath/RF/bus_reg_dataout[1996] ), .ZN(n5697) );
  AOI22_X1 U13063 ( .A1(\DataPath/RF/bus_reg_dataout[1997] ), .A2(n10923), 
        .B1(n10922), .B2(n10965), .ZN(n5696) );
  AOI22_X1 U13064 ( .A1(\DataPath/RF/bus_reg_dataout[1998] ), .A2(n8364), .B1(
        n10922), .B2(n10990), .ZN(n5695) );
  AOI22_X1 U13065 ( .A1(n11019), .A2(n10921), .B1(n8364), .B2(
        \DataPath/RF/bus_reg_dataout[1999] ), .ZN(n5694) );
  AOI22_X1 U13066 ( .A1(\DataPath/RF/bus_reg_dataout[2000] ), .A2(n8364), .B1(
        n10922), .B2(n10966), .ZN(n5693) );
  AOI22_X1 U13067 ( .A1(\DataPath/RF/bus_reg_dataout[2001] ), .A2(n10923), 
        .B1(n10922), .B2(n10967), .ZN(n5692) );
  AOI22_X1 U13068 ( .A1(\DataPath/RF/bus_reg_dataout[2002] ), .A2(n8364), .B1(
        n10922), .B2(n10968), .ZN(n5691) );
  AOI22_X1 U13069 ( .A1(\DataPath/RF/bus_reg_dataout[2003] ), .A2(n10923), 
        .B1(n10922), .B2(n10983), .ZN(n5690) );
  AOI22_X1 U13070 ( .A1(\DataPath/RF/bus_reg_dataout[2004] ), .A2(n8364), .B1(
        n10922), .B2(n10969), .ZN(n5689) );
  AOI22_X1 U13071 ( .A1(n11025), .A2(n10921), .B1(n10923), .B2(
        \DataPath/RF/bus_reg_dataout[2005] ), .ZN(n5688) );
  AOI22_X1 U13072 ( .A1(n11026), .A2(n10921), .B1(n10923), .B2(
        \DataPath/RF/bus_reg_dataout[2006] ), .ZN(n5687) );
  AOI22_X1 U13073 ( .A1(\DataPath/RF/bus_reg_dataout[2007] ), .A2(n8364), .B1(
        n10922), .B2(n10971), .ZN(n5686) );
  AOI22_X1 U13074 ( .A1(n11028), .A2(n10921), .B1(n8364), .B2(
        \DataPath/RF/bus_reg_dataout[2008] ), .ZN(n5685) );
  AOI22_X1 U13075 ( .A1(\DataPath/RF/bus_reg_dataout[2009] ), .A2(n8364), .B1(
        n10922), .B2(n10985), .ZN(n5684) );
  AOI22_X1 U13076 ( .A1(n11030), .A2(n10921), .B1(n8364), .B2(
        \DataPath/RF/bus_reg_dataout[2010] ), .ZN(n5683) );
  AOI22_X1 U13077 ( .A1(n11031), .A2(n10921), .B1(n8364), .B2(
        \DataPath/RF/bus_reg_dataout[2011] ), .ZN(n5682) );
  AOI22_X1 U13078 ( .A1(\DataPath/RF/bus_reg_dataout[2012] ), .A2(n8364), .B1(
        n10922), .B2(n10993), .ZN(n5681) );
  AOI22_X1 U13079 ( .A1(\DataPath/RF/bus_reg_dataout[2013] ), .A2(n8364), .B1(
        n10922), .B2(n10975), .ZN(n5680) );
  AOI22_X1 U13080 ( .A1(n11034), .A2(n10921), .B1(n10923), .B2(
        \DataPath/RF/bus_reg_dataout[2014] ), .ZN(n5679) );
  AOI22_X1 U13081 ( .A1(\DataPath/RF/bus_reg_dataout[2015] ), .A2(n10923), 
        .B1(n10922), .B2(n10995), .ZN(n5676) );
  NAND2_X1 U13082 ( .A1(n10932), .A2(n11460), .ZN(n11745) );
  INV_X1 U13083 ( .A(n10924), .ZN(n10925) );
  OAI22_X1 U13084 ( .A1(n11004), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1952] ), .B2(n8365), .ZN(n5672) );
  OAI22_X1 U13085 ( .A1(n11005), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1953] ), .B2(n10926), .ZN(n5671) );
  OAI22_X1 U13086 ( .A1(n11006), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1954] ), .B2(n8365), .ZN(n5670) );
  OAI22_X1 U13087 ( .A1(n11007), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1955] ), .B2(n10926), .ZN(n5669) );
  OAI22_X1 U13088 ( .A1(n11008), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1956] ), .B2(n8365), .ZN(n5668) );
  OAI22_X1 U13089 ( .A1(n11009), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1957] ), .B2(n10926), .ZN(n5667) );
  OAI22_X1 U13090 ( .A1(n11010), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1958] ), .B2(n8365), .ZN(n5666) );
  OAI22_X1 U13091 ( .A1(n11011), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1959] ), .B2(n8365), .ZN(n5665) );
  OAI22_X1 U13092 ( .A1(n11012), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1960] ), .B2(n8365), .ZN(n5664) );
  OAI22_X1 U13093 ( .A1(n11013), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1961] ), .B2(n8365), .ZN(n5663) );
  OAI22_X1 U13094 ( .A1(n11014), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1962] ), .B2(n10926), .ZN(n5662) );
  OAI22_X1 U13095 ( .A1(n11015), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1963] ), .B2(n8365), .ZN(n5661) );
  OAI22_X1 U13096 ( .A1(n11016), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1964] ), .B2(n10926), .ZN(n5660) );
  OAI22_X1 U13097 ( .A1(n11017), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1965] ), .B2(n8365), .ZN(n5659) );
  OAI22_X1 U13098 ( .A1(n11018), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1966] ), .B2(n10926), .ZN(n5658) );
  OAI22_X1 U13099 ( .A1(n11019), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1967] ), .B2(n8365), .ZN(n5657) );
  OAI22_X1 U13100 ( .A1(n11020), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1968] ), .B2(n8365), .ZN(n5656) );
  OAI22_X1 U13101 ( .A1(n11021), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1969] ), .B2(n8365), .ZN(n5655) );
  AOI22_X1 U13102 ( .A1(n11022), .A2(n8365), .B1(n8366), .B2(
        \DataPath/RF/bus_reg_dataout[1970] ), .ZN(n5654) );
  OAI22_X1 U13103 ( .A1(n11023), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1971] ), .B2(n8365), .ZN(n5653) );
  OAI22_X1 U13104 ( .A1(n11024), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1972] ), .B2(n10926), .ZN(n5652) );
  OAI22_X1 U13105 ( .A1(n11025), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1973] ), .B2(n8365), .ZN(n5651) );
  OAI22_X1 U13106 ( .A1(n11026), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1974] ), .B2(n10926), .ZN(n5650) );
  OAI22_X1 U13107 ( .A1(n11027), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1975] ), .B2(n8365), .ZN(n5649) );
  OAI22_X1 U13108 ( .A1(n11028), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1976] ), .B2(n8365), .ZN(n5648) );
  OAI22_X1 U13109 ( .A1(n11029), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1977] ), .B2(n8365), .ZN(n5647) );
  OAI22_X1 U13110 ( .A1(n11030), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1978] ), .B2(n8365), .ZN(n5646) );
  OAI22_X1 U13111 ( .A1(n11031), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1979] ), .B2(n8365), .ZN(n5645) );
  OAI22_X1 U13112 ( .A1(n11032), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1980] ), .B2(n8365), .ZN(n5644) );
  OAI22_X1 U13113 ( .A1(n11033), .A2(n8366), .B1(
        \DataPath/RF/bus_reg_dataout[1981] ), .B2(n8365), .ZN(n5643) );
  AOI22_X1 U13114 ( .A1(n11034), .A2(n8365), .B1(n8366), .B2(
        \DataPath/RF/bus_reg_dataout[1982] ), .ZN(n5642) );
  OAI22_X1 U13115 ( .A1(n11036), .A2(n10927), .B1(
        \DataPath/RF/bus_reg_dataout[1983] ), .B2(n10926), .ZN(n5639) );
  NAND2_X1 U13116 ( .A1(n10932), .A2(n11464), .ZN(n11758) );
  INV_X1 U13117 ( .A(n10928), .ZN(n10929) );
  AOI22_X1 U13118 ( .A1(n11004), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1920] ), .ZN(n5635) );
  AOI22_X1 U13119 ( .A1(n11005), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1921] ), .ZN(n5634) );
  AOI22_X1 U13120 ( .A1(n11006), .A2(n10931), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1922] ), .ZN(n5633) );
  AOI22_X1 U13121 ( .A1(n11007), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1923] ), .ZN(n5632) );
  AOI22_X1 U13122 ( .A1(n11008), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1924] ), .ZN(n5631) );
  AOI22_X1 U13123 ( .A1(n11009), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1925] ), .ZN(n5630) );
  AOI22_X1 U13124 ( .A1(n11010), .A2(n10931), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1926] ), .ZN(n5629) );
  AOI22_X1 U13125 ( .A1(n11011), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1927] ), .ZN(n5628) );
  AOI22_X1 U13126 ( .A1(n11012), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1928] ), .ZN(n5627) );
  AOI22_X1 U13127 ( .A1(n11013), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1929] ), .ZN(n5626) );
  AOI22_X1 U13128 ( .A1(n11014), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1930] ), .ZN(n5625) );
  AOI22_X1 U13129 ( .A1(n11015), .A2(n10931), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1931] ), .ZN(n5624) );
  AOI22_X1 U13130 ( .A1(n11016), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1932] ), .ZN(n5623) );
  AOI22_X1 U13131 ( .A1(n11017), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1933] ), .ZN(n5622) );
  AOI22_X1 U13132 ( .A1(n11018), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1934] ), .ZN(n5621) );
  AOI22_X1 U13133 ( .A1(n11019), .A2(n10931), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1935] ), .ZN(n5620) );
  AOI22_X1 U13134 ( .A1(n11020), .A2(n10931), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1936] ), .ZN(n5619) );
  AOI22_X1 U13135 ( .A1(n11021), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1937] ), .ZN(n5618) );
  OAI22_X1 U13136 ( .A1(n11022), .A2(n8368), .B1(
        \DataPath/RF/bus_reg_dataout[1938] ), .B2(n8367), .ZN(n5617) );
  AOI22_X1 U13137 ( .A1(n11023), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1939] ), .ZN(n5616) );
  AOI22_X1 U13138 ( .A1(n11024), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1940] ), .ZN(n5615) );
  AOI22_X1 U13139 ( .A1(n11025), .A2(n10931), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1941] ), .ZN(n5614) );
  AOI22_X1 U13140 ( .A1(n11026), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1942] ), .ZN(n5613) );
  AOI22_X1 U13141 ( .A1(n11027), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1943] ), .ZN(n5612) );
  AOI22_X1 U13142 ( .A1(n11028), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1944] ), .ZN(n5611) );
  AOI22_X1 U13143 ( .A1(n11029), .A2(n10931), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1945] ), .ZN(n5610) );
  AOI22_X1 U13144 ( .A1(n11030), .A2(n10931), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1946] ), .ZN(n5609) );
  AOI22_X1 U13145 ( .A1(n11031), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1947] ), .ZN(n5608) );
  AOI22_X1 U13146 ( .A1(n11032), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1948] ), .ZN(n5607) );
  AOI22_X1 U13147 ( .A1(n11033), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1949] ), .ZN(n5606) );
  AOI22_X1 U13148 ( .A1(n11034), .A2(n8367), .B1(n8368), .B2(
        \DataPath/RF/bus_reg_dataout[1950] ), .ZN(n5605) );
  AOI22_X1 U13149 ( .A1(n11036), .A2(n8367), .B1(n10930), .B2(
        \DataPath/RF/bus_reg_dataout[1951] ), .ZN(n5602) );
  NAND2_X1 U13150 ( .A1(n10932), .A2(n11468), .ZN(n11773) );
  INV_X1 U13151 ( .A(n10933), .ZN(n10935) );
  AOI22_X1 U13152 ( .A1(\DataPath/RF/bus_reg_dataout[1888] ), .A2(n8369), .B1(
        n10937), .B2(n10956), .ZN(n5596) );
  AOI22_X1 U13153 ( .A1(\DataPath/RF/bus_reg_dataout[1889] ), .A2(n8369), .B1(
        n10937), .B2(n10980), .ZN(n5595) );
  AOI22_X1 U13154 ( .A1(\DataPath/RF/bus_reg_dataout[1890] ), .A2(n8369), .B1(
        n10937), .B2(n10981), .ZN(n5594) );
  AOI22_X1 U13155 ( .A1(\DataPath/RF/bus_reg_dataout[1891] ), .A2(n8369), .B1(
        n10937), .B2(n10957), .ZN(n5593) );
  AOI22_X1 U13156 ( .A1(\DataPath/RF/bus_reg_dataout[1892] ), .A2(n10938), 
        .B1(n10937), .B2(n10958), .ZN(n5592) );
  AOI22_X1 U13157 ( .A1(\DataPath/RF/bus_reg_dataout[1893] ), .A2(n8369), .B1(
        n10937), .B2(n10959), .ZN(n5591) );
  AOI22_X1 U13158 ( .A1(n11010), .A2(n10936), .B1(n8369), .B2(
        \DataPath/RF/bus_reg_dataout[1894] ), .ZN(n5590) );
  AOI22_X1 U13159 ( .A1(\DataPath/RF/bus_reg_dataout[1895] ), .A2(n10938), 
        .B1(n10937), .B2(n10960), .ZN(n5589) );
  AOI22_X1 U13160 ( .A1(\DataPath/RF/bus_reg_dataout[1896] ), .A2(n8369), .B1(
        n10937), .B2(n10961), .ZN(n5588) );
  AOI22_X1 U13161 ( .A1(n11013), .A2(n10936), .B1(n8369), .B2(
        \DataPath/RF/bus_reg_dataout[1897] ), .ZN(n5587) );
  AOI22_X1 U13162 ( .A1(\DataPath/RF/bus_reg_dataout[1898] ), .A2(n10938), 
        .B1(n10937), .B2(n10962), .ZN(n5586) );
  AOI22_X1 U13163 ( .A1(\DataPath/RF/bus_reg_dataout[1899] ), .A2(n8369), .B1(
        n10937), .B2(n10963), .ZN(n5585) );
  AOI22_X1 U13164 ( .A1(\DataPath/RF/bus_reg_dataout[1900] ), .A2(n8369), .B1(
        n10937), .B2(n10964), .ZN(n5584) );
  AOI22_X1 U13165 ( .A1(\DataPath/RF/bus_reg_dataout[1901] ), .A2(n8369), .B1(
        n10937), .B2(n10965), .ZN(n5583) );
  AOI22_X1 U13166 ( .A1(\DataPath/RF/bus_reg_dataout[1902] ), .A2(n8369), .B1(
        n10937), .B2(n10990), .ZN(n5582) );
  AOI22_X1 U13167 ( .A1(\DataPath/RF/bus_reg_dataout[1903] ), .A2(n10938), 
        .B1(n10937), .B2(n10991), .ZN(n5581) );
  AOI22_X1 U13168 ( .A1(n11020), .A2(n10936), .B1(n10938), .B2(
        \DataPath/RF/bus_reg_dataout[1904] ), .ZN(n5580) );
  AOI22_X1 U13169 ( .A1(\DataPath/RF/bus_reg_dataout[1905] ), .A2(n8369), .B1(
        n10937), .B2(n10967), .ZN(n5579) );
  AOI22_X1 U13170 ( .A1(\DataPath/RF/bus_reg_dataout[1906] ), .A2(n8369), .B1(
        n10937), .B2(n10968), .ZN(n5578) );
  AOI22_X1 U13171 ( .A1(\DataPath/RF/bus_reg_dataout[1907] ), .A2(n8369), .B1(
        n10937), .B2(n10983), .ZN(n5577) );
  AOI22_X1 U13172 ( .A1(\DataPath/RF/bus_reg_dataout[1908] ), .A2(n10938), 
        .B1(n10937), .B2(n10969), .ZN(n5576) );
  AOI22_X1 U13173 ( .A1(n11025), .A2(n10936), .B1(n8369), .B2(
        \DataPath/RF/bus_reg_dataout[1909] ), .ZN(n5575) );
  AOI22_X1 U13174 ( .A1(\DataPath/RF/bus_reg_dataout[1910] ), .A2(n10938), 
        .B1(n10937), .B2(n10984), .ZN(n5574) );
  AOI22_X1 U13175 ( .A1(\DataPath/RF/bus_reg_dataout[1911] ), .A2(n8369), .B1(
        n10937), .B2(n10971), .ZN(n5573) );
  AOI22_X1 U13176 ( .A1(n11028), .A2(n10936), .B1(n10938), .B2(
        \DataPath/RF/bus_reg_dataout[1912] ), .ZN(n5572) );
  AOI22_X1 U13177 ( .A1(n11029), .A2(n10936), .B1(n8369), .B2(
        \DataPath/RF/bus_reg_dataout[1913] ), .ZN(n5571) );
  AOI22_X1 U13178 ( .A1(\DataPath/RF/bus_reg_dataout[1914] ), .A2(n10938), 
        .B1(n10937), .B2(n10992), .ZN(n5570) );
  AOI22_X1 U13179 ( .A1(\DataPath/RF/bus_reg_dataout[1915] ), .A2(n8369), .B1(
        n10937), .B2(n10974), .ZN(n5569) );
  AOI22_X1 U13180 ( .A1(\DataPath/RF/bus_reg_dataout[1916] ), .A2(n8369), .B1(
        n10937), .B2(n10993), .ZN(n5568) );
  AOI22_X1 U13181 ( .A1(n11033), .A2(n10936), .B1(n10938), .B2(
        \DataPath/RF/bus_reg_dataout[1917] ), .ZN(n5567) );
  AOI22_X1 U13182 ( .A1(\DataPath/RF/bus_reg_dataout[1918] ), .A2(n8369), .B1(
        n10937), .B2(n10976), .ZN(n5566) );
  AOI22_X1 U13183 ( .A1(\DataPath/RF/bus_reg_dataout[1919] ), .A2(n8369), .B1(
        n10937), .B2(n10995), .ZN(n5563) );
  OAI22_X1 U13184 ( .A1(n8293), .A2(n11322), .B1(n11321), .B2(n10999), .ZN(
        n10939) );
  AOI22_X1 U13185 ( .A1(\DataPath/RF/bus_reg_dataout[1856] ), .A2(n8370), .B1(
        n10940), .B2(n10956), .ZN(n5561) );
  AOI22_X1 U13186 ( .A1(\DataPath/RF/bus_reg_dataout[1857] ), .A2(n8370), .B1(
        n10940), .B2(n10980), .ZN(n5560) );
  AOI22_X1 U13187 ( .A1(\DataPath/RF/bus_reg_dataout[1858] ), .A2(n8370), .B1(
        n10940), .B2(n10981), .ZN(n5559) );
  AOI22_X1 U13188 ( .A1(\DataPath/RF/bus_reg_dataout[1859] ), .A2(n10941), 
        .B1(n10940), .B2(n10957), .ZN(n5558) );
  AOI22_X1 U13189 ( .A1(\DataPath/RF/bus_reg_dataout[1860] ), .A2(n8370), .B1(
        n10940), .B2(n10958), .ZN(n5557) );
  AOI22_X1 U13190 ( .A1(\DataPath/RF/bus_reg_dataout[1861] ), .A2(n10941), 
        .B1(n10940), .B2(n10959), .ZN(n5556) );
  AOI22_X1 U13191 ( .A1(\DataPath/RF/bus_reg_dataout[1862] ), .A2(n8370), .B1(
        n10940), .B2(n10989), .ZN(n5555) );
  AOI22_X1 U13192 ( .A1(\DataPath/RF/bus_reg_dataout[1863] ), .A2(n10941), 
        .B1(n10940), .B2(n10960), .ZN(n5554) );
  AOI22_X1 U13193 ( .A1(\DataPath/RF/bus_reg_dataout[1864] ), .A2(n8370), .B1(
        n10940), .B2(n10961), .ZN(n5553) );
  AOI22_X1 U13194 ( .A1(\DataPath/RF/bus_reg_dataout[1865] ), .A2(n8370), .B1(
        n10940), .B2(n10982), .ZN(n5552) );
  AOI22_X1 U13195 ( .A1(\DataPath/RF/bus_reg_dataout[1866] ), .A2(n8370), .B1(
        n10940), .B2(n10962), .ZN(n5551) );
  AOI22_X1 U13196 ( .A1(\DataPath/RF/bus_reg_dataout[1867] ), .A2(n8370), .B1(
        n10940), .B2(n10963), .ZN(n5550) );
  AOI22_X1 U13197 ( .A1(\DataPath/RF/bus_reg_dataout[1868] ), .A2(n10941), 
        .B1(n10940), .B2(n10964), .ZN(n5549) );
  AOI22_X1 U13198 ( .A1(\DataPath/RF/bus_reg_dataout[1869] ), .A2(n8370), .B1(
        n10940), .B2(n10965), .ZN(n5548) );
  AOI22_X1 U13199 ( .A1(\DataPath/RF/bus_reg_dataout[1870] ), .A2(n8370), .B1(
        n10940), .B2(n10990), .ZN(n5547) );
  AOI22_X1 U13200 ( .A1(\DataPath/RF/bus_reg_dataout[1871] ), .A2(n8370), .B1(
        n10940), .B2(n10991), .ZN(n5546) );
  AOI22_X1 U13201 ( .A1(\DataPath/RF/bus_reg_dataout[1872] ), .A2(n10941), 
        .B1(n10940), .B2(n10966), .ZN(n5545) );
  AOI22_X1 U13202 ( .A1(\DataPath/RF/bus_reg_dataout[1873] ), .A2(n10941), 
        .B1(n10940), .B2(n10967), .ZN(n5544) );
  AOI22_X1 U13203 ( .A1(\DataPath/RF/bus_reg_dataout[1874] ), .A2(n8370), .B1(
        n10940), .B2(n10968), .ZN(n5543) );
  AOI22_X1 U13204 ( .A1(\DataPath/RF/bus_reg_dataout[1875] ), .A2(n8370), .B1(
        n10940), .B2(n10983), .ZN(n5542) );
  AOI22_X1 U13205 ( .A1(\DataPath/RF/bus_reg_dataout[1876] ), .A2(n8370), .B1(
        n10940), .B2(n10969), .ZN(n5541) );
  AOI22_X1 U13206 ( .A1(\DataPath/RF/bus_reg_dataout[1877] ), .A2(n10941), 
        .B1(n10940), .B2(n10970), .ZN(n5540) );
  AOI22_X1 U13207 ( .A1(\DataPath/RF/bus_reg_dataout[1878] ), .A2(n8370), .B1(
        n10940), .B2(n10984), .ZN(n5539) );
  AOI22_X1 U13208 ( .A1(\DataPath/RF/bus_reg_dataout[1879] ), .A2(n10941), 
        .B1(n10940), .B2(n10971), .ZN(n5538) );
  AOI22_X1 U13209 ( .A1(\DataPath/RF/bus_reg_dataout[1880] ), .A2(n8370), .B1(
        n10940), .B2(n10972), .ZN(n5537) );
  AOI22_X1 U13210 ( .A1(\DataPath/RF/bus_reg_dataout[1881] ), .A2(n8370), .B1(
        n10940), .B2(n10985), .ZN(n5536) );
  AOI22_X1 U13211 ( .A1(\DataPath/RF/bus_reg_dataout[1882] ), .A2(n8370), .B1(
        n10940), .B2(n10992), .ZN(n5535) );
  AOI22_X1 U13212 ( .A1(\DataPath/RF/bus_reg_dataout[1883] ), .A2(n8370), .B1(
        n10940), .B2(n10974), .ZN(n5534) );
  AOI22_X1 U13213 ( .A1(\DataPath/RF/bus_reg_dataout[1884] ), .A2(n8370), .B1(
        n10940), .B2(n10993), .ZN(n5533) );
  AOI22_X1 U13214 ( .A1(\DataPath/RF/bus_reg_dataout[1885] ), .A2(n8370), .B1(
        n10940), .B2(n10975), .ZN(n5532) );
  AOI22_X1 U13215 ( .A1(\DataPath/RF/bus_reg_dataout[1886] ), .A2(n10941), 
        .B1(n10940), .B2(n10976), .ZN(n5531) );
  AOI22_X1 U13216 ( .A1(\DataPath/RF/bus_reg_dataout[1887] ), .A2(n10941), 
        .B1(n10940), .B2(n10995), .ZN(n5528) );
  OAI22_X1 U13217 ( .A1(n8293), .A2(n11327), .B1(n11326), .B2(n10999), .ZN(
        n10942) );
  AOI22_X1 U13218 ( .A1(\DataPath/RF/bus_reg_dataout[1824] ), .A2(n8371), .B1(
        n10943), .B2(n10956), .ZN(n5526) );
  AOI22_X1 U13219 ( .A1(\DataPath/RF/bus_reg_dataout[1825] ), .A2(n8371), .B1(
        n10943), .B2(n10980), .ZN(n5525) );
  AOI22_X1 U13220 ( .A1(\DataPath/RF/bus_reg_dataout[1826] ), .A2(n8371), .B1(
        n10943), .B2(n10981), .ZN(n5524) );
  AOI22_X1 U13221 ( .A1(\DataPath/RF/bus_reg_dataout[1827] ), .A2(n10944), 
        .B1(n10943), .B2(n10957), .ZN(n5523) );
  AOI22_X1 U13222 ( .A1(\DataPath/RF/bus_reg_dataout[1828] ), .A2(n8371), .B1(
        n10943), .B2(n10958), .ZN(n5522) );
  AOI22_X1 U13223 ( .A1(\DataPath/RF/bus_reg_dataout[1829] ), .A2(n10944), 
        .B1(n10943), .B2(n10959), .ZN(n5521) );
  AOI22_X1 U13224 ( .A1(\DataPath/RF/bus_reg_dataout[1830] ), .A2(n8371), .B1(
        n10943), .B2(n10989), .ZN(n5520) );
  AOI22_X1 U13225 ( .A1(\DataPath/RF/bus_reg_dataout[1831] ), .A2(n10944), 
        .B1(n10943), .B2(n10960), .ZN(n5519) );
  AOI22_X1 U13226 ( .A1(\DataPath/RF/bus_reg_dataout[1832] ), .A2(n8371), .B1(
        n10943), .B2(n10961), .ZN(n5518) );
  AOI22_X1 U13227 ( .A1(\DataPath/RF/bus_reg_dataout[1833] ), .A2(n8371), .B1(
        n10943), .B2(n10982), .ZN(n5517) );
  AOI22_X1 U13228 ( .A1(\DataPath/RF/bus_reg_dataout[1834] ), .A2(n8371), .B1(
        n10943), .B2(n10962), .ZN(n5516) );
  AOI22_X1 U13229 ( .A1(\DataPath/RF/bus_reg_dataout[1835] ), .A2(n8371), .B1(
        n10943), .B2(n10963), .ZN(n5515) );
  AOI22_X1 U13230 ( .A1(\DataPath/RF/bus_reg_dataout[1836] ), .A2(n10944), 
        .B1(n10943), .B2(n10964), .ZN(n5514) );
  AOI22_X1 U13231 ( .A1(\DataPath/RF/bus_reg_dataout[1837] ), .A2(n8371), .B1(
        n10943), .B2(n10965), .ZN(n5513) );
  AOI22_X1 U13232 ( .A1(\DataPath/RF/bus_reg_dataout[1838] ), .A2(n8371), .B1(
        n10943), .B2(n10990), .ZN(n5512) );
  AOI22_X1 U13233 ( .A1(\DataPath/RF/bus_reg_dataout[1839] ), .A2(n8371), .B1(
        n10943), .B2(n10991), .ZN(n5511) );
  AOI22_X1 U13234 ( .A1(\DataPath/RF/bus_reg_dataout[1840] ), .A2(n10944), 
        .B1(n10943), .B2(n10966), .ZN(n5510) );
  AOI22_X1 U13235 ( .A1(\DataPath/RF/bus_reg_dataout[1841] ), .A2(n10944), 
        .B1(n10943), .B2(n10967), .ZN(n5509) );
  AOI22_X1 U13236 ( .A1(\DataPath/RF/bus_reg_dataout[1842] ), .A2(n8371), .B1(
        n10943), .B2(n10968), .ZN(n5508) );
  AOI22_X1 U13237 ( .A1(\DataPath/RF/bus_reg_dataout[1843] ), .A2(n8371), .B1(
        n10943), .B2(n10983), .ZN(n5507) );
  AOI22_X1 U13238 ( .A1(\DataPath/RF/bus_reg_dataout[1844] ), .A2(n8371), .B1(
        n10943), .B2(n10969), .ZN(n5506) );
  AOI22_X1 U13239 ( .A1(\DataPath/RF/bus_reg_dataout[1845] ), .A2(n10944), 
        .B1(n10943), .B2(n10970), .ZN(n5505) );
  AOI22_X1 U13240 ( .A1(\DataPath/RF/bus_reg_dataout[1846] ), .A2(n8371), .B1(
        n10943), .B2(n10984), .ZN(n5504) );
  AOI22_X1 U13241 ( .A1(\DataPath/RF/bus_reg_dataout[1847] ), .A2(n10944), 
        .B1(n10943), .B2(n10971), .ZN(n5503) );
  AOI22_X1 U13242 ( .A1(\DataPath/RF/bus_reg_dataout[1848] ), .A2(n8371), .B1(
        n10943), .B2(n10972), .ZN(n5502) );
  AOI22_X1 U13243 ( .A1(\DataPath/RF/bus_reg_dataout[1849] ), .A2(n8371), .B1(
        n10943), .B2(n10985), .ZN(n5501) );
  AOI22_X1 U13244 ( .A1(\DataPath/RF/bus_reg_dataout[1850] ), .A2(n8371), .B1(
        n10943), .B2(n10992), .ZN(n5500) );
  AOI22_X1 U13245 ( .A1(\DataPath/RF/bus_reg_dataout[1851] ), .A2(n8371), .B1(
        n10943), .B2(n10974), .ZN(n5499) );
  AOI22_X1 U13246 ( .A1(\DataPath/RF/bus_reg_dataout[1852] ), .A2(n8371), .B1(
        n10943), .B2(n10993), .ZN(n5498) );
  AOI22_X1 U13247 ( .A1(\DataPath/RF/bus_reg_dataout[1853] ), .A2(n8371), .B1(
        n10943), .B2(n10975), .ZN(n5497) );
  AOI22_X1 U13248 ( .A1(\DataPath/RF/bus_reg_dataout[1854] ), .A2(n10944), 
        .B1(n10943), .B2(n10976), .ZN(n5496) );
  AOI22_X1 U13249 ( .A1(\DataPath/RF/bus_reg_dataout[1855] ), .A2(n10944), 
        .B1(n10943), .B2(n10995), .ZN(n5493) );
  OAI22_X1 U13250 ( .A1(n11004), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1792] ), .B2(n8372), .ZN(n5491) );
  OAI22_X1 U13251 ( .A1(n11005), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1793] ), .B2(n8372), .ZN(n5490) );
  OAI22_X1 U13252 ( .A1(n11006), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1794] ), .B2(n10945), .ZN(n5489) );
  OAI22_X1 U13253 ( .A1(n11007), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1795] ), .B2(n10945), .ZN(n5488) );
  OAI22_X1 U13254 ( .A1(n11008), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1796] ), .B2(n8372), .ZN(n5487) );
  OAI22_X1 U13255 ( .A1(n11009), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1797] ), .B2(n8372), .ZN(n5486) );
  OAI22_X1 U13256 ( .A1(n11010), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1798] ), .B2(n8372), .ZN(n5485) );
  OAI22_X1 U13257 ( .A1(n11011), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1799] ), .B2(n10945), .ZN(n5484) );
  OAI22_X1 U13258 ( .A1(n11012), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1800] ), .B2(n8372), .ZN(n5483) );
  OAI22_X1 U13259 ( .A1(n11013), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1801] ), .B2(n8372), .ZN(n5482) );
  OAI22_X1 U13260 ( .A1(n11014), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1802] ), .B2(n8372), .ZN(n5481) );
  OAI22_X1 U13261 ( .A1(n11015), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1803] ), .B2(n10945), .ZN(n5480) );
  OAI22_X1 U13262 ( .A1(n11016), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1804] ), .B2(n10945), .ZN(n5479) );
  OAI22_X1 U13263 ( .A1(n11017), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1805] ), .B2(n8372), .ZN(n5478) );
  OAI22_X1 U13264 ( .A1(n11018), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1806] ), .B2(n8372), .ZN(n5477) );
  OAI22_X1 U13265 ( .A1(n11019), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1807] ), .B2(n8372), .ZN(n5476) );
  OAI22_X1 U13266 ( .A1(n11020), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1808] ), .B2(n10945), .ZN(n5475) );
  OAI22_X1 U13267 ( .A1(n11021), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1809] ), .B2(n8372), .ZN(n5474) );
  AOI22_X1 U13268 ( .A1(n11022), .A2(n8372), .B1(n8373), .B2(
        \DataPath/RF/bus_reg_dataout[1810] ), .ZN(n5473) );
  OAI22_X1 U13269 ( .A1(n11023), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1811] ), .B2(n8372), .ZN(n5472) );
  OAI22_X1 U13270 ( .A1(n11024), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1812] ), .B2(n8372), .ZN(n5471) );
  OAI22_X1 U13271 ( .A1(n11025), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1813] ), .B2(n10945), .ZN(n5470) );
  OAI22_X1 U13272 ( .A1(n11026), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1814] ), .B2(n10945), .ZN(n5469) );
  OAI22_X1 U13273 ( .A1(n11027), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1815] ), .B2(n8372), .ZN(n5468) );
  OAI22_X1 U13274 ( .A1(n11028), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1816] ), .B2(n8372), .ZN(n5467) );
  OAI22_X1 U13275 ( .A1(n11029), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1817] ), .B2(n8372), .ZN(n5466) );
  OAI22_X1 U13276 ( .A1(n11030), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1818] ), .B2(n10945), .ZN(n5465) );
  OAI22_X1 U13277 ( .A1(n11031), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1819] ), .B2(n8372), .ZN(n5464) );
  OAI22_X1 U13278 ( .A1(n11032), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1820] ), .B2(n8372), .ZN(n5463) );
  OAI22_X1 U13279 ( .A1(n11033), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1821] ), .B2(n8372), .ZN(n5462) );
  OAI22_X1 U13280 ( .A1(n11034), .A2(n10946), .B1(
        \DataPath/RF/bus_reg_dataout[1822] ), .B2(n8372), .ZN(n5461) );
  OAI22_X1 U13281 ( .A1(n11036), .A2(n8373), .B1(
        \DataPath/RF/bus_reg_dataout[1823] ), .B2(n8372), .ZN(n5458) );
  OAI22_X1 U13282 ( .A1(n8271), .A2(n11339), .B1(n8293), .B2(n11338), .ZN(
        n10947) );
  AOI22_X1 U13283 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1760] ), 
        .B1(n11004), .B2(n10948), .ZN(n5456) );
  AOI22_X1 U13284 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1761] ), 
        .B1(n11005), .B2(n10948), .ZN(n5455) );
  AOI22_X1 U13285 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1762] ), 
        .B1(n11006), .B2(n10948), .ZN(n5454) );
  AOI22_X1 U13286 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1763] ), 
        .B1(n11007), .B2(n10948), .ZN(n5453) );
  AOI22_X1 U13287 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1764] ), 
        .B1(n11008), .B2(n10948), .ZN(n5452) );
  AOI22_X1 U13288 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1765] ), 
        .B1(n11009), .B2(n10948), .ZN(n5451) );
  AOI22_X1 U13289 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1766] ), 
        .B1(n11010), .B2(n10948), .ZN(n5450) );
  AOI22_X1 U13290 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1767] ), 
        .B1(n11011), .B2(n10948), .ZN(n5449) );
  AOI22_X1 U13291 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1768] ), 
        .B1(n11012), .B2(n10948), .ZN(n5448) );
  AOI22_X1 U13292 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1769] ), 
        .B1(n11013), .B2(n10948), .ZN(n5447) );
  AOI22_X1 U13293 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1770] ), 
        .B1(n11014), .B2(n10948), .ZN(n5446) );
  AOI22_X1 U13294 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1771] ), 
        .B1(n11015), .B2(n10948), .ZN(n5445) );
  AOI22_X1 U13295 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1772] ), 
        .B1(n11016), .B2(n10948), .ZN(n5444) );
  AOI22_X1 U13296 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1773] ), 
        .B1(n11017), .B2(n10948), .ZN(n5443) );
  AOI22_X1 U13297 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1774] ), 
        .B1(n11018), .B2(n10948), .ZN(n5442) );
  AOI22_X1 U13298 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1775] ), 
        .B1(n11019), .B2(n10948), .ZN(n5441) );
  AOI22_X1 U13299 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1776] ), 
        .B1(n11020), .B2(n10948), .ZN(n5440) );
  AOI22_X1 U13300 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1777] ), 
        .B1(n11021), .B2(n10948), .ZN(n5439) );
  AOI22_X1 U13301 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1778] ), 
        .B1(n11022), .B2(n10948), .ZN(n5438) );
  AOI22_X1 U13302 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1779] ), 
        .B1(n11023), .B2(n10948), .ZN(n5437) );
  AOI22_X1 U13303 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1780] ), 
        .B1(n11024), .B2(n10948), .ZN(n5436) );
  AOI22_X1 U13304 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1781] ), 
        .B1(n11025), .B2(n10948), .ZN(n5435) );
  AOI22_X1 U13305 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1782] ), 
        .B1(n11026), .B2(n10948), .ZN(n5434) );
  AOI22_X1 U13306 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1783] ), 
        .B1(n11027), .B2(n10948), .ZN(n5433) );
  AOI22_X1 U13307 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1784] ), 
        .B1(n11028), .B2(n10948), .ZN(n5432) );
  AOI22_X1 U13308 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1785] ), 
        .B1(n11029), .B2(n10948), .ZN(n5431) );
  AOI22_X1 U13309 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1786] ), 
        .B1(n11030), .B2(n10948), .ZN(n5430) );
  AOI22_X1 U13310 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1787] ), 
        .B1(n11031), .B2(n10948), .ZN(n5429) );
  AOI22_X1 U13311 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1788] ), 
        .B1(n11032), .B2(n10948), .ZN(n5428) );
  AOI22_X1 U13312 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1789] ), 
        .B1(n11033), .B2(n10948), .ZN(n5427) );
  AOI22_X1 U13313 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1790] ), 
        .B1(n11034), .B2(n10948), .ZN(n5426) );
  AOI22_X1 U13314 ( .A1(n10949), .A2(\DataPath/RF/bus_reg_dataout[1791] ), 
        .B1(n11036), .B2(n10948), .ZN(n5423) );
  OAI22_X1 U13315 ( .A1(n8271), .A2(n11346), .B1(n11345), .B2(n10999), .ZN(
        n10950) );
  AOI22_X1 U13316 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1728] ), .B1(
        n11004), .B2(n7754), .ZN(n5421) );
  AOI22_X1 U13317 ( .A1(\DataPath/RF/bus_reg_dataout[1729] ), .A2(n8262), .B1(
        n10951), .B2(n10980), .ZN(n5420) );
  AOI22_X1 U13318 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1730] ), .B1(
        n11006), .B2(n7754), .ZN(n5419) );
  AOI22_X1 U13319 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1731] ), .B1(
        n11007), .B2(n7754), .ZN(n5418) );
  AOI22_X1 U13320 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1732] ), .B1(
        n11008), .B2(n7754), .ZN(n5417) );
  AOI22_X1 U13321 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1733] ), .B1(
        n11009), .B2(n7754), .ZN(n5416) );
  AOI22_X1 U13322 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1734] ), .B1(
        n11010), .B2(n7754), .ZN(n5415) );
  AOI22_X1 U13323 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1735] ), .B1(
        n11011), .B2(n7754), .ZN(n5414) );
  AOI22_X1 U13324 ( .A1(\DataPath/RF/bus_reg_dataout[1736] ), .A2(n8262), .B1(
        n10951), .B2(n10961), .ZN(n5413) );
  AOI22_X1 U13325 ( .A1(\DataPath/RF/bus_reg_dataout[1737] ), .A2(n8262), .B1(
        n10951), .B2(n10982), .ZN(n5412) );
  AOI22_X1 U13326 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1738] ), .B1(
        n11014), .B2(n7754), .ZN(n5411) );
  AOI22_X1 U13327 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1739] ), .B1(
        n11015), .B2(n7754), .ZN(n5410) );
  AOI22_X1 U13328 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1740] ), .B1(
        n11016), .B2(n7754), .ZN(n5409) );
  AOI22_X1 U13329 ( .A1(\DataPath/RF/bus_reg_dataout[1741] ), .A2(n8262), .B1(
        n10951), .B2(n10965), .ZN(n5408) );
  AOI22_X1 U13330 ( .A1(n8263), .A2(\DataPath/RF/bus_reg_dataout[1742] ), .B1(
        n11018), .B2(n7754), .ZN(n5407) );
  AOI22_X1 U13331 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1743] ), .B1(
        n11019), .B2(n7754), .ZN(n5406) );
  AOI22_X1 U13332 ( .A1(\DataPath/RF/bus_reg_dataout[1744] ), .A2(n8262), .B1(
        n10951), .B2(n10966), .ZN(n5405) );
  AOI22_X1 U13333 ( .A1(\DataPath/RF/bus_reg_dataout[1745] ), .A2(n8262), .B1(
        n10951), .B2(n10967), .ZN(n5404) );
  AOI22_X1 U13334 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1746] ), .B1(
        n11022), .B2(n7754), .ZN(n5403) );
  AOI22_X1 U13335 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1747] ), .B1(
        n11023), .B2(n7754), .ZN(n5402) );
  AOI22_X1 U13336 ( .A1(\DataPath/RF/bus_reg_dataout[1748] ), .A2(n8262), .B1(
        n10951), .B2(n10969), .ZN(n5401) );
  AOI22_X1 U13337 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1749] ), .B1(
        n11025), .B2(n7754), .ZN(n5400) );
  AOI22_X1 U13338 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1750] ), .B1(
        n11026), .B2(n7754), .ZN(n5399) );
  AOI22_X1 U13339 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1751] ), .B1(
        n11027), .B2(n7754), .ZN(n5398) );
  AOI22_X1 U13340 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1752] ), .B1(
        n11028), .B2(n7754), .ZN(n5397) );
  AOI22_X1 U13341 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1753] ), .B1(
        n11029), .B2(n7754), .ZN(n5396) );
  AOI22_X1 U13342 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1754] ), .B1(
        n11030), .B2(n7754), .ZN(n5395) );
  AOI22_X1 U13343 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1755] ), .B1(
        n11031), .B2(n7754), .ZN(n5394) );
  AOI22_X1 U13344 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1756] ), .B1(
        n11032), .B2(n7754), .ZN(n5393) );
  AOI22_X1 U13345 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1757] ), .B1(
        n11033), .B2(n7754), .ZN(n5392) );
  AOI22_X1 U13346 ( .A1(n8262), .A2(\DataPath/RF/bus_reg_dataout[1758] ), .B1(
        n11034), .B2(n7754), .ZN(n5391) );
  AOI22_X1 U13347 ( .A1(\DataPath/RF/bus_reg_dataout[1759] ), .A2(n8262), .B1(
        n10951), .B2(n10995), .ZN(n5388) );
  OAI22_X1 U13348 ( .A1(n8271), .A2(n11353), .B1(n11352), .B2(n10999), .ZN(
        n10953) );
  AOI22_X1 U13349 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1696] ), .B1(
        n11004), .B2(n8266), .ZN(n5386) );
  AOI22_X1 U13350 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1697] ), .B1(
        n11005), .B2(n8266), .ZN(n5385) );
  AOI22_X1 U13351 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1698] ), .B1(
        n11006), .B2(n8266), .ZN(n5384) );
  AOI22_X1 U13352 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1699] ), .B1(
        n11007), .B2(n8266), .ZN(n5383) );
  NOR2_X1 U13353 ( .A1(RST), .A2(n8265), .ZN(n10954) );
  AOI22_X1 U13354 ( .A1(\DataPath/RF/bus_reg_dataout[1700] ), .A2(n8264), .B1(
        n10954), .B2(n10958), .ZN(n5382) );
  AOI22_X1 U13355 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1701] ), .B1(
        n11009), .B2(n8266), .ZN(n5381) );
  AOI22_X1 U13356 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1702] ), .B1(
        n11010), .B2(n8266), .ZN(n5380) );
  AOI22_X1 U13357 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1703] ), .B1(
        n11011), .B2(n8266), .ZN(n5379) );
  AOI22_X1 U13358 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1704] ), .B1(
        n11012), .B2(n8266), .ZN(n5378) );
  AOI22_X1 U13359 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1705] ), .B1(
        n11013), .B2(n8266), .ZN(n5377) );
  AOI22_X1 U13360 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1706] ), .B1(
        n11014), .B2(n8266), .ZN(n5376) );
  AOI22_X1 U13361 ( .A1(n8265), .A2(\DataPath/RF/bus_reg_dataout[1707] ), .B1(
        n11015), .B2(n8266), .ZN(n5375) );
  AOI22_X1 U13362 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1708] ), .B1(
        n11016), .B2(n8266), .ZN(n5374) );
  AOI22_X1 U13363 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1709] ), .B1(
        n11017), .B2(n8266), .ZN(n5373) );
  AOI22_X1 U13364 ( .A1(\DataPath/RF/bus_reg_dataout[1710] ), .A2(n8264), .B1(
        n10954), .B2(n10990), .ZN(n5372) );
  AOI22_X1 U13365 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1711] ), .B1(
        n11019), .B2(n8266), .ZN(n5371) );
  AOI22_X1 U13366 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1712] ), .B1(
        n11020), .B2(n8266), .ZN(n5370) );
  AOI22_X1 U13367 ( .A1(\DataPath/RF/bus_reg_dataout[1713] ), .A2(n8264), .B1(
        n10954), .B2(n10967), .ZN(n5369) );
  AOI22_X1 U13368 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1714] ), .B1(
        n11022), .B2(n8266), .ZN(n5368) );
  AOI22_X1 U13369 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1715] ), .B1(
        n11023), .B2(n8266), .ZN(n5367) );
  AOI22_X1 U13370 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1716] ), .B1(
        n11024), .B2(n8266), .ZN(n5366) );
  AOI22_X1 U13371 ( .A1(\DataPath/RF/bus_reg_dataout[1717] ), .A2(n8264), .B1(
        n10954), .B2(n10970), .ZN(n5365) );
  AOI22_X1 U13372 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1718] ), .B1(
        n11026), .B2(n8266), .ZN(n5364) );
  AOI22_X1 U13373 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1719] ), .B1(
        n11027), .B2(n8266), .ZN(n5363) );
  AOI22_X1 U13374 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1720] ), .B1(
        n11028), .B2(n8266), .ZN(n5362) );
  AOI22_X1 U13375 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1721] ), .B1(
        n11029), .B2(n8266), .ZN(n5361) );
  AOI22_X1 U13376 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1722] ), .B1(
        n11030), .B2(n8266), .ZN(n5360) );
  AOI22_X1 U13377 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1723] ), .B1(
        n11031), .B2(n8266), .ZN(n5359) );
  AOI22_X1 U13378 ( .A1(\DataPath/RF/bus_reg_dataout[1724] ), .A2(n8264), .B1(
        n10954), .B2(n10993), .ZN(n5358) );
  AOI22_X1 U13379 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1725] ), .B1(
        n11033), .B2(n8266), .ZN(n5357) );
  AOI22_X1 U13380 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1726] ), .B1(
        n11034), .B2(n8266), .ZN(n5356) );
  AOI22_X1 U13381 ( .A1(n8264), .A2(\DataPath/RF/bus_reg_dataout[1727] ), .B1(
        n11036), .B2(n8266), .ZN(n5353) );
  OAI222_X1 U13382 ( .A1(n10999), .A2(n11361), .B1(n11360), .B2(n8271), .C1(
        n11359), .C2(n8293), .ZN(n10973) );
  AOI22_X1 U13383 ( .A1(\DataPath/RF/bus_reg_dataout[1664] ), .A2(n8374), .B1(
        n10977), .B2(n10956), .ZN(n5351) );
  AOI22_X1 U13384 ( .A1(\DataPath/RF/bus_reg_dataout[1665] ), .A2(n10978), 
        .B1(n10977), .B2(n10980), .ZN(n5350) );
  AOI22_X1 U13385 ( .A1(\DataPath/RF/bus_reg_dataout[1666] ), .A2(n8374), .B1(
        n10977), .B2(n10981), .ZN(n5349) );
  AOI22_X1 U13386 ( .A1(\DataPath/RF/bus_reg_dataout[1667] ), .A2(n8374), .B1(
        n10977), .B2(n10957), .ZN(n5348) );
  AOI22_X1 U13387 ( .A1(\DataPath/RF/bus_reg_dataout[1668] ), .A2(n10978), 
        .B1(n10977), .B2(n10958), .ZN(n5347) );
  AOI22_X1 U13388 ( .A1(\DataPath/RF/bus_reg_dataout[1669] ), .A2(n8374), .B1(
        n10977), .B2(n10959), .ZN(n5346) );
  AOI22_X1 U13389 ( .A1(\DataPath/RF/bus_reg_dataout[1670] ), .A2(n8374), .B1(
        n10977), .B2(n10989), .ZN(n5345) );
  AOI22_X1 U13390 ( .A1(\DataPath/RF/bus_reg_dataout[1671] ), .A2(n8374), .B1(
        n10977), .B2(n10960), .ZN(n5344) );
  AOI22_X1 U13391 ( .A1(\DataPath/RF/bus_reg_dataout[1672] ), .A2(n8374), .B1(
        n10977), .B2(n10961), .ZN(n5343) );
  AOI22_X1 U13392 ( .A1(\DataPath/RF/bus_reg_dataout[1673] ), .A2(n8374), .B1(
        n10977), .B2(n10982), .ZN(n5342) );
  AOI22_X1 U13393 ( .A1(\DataPath/RF/bus_reg_dataout[1674] ), .A2(n8374), .B1(
        n10977), .B2(n10962), .ZN(n5341) );
  AOI22_X1 U13394 ( .A1(\DataPath/RF/bus_reg_dataout[1675] ), .A2(n10978), 
        .B1(n10977), .B2(n10963), .ZN(n5340) );
  AOI22_X1 U13395 ( .A1(\DataPath/RF/bus_reg_dataout[1676] ), .A2(n8374), .B1(
        n10977), .B2(n10964), .ZN(n5339) );
  AOI22_X1 U13396 ( .A1(\DataPath/RF/bus_reg_dataout[1677] ), .A2(n8374), .B1(
        n10977), .B2(n10965), .ZN(n5338) );
  AOI22_X1 U13397 ( .A1(\DataPath/RF/bus_reg_dataout[1678] ), .A2(n8374), .B1(
        n10977), .B2(n10990), .ZN(n5337) );
  AOI22_X1 U13398 ( .A1(\DataPath/RF/bus_reg_dataout[1679] ), .A2(n10978), 
        .B1(n10977), .B2(n10991), .ZN(n5336) );
  AOI22_X1 U13399 ( .A1(\DataPath/RF/bus_reg_dataout[1680] ), .A2(n8374), .B1(
        n10977), .B2(n10966), .ZN(n5335) );
  AOI22_X1 U13400 ( .A1(\DataPath/RF/bus_reg_dataout[1681] ), .A2(n10978), 
        .B1(n10977), .B2(n10967), .ZN(n5334) );
  AOI22_X1 U13401 ( .A1(\DataPath/RF/bus_reg_dataout[1682] ), .A2(n8374), .B1(
        n10977), .B2(n10968), .ZN(n5333) );
  AOI22_X1 U13402 ( .A1(\DataPath/RF/bus_reg_dataout[1683] ), .A2(n10978), 
        .B1(n10977), .B2(n10983), .ZN(n5332) );
  AOI22_X1 U13403 ( .A1(\DataPath/RF/bus_reg_dataout[1684] ), .A2(n8374), .B1(
        n10977), .B2(n10969), .ZN(n5331) );
  AOI22_X1 U13404 ( .A1(\DataPath/RF/bus_reg_dataout[1685] ), .A2(n8374), .B1(
        n10977), .B2(n10970), .ZN(n5330) );
  AOI22_X1 U13405 ( .A1(\DataPath/RF/bus_reg_dataout[1686] ), .A2(n10978), 
        .B1(n10977), .B2(n10984), .ZN(n5329) );
  AOI22_X1 U13406 ( .A1(\DataPath/RF/bus_reg_dataout[1687] ), .A2(n8374), .B1(
        n10977), .B2(n10971), .ZN(n5328) );
  AOI22_X1 U13407 ( .A1(\DataPath/RF/bus_reg_dataout[1688] ), .A2(n10978), 
        .B1(n10977), .B2(n10972), .ZN(n5327) );
  AOI22_X1 U13408 ( .A1(\DataPath/RF/bus_reg_dataout[1689] ), .A2(n8374), .B1(
        n10977), .B2(n10985), .ZN(n5326) );
  AOI22_X1 U13409 ( .A1(n11030), .A2(n10973), .B1(n8374), .B2(
        \DataPath/RF/bus_reg_dataout[1690] ), .ZN(n5325) );
  AOI22_X1 U13410 ( .A1(\DataPath/RF/bus_reg_dataout[1691] ), .A2(n8374), .B1(
        n10977), .B2(n10974), .ZN(n5324) );
  AOI22_X1 U13411 ( .A1(\DataPath/RF/bus_reg_dataout[1692] ), .A2(n8374), .B1(
        n10977), .B2(n10993), .ZN(n5323) );
  AOI22_X1 U13412 ( .A1(\DataPath/RF/bus_reg_dataout[1693] ), .A2(n8374), .B1(
        n10977), .B2(n10975), .ZN(n5322) );
  AOI22_X1 U13413 ( .A1(\DataPath/RF/bus_reg_dataout[1694] ), .A2(n10978), 
        .B1(n10977), .B2(n10976), .ZN(n5321) );
  AOI22_X1 U13414 ( .A1(\DataPath/RF/bus_reg_dataout[1695] ), .A2(n10978), 
        .B1(n10977), .B2(n10995), .ZN(n5318) );
  OAI22_X1 U13415 ( .A1(n8271), .A2(n11367), .B1(n11366), .B2(n10999), .ZN(
        n10979) );
  AOI22_X1 U13416 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1632] ), .B1(
        n11004), .B2(n7755), .ZN(n5316) );
  AOI22_X1 U13417 ( .A1(\DataPath/RF/bus_reg_dataout[1633] ), .A2(n8267), .B1(
        n10986), .B2(n10980), .ZN(n5315) );
  AOI22_X1 U13418 ( .A1(\DataPath/RF/bus_reg_dataout[1634] ), .A2(n8267), .B1(
        n10986), .B2(n10981), .ZN(n5314) );
  AOI22_X1 U13419 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1635] ), .B1(
        n11007), .B2(n7755), .ZN(n5313) );
  AOI22_X1 U13420 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1636] ), .B1(
        n11008), .B2(n7755), .ZN(n5312) );
  AOI22_X1 U13421 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1637] ), .B1(
        n11009), .B2(n7755), .ZN(n5311) );
  AOI22_X1 U13422 ( .A1(\DataPath/RF/bus_reg_dataout[1638] ), .A2(n8267), .B1(
        n10986), .B2(n10989), .ZN(n5310) );
  AOI22_X1 U13423 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1639] ), .B1(
        n11011), .B2(n7755), .ZN(n5309) );
  AOI22_X1 U13424 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1640] ), .B1(
        n11012), .B2(n7755), .ZN(n5308) );
  AOI22_X1 U13425 ( .A1(\DataPath/RF/bus_reg_dataout[1641] ), .A2(n8267), .B1(
        n10986), .B2(n10982), .ZN(n5307) );
  AOI22_X1 U13426 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1642] ), .B1(
        n11014), .B2(n7755), .ZN(n5306) );
  AOI22_X1 U13427 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1643] ), .B1(
        n11015), .B2(n7755), .ZN(n5305) );
  AOI22_X1 U13428 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1644] ), .B1(
        n11016), .B2(n7755), .ZN(n5304) );
  AOI22_X1 U13429 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1645] ), .B1(
        n11017), .B2(n7755), .ZN(n5303) );
  AOI22_X1 U13430 ( .A1(n8268), .A2(\DataPath/RF/bus_reg_dataout[1646] ), .B1(
        n11018), .B2(n7755), .ZN(n5302) );
  AOI22_X1 U13431 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1647] ), .B1(
        n11019), .B2(n7755), .ZN(n5301) );
  AOI22_X1 U13432 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1648] ), .B1(
        n11020), .B2(n7755), .ZN(n5300) );
  AOI22_X1 U13433 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1649] ), .B1(
        n11021), .B2(n7755), .ZN(n5299) );
  AOI22_X1 U13434 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1650] ), .B1(
        n11022), .B2(n7755), .ZN(n5298) );
  AOI22_X1 U13435 ( .A1(\DataPath/RF/bus_reg_dataout[1651] ), .A2(n8267), .B1(
        n10986), .B2(n10983), .ZN(n5297) );
  AOI22_X1 U13436 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1652] ), .B1(
        n11024), .B2(n7755), .ZN(n5296) );
  AOI22_X1 U13437 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1653] ), .B1(
        n11025), .B2(n7755), .ZN(n5295) );
  AOI22_X1 U13438 ( .A1(\DataPath/RF/bus_reg_dataout[1654] ), .A2(n8267), .B1(
        n10986), .B2(n10984), .ZN(n5294) );
  AOI22_X1 U13439 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1655] ), .B1(
        n11027), .B2(n7755), .ZN(n5293) );
  AOI22_X1 U13440 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1656] ), .B1(
        n11028), .B2(n7755), .ZN(n5292) );
  AOI22_X1 U13441 ( .A1(\DataPath/RF/bus_reg_dataout[1657] ), .A2(n8267), .B1(
        n10986), .B2(n10985), .ZN(n5291) );
  AOI22_X1 U13442 ( .A1(\DataPath/RF/bus_reg_dataout[1658] ), .A2(n8267), .B1(
        n10986), .B2(n10992), .ZN(n5290) );
  AOI22_X1 U13443 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1659] ), .B1(
        n11031), .B2(n7755), .ZN(n5289) );
  AOI22_X1 U13444 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1660] ), .B1(
        n11032), .B2(n7755), .ZN(n5288) );
  AOI22_X1 U13445 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1661] ), .B1(
        n11033), .B2(n7755), .ZN(n5287) );
  AOI22_X1 U13446 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1662] ), .B1(
        n11034), .B2(n7755), .ZN(n5286) );
  AOI22_X1 U13447 ( .A1(n8267), .A2(\DataPath/RF/bus_reg_dataout[1663] ), .B1(
        n11036), .B2(n7755), .ZN(n5283) );
  OAI22_X1 U13448 ( .A1(n8271), .A2(n11375), .B1(n8293), .B2(n11374), .ZN(
        n10988) );
  AOI22_X1 U13449 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1600] ), 
        .B1(n11004), .B2(n10994), .ZN(n5281) );
  AOI22_X1 U13450 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1601] ), 
        .B1(n11005), .B2(n10994), .ZN(n5280) );
  AOI22_X1 U13451 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1602] ), 
        .B1(n11006), .B2(n10994), .ZN(n5279) );
  AOI22_X1 U13452 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1603] ), 
        .B1(n11007), .B2(n10994), .ZN(n5278) );
  AOI22_X1 U13453 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1604] ), 
        .B1(n11008), .B2(n10994), .ZN(n5277) );
  AOI22_X1 U13454 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1605] ), 
        .B1(n11009), .B2(n10994), .ZN(n5276) );
  NOR2_X1 U13455 ( .A1(RST), .A2(n10997), .ZN(n10996) );
  AOI22_X1 U13456 ( .A1(\DataPath/RF/bus_reg_dataout[1606] ), .A2(n10997), 
        .B1(n10996), .B2(n10989), .ZN(n5275) );
  AOI22_X1 U13457 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1607] ), 
        .B1(n11011), .B2(n10994), .ZN(n5274) );
  AOI22_X1 U13458 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1608] ), 
        .B1(n11012), .B2(n10994), .ZN(n5273) );
  AOI22_X1 U13459 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1609] ), 
        .B1(n11013), .B2(n10994), .ZN(n5272) );
  AOI22_X1 U13460 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1610] ), 
        .B1(n11014), .B2(n10994), .ZN(n5271) );
  AOI22_X1 U13461 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1611] ), 
        .B1(n11015), .B2(n10994), .ZN(n5270) );
  AOI22_X1 U13462 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1612] ), 
        .B1(n11016), .B2(n10994), .ZN(n5269) );
  AOI22_X1 U13463 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1613] ), 
        .B1(n11017), .B2(n10994), .ZN(n5268) );
  AOI22_X1 U13464 ( .A1(\DataPath/RF/bus_reg_dataout[1614] ), .A2(n10997), 
        .B1(n10996), .B2(n10990), .ZN(n5267) );
  AOI22_X1 U13465 ( .A1(\DataPath/RF/bus_reg_dataout[1615] ), .A2(n10997), 
        .B1(n10996), .B2(n10991), .ZN(n5266) );
  AOI22_X1 U13466 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1616] ), 
        .B1(n11020), .B2(n10994), .ZN(n5265) );
  AOI22_X1 U13467 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1617] ), 
        .B1(n11021), .B2(n10994), .ZN(n5264) );
  AOI22_X1 U13468 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1618] ), 
        .B1(n11022), .B2(n10994), .ZN(n5263) );
  AOI22_X1 U13469 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1619] ), 
        .B1(n11023), .B2(n10994), .ZN(n5262) );
  AOI22_X1 U13470 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1620] ), 
        .B1(n11024), .B2(n10994), .ZN(n5261) );
  AOI22_X1 U13471 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1621] ), 
        .B1(n11025), .B2(n10994), .ZN(n5260) );
  AOI22_X1 U13472 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1622] ), 
        .B1(n11026), .B2(n10994), .ZN(n5259) );
  AOI22_X1 U13473 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1623] ), 
        .B1(n11027), .B2(n10994), .ZN(n5258) );
  AOI22_X1 U13474 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1624] ), 
        .B1(n11028), .B2(n10994), .ZN(n5257) );
  AOI22_X1 U13475 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1625] ), 
        .B1(n11029), .B2(n10994), .ZN(n5256) );
  AOI22_X1 U13476 ( .A1(\DataPath/RF/bus_reg_dataout[1626] ), .A2(n10997), 
        .B1(n10996), .B2(n10992), .ZN(n5255) );
  AOI22_X1 U13477 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1627] ), 
        .B1(n11031), .B2(n10994), .ZN(n5254) );
  AOI22_X1 U13478 ( .A1(\DataPath/RF/bus_reg_dataout[1628] ), .A2(n10997), 
        .B1(n10996), .B2(n10993), .ZN(n5253) );
  AOI22_X1 U13479 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1629] ), 
        .B1(n11033), .B2(n10994), .ZN(n5252) );
  AOI22_X1 U13480 ( .A1(n10997), .A2(\DataPath/RF/bus_reg_dataout[1630] ), 
        .B1(n11034), .B2(n10994), .ZN(n5251) );
  AOI22_X1 U13481 ( .A1(\DataPath/RF/bus_reg_dataout[1631] ), .A2(n10997), 
        .B1(n10996), .B2(n10995), .ZN(n5248) );
  AOI22_X1 U13482 ( .A1(n11004), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1568] ), .ZN(n5245) );
  OAI22_X1 U13483 ( .A1(n11005), .A2(n11000), .B1(
        \DataPath/RF/bus_reg_dataout[1569] ), .B2(n8269), .ZN(n5244) );
  AOI22_X1 U13484 ( .A1(n11006), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1570] ), .ZN(n5243) );
  AOI22_X1 U13485 ( .A1(n11007), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1571] ), .ZN(n5242) );
  AOI22_X1 U13486 ( .A1(n11008), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1572] ), .ZN(n5241) );
  AOI22_X1 U13487 ( .A1(n11009), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1573] ), .ZN(n5240) );
  AOI22_X1 U13488 ( .A1(n11010), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1574] ), .ZN(n5239) );
  AOI22_X1 U13489 ( .A1(n11011), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1575] ), .ZN(n5238) );
  AOI22_X1 U13490 ( .A1(n11012), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1576] ), .ZN(n5237) );
  AOI22_X1 U13491 ( .A1(n11013), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1577] ), .ZN(n5236) );
  AOI22_X1 U13492 ( .A1(n11014), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1578] ), .ZN(n5235) );
  AOI22_X1 U13493 ( .A1(n11015), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1579] ), .ZN(n5234) );
  AOI22_X1 U13494 ( .A1(n11016), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1580] ), .ZN(n5233) );
  AOI22_X1 U13495 ( .A1(n11017), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1581] ), .ZN(n5232) );
  AOI22_X1 U13496 ( .A1(n11018), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1582] ), .ZN(n5231) );
  AOI22_X1 U13497 ( .A1(n11019), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1583] ), .ZN(n5230) );
  AOI22_X1 U13498 ( .A1(n11020), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1584] ), .ZN(n5229) );
  AOI22_X1 U13499 ( .A1(n11021), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1585] ), .ZN(n5228) );
  OAI22_X1 U13500 ( .A1(n11022), .A2(n8375), .B1(
        \DataPath/RF/bus_reg_dataout[1586] ), .B2(n8269), .ZN(n5227) );
  AOI22_X1 U13501 ( .A1(n11023), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1587] ), .ZN(n5226) );
  AOI22_X1 U13502 ( .A1(n11024), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1588] ), .ZN(n5225) );
  AOI22_X1 U13503 ( .A1(n11025), .A2(n8269), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1589] ), .ZN(n5224) );
  AOI22_X1 U13504 ( .A1(n11026), .A2(n11001), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1590] ), .ZN(n5223) );
  AOI22_X1 U13505 ( .A1(n11027), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1591] ), .ZN(n5222) );
  AOI22_X1 U13506 ( .A1(n11028), .A2(n11001), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1592] ), .ZN(n5221) );
  AOI22_X1 U13507 ( .A1(n11029), .A2(n11001), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1593] ), .ZN(n5220) );
  AOI22_X1 U13508 ( .A1(n11030), .A2(n11001), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1594] ), .ZN(n5219) );
  AOI22_X1 U13509 ( .A1(n11031), .A2(n11001), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1595] ), .ZN(n5218) );
  AOI22_X1 U13510 ( .A1(n11032), .A2(n11001), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1596] ), .ZN(n5217) );
  AOI22_X1 U13511 ( .A1(n11033), .A2(n11001), .B1(n8375), .B2(
        \DataPath/RF/bus_reg_dataout[1597] ), .ZN(n5216) );
  AOI22_X1 U13512 ( .A1(n11034), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1598] ), .ZN(n5215) );
  AOI22_X1 U13513 ( .A1(n11036), .A2(n8269), .B1(n11000), .B2(
        \DataPath/RF/bus_reg_dataout[1599] ), .ZN(n5212) );
  OAI22_X1 U13514 ( .A1(n8271), .A2(n11416), .B1(n8293), .B2(n11414), .ZN(
        n11002) );
  AOI22_X1 U13515 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1536] ), 
        .B1(n11004), .B2(n11035), .ZN(n5209) );
  AOI22_X1 U13516 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1537] ), 
        .B1(n11005), .B2(n11035), .ZN(n5207) );
  AOI22_X1 U13517 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1538] ), 
        .B1(n11006), .B2(n11035), .ZN(n5205) );
  AOI22_X1 U13518 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1539] ), 
        .B1(n11007), .B2(n11035), .ZN(n5203) );
  AOI22_X1 U13519 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1540] ), 
        .B1(n11008), .B2(n11035), .ZN(n5201) );
  AOI22_X1 U13520 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1541] ), 
        .B1(n11009), .B2(n11035), .ZN(n5199) );
  AOI22_X1 U13521 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1542] ), 
        .B1(n11010), .B2(n11035), .ZN(n5197) );
  AOI22_X1 U13522 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1543] ), 
        .B1(n11011), .B2(n11035), .ZN(n5195) );
  AOI22_X1 U13523 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1544] ), 
        .B1(n11012), .B2(n11035), .ZN(n5193) );
  AOI22_X1 U13524 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1545] ), 
        .B1(n11013), .B2(n11035), .ZN(n5191) );
  AOI22_X1 U13525 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1546] ), 
        .B1(n11014), .B2(n11035), .ZN(n5189) );
  AOI22_X1 U13526 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1547] ), 
        .B1(n11015), .B2(n11035), .ZN(n5187) );
  AOI22_X1 U13527 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1548] ), 
        .B1(n11016), .B2(n11035), .ZN(n5185) );
  AOI22_X1 U13528 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1549] ), 
        .B1(n11017), .B2(n11035), .ZN(n5183) );
  AOI22_X1 U13529 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1550] ), 
        .B1(n11018), .B2(n11035), .ZN(n5181) );
  AOI22_X1 U13530 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1551] ), 
        .B1(n11019), .B2(n11035), .ZN(n5179) );
  AOI22_X1 U13531 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1552] ), 
        .B1(n11020), .B2(n11035), .ZN(n5177) );
  AOI22_X1 U13532 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1553] ), 
        .B1(n11021), .B2(n11035), .ZN(n5175) );
  AOI22_X1 U13533 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1554] ), 
        .B1(n11022), .B2(n11035), .ZN(n5173) );
  AOI22_X1 U13534 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1555] ), 
        .B1(n11023), .B2(n11035), .ZN(n5171) );
  AOI22_X1 U13535 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1556] ), 
        .B1(n11024), .B2(n11035), .ZN(n5169) );
  AOI22_X1 U13536 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1557] ), 
        .B1(n11025), .B2(n11035), .ZN(n5167) );
  AOI22_X1 U13537 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1558] ), 
        .B1(n11026), .B2(n11035), .ZN(n5165) );
  AOI22_X1 U13538 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1559] ), 
        .B1(n11027), .B2(n11035), .ZN(n5163) );
  AOI22_X1 U13539 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1560] ), 
        .B1(n11028), .B2(n11035), .ZN(n5161) );
  AOI22_X1 U13540 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1561] ), 
        .B1(n11029), .B2(n11035), .ZN(n5159) );
  AOI22_X1 U13541 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1562] ), 
        .B1(n11030), .B2(n11035), .ZN(n5157) );
  AOI22_X1 U13542 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1563] ), 
        .B1(n11031), .B2(n11035), .ZN(n5155) );
  AOI22_X1 U13543 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1564] ), 
        .B1(n11032), .B2(n11035), .ZN(n5153) );
  AOI22_X1 U13544 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1565] ), 
        .B1(n11033), .B2(n11035), .ZN(n5151) );
  AOI22_X1 U13545 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1566] ), 
        .B1(n11034), .B2(n11035), .ZN(n5149) );
  AOI22_X1 U13546 ( .A1(n11037), .A2(\DataPath/RF/bus_reg_dataout[1567] ), 
        .B1(n11036), .B2(n11035), .ZN(n5145) );
  AOI22_X1 U13547 ( .A1(n7762), .A2(n11272), .B1(n11479), .B2(n11102), .ZN(
        n11071) );
  AOI22_X1 U13548 ( .A1(n11040), .A2(\DataPath/RF/bus_reg_dataout[1504] ), 
        .B1(n11038), .B2(n11071), .ZN(n5143) );
  AOI22_X1 U13549 ( .A1(n7762), .A2(n11273), .B1(n11480), .B2(n11102), .ZN(
        n11072) );
  AOI22_X1 U13550 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1505] ), .B1(
        n11038), .B2(n11072), .ZN(n5142) );
  AOI22_X1 U13551 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1506] ), .B1(
        n11038), .B2(n7779), .ZN(n5141) );
  AOI22_X1 U13552 ( .A1(n7762), .A2(n11275), .B1(n11482), .B2(n11102), .ZN(
        n11107) );
  AOI22_X1 U13553 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1507] ), .B1(
        n11038), .B2(n11107), .ZN(n5140) );
  OAI22_X1 U13554 ( .A1(n11102), .A2(n11276), .B1(n11483), .B2(n7762), .ZN(
        n11074) );
  AOI22_X1 U13555 ( .A1(\DataPath/RF/bus_reg_dataout[1508] ), .A2(n8376), .B1(
        n11124), .B2(n11039), .ZN(n5139) );
  OAI22_X1 U13556 ( .A1(n11102), .A2(n11277), .B1(n11484), .B2(n7762), .ZN(
        n11075) );
  AOI22_X1 U13557 ( .A1(\DataPath/RF/bus_reg_dataout[1509] ), .A2(n11040), 
        .B1(n11125), .B2(n11039), .ZN(n5138) );
  OAI22_X1 U13558 ( .A1(n11102), .A2(n11278), .B1(n11485), .B2(n7762), .ZN(
        n11076) );
  AOI22_X1 U13559 ( .A1(\DataPath/RF/bus_reg_dataout[1510] ), .A2(n8376), .B1(
        n11126), .B2(n11039), .ZN(n5137) );
  OAI22_X1 U13560 ( .A1(n11102), .A2(n11279), .B1(n11486), .B2(n7762), .ZN(
        n11108) );
  AOI22_X1 U13561 ( .A1(\DataPath/RF/bus_reg_dataout[1511] ), .A2(n8376), .B1(
        n11127), .B2(n11039), .ZN(n5136) );
  AOI22_X1 U13562 ( .A1(n7762), .A2(n11280), .B1(n11487), .B2(n11102), .ZN(
        n11077) );
  AOI22_X1 U13563 ( .A1(n11040), .A2(\DataPath/RF/bus_reg_dataout[1512] ), 
        .B1(n11038), .B2(n11077), .ZN(n5135) );
  AOI22_X1 U13564 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1513] ), .B1(
        n11038), .B2(n11078), .ZN(n5134) );
  AOI22_X1 U13565 ( .A1(n7762), .A2(n11282), .B1(n11489), .B2(n11102), .ZN(
        n11079) );
  AOI22_X1 U13566 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1514] ), .B1(
        n11038), .B2(n11079), .ZN(n5133) );
  AOI22_X1 U13567 ( .A1(n7762), .A2(n11283), .B1(n11490), .B2(n11102), .ZN(
        n11080) );
  AOI22_X1 U13568 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1515] ), .B1(
        n11038), .B2(n11080), .ZN(n5132) );
  AOI22_X1 U13569 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1516] ), .B1(
        n11038), .B2(n7781), .ZN(n5131) );
  AOI22_X1 U13570 ( .A1(n7762), .A2(n11285), .B1(n11492), .B2(n11102), .ZN(
        n11082) );
  AOI22_X1 U13571 ( .A1(n11040), .A2(\DataPath/RF/bus_reg_dataout[1517] ), 
        .B1(n11038), .B2(n11082), .ZN(n5130) );
  OAI22_X1 U13572 ( .A1(n11102), .A2(n11286), .B1(n11493), .B2(n7762), .ZN(
        n11109) );
  AOI22_X1 U13573 ( .A1(\DataPath/RF/bus_reg_dataout[1518] ), .A2(n8376), .B1(
        n11134), .B2(n11039), .ZN(n5129) );
  AOI22_X1 U13574 ( .A1(n11040), .A2(\DataPath/RF/bus_reg_dataout[1519] ), 
        .B1(n11038), .B2(n7778), .ZN(n5128) );
  OAI22_X1 U13575 ( .A1(n11102), .A2(n11288), .B1(n11495), .B2(n7762), .ZN(
        n11083) );
  AOI22_X1 U13576 ( .A1(\DataPath/RF/bus_reg_dataout[1520] ), .A2(n11040), 
        .B1(n11136), .B2(n11039), .ZN(n5127) );
  AOI22_X1 U13577 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1521] ), .B1(
        n11038), .B2(n7780), .ZN(n5126) );
  AOI22_X1 U13578 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1522] ), .B1(
        n11038), .B2(n11085), .ZN(n5125) );
  AOI22_X1 U13579 ( .A1(n7762), .A2(n11291), .B1(n11498), .B2(n11102), .ZN(
        n11086) );
  AOI22_X1 U13580 ( .A1(n11040), .A2(\DataPath/RF/bus_reg_dataout[1523] ), 
        .B1(n11038), .B2(n11086), .ZN(n5124) );
  AOI22_X1 U13581 ( .A1(n7762), .A2(n11292), .B1(n11499), .B2(n11102), .ZN(
        n11087) );
  AOI22_X1 U13582 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1524] ), .B1(
        n11038), .B2(n11087), .ZN(n5123) );
  AOI22_X1 U13583 ( .A1(n7762), .A2(n11293), .B1(n11500), .B2(n11102), .ZN(
        n11088) );
  AOI22_X1 U13584 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1525] ), .B1(
        n11038), .B2(n11088), .ZN(n5122) );
  AOI22_X1 U13585 ( .A1(n7762), .A2(n11294), .B1(n11501), .B2(n11102), .ZN(
        n11089) );
  AOI22_X1 U13586 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1526] ), .B1(
        n11038), .B2(n11089), .ZN(n5121) );
  OAI22_X1 U13587 ( .A1(n11102), .A2(n11295), .B1(n11502), .B2(n7762), .ZN(
        n11090) );
  AOI22_X1 U13588 ( .A1(\DataPath/RF/bus_reg_dataout[1527] ), .A2(n11040), 
        .B1(n11143), .B2(n11039), .ZN(n5120) );
  AOI22_X1 U13589 ( .A1(n7762), .A2(n11296), .B1(n11503), .B2(n11102), .ZN(
        n11055) );
  AOI22_X1 U13590 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1528] ), .B1(
        n11038), .B2(n11055), .ZN(n5119) );
  OAI22_X1 U13591 ( .A1(n11102), .A2(n11297), .B1(n11504), .B2(n7762), .ZN(
        n11111) );
  AOI22_X1 U13592 ( .A1(\DataPath/RF/bus_reg_dataout[1529] ), .A2(n8376), .B1(
        n11145), .B2(n11039), .ZN(n5118) );
  OAI22_X1 U13593 ( .A1(n11102), .A2(n11298), .B1(n11505), .B2(n7762), .ZN(
        n11091) );
  AOI22_X1 U13594 ( .A1(\DataPath/RF/bus_reg_dataout[1530] ), .A2(n8376), .B1(
        n11146), .B2(n11039), .ZN(n5117) );
  AOI22_X1 U13595 ( .A1(n7762), .A2(n11299), .B1(n11506), .B2(n11102), .ZN(
        n11092) );
  AOI22_X1 U13596 ( .A1(n11040), .A2(\DataPath/RF/bus_reg_dataout[1531] ), 
        .B1(n11038), .B2(n11092), .ZN(n5116) );
  AOI22_X1 U13597 ( .A1(n7762), .A2(n11300), .B1(n11507), .B2(n11102), .ZN(
        n11093) );
  AOI22_X1 U13598 ( .A1(n8376), .A2(\DataPath/RF/bus_reg_dataout[1532] ), .B1(
        n11038), .B2(n11093), .ZN(n5115) );
  OAI22_X1 U13599 ( .A1(n11102), .A2(n11301), .B1(n11508), .B2(n7762), .ZN(
        n11067) );
  AOI22_X1 U13600 ( .A1(\DataPath/RF/bus_reg_dataout[1533] ), .A2(n8376), .B1(
        n11149), .B2(n11039), .ZN(n5114) );
  OAI22_X1 U13601 ( .A1(n11102), .A2(n11302), .B1(n11509), .B2(n7762), .ZN(
        n11095) );
  AOI22_X1 U13602 ( .A1(\DataPath/RF/bus_reg_dataout[1534] ), .A2(n11040), 
        .B1(n11150), .B2(n11039), .ZN(n5113) );
  OAI22_X1 U13603 ( .A1(n11102), .A2(n11304), .B1(n11512), .B2(n7762), .ZN(
        n11096) );
  AOI22_X1 U13604 ( .A1(\DataPath/RF/bus_reg_dataout[1535] ), .A2(n8376), .B1(
        n11152), .B2(n11039), .ZN(n5110) );
  AOI22_X1 U13605 ( .A1(\DataPath/RF/bus_reg_dataout[1472] ), .A2(n8377), .B1(
        n11041), .B2(n11071), .ZN(n5108) );
  AOI22_X1 U13606 ( .A1(\DataPath/RF/bus_reg_dataout[1473] ), .A2(n8377), .B1(
        n11041), .B2(n11072), .ZN(n5107) );
  AOI22_X1 U13607 ( .A1(\DataPath/RF/bus_reg_dataout[1474] ), .A2(n11042), 
        .B1(n11041), .B2(n7779), .ZN(n5106) );
  AOI22_X1 U13608 ( .A1(\DataPath/RF/bus_reg_dataout[1475] ), .A2(n11042), 
        .B1(n11041), .B2(n11107), .ZN(n5105) );
  AOI22_X1 U13609 ( .A1(\DataPath/RF/bus_reg_dataout[1476] ), .A2(n11042), 
        .B1(n11041), .B2(n11074), .ZN(n5104) );
  AOI22_X1 U13610 ( .A1(\DataPath/RF/bus_reg_dataout[1477] ), .A2(n8377), .B1(
        n11041), .B2(n11075), .ZN(n5103) );
  AOI22_X1 U13611 ( .A1(n11126), .A2(n11043), .B1(n8377), .B2(
        \DataPath/RF/bus_reg_dataout[1478] ), .ZN(n5102) );
  AOI22_X1 U13612 ( .A1(\DataPath/RF/bus_reg_dataout[1479] ), .A2(n8377), .B1(
        n11041), .B2(n11108), .ZN(n5101) );
  AOI22_X1 U13613 ( .A1(\DataPath/RF/bus_reg_dataout[1480] ), .A2(n8377), .B1(
        n11041), .B2(n11077), .ZN(n5100) );
  AOI22_X1 U13614 ( .A1(\DataPath/RF/bus_reg_dataout[1481] ), .A2(n8377), .B1(
        n11041), .B2(n11078), .ZN(n5099) );
  AOI22_X1 U13615 ( .A1(\DataPath/RF/bus_reg_dataout[1482] ), .A2(n8377), .B1(
        n11041), .B2(n11079), .ZN(n5098) );
  AOI22_X1 U13616 ( .A1(\DataPath/RF/bus_reg_dataout[1483] ), .A2(n8377), .B1(
        n11041), .B2(n11080), .ZN(n5097) );
  AOI22_X1 U13617 ( .A1(\DataPath/RF/bus_reg_dataout[1484] ), .A2(n11042), 
        .B1(n11041), .B2(n7781), .ZN(n5096) );
  AOI22_X1 U13618 ( .A1(\DataPath/RF/bus_reg_dataout[1485] ), .A2(n11042), 
        .B1(n11041), .B2(n11082), .ZN(n5095) );
  AOI22_X1 U13619 ( .A1(\DataPath/RF/bus_reg_dataout[1486] ), .A2(n8377), .B1(
        n11041), .B2(n11109), .ZN(n5094) );
  AOI22_X1 U13620 ( .A1(\DataPath/RF/bus_reg_dataout[1487] ), .A2(n8377), .B1(
        n11041), .B2(n7778), .ZN(n5093) );
  AOI22_X1 U13621 ( .A1(\DataPath/RF/bus_reg_dataout[1488] ), .A2(n8377), .B1(
        n11041), .B2(n11083), .ZN(n5092) );
  AOI22_X1 U13622 ( .A1(\DataPath/RF/bus_reg_dataout[1489] ), .A2(n11042), 
        .B1(n11041), .B2(n7780), .ZN(n5091) );
  AOI22_X1 U13623 ( .A1(\DataPath/RF/bus_reg_dataout[1490] ), .A2(n11042), 
        .B1(n11041), .B2(n11085), .ZN(n5090) );
  AOI22_X1 U13624 ( .A1(\DataPath/RF/bus_reg_dataout[1491] ), .A2(n8377), .B1(
        n11139), .B2(n11043), .ZN(n5089) );
  AOI22_X1 U13625 ( .A1(\DataPath/RF/bus_reg_dataout[1492] ), .A2(n8377), .B1(
        n11041), .B2(n11087), .ZN(n5088) );
  AOI22_X1 U13626 ( .A1(\DataPath/RF/bus_reg_dataout[1493] ), .A2(n8377), .B1(
        n11041), .B2(n11088), .ZN(n5087) );
  AOI22_X1 U13627 ( .A1(\DataPath/RF/bus_reg_dataout[1494] ), .A2(n11042), 
        .B1(n11041), .B2(n11089), .ZN(n5086) );
  AOI22_X1 U13628 ( .A1(\DataPath/RF/bus_reg_dataout[1495] ), .A2(n11042), 
        .B1(n11041), .B2(n11090), .ZN(n5085) );
  AOI22_X1 U13629 ( .A1(\DataPath/RF/bus_reg_dataout[1496] ), .A2(n8377), .B1(
        n11041), .B2(n11055), .ZN(n5084) );
  AOI22_X1 U13630 ( .A1(\DataPath/RF/bus_reg_dataout[1497] ), .A2(n8377), .B1(
        n11041), .B2(n11111), .ZN(n5083) );
  AOI22_X1 U13631 ( .A1(\DataPath/RF/bus_reg_dataout[1498] ), .A2(n8377), .B1(
        n11041), .B2(n11091), .ZN(n5082) );
  AOI22_X1 U13632 ( .A1(\DataPath/RF/bus_reg_dataout[1499] ), .A2(n11042), 
        .B1(n11041), .B2(n11092), .ZN(n5081) );
  AOI22_X1 U13633 ( .A1(\DataPath/RF/bus_reg_dataout[1500] ), .A2(n8377), .B1(
        n11041), .B2(n11093), .ZN(n5080) );
  AOI22_X1 U13634 ( .A1(\DataPath/RF/bus_reg_dataout[1501] ), .A2(n8377), .B1(
        n11041), .B2(n11067), .ZN(n5079) );
  AOI22_X1 U13635 ( .A1(\DataPath/RF/bus_reg_dataout[1502] ), .A2(n8377), .B1(
        n11041), .B2(n11095), .ZN(n5078) );
  AOI22_X1 U13636 ( .A1(n11152), .A2(n11043), .B1(n8377), .B2(
        \DataPath/RF/bus_reg_dataout[1503] ), .ZN(n5075) );
  OAI22_X1 U13637 ( .A1(n11120), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1440] ), .B2(n11044), .ZN(n5073) );
  OAI22_X1 U13638 ( .A1(n8379), .A2(n11121), .B1(
        \DataPath/RF/bus_reg_dataout[1441] ), .B2(n8378), .ZN(n5072) );
  OAI22_X1 U13639 ( .A1(n8379), .A2(n11122), .B1(
        \DataPath/RF/bus_reg_dataout[1442] ), .B2(n8378), .ZN(n5071) );
  OAI22_X1 U13640 ( .A1(n8379), .A2(n11123), .B1(
        \DataPath/RF/bus_reg_dataout[1443] ), .B2(n8378), .ZN(n5070) );
  OAI22_X1 U13641 ( .A1(n11124), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1444] ), .B2(n11044), .ZN(n5069) );
  OAI22_X1 U13642 ( .A1(n11125), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1445] ), .B2(n11044), .ZN(n5068) );
  OAI22_X1 U13643 ( .A1(n11126), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1446] ), .B2(n8378), .ZN(n5067) );
  OAI22_X1 U13644 ( .A1(n11127), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1447] ), .B2(n8378), .ZN(n5066) );
  OAI22_X1 U13645 ( .A1(n11045), .A2(n11128), .B1(
        \DataPath/RF/bus_reg_dataout[1448] ), .B2(n8378), .ZN(n5065) );
  OAI22_X1 U13646 ( .A1(n11045), .A2(n11129), .B1(
        \DataPath/RF/bus_reg_dataout[1449] ), .B2(n11044), .ZN(n5064) );
  OAI22_X1 U13647 ( .A1(n8379), .A2(n11130), .B1(
        \DataPath/RF/bus_reg_dataout[1450] ), .B2(n8378), .ZN(n5063) );
  OAI22_X1 U13648 ( .A1(n8379), .A2(n11131), .B1(
        \DataPath/RF/bus_reg_dataout[1451] ), .B2(n8378), .ZN(n5062) );
  OAI22_X1 U13649 ( .A1(n8379), .A2(n11132), .B1(
        \DataPath/RF/bus_reg_dataout[1452] ), .B2(n11044), .ZN(n5061) );
  OAI22_X1 U13650 ( .A1(n11045), .A2(n11133), .B1(
        \DataPath/RF/bus_reg_dataout[1453] ), .B2(n11044), .ZN(n5060) );
  OAI22_X1 U13651 ( .A1(n11134), .A2(n11045), .B1(
        \DataPath/RF/bus_reg_dataout[1454] ), .B2(n11044), .ZN(n5059) );
  OAI22_X1 U13652 ( .A1(n8379), .A2(n11135), .B1(
        \DataPath/RF/bus_reg_dataout[1455] ), .B2(n8378), .ZN(n5058) );
  OAI22_X1 U13653 ( .A1(n11136), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1456] ), .B2(n8378), .ZN(n5057) );
  OAI22_X1 U13654 ( .A1(n8379), .A2(n11137), .B1(
        \DataPath/RF/bus_reg_dataout[1457] ), .B2(n8378), .ZN(n5056) );
  OAI22_X1 U13655 ( .A1(n8379), .A2(n11138), .B1(
        \DataPath/RF/bus_reg_dataout[1458] ), .B2(n11044), .ZN(n5055) );
  OAI22_X1 U13656 ( .A1(n11139), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1459] ), .B2(n8378), .ZN(n5054) );
  OAI22_X1 U13657 ( .A1(n11045), .A2(n11140), .B1(
        \DataPath/RF/bus_reg_dataout[1460] ), .B2(n8378), .ZN(n5053) );
  OAI22_X1 U13658 ( .A1(n11045), .A2(n11141), .B1(
        \DataPath/RF/bus_reg_dataout[1461] ), .B2(n8378), .ZN(n5052) );
  OAI22_X1 U13659 ( .A1(n8379), .A2(n11142), .B1(
        \DataPath/RF/bus_reg_dataout[1462] ), .B2(n11044), .ZN(n5051) );
  OAI22_X1 U13660 ( .A1(n11143), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1463] ), .B2(n8378), .ZN(n5050) );
  OAI22_X1 U13661 ( .A1(n8379), .A2(n11144), .B1(
        \DataPath/RF/bus_reg_dataout[1464] ), .B2(n8378), .ZN(n5049) );
  OAI22_X1 U13662 ( .A1(n11145), .A2(n11045), .B1(
        \DataPath/RF/bus_reg_dataout[1465] ), .B2(n8378), .ZN(n5048) );
  OAI22_X1 U13663 ( .A1(n11146), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1466] ), .B2(n8378), .ZN(n5047) );
  OAI22_X1 U13664 ( .A1(n8379), .A2(n11147), .B1(
        \DataPath/RF/bus_reg_dataout[1467] ), .B2(n8378), .ZN(n5046) );
  OAI22_X1 U13665 ( .A1(n11045), .A2(n11148), .B1(
        \DataPath/RF/bus_reg_dataout[1468] ), .B2(n8378), .ZN(n5045) );
  OAI22_X1 U13666 ( .A1(n11149), .A2(n8379), .B1(
        \DataPath/RF/bus_reg_dataout[1469] ), .B2(n8378), .ZN(n5044) );
  OAI22_X1 U13667 ( .A1(n11150), .A2(n11045), .B1(
        \DataPath/RF/bus_reg_dataout[1470] ), .B2(n8378), .ZN(n5043) );
  OAI22_X1 U13668 ( .A1(n11152), .A2(n11045), .B1(
        \DataPath/RF/bus_reg_dataout[1471] ), .B2(n8378), .ZN(n5040) );
  AOI22_X1 U13669 ( .A1(\DataPath/RF/bus_reg_dataout[1408] ), .A2(n8380), .B1(
        n11046), .B2(n11071), .ZN(n5038) );
  AOI22_X1 U13670 ( .A1(\DataPath/RF/bus_reg_dataout[1409] ), .A2(n8380), .B1(
        n11046), .B2(n11072), .ZN(n5037) );
  AOI22_X1 U13671 ( .A1(\DataPath/RF/bus_reg_dataout[1410] ), .A2(n8380), .B1(
        n11046), .B2(n7779), .ZN(n5036) );
  AOI22_X1 U13672 ( .A1(\DataPath/RF/bus_reg_dataout[1411] ), .A2(n11047), 
        .B1(n11046), .B2(n11107), .ZN(n5035) );
  AOI22_X1 U13673 ( .A1(\DataPath/RF/bus_reg_dataout[1412] ), .A2(n8380), .B1(
        n11046), .B2(n11074), .ZN(n5034) );
  AOI22_X1 U13674 ( .A1(\DataPath/RF/bus_reg_dataout[1413] ), .A2(n11047), 
        .B1(n11046), .B2(n11075), .ZN(n5033) );
  AOI22_X1 U13675 ( .A1(\DataPath/RF/bus_reg_dataout[1414] ), .A2(n8380), .B1(
        n11046), .B2(n11076), .ZN(n5032) );
  AOI22_X1 U13676 ( .A1(\DataPath/RF/bus_reg_dataout[1415] ), .A2(n11047), 
        .B1(n11046), .B2(n11108), .ZN(n5031) );
  AOI22_X1 U13677 ( .A1(\DataPath/RF/bus_reg_dataout[1416] ), .A2(n8380), .B1(
        n11046), .B2(n11077), .ZN(n5030) );
  AOI22_X1 U13678 ( .A1(\DataPath/RF/bus_reg_dataout[1417] ), .A2(n11047), 
        .B1(n11046), .B2(n11078), .ZN(n5029) );
  AOI22_X1 U13679 ( .A1(\DataPath/RF/bus_reg_dataout[1418] ), .A2(n8380), .B1(
        n11046), .B2(n11079), .ZN(n5028) );
  AOI22_X1 U13680 ( .A1(\DataPath/RF/bus_reg_dataout[1419] ), .A2(n8380), .B1(
        n11046), .B2(n11080), .ZN(n5027) );
  AOI22_X1 U13681 ( .A1(\DataPath/RF/bus_reg_dataout[1420] ), .A2(n8380), .B1(
        n11046), .B2(n7781), .ZN(n5026) );
  AOI22_X1 U13682 ( .A1(\DataPath/RF/bus_reg_dataout[1421] ), .A2(n8380), .B1(
        n11046), .B2(n11082), .ZN(n5025) );
  AOI22_X1 U13683 ( .A1(\DataPath/RF/bus_reg_dataout[1422] ), .A2(n8380), .B1(
        n11046), .B2(n11109), .ZN(n5024) );
  AOI22_X1 U13684 ( .A1(\DataPath/RF/bus_reg_dataout[1423] ), .A2(n8380), .B1(
        n11046), .B2(n7778), .ZN(n5023) );
  AOI22_X1 U13685 ( .A1(\DataPath/RF/bus_reg_dataout[1424] ), .A2(n11047), 
        .B1(n11046), .B2(n11083), .ZN(n5022) );
  AOI22_X1 U13686 ( .A1(\DataPath/RF/bus_reg_dataout[1425] ), .A2(n11047), 
        .B1(n11046), .B2(n7780), .ZN(n5021) );
  AOI22_X1 U13687 ( .A1(\DataPath/RF/bus_reg_dataout[1426] ), .A2(n11047), 
        .B1(n11046), .B2(n11085), .ZN(n5020) );
  AOI22_X1 U13688 ( .A1(\DataPath/RF/bus_reg_dataout[1427] ), .A2(n8380), .B1(
        n11046), .B2(n11086), .ZN(n5019) );
  AOI22_X1 U13689 ( .A1(\DataPath/RF/bus_reg_dataout[1428] ), .A2(n8380), .B1(
        n11046), .B2(n11087), .ZN(n5018) );
  AOI22_X1 U13690 ( .A1(\DataPath/RF/bus_reg_dataout[1429] ), .A2(n11047), 
        .B1(n11046), .B2(n11088), .ZN(n5017) );
  AOI22_X1 U13691 ( .A1(\DataPath/RF/bus_reg_dataout[1430] ), .A2(n8380), .B1(
        n11046), .B2(n11089), .ZN(n5016) );
  AOI22_X1 U13692 ( .A1(\DataPath/RF/bus_reg_dataout[1431] ), .A2(n8380), .B1(
        n11046), .B2(n11090), .ZN(n5015) );
  AOI22_X1 U13693 ( .A1(\DataPath/RF/bus_reg_dataout[1432] ), .A2(n8380), .B1(
        n11046), .B2(n11055), .ZN(n5014) );
  AOI22_X1 U13694 ( .A1(\DataPath/RF/bus_reg_dataout[1433] ), .A2(n11047), 
        .B1(n11046), .B2(n11111), .ZN(n5013) );
  AOI22_X1 U13695 ( .A1(\DataPath/RF/bus_reg_dataout[1434] ), .A2(n8380), .B1(
        n11046), .B2(n11091), .ZN(n5012) );
  AOI22_X1 U13696 ( .A1(\DataPath/RF/bus_reg_dataout[1435] ), .A2(n8380), .B1(
        n11046), .B2(n11092), .ZN(n5011) );
  AOI22_X1 U13697 ( .A1(n11148), .A2(n11048), .B1(n8380), .B2(
        \DataPath/RF/bus_reg_dataout[1436] ), .ZN(n5010) );
  AOI22_X1 U13698 ( .A1(\DataPath/RF/bus_reg_dataout[1437] ), .A2(n8380), .B1(
        n11046), .B2(n11067), .ZN(n5009) );
  AOI22_X1 U13699 ( .A1(n11150), .A2(n11048), .B1(n11047), .B2(
        \DataPath/RF/bus_reg_dataout[1438] ), .ZN(n5008) );
  AOI22_X1 U13700 ( .A1(n11152), .A2(n11048), .B1(n8380), .B2(
        \DataPath/RF/bus_reg_dataout[1439] ), .ZN(n5005) );
  OAI22_X1 U13701 ( .A1(n8271), .A2(n11773), .B1(n11772), .B2(n11102), .ZN(
        n11049) );
  AOI22_X1 U13702 ( .A1(\DataPath/RF/bus_reg_dataout[1376] ), .A2(n8381), .B1(
        n11050), .B2(n11071), .ZN(n5003) );
  AOI22_X1 U13703 ( .A1(\DataPath/RF/bus_reg_dataout[1377] ), .A2(n8381), .B1(
        n11050), .B2(n11072), .ZN(n5002) );
  AOI22_X1 U13704 ( .A1(\DataPath/RF/bus_reg_dataout[1378] ), .A2(n8381), .B1(
        n11050), .B2(n7779), .ZN(n5001) );
  AOI22_X1 U13705 ( .A1(\DataPath/RF/bus_reg_dataout[1379] ), .A2(n8381), .B1(
        n11050), .B2(n11107), .ZN(n5000) );
  AOI22_X1 U13706 ( .A1(\DataPath/RF/bus_reg_dataout[1380] ), .A2(n8381), .B1(
        n11050), .B2(n11074), .ZN(n4999) );
  AOI22_X1 U13707 ( .A1(\DataPath/RF/bus_reg_dataout[1381] ), .A2(n11051), 
        .B1(n11050), .B2(n11075), .ZN(n4998) );
  AOI22_X1 U13708 ( .A1(\DataPath/RF/bus_reg_dataout[1382] ), .A2(n8381), .B1(
        n11050), .B2(n11076), .ZN(n4997) );
  AOI22_X1 U13709 ( .A1(\DataPath/RF/bus_reg_dataout[1383] ), .A2(n11051), 
        .B1(n11050), .B2(n11108), .ZN(n4996) );
  AOI22_X1 U13710 ( .A1(\DataPath/RF/bus_reg_dataout[1384] ), .A2(n8381), .B1(
        n11050), .B2(n11077), .ZN(n4995) );
  AOI22_X1 U13711 ( .A1(\DataPath/RF/bus_reg_dataout[1385] ), .A2(n8381), .B1(
        n11050), .B2(n11078), .ZN(n4994) );
  AOI22_X1 U13712 ( .A1(\DataPath/RF/bus_reg_dataout[1386] ), .A2(n8381), .B1(
        n11050), .B2(n11079), .ZN(n4993) );
  AOI22_X1 U13713 ( .A1(\DataPath/RF/bus_reg_dataout[1387] ), .A2(n8381), .B1(
        n11050), .B2(n11080), .ZN(n4992) );
  AOI22_X1 U13714 ( .A1(\DataPath/RF/bus_reg_dataout[1388] ), .A2(n8381), .B1(
        n11050), .B2(n7781), .ZN(n4991) );
  AOI22_X1 U13715 ( .A1(\DataPath/RF/bus_reg_dataout[1389] ), .A2(n8381), .B1(
        n11050), .B2(n11082), .ZN(n4990) );
  AOI22_X1 U13716 ( .A1(\DataPath/RF/bus_reg_dataout[1390] ), .A2(n11051), 
        .B1(n11050), .B2(n11109), .ZN(n4989) );
  AOI22_X1 U13717 ( .A1(\DataPath/RF/bus_reg_dataout[1391] ), .A2(n8381), .B1(
        n11050), .B2(n7778), .ZN(n4988) );
  AOI22_X1 U13718 ( .A1(\DataPath/RF/bus_reg_dataout[1392] ), .A2(n11051), 
        .B1(n11050), .B2(n11083), .ZN(n4987) );
  AOI22_X1 U13719 ( .A1(\DataPath/RF/bus_reg_dataout[1393] ), .A2(n11051), 
        .B1(n11050), .B2(n7780), .ZN(n4986) );
  AOI22_X1 U13720 ( .A1(\DataPath/RF/bus_reg_dataout[1394] ), .A2(n11051), 
        .B1(n11050), .B2(n11085), .ZN(n4985) );
  AOI22_X1 U13721 ( .A1(\DataPath/RF/bus_reg_dataout[1395] ), .A2(n8381), .B1(
        n11050), .B2(n11086), .ZN(n4984) );
  AOI22_X1 U13722 ( .A1(\DataPath/RF/bus_reg_dataout[1396] ), .A2(n8381), .B1(
        n11050), .B2(n11087), .ZN(n4983) );
  AOI22_X1 U13723 ( .A1(\DataPath/RF/bus_reg_dataout[1397] ), .A2(n11051), 
        .B1(n11050), .B2(n11088), .ZN(n4982) );
  AOI22_X1 U13724 ( .A1(\DataPath/RF/bus_reg_dataout[1398] ), .A2(n8381), .B1(
        n11050), .B2(n11089), .ZN(n4981) );
  AOI22_X1 U13725 ( .A1(\DataPath/RF/bus_reg_dataout[1399] ), .A2(n11051), 
        .B1(n11050), .B2(n11090), .ZN(n4980) );
  AOI22_X1 U13726 ( .A1(\DataPath/RF/bus_reg_dataout[1400] ), .A2(n8381), .B1(
        n11050), .B2(n11055), .ZN(n4979) );
  AOI22_X1 U13727 ( .A1(\DataPath/RF/bus_reg_dataout[1401] ), .A2(n11051), 
        .B1(n11050), .B2(n11111), .ZN(n4978) );
  AOI22_X1 U13728 ( .A1(\DataPath/RF/bus_reg_dataout[1402] ), .A2(n8381), .B1(
        n11050), .B2(n11091), .ZN(n4977) );
  AOI22_X1 U13729 ( .A1(\DataPath/RF/bus_reg_dataout[1403] ), .A2(n8381), .B1(
        n11050), .B2(n11092), .ZN(n4976) );
  AOI22_X1 U13730 ( .A1(\DataPath/RF/bus_reg_dataout[1404] ), .A2(n8381), .B1(
        n11050), .B2(n11093), .ZN(n4975) );
  AOI22_X1 U13731 ( .A1(\DataPath/RF/bus_reg_dataout[1405] ), .A2(n8381), .B1(
        n11050), .B2(n11067), .ZN(n4974) );
  AOI22_X1 U13732 ( .A1(\DataPath/RF/bus_reg_dataout[1406] ), .A2(n11051), 
        .B1(n11050), .B2(n11095), .ZN(n4973) );
  AOI22_X1 U13733 ( .A1(\DataPath/RF/bus_reg_dataout[1407] ), .A2(n8381), .B1(
        n11050), .B2(n11096), .ZN(n4970) );
  OAI22_X1 U13734 ( .A1(n8271), .A2(n11322), .B1(n11321), .B2(n11102), .ZN(
        n11052) );
  AOI22_X1 U13735 ( .A1(\DataPath/RF/bus_reg_dataout[1344] ), .A2(n8382), .B1(
        n11053), .B2(n11071), .ZN(n4968) );
  AOI22_X1 U13736 ( .A1(\DataPath/RF/bus_reg_dataout[1345] ), .A2(n8382), .B1(
        n11053), .B2(n11072), .ZN(n4967) );
  AOI22_X1 U13737 ( .A1(\DataPath/RF/bus_reg_dataout[1346] ), .A2(n11054), 
        .B1(n11053), .B2(n7779), .ZN(n4966) );
  AOI22_X1 U13738 ( .A1(\DataPath/RF/bus_reg_dataout[1347] ), .A2(n11054), 
        .B1(n11053), .B2(n11107), .ZN(n4965) );
  AOI22_X1 U13739 ( .A1(\DataPath/RF/bus_reg_dataout[1348] ), .A2(n11054), 
        .B1(n11053), .B2(n11074), .ZN(n4964) );
  AOI22_X1 U13740 ( .A1(\DataPath/RF/bus_reg_dataout[1349] ), .A2(n8382), .B1(
        n11053), .B2(n11075), .ZN(n4963) );
  AOI22_X1 U13741 ( .A1(\DataPath/RF/bus_reg_dataout[1350] ), .A2(n8382), .B1(
        n11053), .B2(n11076), .ZN(n4962) );
  AOI22_X1 U13742 ( .A1(\DataPath/RF/bus_reg_dataout[1351] ), .A2(n8382), .B1(
        n11053), .B2(n11108), .ZN(n4961) );
  AOI22_X1 U13743 ( .A1(\DataPath/RF/bus_reg_dataout[1352] ), .A2(n11054), 
        .B1(n11053), .B2(n11077), .ZN(n4960) );
  AOI22_X1 U13744 ( .A1(\DataPath/RF/bus_reg_dataout[1353] ), .A2(n11054), 
        .B1(n11053), .B2(n11078), .ZN(n4959) );
  AOI22_X1 U13745 ( .A1(\DataPath/RF/bus_reg_dataout[1354] ), .A2(n8382), .B1(
        n11053), .B2(n11079), .ZN(n4958) );
  AOI22_X1 U13746 ( .A1(\DataPath/RF/bus_reg_dataout[1355] ), .A2(n8382), .B1(
        n11053), .B2(n11080), .ZN(n4957) );
  AOI22_X1 U13747 ( .A1(\DataPath/RF/bus_reg_dataout[1356] ), .A2(n11054), 
        .B1(n11053), .B2(n7781), .ZN(n4956) );
  AOI22_X1 U13748 ( .A1(\DataPath/RF/bus_reg_dataout[1357] ), .A2(n11054), 
        .B1(n11053), .B2(n11082), .ZN(n4955) );
  AOI22_X1 U13749 ( .A1(\DataPath/RF/bus_reg_dataout[1358] ), .A2(n8382), .B1(
        n11053), .B2(n11109), .ZN(n4954) );
  AOI22_X1 U13750 ( .A1(\DataPath/RF/bus_reg_dataout[1359] ), .A2(n8382), .B1(
        n11053), .B2(n7778), .ZN(n4953) );
  AOI22_X1 U13751 ( .A1(\DataPath/RF/bus_reg_dataout[1360] ), .A2(n8382), .B1(
        n11053), .B2(n11083), .ZN(n4952) );
  AOI22_X1 U13752 ( .A1(\DataPath/RF/bus_reg_dataout[1361] ), .A2(n8382), .B1(
        n11053), .B2(n7780), .ZN(n4951) );
  AOI22_X1 U13753 ( .A1(\DataPath/RF/bus_reg_dataout[1362] ), .A2(n11054), 
        .B1(n11053), .B2(n11085), .ZN(n4950) );
  AOI22_X1 U13754 ( .A1(\DataPath/RF/bus_reg_dataout[1363] ), .A2(n8382), .B1(
        n11053), .B2(n11086), .ZN(n4949) );
  AOI22_X1 U13755 ( .A1(\DataPath/RF/bus_reg_dataout[1364] ), .A2(n8382), .B1(
        n11053), .B2(n11087), .ZN(n4948) );
  AOI22_X1 U13756 ( .A1(\DataPath/RF/bus_reg_dataout[1365] ), .A2(n11054), 
        .B1(n11053), .B2(n11088), .ZN(n4947) );
  AOI22_X1 U13757 ( .A1(\DataPath/RF/bus_reg_dataout[1366] ), .A2(n8382), .B1(
        n11053), .B2(n11089), .ZN(n4946) );
  AOI22_X1 U13758 ( .A1(\DataPath/RF/bus_reg_dataout[1367] ), .A2(n8382), .B1(
        n11053), .B2(n11090), .ZN(n4945) );
  AOI22_X1 U13759 ( .A1(\DataPath/RF/bus_reg_dataout[1368] ), .A2(n8382), .B1(
        n11053), .B2(n11055), .ZN(n4944) );
  AOI22_X1 U13760 ( .A1(\DataPath/RF/bus_reg_dataout[1369] ), .A2(n8382), .B1(
        n11053), .B2(n11111), .ZN(n4943) );
  AOI22_X1 U13761 ( .A1(\DataPath/RF/bus_reg_dataout[1370] ), .A2(n11054), 
        .B1(n11053), .B2(n11091), .ZN(n4942) );
  AOI22_X1 U13762 ( .A1(\DataPath/RF/bus_reg_dataout[1371] ), .A2(n8382), .B1(
        n11053), .B2(n11092), .ZN(n4941) );
  AOI22_X1 U13763 ( .A1(\DataPath/RF/bus_reg_dataout[1372] ), .A2(n8382), .B1(
        n11053), .B2(n11093), .ZN(n4940) );
  AOI22_X1 U13764 ( .A1(n11149), .A2(n11052), .B1(n8382), .B2(
        \DataPath/RF/bus_reg_dataout[1373] ), .ZN(n4939) );
  AOI22_X1 U13765 ( .A1(n11150), .A2(n11052), .B1(n8382), .B2(
        \DataPath/RF/bus_reg_dataout[1374] ), .ZN(n4938) );
  AOI22_X1 U13766 ( .A1(\DataPath/RF/bus_reg_dataout[1375] ), .A2(n8382), .B1(
        n11053), .B2(n11096), .ZN(n4935) );
  OAI22_X1 U13767 ( .A1(n8271), .A2(n11327), .B1(n11326), .B2(n11102), .ZN(
        n11056) );
  AOI22_X1 U13768 ( .A1(\DataPath/RF/bus_reg_dataout[1312] ), .A2(n8383), .B1(
        n11057), .B2(n11071), .ZN(n4933) );
  AOI22_X1 U13769 ( .A1(\DataPath/RF/bus_reg_dataout[1313] ), .A2(n8383), .B1(
        n11057), .B2(n11072), .ZN(n4932) );
  AOI22_X1 U13770 ( .A1(\DataPath/RF/bus_reg_dataout[1314] ), .A2(n11058), 
        .B1(n11057), .B2(n7779), .ZN(n4931) );
  AOI22_X1 U13771 ( .A1(\DataPath/RF/bus_reg_dataout[1315] ), .A2(n11058), 
        .B1(n11057), .B2(n11107), .ZN(n4930) );
  AOI22_X1 U13772 ( .A1(\DataPath/RF/bus_reg_dataout[1316] ), .A2(n11058), 
        .B1(n11057), .B2(n11074), .ZN(n4929) );
  AOI22_X1 U13773 ( .A1(\DataPath/RF/bus_reg_dataout[1317] ), .A2(n8383), .B1(
        n11057), .B2(n11075), .ZN(n4928) );
  AOI22_X1 U13774 ( .A1(\DataPath/RF/bus_reg_dataout[1318] ), .A2(n8383), .B1(
        n11057), .B2(n11076), .ZN(n4927) );
  AOI22_X1 U13775 ( .A1(\DataPath/RF/bus_reg_dataout[1319] ), .A2(n8383), .B1(
        n11057), .B2(n11108), .ZN(n4926) );
  AOI22_X1 U13776 ( .A1(\DataPath/RF/bus_reg_dataout[1320] ), .A2(n11058), 
        .B1(n11057), .B2(n11077), .ZN(n4925) );
  AOI22_X1 U13777 ( .A1(\DataPath/RF/bus_reg_dataout[1321] ), .A2(n11058), 
        .B1(n11057), .B2(n11078), .ZN(n4924) );
  AOI22_X1 U13778 ( .A1(\DataPath/RF/bus_reg_dataout[1322] ), .A2(n8383), .B1(
        n11057), .B2(n11079), .ZN(n4923) );
  AOI22_X1 U13779 ( .A1(\DataPath/RF/bus_reg_dataout[1323] ), .A2(n8383), .B1(
        n11057), .B2(n11080), .ZN(n4922) );
  AOI22_X1 U13780 ( .A1(\DataPath/RF/bus_reg_dataout[1324] ), .A2(n11058), 
        .B1(n11057), .B2(n7781), .ZN(n4921) );
  AOI22_X1 U13781 ( .A1(\DataPath/RF/bus_reg_dataout[1325] ), .A2(n11058), 
        .B1(n11057), .B2(n11082), .ZN(n4920) );
  AOI22_X1 U13782 ( .A1(\DataPath/RF/bus_reg_dataout[1326] ), .A2(n8383), .B1(
        n11057), .B2(n11109), .ZN(n4919) );
  AOI22_X1 U13783 ( .A1(\DataPath/RF/bus_reg_dataout[1327] ), .A2(n8383), .B1(
        n11057), .B2(n7778), .ZN(n4918) );
  AOI22_X1 U13784 ( .A1(\DataPath/RF/bus_reg_dataout[1328] ), .A2(n8383), .B1(
        n11057), .B2(n11083), .ZN(n4917) );
  AOI22_X1 U13785 ( .A1(\DataPath/RF/bus_reg_dataout[1329] ), .A2(n8383), .B1(
        n11057), .B2(n7780), .ZN(n4916) );
  AOI22_X1 U13786 ( .A1(\DataPath/RF/bus_reg_dataout[1330] ), .A2(n11058), 
        .B1(n11057), .B2(n11085), .ZN(n4915) );
  AOI22_X1 U13787 ( .A1(\DataPath/RF/bus_reg_dataout[1331] ), .A2(n8383), .B1(
        n11057), .B2(n11086), .ZN(n4914) );
  AOI22_X1 U13788 ( .A1(\DataPath/RF/bus_reg_dataout[1332] ), .A2(n8383), .B1(
        n11057), .B2(n11087), .ZN(n4913) );
  AOI22_X1 U13789 ( .A1(\DataPath/RF/bus_reg_dataout[1333] ), .A2(n11058), 
        .B1(n11057), .B2(n11088), .ZN(n4912) );
  AOI22_X1 U13790 ( .A1(\DataPath/RF/bus_reg_dataout[1334] ), .A2(n8383), .B1(
        n11057), .B2(n11089), .ZN(n4911) );
  AOI22_X1 U13791 ( .A1(\DataPath/RF/bus_reg_dataout[1335] ), .A2(n8383), .B1(
        n11057), .B2(n11090), .ZN(n4910) );
  AOI22_X1 U13792 ( .A1(\DataPath/RF/bus_reg_dataout[1336] ), .A2(n8383), .B1(
        n11057), .B2(n11055), .ZN(n4909) );
  AOI22_X1 U13793 ( .A1(n11145), .A2(n11056), .B1(n8383), .B2(
        \DataPath/RF/bus_reg_dataout[1337] ), .ZN(n4908) );
  AOI22_X1 U13794 ( .A1(\DataPath/RF/bus_reg_dataout[1338] ), .A2(n8383), .B1(
        n11057), .B2(n11091), .ZN(n4907) );
  AOI22_X1 U13795 ( .A1(\DataPath/RF/bus_reg_dataout[1339] ), .A2(n11058), 
        .B1(n11057), .B2(n11092), .ZN(n4906) );
  AOI22_X1 U13796 ( .A1(n11148), .A2(n11056), .B1(n8383), .B2(
        \DataPath/RF/bus_reg_dataout[1340] ), .ZN(n4905) );
  AOI22_X1 U13797 ( .A1(\DataPath/RF/bus_reg_dataout[1341] ), .A2(n8383), .B1(
        n11057), .B2(n11067), .ZN(n4904) );
  AOI22_X1 U13798 ( .A1(\DataPath/RF/bus_reg_dataout[1342] ), .A2(n8383), .B1(
        n11057), .B2(n11095), .ZN(n4903) );
  AOI22_X1 U13799 ( .A1(\DataPath/RF/bus_reg_dataout[1343] ), .A2(n8383), .B1(
        n11057), .B2(n11096), .ZN(n4900) );
  AOI22_X1 U13800 ( .A1(\DataPath/RF/bus_reg_dataout[1280] ), .A2(n8384), .B1(
        n11060), .B2(n11071), .ZN(n4898) );
  AOI22_X1 U13801 ( .A1(\DataPath/RF/bus_reg_dataout[1281] ), .A2(n8384), .B1(
        n11060), .B2(n11072), .ZN(n4897) );
  AOI22_X1 U13802 ( .A1(\DataPath/RF/bus_reg_dataout[1282] ), .A2(n8384), .B1(
        n11060), .B2(n7779), .ZN(n4896) );
  AOI22_X1 U13803 ( .A1(n11123), .A2(n11059), .B1(n11061), .B2(
        \DataPath/RF/bus_reg_dataout[1283] ), .ZN(n4895) );
  AOI22_X1 U13804 ( .A1(\DataPath/RF/bus_reg_dataout[1284] ), .A2(n11061), 
        .B1(n11060), .B2(n11074), .ZN(n4894) );
  AOI22_X1 U13805 ( .A1(\DataPath/RF/bus_reg_dataout[1285] ), .A2(n11061), 
        .B1(n11060), .B2(n11075), .ZN(n4893) );
  AOI22_X1 U13806 ( .A1(\DataPath/RF/bus_reg_dataout[1286] ), .A2(n8384), .B1(
        n11060), .B2(n11076), .ZN(n4892) );
  AOI22_X1 U13807 ( .A1(\DataPath/RF/bus_reg_dataout[1287] ), .A2(n8384), .B1(
        n11060), .B2(n11108), .ZN(n4891) );
  AOI22_X1 U13808 ( .A1(\DataPath/RF/bus_reg_dataout[1288] ), .A2(n8384), .B1(
        n11060), .B2(n11077), .ZN(n4890) );
  AOI22_X1 U13809 ( .A1(\DataPath/RF/bus_reg_dataout[1289] ), .A2(n8384), .B1(
        n11060), .B2(n11078), .ZN(n4889) );
  AOI22_X1 U13810 ( .A1(n11130), .A2(n11059), .B1(n8384), .B2(
        \DataPath/RF/bus_reg_dataout[1290] ), .ZN(n4888) );
  AOI22_X1 U13811 ( .A1(\DataPath/RF/bus_reg_dataout[1291] ), .A2(n8384), .B1(
        n11060), .B2(n11080), .ZN(n4887) );
  AOI22_X1 U13812 ( .A1(\DataPath/RF/bus_reg_dataout[1292] ), .A2(n8384), .B1(
        n11060), .B2(n7781), .ZN(n4886) );
  AOI22_X1 U13813 ( .A1(\DataPath/RF/bus_reg_dataout[1293] ), .A2(n8384), .B1(
        n11060), .B2(n11082), .ZN(n4885) );
  AOI22_X1 U13814 ( .A1(\DataPath/RF/bus_reg_dataout[1294] ), .A2(n8384), .B1(
        n11060), .B2(n11109), .ZN(n4884) );
  AOI22_X1 U13815 ( .A1(\DataPath/RF/bus_reg_dataout[1295] ), .A2(n11061), 
        .B1(n11060), .B2(n7778), .ZN(n4883) );
  AOI22_X1 U13816 ( .A1(n11136), .A2(n11059), .B1(n8384), .B2(
        \DataPath/RF/bus_reg_dataout[1296] ), .ZN(n4882) );
  AOI22_X1 U13817 ( .A1(\DataPath/RF/bus_reg_dataout[1297] ), .A2(n8384), .B1(
        n11060), .B2(n7780), .ZN(n4881) );
  AOI22_X1 U13818 ( .A1(\DataPath/RF/bus_reg_dataout[1298] ), .A2(n11061), 
        .B1(n11060), .B2(n11085), .ZN(n4880) );
  AOI22_X1 U13819 ( .A1(\DataPath/RF/bus_reg_dataout[1299] ), .A2(n8384), .B1(
        n11060), .B2(n11086), .ZN(n4879) );
  AOI22_X1 U13820 ( .A1(\DataPath/RF/bus_reg_dataout[1300] ), .A2(n11061), 
        .B1(n11060), .B2(n11087), .ZN(n4878) );
  AOI22_X1 U13821 ( .A1(\DataPath/RF/bus_reg_dataout[1301] ), .A2(n8384), .B1(
        n11060), .B2(n11088), .ZN(n4877) );
  AOI22_X1 U13822 ( .A1(\DataPath/RF/bus_reg_dataout[1302] ), .A2(n8384), .B1(
        n11060), .B2(n11089), .ZN(n4876) );
  AOI22_X1 U13823 ( .A1(\DataPath/RF/bus_reg_dataout[1303] ), .A2(n8384), .B1(
        n11060), .B2(n11090), .ZN(n4875) );
  AOI22_X1 U13824 ( .A1(n11144), .A2(n11059), .B1(n8384), .B2(
        \DataPath/RF/bus_reg_dataout[1304] ), .ZN(n4874) );
  AOI22_X1 U13825 ( .A1(n11145), .A2(n11059), .B1(n11061), .B2(
        \DataPath/RF/bus_reg_dataout[1305] ), .ZN(n4873) );
  AOI22_X1 U13826 ( .A1(\DataPath/RF/bus_reg_dataout[1306] ), .A2(n11061), 
        .B1(n11060), .B2(n11091), .ZN(n4872) );
  AOI22_X1 U13827 ( .A1(\DataPath/RF/bus_reg_dataout[1307] ), .A2(n11061), 
        .B1(n11060), .B2(n11092), .ZN(n4871) );
  AOI22_X1 U13828 ( .A1(\DataPath/RF/bus_reg_dataout[1308] ), .A2(n8384), .B1(
        n11060), .B2(n11093), .ZN(n4870) );
  AOI22_X1 U13829 ( .A1(\DataPath/RF/bus_reg_dataout[1309] ), .A2(n8384), .B1(
        n11060), .B2(n11067), .ZN(n4869) );
  AOI22_X1 U13830 ( .A1(\DataPath/RF/bus_reg_dataout[1310] ), .A2(n8384), .B1(
        n11060), .B2(n11095), .ZN(n4868) );
  AOI22_X1 U13831 ( .A1(\DataPath/RF/bus_reg_dataout[1311] ), .A2(n11061), 
        .B1(n11060), .B2(n11096), .ZN(n4865) );
  OAI22_X1 U13832 ( .A1(n8271), .A2(n11338), .B1(n11339), .B2(n11640), .ZN(
        n11062) );
  AOI22_X1 U13833 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1248] ), 
        .B1(n11120), .B2(n11064), .ZN(n4863) );
  AOI22_X1 U13834 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1249] ), 
        .B1(n11121), .B2(n11064), .ZN(n4862) );
  NOR2_X1 U13835 ( .A1(RST), .A2(n11065), .ZN(n11063) );
  AOI22_X1 U13836 ( .A1(\DataPath/RF/bus_reg_dataout[1250] ), .A2(n11065), 
        .B1(n11063), .B2(n7779), .ZN(n4861) );
  AOI22_X1 U13837 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1251] ), 
        .B1(n11123), .B2(n11064), .ZN(n4860) );
  AOI22_X1 U13838 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1252] ), 
        .B1(n11124), .B2(n11064), .ZN(n4859) );
  AOI22_X1 U13839 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1253] ), 
        .B1(n11125), .B2(n11064), .ZN(n4858) );
  AOI22_X1 U13840 ( .A1(\DataPath/RF/bus_reg_dataout[1254] ), .A2(n11065), 
        .B1(n11063), .B2(n11076), .ZN(n4857) );
  AOI22_X1 U13841 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1255] ), 
        .B1(n11127), .B2(n11064), .ZN(n4856) );
  AOI22_X1 U13842 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1256] ), 
        .B1(n11128), .B2(n11064), .ZN(n4855) );
  AOI22_X1 U13843 ( .A1(\DataPath/RF/bus_reg_dataout[1257] ), .A2(n11065), 
        .B1(n11063), .B2(n11078), .ZN(n4854) );
  AOI22_X1 U13844 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1258] ), 
        .B1(n11130), .B2(n11064), .ZN(n4853) );
  AOI22_X1 U13845 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1259] ), 
        .B1(n11131), .B2(n11064), .ZN(n4852) );
  AOI22_X1 U13846 ( .A1(\DataPath/RF/bus_reg_dataout[1260] ), .A2(n11065), 
        .B1(n11063), .B2(n7781), .ZN(n4851) );
  AOI22_X1 U13847 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1261] ), 
        .B1(n11133), .B2(n11064), .ZN(n4850) );
  AOI22_X1 U13848 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1262] ), 
        .B1(n11134), .B2(n11064), .ZN(n4849) );
  AOI22_X1 U13849 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1263] ), 
        .B1(n11135), .B2(n11064), .ZN(n4848) );
  AOI22_X1 U13850 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1264] ), 
        .B1(n11136), .B2(n11064), .ZN(n4847) );
  AOI22_X1 U13851 ( .A1(\DataPath/RF/bus_reg_dataout[1265] ), .A2(n11065), 
        .B1(n11063), .B2(n7780), .ZN(n4846) );
  AOI22_X1 U13852 ( .A1(\DataPath/RF/bus_reg_dataout[1266] ), .A2(n11065), 
        .B1(n11063), .B2(n11085), .ZN(n4845) );
  AOI22_X1 U13853 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1267] ), 
        .B1(n11139), .B2(n11064), .ZN(n4844) );
  AOI22_X1 U13854 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1268] ), 
        .B1(n11140), .B2(n11064), .ZN(n4843) );
  AOI22_X1 U13855 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1269] ), 
        .B1(n11141), .B2(n11064), .ZN(n4842) );
  AOI22_X1 U13856 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1270] ), 
        .B1(n11142), .B2(n11064), .ZN(n4841) );
  AOI22_X1 U13857 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1271] ), 
        .B1(n11143), .B2(n11064), .ZN(n4840) );
  AOI22_X1 U13858 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1272] ), 
        .B1(n11144), .B2(n11064), .ZN(n4839) );
  AOI22_X1 U13859 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1273] ), 
        .B1(n11145), .B2(n11064), .ZN(n4838) );
  AOI22_X1 U13860 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1274] ), 
        .B1(n11146), .B2(n11064), .ZN(n4837) );
  AOI22_X1 U13861 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1275] ), 
        .B1(n11147), .B2(n11064), .ZN(n4836) );
  AOI22_X1 U13862 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1276] ), 
        .B1(n11148), .B2(n11064), .ZN(n4835) );
  AOI22_X1 U13863 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1277] ), 
        .B1(n11149), .B2(n11064), .ZN(n4834) );
  AOI22_X1 U13864 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1278] ), 
        .B1(n11150), .B2(n11064), .ZN(n4833) );
  AOI22_X1 U13865 ( .A1(n11065), .A2(\DataPath/RF/bus_reg_dataout[1279] ), 
        .B1(n11152), .B2(n11064), .ZN(n4830) );
  AOI22_X1 U13866 ( .A1(\DataPath/RF/bus_reg_dataout[1216] ), .A2(n8385), .B1(
        n11068), .B2(n11071), .ZN(n4828) );
  AOI22_X1 U13867 ( .A1(\DataPath/RF/bus_reg_dataout[1217] ), .A2(n8385), .B1(
        n11068), .B2(n11072), .ZN(n4827) );
  AOI22_X1 U13868 ( .A1(\DataPath/RF/bus_reg_dataout[1218] ), .A2(n11069), 
        .B1(n11068), .B2(n7779), .ZN(n4826) );
  AOI22_X1 U13869 ( .A1(\DataPath/RF/bus_reg_dataout[1219] ), .A2(n8385), .B1(
        n11068), .B2(n11107), .ZN(n4825) );
  AOI22_X1 U13870 ( .A1(\DataPath/RF/bus_reg_dataout[1220] ), .A2(n11069), 
        .B1(n11068), .B2(n11074), .ZN(n4824) );
  AOI22_X1 U13871 ( .A1(\DataPath/RF/bus_reg_dataout[1221] ), .A2(n8385), .B1(
        n11068), .B2(n11075), .ZN(n4823) );
  AOI22_X1 U13872 ( .A1(\DataPath/RF/bus_reg_dataout[1222] ), .A2(n8385), .B1(
        n11068), .B2(n11076), .ZN(n4822) );
  AOI22_X1 U13873 ( .A1(n11127), .A2(n11066), .B1(n8385), .B2(
        \DataPath/RF/bus_reg_dataout[1223] ), .ZN(n4821) );
  AOI22_X1 U13874 ( .A1(\DataPath/RF/bus_reg_dataout[1224] ), .A2(n8385), .B1(
        n11068), .B2(n11077), .ZN(n4820) );
  AOI22_X1 U13875 ( .A1(\DataPath/RF/bus_reg_dataout[1225] ), .A2(n11069), 
        .B1(n11068), .B2(n11078), .ZN(n4819) );
  AOI22_X1 U13876 ( .A1(\DataPath/RF/bus_reg_dataout[1226] ), .A2(n8385), .B1(
        n11068), .B2(n11079), .ZN(n4818) );
  AOI22_X1 U13877 ( .A1(n11131), .A2(n11066), .B1(n8385), .B2(
        \DataPath/RF/bus_reg_dataout[1227] ), .ZN(n4817) );
  AOI22_X1 U13878 ( .A1(\DataPath/RF/bus_reg_dataout[1228] ), .A2(n8385), .B1(
        n11068), .B2(n7781), .ZN(n4816) );
  AOI22_X1 U13879 ( .A1(\DataPath/RF/bus_reg_dataout[1229] ), .A2(n8385), .B1(
        n11068), .B2(n11082), .ZN(n4815) );
  AOI22_X1 U13880 ( .A1(\DataPath/RF/bus_reg_dataout[1230] ), .A2(n8385), .B1(
        n11068), .B2(n11109), .ZN(n4814) );
  AOI22_X1 U13881 ( .A1(\DataPath/RF/bus_reg_dataout[1231] ), .A2(n8385), .B1(
        n11068), .B2(n7778), .ZN(n4813) );
  AOI22_X1 U13882 ( .A1(n11136), .A2(n11066), .B1(n11069), .B2(
        \DataPath/RF/bus_reg_dataout[1232] ), .ZN(n4812) );
  AOI22_X1 U13883 ( .A1(\DataPath/RF/bus_reg_dataout[1233] ), .A2(n8385), .B1(
        n11068), .B2(n7780), .ZN(n4811) );
  AOI22_X1 U13884 ( .A1(\DataPath/RF/bus_reg_dataout[1234] ), .A2(n8385), .B1(
        n11068), .B2(n11085), .ZN(n4810) );
  AOI22_X1 U13885 ( .A1(\DataPath/RF/bus_reg_dataout[1235] ), .A2(n8385), .B1(
        n11068), .B2(n11086), .ZN(n4809) );
  AOI22_X1 U13886 ( .A1(n11140), .A2(n11066), .B1(n8385), .B2(
        \DataPath/RF/bus_reg_dataout[1236] ), .ZN(n4808) );
  AOI22_X1 U13887 ( .A1(n11141), .A2(n11066), .B1(n11069), .B2(
        \DataPath/RF/bus_reg_dataout[1237] ), .ZN(n4807) );
  AOI22_X1 U13888 ( .A1(\DataPath/RF/bus_reg_dataout[1238] ), .A2(n11069), 
        .B1(n11068), .B2(n11089), .ZN(n4806) );
  AOI22_X1 U13889 ( .A1(\DataPath/RF/bus_reg_dataout[1239] ), .A2(n8385), .B1(
        n11068), .B2(n11090), .ZN(n4805) );
  AOI22_X1 U13890 ( .A1(n11144), .A2(n11066), .B1(n8385), .B2(
        \DataPath/RF/bus_reg_dataout[1240] ), .ZN(n4804) );
  AOI22_X1 U13891 ( .A1(\DataPath/RF/bus_reg_dataout[1241] ), .A2(n8385), .B1(
        n11068), .B2(n11111), .ZN(n4803) );
  AOI22_X1 U13892 ( .A1(\DataPath/RF/bus_reg_dataout[1242] ), .A2(n11069), 
        .B1(n11068), .B2(n11091), .ZN(n4802) );
  AOI22_X1 U13893 ( .A1(n11147), .A2(n11066), .B1(n11069), .B2(
        \DataPath/RF/bus_reg_dataout[1243] ), .ZN(n4801) );
  AOI22_X1 U13894 ( .A1(\DataPath/RF/bus_reg_dataout[1244] ), .A2(n8385), .B1(
        n11068), .B2(n11093), .ZN(n4800) );
  AOI22_X1 U13895 ( .A1(\DataPath/RF/bus_reg_dataout[1245] ), .A2(n11069), 
        .B1(n11068), .B2(n11067), .ZN(n4799) );
  AOI22_X1 U13896 ( .A1(\DataPath/RF/bus_reg_dataout[1246] ), .A2(n8385), .B1(
        n11068), .B2(n11095), .ZN(n4798) );
  AOI22_X1 U13897 ( .A1(\DataPath/RF/bus_reg_dataout[1247] ), .A2(n11069), 
        .B1(n11068), .B2(n11096), .ZN(n4795) );
  OAI222_X1 U13898 ( .A1(n11352), .A2(n11102), .B1(n11070), .B2(n8271), .C1(
        n11353), .C2(n11640), .ZN(n11094) );
  AOI22_X1 U13899 ( .A1(\DataPath/RF/bus_reg_dataout[1184] ), .A2(n8386), .B1(
        n11097), .B2(n11071), .ZN(n4793) );
  AOI22_X1 U13900 ( .A1(\DataPath/RF/bus_reg_dataout[1185] ), .A2(n8386), .B1(
        n11097), .B2(n11072), .ZN(n4792) );
  AOI22_X1 U13901 ( .A1(\DataPath/RF/bus_reg_dataout[1186] ), .A2(n11098), 
        .B1(n11097), .B2(n7779), .ZN(n4791) );
  AOI22_X1 U13902 ( .A1(\DataPath/RF/bus_reg_dataout[1187] ), .A2(n11098), 
        .B1(n11097), .B2(n11107), .ZN(n4790) );
  AOI22_X1 U13903 ( .A1(\DataPath/RF/bus_reg_dataout[1188] ), .A2(n11098), 
        .B1(n11097), .B2(n11074), .ZN(n4789) );
  AOI22_X1 U13904 ( .A1(\DataPath/RF/bus_reg_dataout[1189] ), .A2(n8386), .B1(
        n11097), .B2(n11075), .ZN(n4788) );
  AOI22_X1 U13905 ( .A1(\DataPath/RF/bus_reg_dataout[1190] ), .A2(n8386), .B1(
        n11097), .B2(n11076), .ZN(n4787) );
  AOI22_X1 U13906 ( .A1(\DataPath/RF/bus_reg_dataout[1191] ), .A2(n8386), .B1(
        n11097), .B2(n11108), .ZN(n4786) );
  AOI22_X1 U13907 ( .A1(\DataPath/RF/bus_reg_dataout[1192] ), .A2(n11098), 
        .B1(n11097), .B2(n11077), .ZN(n4785) );
  AOI22_X1 U13908 ( .A1(\DataPath/RF/bus_reg_dataout[1193] ), .A2(n11098), 
        .B1(n11097), .B2(n11078), .ZN(n4784) );
  AOI22_X1 U13909 ( .A1(\DataPath/RF/bus_reg_dataout[1194] ), .A2(n8386), .B1(
        n11097), .B2(n11079), .ZN(n4783) );
  AOI22_X1 U13910 ( .A1(\DataPath/RF/bus_reg_dataout[1195] ), .A2(n8386), .B1(
        n11097), .B2(n11080), .ZN(n4782) );
  AOI22_X1 U13911 ( .A1(\DataPath/RF/bus_reg_dataout[1196] ), .A2(n11098), 
        .B1(n11097), .B2(n7781), .ZN(n4781) );
  AOI22_X1 U13912 ( .A1(\DataPath/RF/bus_reg_dataout[1197] ), .A2(n11098), 
        .B1(n11097), .B2(n11082), .ZN(n4780) );
  AOI22_X1 U13913 ( .A1(\DataPath/RF/bus_reg_dataout[1198] ), .A2(n8386), .B1(
        n11097), .B2(n11109), .ZN(n4779) );
  AOI22_X1 U13914 ( .A1(\DataPath/RF/bus_reg_dataout[1199] ), .A2(n8386), .B1(
        n11097), .B2(n7778), .ZN(n4778) );
  AOI22_X1 U13915 ( .A1(\DataPath/RF/bus_reg_dataout[1200] ), .A2(n8386), .B1(
        n11097), .B2(n11083), .ZN(n4777) );
  AOI22_X1 U13916 ( .A1(\DataPath/RF/bus_reg_dataout[1201] ), .A2(n8386), .B1(
        n11097), .B2(n7780), .ZN(n4776) );
  AOI22_X1 U13917 ( .A1(\DataPath/RF/bus_reg_dataout[1202] ), .A2(n11098), 
        .B1(n11097), .B2(n11085), .ZN(n4775) );
  AOI22_X1 U13918 ( .A1(\DataPath/RF/bus_reg_dataout[1203] ), .A2(n8386), .B1(
        n11097), .B2(n11086), .ZN(n4774) );
  AOI22_X1 U13919 ( .A1(\DataPath/RF/bus_reg_dataout[1204] ), .A2(n8386), .B1(
        n11097), .B2(n11087), .ZN(n4773) );
  AOI22_X1 U13920 ( .A1(\DataPath/RF/bus_reg_dataout[1205] ), .A2(n11098), 
        .B1(n11097), .B2(n11088), .ZN(n4772) );
  AOI22_X1 U13921 ( .A1(\DataPath/RF/bus_reg_dataout[1206] ), .A2(n8386), .B1(
        n11097), .B2(n11089), .ZN(n4771) );
  AOI22_X1 U13922 ( .A1(\DataPath/RF/bus_reg_dataout[1207] ), .A2(n8386), .B1(
        n11097), .B2(n11090), .ZN(n4770) );
  AOI22_X1 U13923 ( .A1(n11144), .A2(n11094), .B1(n8386), .B2(
        \DataPath/RF/bus_reg_dataout[1208] ), .ZN(n4769) );
  AOI22_X1 U13924 ( .A1(\DataPath/RF/bus_reg_dataout[1209] ), .A2(n8386), .B1(
        n11097), .B2(n11111), .ZN(n4768) );
  AOI22_X1 U13925 ( .A1(\DataPath/RF/bus_reg_dataout[1210] ), .A2(n8386), .B1(
        n11097), .B2(n11091), .ZN(n4767) );
  AOI22_X1 U13926 ( .A1(\DataPath/RF/bus_reg_dataout[1211] ), .A2(n11098), 
        .B1(n11097), .B2(n11092), .ZN(n4766) );
  AOI22_X1 U13927 ( .A1(\DataPath/RF/bus_reg_dataout[1212] ), .A2(n8386), .B1(
        n11097), .B2(n11093), .ZN(n4765) );
  AOI22_X1 U13928 ( .A1(n11149), .A2(n11094), .B1(n8386), .B2(
        \DataPath/RF/bus_reg_dataout[1213] ), .ZN(n4764) );
  AOI22_X1 U13929 ( .A1(\DataPath/RF/bus_reg_dataout[1214] ), .A2(n8386), .B1(
        n11097), .B2(n11095), .ZN(n4763) );
  AOI22_X1 U13930 ( .A1(\DataPath/RF/bus_reg_dataout[1215] ), .A2(n8386), .B1(
        n11097), .B2(n11096), .ZN(n4760) );
  OAI22_X1 U13931 ( .A1(n11640), .A2(n11360), .B1(n11102), .B2(n11361), .ZN(
        n11099) );
  AOI22_X1 U13932 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1152] ), 
        .B1(n11120), .B2(n11100), .ZN(n4758) );
  AOI22_X1 U13933 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1153] ), 
        .B1(n11121), .B2(n11100), .ZN(n4757) );
  AOI22_X1 U13934 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1154] ), 
        .B1(n11122), .B2(n11100), .ZN(n4756) );
  AOI22_X1 U13935 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1155] ), 
        .B1(n11123), .B2(n11100), .ZN(n4755) );
  AOI22_X1 U13936 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1156] ), 
        .B1(n11124), .B2(n11100), .ZN(n4754) );
  AOI22_X1 U13937 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1157] ), 
        .B1(n11125), .B2(n11100), .ZN(n4753) );
  AOI22_X1 U13938 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1158] ), 
        .B1(n11126), .B2(n11100), .ZN(n4752) );
  AOI22_X1 U13939 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1159] ), 
        .B1(n11127), .B2(n11100), .ZN(n4751) );
  AOI22_X1 U13940 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1160] ), 
        .B1(n11128), .B2(n11100), .ZN(n4750) );
  AOI22_X1 U13941 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1161] ), 
        .B1(n11129), .B2(n11100), .ZN(n4749) );
  AOI22_X1 U13942 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1162] ), 
        .B1(n11130), .B2(n11100), .ZN(n4748) );
  AOI22_X1 U13943 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1163] ), 
        .B1(n11131), .B2(n11100), .ZN(n4747) );
  AOI22_X1 U13944 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1164] ), 
        .B1(n11132), .B2(n11100), .ZN(n4746) );
  AOI22_X1 U13945 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1165] ), 
        .B1(n11133), .B2(n11100), .ZN(n4745) );
  AOI22_X1 U13946 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1166] ), 
        .B1(n11134), .B2(n11100), .ZN(n4744) );
  AOI22_X1 U13947 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1167] ), 
        .B1(n11135), .B2(n11100), .ZN(n4743) );
  AOI22_X1 U13948 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1168] ), 
        .B1(n11136), .B2(n11100), .ZN(n4742) );
  AOI22_X1 U13949 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1169] ), 
        .B1(n11137), .B2(n11100), .ZN(n4741) );
  AOI22_X1 U13950 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1170] ), 
        .B1(n11138), .B2(n11100), .ZN(n4740) );
  AOI22_X1 U13951 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1171] ), 
        .B1(n11139), .B2(n11100), .ZN(n4739) );
  AOI22_X1 U13952 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1172] ), 
        .B1(n11140), .B2(n11100), .ZN(n4738) );
  AOI22_X1 U13953 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1173] ), 
        .B1(n11141), .B2(n11100), .ZN(n4737) );
  AOI22_X1 U13954 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1174] ), 
        .B1(n11142), .B2(n11100), .ZN(n4736) );
  AOI22_X1 U13955 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1175] ), 
        .B1(n11143), .B2(n11100), .ZN(n4735) );
  AOI22_X1 U13956 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1176] ), 
        .B1(n11144), .B2(n11100), .ZN(n4734) );
  AOI22_X1 U13957 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1177] ), 
        .B1(n11145), .B2(n11100), .ZN(n4733) );
  AOI22_X1 U13958 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1178] ), 
        .B1(n11146), .B2(n11100), .ZN(n4732) );
  AOI22_X1 U13959 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1179] ), 
        .B1(n11147), .B2(n11100), .ZN(n4731) );
  AOI22_X1 U13960 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1180] ), 
        .B1(n11148), .B2(n11100), .ZN(n4730) );
  AOI22_X1 U13961 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1181] ), 
        .B1(n11149), .B2(n11100), .ZN(n4729) );
  AOI22_X1 U13962 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1182] ), 
        .B1(n11150), .B2(n11100), .ZN(n4728) );
  AOI22_X1 U13963 ( .A1(n11101), .A2(\DataPath/RF/bus_reg_dataout[1183] ), 
        .B1(n11152), .B2(n11100), .ZN(n4725) );
  OAI22_X1 U13964 ( .A1(n11640), .A2(n11367), .B1(n11102), .B2(n11366), .ZN(
        n11103) );
  AOI22_X1 U13965 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1120] ), 
        .B1(n11120), .B2(n11104), .ZN(n4723) );
  AOI22_X1 U13966 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1121] ), 
        .B1(n11121), .B2(n11104), .ZN(n4722) );
  AOI22_X1 U13967 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1122] ), 
        .B1(n11122), .B2(n11104), .ZN(n4721) );
  AOI22_X1 U13968 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1123] ), 
        .B1(n11123), .B2(n11104), .ZN(n4720) );
  AOI22_X1 U13969 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1124] ), 
        .B1(n11124), .B2(n11104), .ZN(n4719) );
  AOI22_X1 U13970 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1125] ), 
        .B1(n11125), .B2(n11104), .ZN(n4718) );
  AOI22_X1 U13971 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1126] ), 
        .B1(n11126), .B2(n11104), .ZN(n4717) );
  AOI22_X1 U13972 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1127] ), 
        .B1(n11127), .B2(n11104), .ZN(n4716) );
  AOI22_X1 U13973 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1128] ), 
        .B1(n11128), .B2(n11104), .ZN(n4715) );
  AOI22_X1 U13974 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1129] ), 
        .B1(n11129), .B2(n11104), .ZN(n4714) );
  AOI22_X1 U13975 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1130] ), 
        .B1(n11130), .B2(n11104), .ZN(n4713) );
  AOI22_X1 U13976 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1131] ), 
        .B1(n11131), .B2(n11104), .ZN(n4712) );
  AOI22_X1 U13977 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1132] ), 
        .B1(n11132), .B2(n11104), .ZN(n4711) );
  AOI22_X1 U13978 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1133] ), 
        .B1(n11133), .B2(n11104), .ZN(n4710) );
  AOI22_X1 U13979 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1134] ), 
        .B1(n11134), .B2(n11104), .ZN(n4709) );
  AOI22_X1 U13980 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1135] ), 
        .B1(n11135), .B2(n11104), .ZN(n4708) );
  AOI22_X1 U13981 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1136] ), 
        .B1(n11136), .B2(n11104), .ZN(n4707) );
  AOI22_X1 U13982 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1137] ), 
        .B1(n11137), .B2(n11104), .ZN(n4706) );
  AOI22_X1 U13983 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1138] ), 
        .B1(n11138), .B2(n11104), .ZN(n4705) );
  AOI22_X1 U13984 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1139] ), 
        .B1(n11139), .B2(n11104), .ZN(n4704) );
  AOI22_X1 U13985 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1140] ), 
        .B1(n11140), .B2(n11104), .ZN(n4703) );
  AOI22_X1 U13986 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1141] ), 
        .B1(n11141), .B2(n11104), .ZN(n4702) );
  AOI22_X1 U13987 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1142] ), 
        .B1(n11142), .B2(n11104), .ZN(n4701) );
  AOI22_X1 U13988 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1143] ), 
        .B1(n11143), .B2(n11104), .ZN(n4700) );
  AOI22_X1 U13989 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1144] ), 
        .B1(n11144), .B2(n11104), .ZN(n4699) );
  AOI22_X1 U13990 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1145] ), 
        .B1(n11145), .B2(n11104), .ZN(n4698) );
  AOI22_X1 U13991 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1146] ), 
        .B1(n11146), .B2(n11104), .ZN(n4697) );
  AOI22_X1 U13992 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1147] ), 
        .B1(n11147), .B2(n11104), .ZN(n4696) );
  AOI22_X1 U13993 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1148] ), 
        .B1(n11148), .B2(n11104), .ZN(n4695) );
  AOI22_X1 U13994 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1149] ), 
        .B1(n11149), .B2(n11104), .ZN(n4694) );
  AOI22_X1 U13995 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1150] ), 
        .B1(n11150), .B2(n11104), .ZN(n4693) );
  AOI22_X1 U13996 ( .A1(n11105), .A2(\DataPath/RF/bus_reg_dataout[1151] ), 
        .B1(n11152), .B2(n11104), .ZN(n4690) );
  OAI22_X1 U13997 ( .A1(n8271), .A2(n11374), .B1(n11375), .B2(n11640), .ZN(
        n11106) );
  AOI22_X1 U13998 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1088] ), 
        .B1(n11120), .B2(n11113), .ZN(n4688) );
  AOI22_X1 U13999 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1089] ), 
        .B1(n11121), .B2(n11113), .ZN(n4687) );
  AOI22_X1 U14000 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1090] ), 
        .B1(n11122), .B2(n11113), .ZN(n4686) );
  NOR2_X1 U14001 ( .A1(RST), .A2(n11114), .ZN(n11112) );
  AOI22_X1 U14002 ( .A1(\DataPath/RF/bus_reg_dataout[1091] ), .A2(n11114), 
        .B1(n11112), .B2(n11107), .ZN(n4685) );
  AOI22_X1 U14003 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1092] ), 
        .B1(n11124), .B2(n11113), .ZN(n4684) );
  AOI22_X1 U14004 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1093] ), 
        .B1(n11125), .B2(n11113), .ZN(n4683) );
  AOI22_X1 U14005 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1094] ), 
        .B1(n11126), .B2(n11113), .ZN(n4682) );
  AOI22_X1 U14006 ( .A1(\DataPath/RF/bus_reg_dataout[1095] ), .A2(n11114), 
        .B1(n11112), .B2(n11108), .ZN(n4681) );
  AOI22_X1 U14007 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1096] ), 
        .B1(n11128), .B2(n11113), .ZN(n4680) );
  AOI22_X1 U14008 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1097] ), 
        .B1(n11129), .B2(n11113), .ZN(n4679) );
  AOI22_X1 U14009 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1098] ), 
        .B1(n11130), .B2(n11113), .ZN(n4678) );
  AOI22_X1 U14010 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1099] ), 
        .B1(n11131), .B2(n11113), .ZN(n4677) );
  AOI22_X1 U14011 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1100] ), 
        .B1(n11132), .B2(n11113), .ZN(n4676) );
  AOI22_X1 U14012 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1101] ), 
        .B1(n11133), .B2(n11113), .ZN(n4675) );
  AOI22_X1 U14013 ( .A1(\DataPath/RF/bus_reg_dataout[1102] ), .A2(n11114), 
        .B1(n11112), .B2(n11109), .ZN(n4674) );
  AOI22_X1 U14014 ( .A1(\DataPath/RF/bus_reg_dataout[1103] ), .A2(n11114), 
        .B1(n11112), .B2(n7778), .ZN(n4673) );
  AOI22_X1 U14015 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1104] ), 
        .B1(n11136), .B2(n11113), .ZN(n4672) );
  AOI22_X1 U14016 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1105] ), 
        .B1(n11137), .B2(n11113), .ZN(n4671) );
  AOI22_X1 U14017 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1106] ), 
        .B1(n11138), .B2(n11113), .ZN(n4670) );
  AOI22_X1 U14018 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1107] ), 
        .B1(n11139), .B2(n11113), .ZN(n4669) );
  AOI22_X1 U14019 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1108] ), 
        .B1(n11140), .B2(n11113), .ZN(n4668) );
  AOI22_X1 U14020 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1109] ), 
        .B1(n11141), .B2(n11113), .ZN(n4667) );
  AOI22_X1 U14021 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1110] ), 
        .B1(n11142), .B2(n11113), .ZN(n4666) );
  AOI22_X1 U14022 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1111] ), 
        .B1(n11143), .B2(n11113), .ZN(n4665) );
  AOI22_X1 U14023 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1112] ), 
        .B1(n11144), .B2(n11113), .ZN(n4664) );
  AOI22_X1 U14024 ( .A1(\DataPath/RF/bus_reg_dataout[1113] ), .A2(n11114), 
        .B1(n11112), .B2(n11111), .ZN(n4663) );
  AOI22_X1 U14025 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1114] ), 
        .B1(n11146), .B2(n11113), .ZN(n4662) );
  AOI22_X1 U14026 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1115] ), 
        .B1(n11147), .B2(n11113), .ZN(n4661) );
  AOI22_X1 U14027 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1116] ), 
        .B1(n11148), .B2(n11113), .ZN(n4660) );
  AOI22_X1 U14028 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1117] ), 
        .B1(n11149), .B2(n11113), .ZN(n4659) );
  AOI22_X1 U14029 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1118] ), 
        .B1(n11150), .B2(n11113), .ZN(n4658) );
  AOI22_X1 U14030 ( .A1(n11114), .A2(\DataPath/RF/bus_reg_dataout[1119] ), 
        .B1(n11152), .B2(n11113), .ZN(n4655) );
  OAI22_X1 U14031 ( .A1(n8271), .A2(n11406), .B1(n11407), .B2(n11640), .ZN(
        n11115) );
  AOI22_X1 U14032 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1056] ), 
        .B1(n11120), .B2(n11116), .ZN(n4653) );
  AOI22_X1 U14033 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1057] ), 
        .B1(n11121), .B2(n11116), .ZN(n4652) );
  AOI22_X1 U14034 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1058] ), 
        .B1(n11122), .B2(n11116), .ZN(n4651) );
  AOI22_X1 U14035 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1059] ), 
        .B1(n11123), .B2(n11116), .ZN(n4650) );
  AOI22_X1 U14036 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1060] ), 
        .B1(n11124), .B2(n11116), .ZN(n4649) );
  AOI22_X1 U14037 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1061] ), 
        .B1(n11125), .B2(n11116), .ZN(n4648) );
  AOI22_X1 U14038 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1062] ), 
        .B1(n11126), .B2(n11116), .ZN(n4647) );
  AOI22_X1 U14039 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1063] ), 
        .B1(n11127), .B2(n11116), .ZN(n4646) );
  AOI22_X1 U14040 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1064] ), 
        .B1(n11128), .B2(n11116), .ZN(n4645) );
  AOI22_X1 U14041 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1065] ), 
        .B1(n11129), .B2(n11116), .ZN(n4644) );
  AOI22_X1 U14042 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1066] ), 
        .B1(n11130), .B2(n11116), .ZN(n4643) );
  AOI22_X1 U14043 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1067] ), 
        .B1(n11131), .B2(n11116), .ZN(n4642) );
  AOI22_X1 U14044 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1068] ), 
        .B1(n11132), .B2(n11116), .ZN(n4641) );
  AOI22_X1 U14045 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1069] ), 
        .B1(n11133), .B2(n11116), .ZN(n4640) );
  AOI22_X1 U14046 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1070] ), 
        .B1(n11134), .B2(n11116), .ZN(n4639) );
  AOI22_X1 U14047 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1071] ), 
        .B1(n11135), .B2(n11116), .ZN(n4638) );
  AOI22_X1 U14048 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1072] ), 
        .B1(n11136), .B2(n11116), .ZN(n4637) );
  AOI22_X1 U14049 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1073] ), 
        .B1(n11137), .B2(n11116), .ZN(n4636) );
  AOI22_X1 U14050 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1074] ), 
        .B1(n11138), .B2(n11116), .ZN(n4635) );
  AOI22_X1 U14051 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1075] ), 
        .B1(n11139), .B2(n11116), .ZN(n4634) );
  AOI22_X1 U14052 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1076] ), 
        .B1(n11140), .B2(n11116), .ZN(n4633) );
  AOI22_X1 U14053 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1077] ), 
        .B1(n11141), .B2(n11116), .ZN(n4632) );
  AOI22_X1 U14054 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1078] ), 
        .B1(n11142), .B2(n11116), .ZN(n4631) );
  AOI22_X1 U14055 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1079] ), 
        .B1(n11143), .B2(n11116), .ZN(n4630) );
  AOI22_X1 U14056 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1080] ), 
        .B1(n11144), .B2(n11116), .ZN(n4629) );
  AOI22_X1 U14057 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1081] ), 
        .B1(n11145), .B2(n11116), .ZN(n4628) );
  AOI22_X1 U14058 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1082] ), 
        .B1(n11146), .B2(n11116), .ZN(n4627) );
  AOI22_X1 U14059 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1083] ), 
        .B1(n11147), .B2(n11116), .ZN(n4626) );
  AOI22_X1 U14060 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1084] ), 
        .B1(n11148), .B2(n11116), .ZN(n4625) );
  AOI22_X1 U14061 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1085] ), 
        .B1(n11149), .B2(n11116), .ZN(n4624) );
  AOI22_X1 U14062 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1086] ), 
        .B1(n11150), .B2(n11116), .ZN(n4623) );
  AOI22_X1 U14063 ( .A1(n11117), .A2(\DataPath/RF/bus_reg_dataout[1087] ), 
        .B1(n11152), .B2(n11116), .ZN(n4620) );
  OAI22_X1 U14064 ( .A1(n8271), .A2(n11414), .B1(n11416), .B2(n11640), .ZN(
        n11118) );
  AOI22_X1 U14065 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1024] ), 
        .B1(n11120), .B2(n11151), .ZN(n4616) );
  AOI22_X1 U14066 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1025] ), 
        .B1(n11121), .B2(n11151), .ZN(n4614) );
  AOI22_X1 U14067 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1026] ), 
        .B1(n11122), .B2(n11151), .ZN(n4612) );
  AOI22_X1 U14068 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1027] ), 
        .B1(n11123), .B2(n11151), .ZN(n4610) );
  AOI22_X1 U14069 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1028] ), 
        .B1(n11124), .B2(n11151), .ZN(n4608) );
  AOI22_X1 U14070 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1029] ), 
        .B1(n11125), .B2(n11151), .ZN(n4606) );
  AOI22_X1 U14071 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1030] ), 
        .B1(n11126), .B2(n11151), .ZN(n4604) );
  AOI22_X1 U14072 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1031] ), 
        .B1(n11127), .B2(n11151), .ZN(n4602) );
  AOI22_X1 U14073 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1032] ), 
        .B1(n11128), .B2(n11151), .ZN(n4600) );
  AOI22_X1 U14074 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1033] ), 
        .B1(n11129), .B2(n11151), .ZN(n4598) );
  AOI22_X1 U14075 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1034] ), 
        .B1(n11130), .B2(n11151), .ZN(n4596) );
  AOI22_X1 U14076 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1035] ), 
        .B1(n11131), .B2(n11151), .ZN(n4594) );
  AOI22_X1 U14077 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1036] ), 
        .B1(n11132), .B2(n11151), .ZN(n4592) );
  AOI22_X1 U14078 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1037] ), 
        .B1(n11133), .B2(n11151), .ZN(n4590) );
  AOI22_X1 U14079 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1038] ), 
        .B1(n11134), .B2(n11151), .ZN(n4588) );
  AOI22_X1 U14080 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1039] ), 
        .B1(n11135), .B2(n11151), .ZN(n4586) );
  AOI22_X1 U14081 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1040] ), 
        .B1(n11136), .B2(n11151), .ZN(n4584) );
  AOI22_X1 U14082 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1041] ), 
        .B1(n11137), .B2(n11151), .ZN(n4582) );
  AOI22_X1 U14083 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1042] ), 
        .B1(n11138), .B2(n11151), .ZN(n4580) );
  AOI22_X1 U14084 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1043] ), 
        .B1(n11139), .B2(n11151), .ZN(n4578) );
  AOI22_X1 U14085 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1044] ), 
        .B1(n11140), .B2(n11151), .ZN(n4576) );
  AOI22_X1 U14086 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1045] ), 
        .B1(n11141), .B2(n11151), .ZN(n4574) );
  AOI22_X1 U14087 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1046] ), 
        .B1(n11142), .B2(n11151), .ZN(n4572) );
  AOI22_X1 U14088 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1047] ), 
        .B1(n11143), .B2(n11151), .ZN(n4570) );
  AOI22_X1 U14089 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1048] ), 
        .B1(n11144), .B2(n11151), .ZN(n4568) );
  AOI22_X1 U14090 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1049] ), 
        .B1(n11145), .B2(n11151), .ZN(n4566) );
  AOI22_X1 U14091 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1050] ), 
        .B1(n11146), .B2(n11151), .ZN(n4564) );
  AOI22_X1 U14092 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1051] ), 
        .B1(n11147), .B2(n11151), .ZN(n4562) );
  AOI22_X1 U14093 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1052] ), 
        .B1(n11148), .B2(n11151), .ZN(n4560) );
  AOI22_X1 U14094 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1053] ), 
        .B1(n11149), .B2(n11151), .ZN(n4558) );
  AOI22_X1 U14095 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1054] ), 
        .B1(n11150), .B2(n11151), .ZN(n4556) );
  AOI22_X1 U14096 ( .A1(n11153), .A2(\DataPath/RF/bus_reg_dataout[1055] ), 
        .B1(n11152), .B2(n11151), .ZN(n4552) );
  OAI22_X1 U14097 ( .A1(n11640), .A2(n11737), .B1(n11736), .B2(n11211), .ZN(
        n11154) );
  AOI22_X1 U14098 ( .A1(n7761), .A2(n11272), .B1(n11479), .B2(n11211), .ZN(
        n11174) );
  AOI22_X1 U14099 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[992] ), .B1(
        n11155), .B2(n11174), .ZN(n4550) );
  AOI22_X1 U14100 ( .A1(n7761), .A2(n11273), .B1(n11480), .B2(n11211), .ZN(
        n11213) );
  AOI22_X1 U14101 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[993] ), .B1(
        n11155), .B2(n11213), .ZN(n4549) );
  AOI22_X1 U14102 ( .A1(n7761), .A2(n11274), .B1(n11481), .B2(n11211), .ZN(
        n11203) );
  AOI22_X1 U14103 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[994] ), .B1(
        n11155), .B2(n11203), .ZN(n4548) );
  AOI22_X1 U14104 ( .A1(n7761), .A2(n11275), .B1(n11482), .B2(n11211), .ZN(
        n11175) );
  AOI22_X1 U14105 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[995] ), .B1(
        n11155), .B2(n11175), .ZN(n4547) );
  AOI22_X1 U14106 ( .A1(n7761), .A2(n11276), .B1(n11483), .B2(n11211), .ZN(
        n11189) );
  AOI22_X1 U14107 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[996] ), .B1(
        n11155), .B2(n11189), .ZN(n4546) );
  AOI22_X1 U14108 ( .A1(n7761), .A2(n11277), .B1(n11484), .B2(n11211), .ZN(
        n11176) );
  AOI22_X1 U14109 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[997] ), .B1(
        n11155), .B2(n11176), .ZN(n4545) );
  AOI22_X1 U14110 ( .A1(n7761), .A2(n11278), .B1(n11485), .B2(n11211), .ZN(
        n11227) );
  AOI22_X1 U14111 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[998] ), .B1(
        n11155), .B2(n11227), .ZN(n4544) );
  AOI22_X1 U14112 ( .A1(n7761), .A2(n11279), .B1(n11486), .B2(n11211), .ZN(
        n11214) );
  AOI22_X1 U14113 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[999] ), .B1(
        n11155), .B2(n11214), .ZN(n4543) );
  AOI22_X1 U14114 ( .A1(n7761), .A2(n11280), .B1(n11487), .B2(n11211), .ZN(
        n11177) );
  AOI22_X1 U14115 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1000] ), .B1(
        n11155), .B2(n11177), .ZN(n4542) );
  AOI22_X1 U14116 ( .A1(n7761), .A2(n11281), .B1(n11488), .B2(n11211), .ZN(
        n11204) );
  AOI22_X1 U14117 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1001] ), .B1(
        n11155), .B2(n11204), .ZN(n4541) );
  AOI22_X1 U14118 ( .A1(n7761), .A2(n11282), .B1(n11489), .B2(n11211), .ZN(
        n11228) );
  AOI22_X1 U14119 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1002] ), .B1(
        n11155), .B2(n11228), .ZN(n4540) );
  AOI22_X1 U14120 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1003] ), .B1(
        n11155), .B2(n11229), .ZN(n4539) );
  AOI22_X1 U14121 ( .A1(n7761), .A2(n11284), .B1(n11491), .B2(n11211), .ZN(
        n11178) );
  AOI22_X1 U14122 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[1004] ), 
        .B1(n11155), .B2(n11178), .ZN(n4538) );
  AOI22_X1 U14123 ( .A1(n7761), .A2(n11285), .B1(n11492), .B2(n11211), .ZN(
        n11215) );
  AOI22_X1 U14124 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[1005] ), 
        .B1(n11155), .B2(n11215), .ZN(n4537) );
  AOI22_X1 U14125 ( .A1(n7761), .A2(n11286), .B1(n11493), .B2(n11211), .ZN(
        n11216) );
  AOI22_X1 U14126 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1006] ), .B1(
        n11155), .B2(n11216), .ZN(n4536) );
  AOI22_X1 U14127 ( .A1(n7761), .A2(n11287), .B1(n11494), .B2(n11211), .ZN(
        n11179) );
  AOI22_X1 U14128 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1007] ), .B1(
        n11155), .B2(n11179), .ZN(n4535) );
  AOI22_X1 U14129 ( .A1(n7761), .A2(n11288), .B1(n11495), .B2(n11211), .ZN(
        n11205) );
  AOI22_X1 U14130 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[1008] ), 
        .B1(n11155), .B2(n11205), .ZN(n4534) );
  AOI22_X1 U14131 ( .A1(n7761), .A2(n11289), .B1(n11496), .B2(n11211), .ZN(
        n11180) );
  AOI22_X1 U14132 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1009] ), .B1(
        n11155), .B2(n11180), .ZN(n4533) );
  AOI22_X1 U14133 ( .A1(n7761), .A2(n11290), .B1(n11497), .B2(n11211), .ZN(
        n11230) );
  AOI22_X1 U14134 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1010] ), .B1(
        n11155), .B2(n11230), .ZN(n4532) );
  AOI22_X1 U14135 ( .A1(n7761), .A2(n11291), .B1(n11498), .B2(n11211), .ZN(
        n11217) );
  AOI22_X1 U14136 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1011] ), .B1(
        n11155), .B2(n11217), .ZN(n4531) );
  AOI22_X1 U14137 ( .A1(n7761), .A2(n11292), .B1(n11499), .B2(n11211), .ZN(
        n11231) );
  AOI22_X1 U14138 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1012] ), .B1(
        n11155), .B2(n11231), .ZN(n4530) );
  AOI22_X1 U14139 ( .A1(n7761), .A2(n11293), .B1(n11500), .B2(n11211), .ZN(
        n11232) );
  AOI22_X1 U14140 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[1013] ), 
        .B1(n11155), .B2(n11232), .ZN(n4529) );
  AOI22_X1 U14141 ( .A1(n7761), .A2(n11294), .B1(n11501), .B2(n11211), .ZN(
        n11218) );
  AOI22_X1 U14142 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1014] ), .B1(
        n11155), .B2(n11218), .ZN(n4528) );
  AOI22_X1 U14143 ( .A1(n7761), .A2(n11295), .B1(n11502), .B2(n11211), .ZN(
        n11181) );
  AOI22_X1 U14144 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[1015] ), 
        .B1(n11155), .B2(n11181), .ZN(n4527) );
  AOI22_X1 U14145 ( .A1(n7761), .A2(n11296), .B1(n11503), .B2(n11211), .ZN(
        n11206) );
  AOI22_X1 U14146 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1016] ), .B1(
        n11155), .B2(n11206), .ZN(n4526) );
  AOI22_X1 U14147 ( .A1(n7761), .A2(n11297), .B1(n11504), .B2(n11211), .ZN(
        n11182) );
  AOI22_X1 U14148 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[1017] ), 
        .B1(n11155), .B2(n11182), .ZN(n4525) );
  AOI22_X1 U14149 ( .A1(n7761), .A2(n11298), .B1(n11505), .B2(n11211), .ZN(
        n11207) );
  AOI22_X1 U14150 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1018] ), .B1(
        n11155), .B2(n11207), .ZN(n4524) );
  AOI22_X1 U14151 ( .A1(n7761), .A2(n11299), .B1(n11506), .B2(n11211), .ZN(
        n11183) );
  AOI22_X1 U14152 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1019] ), .B1(
        n11155), .B2(n11183), .ZN(n4523) );
  AOI22_X1 U14153 ( .A1(n7761), .A2(n11300), .B1(n11507), .B2(n11211), .ZN(
        n11184) );
  AOI22_X1 U14154 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1020] ), .B1(
        n11155), .B2(n11184), .ZN(n4522) );
  AOI22_X1 U14155 ( .A1(n7761), .A2(n11301), .B1(n11508), .B2(n11211), .ZN(
        n11185) );
  AOI22_X1 U14156 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1021] ), .B1(
        n11155), .B2(n11185), .ZN(n4521) );
  AOI22_X1 U14157 ( .A1(n7761), .A2(n11302), .B1(n11509), .B2(n11211), .ZN(
        n11219) );
  AOI22_X1 U14158 ( .A1(n8387), .A2(\DataPath/RF/bus_reg_dataout[1022] ), .B1(
        n11155), .B2(n11219), .ZN(n4520) );
  AOI22_X1 U14159 ( .A1(n7761), .A2(n11304), .B1(n11512), .B2(n11211), .ZN(
        n11191) );
  AOI22_X1 U14160 ( .A1(n11156), .A2(\DataPath/RF/bus_reg_dataout[1023] ), 
        .B1(n11155), .B2(n11191), .ZN(n4517) );
  AOI22_X1 U14161 ( .A1(n11238), .A2(n8388), .B1(n8389), .B2(
        \DataPath/RF/bus_reg_dataout[960] ), .ZN(n4515) );
  AOI22_X1 U14162 ( .A1(\DataPath/RF/bus_reg_dataout[961] ), .A2(n8389), .B1(
        n11239), .B2(n11157), .ZN(n4514) );
  AOI22_X1 U14163 ( .A1(\DataPath/RF/bus_reg_dataout[962] ), .A2(n8389), .B1(
        n11240), .B2(n8388), .ZN(n4513) );
  AOI22_X1 U14164 ( .A1(\DataPath/RF/bus_reg_dataout[963] ), .A2(n8389), .B1(
        n11241), .B2(n8388), .ZN(n4512) );
  AOI22_X1 U14165 ( .A1(\DataPath/RF/bus_reg_dataout[964] ), .A2(n11158), .B1(
        n11242), .B2(n8388), .ZN(n4511) );
  AOI22_X1 U14166 ( .A1(\DataPath/RF/bus_reg_dataout[965] ), .A2(n8389), .B1(
        n11243), .B2(n8388), .ZN(n4510) );
  AOI22_X1 U14167 ( .A1(\DataPath/RF/bus_reg_dataout[966] ), .A2(n11158), .B1(
        n11244), .B2(n8388), .ZN(n4509) );
  AOI22_X1 U14168 ( .A1(\DataPath/RF/bus_reg_dataout[967] ), .A2(n8389), .B1(
        n11245), .B2(n8388), .ZN(n4508) );
  AOI22_X1 U14169 ( .A1(\DataPath/RF/bus_reg_dataout[968] ), .A2(n11158), .B1(
        n11246), .B2(n11157), .ZN(n4507) );
  AOI22_X1 U14170 ( .A1(\DataPath/RF/bus_reg_dataout[969] ), .A2(n8389), .B1(
        n11247), .B2(n11157), .ZN(n4506) );
  AOI22_X1 U14171 ( .A1(\DataPath/RF/bus_reg_dataout[970] ), .A2(n8389), .B1(
        n11248), .B2(n11157), .ZN(n4505) );
  AOI22_X1 U14172 ( .A1(\DataPath/RF/bus_reg_dataout[971] ), .A2(n8389), .B1(
        n11249), .B2(n8388), .ZN(n4504) );
  AOI22_X1 U14173 ( .A1(\DataPath/RF/bus_reg_dataout[972] ), .A2(n8389), .B1(
        n11250), .B2(n8388), .ZN(n4503) );
  AOI22_X1 U14174 ( .A1(\DataPath/RF/bus_reg_dataout[973] ), .A2(n8389), .B1(
        n11251), .B2(n8388), .ZN(n4502) );
  AOI22_X1 U14175 ( .A1(\DataPath/RF/bus_reg_dataout[974] ), .A2(n8389), .B1(
        n11252), .B2(n8388), .ZN(n4501) );
  AOI22_X1 U14176 ( .A1(\DataPath/RF/bus_reg_dataout[975] ), .A2(n11158), .B1(
        n11253), .B2(n8388), .ZN(n4500) );
  AOI22_X1 U14177 ( .A1(\DataPath/RF/bus_reg_dataout[976] ), .A2(n8389), .B1(
        n11254), .B2(n8388), .ZN(n4499) );
  AOI22_X1 U14178 ( .A1(\DataPath/RF/bus_reg_dataout[977] ), .A2(n11158), .B1(
        n11255), .B2(n11157), .ZN(n4498) );
  AOI22_X1 U14179 ( .A1(\DataPath/RF/bus_reg_dataout[978] ), .A2(n8389), .B1(
        n11256), .B2(n11157), .ZN(n4497) );
  AOI22_X1 U14180 ( .A1(\DataPath/RF/bus_reg_dataout[979] ), .A2(n11158), .B1(
        n11257), .B2(n11157), .ZN(n4496) );
  AOI22_X1 U14181 ( .A1(\DataPath/RF/bus_reg_dataout[980] ), .A2(n8389), .B1(
        n11258), .B2(n8388), .ZN(n4495) );
  AOI22_X1 U14182 ( .A1(\DataPath/RF/bus_reg_dataout[981] ), .A2(n11158), .B1(
        n11259), .B2(n8388), .ZN(n4494) );
  AOI22_X1 U14183 ( .A1(\DataPath/RF/bus_reg_dataout[982] ), .A2(n8389), .B1(
        n11260), .B2(n8388), .ZN(n4493) );
  OAI22_X1 U14184 ( .A1(n11158), .A2(n11261), .B1(
        \DataPath/RF/bus_reg_dataout[983] ), .B2(n11157), .ZN(n4492) );
  OAI22_X1 U14185 ( .A1(n8389), .A2(n11262), .B1(
        \DataPath/RF/bus_reg_dataout[984] ), .B2(n8388), .ZN(n4491) );
  AOI22_X1 U14186 ( .A1(\DataPath/RF/bus_reg_dataout[985] ), .A2(n11158), .B1(
        n11263), .B2(n8388), .ZN(n4490) );
  AOI22_X1 U14187 ( .A1(\DataPath/RF/bus_reg_dataout[986] ), .A2(n8389), .B1(
        n11264), .B2(n8388), .ZN(n4489) );
  AOI22_X1 U14188 ( .A1(\DataPath/RF/bus_reg_dataout[987] ), .A2(n8389), .B1(
        n11265), .B2(n8388), .ZN(n4488) );
  AOI22_X1 U14189 ( .A1(\DataPath/RF/bus_reg_dataout[988] ), .A2(n8389), .B1(
        n11266), .B2(n8388), .ZN(n4487) );
  AOI22_X1 U14190 ( .A1(\DataPath/RF/bus_reg_dataout[989] ), .A2(n8389), .B1(
        n11267), .B2(n8388), .ZN(n4486) );
  AOI22_X1 U14191 ( .A1(\DataPath/RF/bus_reg_dataout[990] ), .A2(n11158), .B1(
        n11268), .B2(n11157), .ZN(n4485) );
  AOI22_X1 U14192 ( .A1(\DataPath/RF/bus_reg_dataout[991] ), .A2(n8389), .B1(
        n11270), .B2(n8388), .ZN(n4482) );
  OAI22_X1 U14193 ( .A1(n11640), .A2(n11745), .B1(n11211), .B2(n11744), .ZN(
        n11159) );
  AOI22_X1 U14194 ( .A1(\DataPath/RF/bus_reg_dataout[928] ), .A2(n8390), .B1(
        n11160), .B2(n11174), .ZN(n4480) );
  AOI22_X1 U14195 ( .A1(\DataPath/RF/bus_reg_dataout[929] ), .A2(n8390), .B1(
        n11160), .B2(n11213), .ZN(n4479) );
  AOI22_X1 U14196 ( .A1(\DataPath/RF/bus_reg_dataout[930] ), .A2(n8390), .B1(
        n11160), .B2(n11203), .ZN(n4478) );
  AOI22_X1 U14197 ( .A1(\DataPath/RF/bus_reg_dataout[931] ), .A2(n11161), .B1(
        n11160), .B2(n11175), .ZN(n4477) );
  AOI22_X1 U14198 ( .A1(\DataPath/RF/bus_reg_dataout[932] ), .A2(n11161), .B1(
        n11160), .B2(n11189), .ZN(n4476) );
  AOI22_X1 U14199 ( .A1(\DataPath/RF/bus_reg_dataout[933] ), .A2(n11161), .B1(
        n11160), .B2(n11176), .ZN(n4475) );
  AOI22_X1 U14200 ( .A1(\DataPath/RF/bus_reg_dataout[934] ), .A2(n8390), .B1(
        n11160), .B2(n11227), .ZN(n4474) );
  AOI22_X1 U14201 ( .A1(\DataPath/RF/bus_reg_dataout[935] ), .A2(n11161), .B1(
        n11160), .B2(n11214), .ZN(n4473) );
  AOI22_X1 U14202 ( .A1(\DataPath/RF/bus_reg_dataout[936] ), .A2(n8390), .B1(
        n11160), .B2(n11177), .ZN(n4472) );
  AOI22_X1 U14203 ( .A1(\DataPath/RF/bus_reg_dataout[937] ), .A2(n8390), .B1(
        n11160), .B2(n11204), .ZN(n4471) );
  AOI22_X1 U14204 ( .A1(\DataPath/RF/bus_reg_dataout[938] ), .A2(n8390), .B1(
        n11160), .B2(n11228), .ZN(n4470) );
  AOI22_X1 U14205 ( .A1(\DataPath/RF/bus_reg_dataout[939] ), .A2(n8390), .B1(
        n11160), .B2(n11229), .ZN(n4469) );
  AOI22_X1 U14206 ( .A1(\DataPath/RF/bus_reg_dataout[940] ), .A2(n8390), .B1(
        n11160), .B2(n11178), .ZN(n4468) );
  AOI22_X1 U14207 ( .A1(\DataPath/RF/bus_reg_dataout[941] ), .A2(n11161), .B1(
        n11160), .B2(n11215), .ZN(n4467) );
  AOI22_X1 U14208 ( .A1(\DataPath/RF/bus_reg_dataout[942] ), .A2(n8390), .B1(
        n11160), .B2(n11216), .ZN(n4466) );
  AOI22_X1 U14209 ( .A1(\DataPath/RF/bus_reg_dataout[943] ), .A2(n8390), .B1(
        n11160), .B2(n11179), .ZN(n4465) );
  AOI22_X1 U14210 ( .A1(\DataPath/RF/bus_reg_dataout[944] ), .A2(n11161), .B1(
        n11160), .B2(n11205), .ZN(n4464) );
  AOI22_X1 U14211 ( .A1(\DataPath/RF/bus_reg_dataout[945] ), .A2(n8390), .B1(
        n11160), .B2(n11180), .ZN(n4463) );
  AOI22_X1 U14212 ( .A1(\DataPath/RF/bus_reg_dataout[946] ), .A2(n8390), .B1(
        n11160), .B2(n11230), .ZN(n4462) );
  AOI22_X1 U14213 ( .A1(\DataPath/RF/bus_reg_dataout[947] ), .A2(n8390), .B1(
        n11160), .B2(n11217), .ZN(n4461) );
  AOI22_X1 U14214 ( .A1(\DataPath/RF/bus_reg_dataout[948] ), .A2(n8390), .B1(
        n11160), .B2(n11231), .ZN(n4460) );
  AOI22_X1 U14215 ( .A1(\DataPath/RF/bus_reg_dataout[949] ), .A2(n8390), .B1(
        n11160), .B2(n11232), .ZN(n4459) );
  AOI22_X1 U14216 ( .A1(\DataPath/RF/bus_reg_dataout[950] ), .A2(n8390), .B1(
        n11160), .B2(n11218), .ZN(n4458) );
  AOI22_X1 U14217 ( .A1(\DataPath/RF/bus_reg_dataout[951] ), .A2(n11161), .B1(
        n11160), .B2(n11181), .ZN(n4457) );
  AOI22_X1 U14218 ( .A1(\DataPath/RF/bus_reg_dataout[952] ), .A2(n8390), .B1(
        n11160), .B2(n11206), .ZN(n4456) );
  AOI22_X1 U14219 ( .A1(\DataPath/RF/bus_reg_dataout[953] ), .A2(n11161), .B1(
        n11160), .B2(n11182), .ZN(n4455) );
  AOI22_X1 U14220 ( .A1(\DataPath/RF/bus_reg_dataout[954] ), .A2(n11161), .B1(
        n11160), .B2(n11207), .ZN(n4454) );
  AOI22_X1 U14221 ( .A1(\DataPath/RF/bus_reg_dataout[955] ), .A2(n8390), .B1(
        n11160), .B2(n11183), .ZN(n4453) );
  AOI22_X1 U14222 ( .A1(\DataPath/RF/bus_reg_dataout[956] ), .A2(n8390), .B1(
        n11160), .B2(n11184), .ZN(n4452) );
  AOI22_X1 U14223 ( .A1(\DataPath/RF/bus_reg_dataout[957] ), .A2(n8390), .B1(
        n11160), .B2(n11185), .ZN(n4451) );
  AOI22_X1 U14224 ( .A1(\DataPath/RF/bus_reg_dataout[958] ), .A2(n8390), .B1(
        n11160), .B2(n11219), .ZN(n4450) );
  AOI22_X1 U14225 ( .A1(\DataPath/RF/bus_reg_dataout[959] ), .A2(n11161), .B1(
        n11160), .B2(n11191), .ZN(n4447) );
  AOI22_X1 U14226 ( .A1(\DataPath/RF/bus_reg_dataout[896] ), .A2(n8391), .B1(
        n11163), .B2(n11174), .ZN(n4445) );
  AOI22_X1 U14227 ( .A1(\DataPath/RF/bus_reg_dataout[897] ), .A2(n8391), .B1(
        n11163), .B2(n11213), .ZN(n4444) );
  AOI22_X1 U14228 ( .A1(\DataPath/RF/bus_reg_dataout[898] ), .A2(n8391), .B1(
        n11163), .B2(n11203), .ZN(n4443) );
  AOI22_X1 U14229 ( .A1(\DataPath/RF/bus_reg_dataout[899] ), .A2(n11164), .B1(
        n11163), .B2(n11175), .ZN(n4442) );
  AOI22_X1 U14230 ( .A1(\DataPath/RF/bus_reg_dataout[900] ), .A2(n8391), .B1(
        n11163), .B2(n11189), .ZN(n4441) );
  AOI22_X1 U14231 ( .A1(n11243), .A2(n11162), .B1(n8391), .B2(
        \DataPath/RF/bus_reg_dataout[901] ), .ZN(n4440) );
  AOI22_X1 U14232 ( .A1(\DataPath/RF/bus_reg_dataout[902] ), .A2(n11164), .B1(
        n11163), .B2(n11227), .ZN(n4439) );
  AOI22_X1 U14233 ( .A1(n11245), .A2(n11162), .B1(n8391), .B2(
        \DataPath/RF/bus_reg_dataout[903] ), .ZN(n4438) );
  AOI22_X1 U14234 ( .A1(\DataPath/RF/bus_reg_dataout[904] ), .A2(n8391), .B1(
        n11163), .B2(n11177), .ZN(n4437) );
  AOI22_X1 U14235 ( .A1(n11247), .A2(n11162), .B1(n8391), .B2(
        \DataPath/RF/bus_reg_dataout[905] ), .ZN(n4436) );
  AOI22_X1 U14236 ( .A1(n11248), .A2(n11162), .B1(n11164), .B2(
        \DataPath/RF/bus_reg_dataout[906] ), .ZN(n4435) );
  AOI22_X1 U14237 ( .A1(n11249), .A2(n11162), .B1(n8391), .B2(
        \DataPath/RF/bus_reg_dataout[907] ), .ZN(n4434) );
  AOI22_X1 U14238 ( .A1(\DataPath/RF/bus_reg_dataout[908] ), .A2(n11164), .B1(
        n11163), .B2(n11178), .ZN(n4433) );
  AOI22_X1 U14239 ( .A1(\DataPath/RF/bus_reg_dataout[909] ), .A2(n11164), .B1(
        n11163), .B2(n11215), .ZN(n4432) );
  AOI22_X1 U14240 ( .A1(\DataPath/RF/bus_reg_dataout[910] ), .A2(n11164), .B1(
        n11163), .B2(n11216), .ZN(n4431) );
  AOI22_X1 U14241 ( .A1(n11253), .A2(n11162), .B1(n11164), .B2(
        \DataPath/RF/bus_reg_dataout[911] ), .ZN(n4430) );
  AOI22_X1 U14242 ( .A1(n11254), .A2(n11162), .B1(n8391), .B2(
        \DataPath/RF/bus_reg_dataout[912] ), .ZN(n4429) );
  AOI22_X1 U14243 ( .A1(\DataPath/RF/bus_reg_dataout[913] ), .A2(n8391), .B1(
        n11163), .B2(n11180), .ZN(n4428) );
  AOI22_X1 U14244 ( .A1(n11256), .A2(n11162), .B1(n11164), .B2(
        \DataPath/RF/bus_reg_dataout[914] ), .ZN(n4427) );
  AOI22_X1 U14245 ( .A1(\DataPath/RF/bus_reg_dataout[915] ), .A2(n8391), .B1(
        n11163), .B2(n11217), .ZN(n4426) );
  AOI22_X1 U14246 ( .A1(\DataPath/RF/bus_reg_dataout[916] ), .A2(n11164), .B1(
        n11163), .B2(n11231), .ZN(n4425) );
  AOI22_X1 U14247 ( .A1(\DataPath/RF/bus_reg_dataout[917] ), .A2(n8391), .B1(
        n11163), .B2(n11232), .ZN(n4424) );
  AOI22_X1 U14248 ( .A1(\DataPath/RF/bus_reg_dataout[918] ), .A2(n8391), .B1(
        n11163), .B2(n11218), .ZN(n4423) );
  AOI22_X1 U14249 ( .A1(n11261), .A2(n11162), .B1(n8391), .B2(
        \DataPath/RF/bus_reg_dataout[919] ), .ZN(n4422) );
  AOI22_X1 U14250 ( .A1(\DataPath/RF/bus_reg_dataout[920] ), .A2(n8391), .B1(
        n11163), .B2(n11206), .ZN(n4421) );
  AOI22_X1 U14251 ( .A1(\DataPath/RF/bus_reg_dataout[921] ), .A2(n11164), .B1(
        n11163), .B2(n11182), .ZN(n4420) );
  AOI22_X1 U14252 ( .A1(\DataPath/RF/bus_reg_dataout[922] ), .A2(n8391), .B1(
        n11163), .B2(n11207), .ZN(n4419) );
  AOI22_X1 U14253 ( .A1(\DataPath/RF/bus_reg_dataout[923] ), .A2(n8391), .B1(
        n11163), .B2(n11183), .ZN(n4418) );
  AOI22_X1 U14254 ( .A1(\DataPath/RF/bus_reg_dataout[924] ), .A2(n8391), .B1(
        n11163), .B2(n11184), .ZN(n4417) );
  AOI22_X1 U14255 ( .A1(\DataPath/RF/bus_reg_dataout[925] ), .A2(n8391), .B1(
        n11163), .B2(n11185), .ZN(n4416) );
  AOI22_X1 U14256 ( .A1(\DataPath/RF/bus_reg_dataout[926] ), .A2(n8391), .B1(
        n11163), .B2(n11219), .ZN(n4415) );
  AOI22_X1 U14257 ( .A1(\DataPath/RF/bus_reg_dataout[927] ), .A2(n8391), .B1(
        n11163), .B2(n11191), .ZN(n4412) );
  AOI22_X1 U14258 ( .A1(\DataPath/RF/bus_reg_dataout[864] ), .A2(n8392), .B1(
        n11166), .B2(n11174), .ZN(n4410) );
  AOI22_X1 U14259 ( .A1(\DataPath/RF/bus_reg_dataout[865] ), .A2(n8392), .B1(
        n11166), .B2(n11213), .ZN(n4409) );
  AOI22_X1 U14260 ( .A1(\DataPath/RF/bus_reg_dataout[866] ), .A2(n8392), .B1(
        n11166), .B2(n11203), .ZN(n4408) );
  AOI22_X1 U14261 ( .A1(\DataPath/RF/bus_reg_dataout[867] ), .A2(n11167), .B1(
        n11166), .B2(n11175), .ZN(n4407) );
  AOI22_X1 U14262 ( .A1(\DataPath/RF/bus_reg_dataout[868] ), .A2(n8392), .B1(
        n11166), .B2(n11189), .ZN(n4406) );
  AOI22_X1 U14263 ( .A1(n11243), .A2(n11165), .B1(n11167), .B2(
        \DataPath/RF/bus_reg_dataout[869] ), .ZN(n4405) );
  AOI22_X1 U14264 ( .A1(\DataPath/RF/bus_reg_dataout[870] ), .A2(n11167), .B1(
        n11166), .B2(n11227), .ZN(n4404) );
  AOI22_X1 U14265 ( .A1(\DataPath/RF/bus_reg_dataout[871] ), .A2(n8392), .B1(
        n11166), .B2(n11214), .ZN(n4403) );
  AOI22_X1 U14266 ( .A1(\DataPath/RF/bus_reg_dataout[872] ), .A2(n11167), .B1(
        n11166), .B2(n11177), .ZN(n4402) );
  AOI22_X1 U14267 ( .A1(\DataPath/RF/bus_reg_dataout[873] ), .A2(n8392), .B1(
        n11166), .B2(n11204), .ZN(n4401) );
  AOI22_X1 U14268 ( .A1(\DataPath/RF/bus_reg_dataout[874] ), .A2(n8392), .B1(
        n11166), .B2(n11228), .ZN(n4400) );
  AOI22_X1 U14269 ( .A1(\DataPath/RF/bus_reg_dataout[875] ), .A2(n8392), .B1(
        n11166), .B2(n11229), .ZN(n4399) );
  AOI22_X1 U14270 ( .A1(\DataPath/RF/bus_reg_dataout[876] ), .A2(n8392), .B1(
        n11166), .B2(n11178), .ZN(n4398) );
  AOI22_X1 U14271 ( .A1(\DataPath/RF/bus_reg_dataout[877] ), .A2(n11167), .B1(
        n11166), .B2(n11215), .ZN(n4397) );
  AOI22_X1 U14272 ( .A1(\DataPath/RF/bus_reg_dataout[878] ), .A2(n8392), .B1(
        n11166), .B2(n11216), .ZN(n4396) );
  AOI22_X1 U14273 ( .A1(n11253), .A2(n11165), .B1(n8392), .B2(
        \DataPath/RF/bus_reg_dataout[879] ), .ZN(n4395) );
  AOI22_X1 U14274 ( .A1(\DataPath/RF/bus_reg_dataout[880] ), .A2(n11167), .B1(
        n11166), .B2(n11205), .ZN(n4394) );
  AOI22_X1 U14275 ( .A1(n11255), .A2(n11165), .B1(n11167), .B2(
        \DataPath/RF/bus_reg_dataout[881] ), .ZN(n4393) );
  AOI22_X1 U14276 ( .A1(\DataPath/RF/bus_reg_dataout[882] ), .A2(n8392), .B1(
        n11166), .B2(n11230), .ZN(n4392) );
  AOI22_X1 U14277 ( .A1(\DataPath/RF/bus_reg_dataout[883] ), .A2(n8392), .B1(
        n11166), .B2(n11217), .ZN(n4391) );
  AOI22_X1 U14278 ( .A1(\DataPath/RF/bus_reg_dataout[884] ), .A2(n8392), .B1(
        n11166), .B2(n11231), .ZN(n4390) );
  AOI22_X1 U14279 ( .A1(\DataPath/RF/bus_reg_dataout[885] ), .A2(n8392), .B1(
        n11166), .B2(n11232), .ZN(n4389) );
  AOI22_X1 U14280 ( .A1(n11260), .A2(n11165), .B1(n8392), .B2(
        \DataPath/RF/bus_reg_dataout[886] ), .ZN(n4388) );
  AOI22_X1 U14281 ( .A1(\DataPath/RF/bus_reg_dataout[887] ), .A2(n8392), .B1(
        n11166), .B2(n11181), .ZN(n4387) );
  AOI22_X1 U14282 ( .A1(\DataPath/RF/bus_reg_dataout[888] ), .A2(n8392), .B1(
        n11166), .B2(n11206), .ZN(n4386) );
  AOI22_X1 U14283 ( .A1(\DataPath/RF/bus_reg_dataout[889] ), .A2(n11167), .B1(
        n11166), .B2(n11182), .ZN(n4385) );
  AOI22_X1 U14284 ( .A1(n11264), .A2(n11165), .B1(n11167), .B2(
        \DataPath/RF/bus_reg_dataout[890] ), .ZN(n4384) );
  AOI22_X1 U14285 ( .A1(\DataPath/RF/bus_reg_dataout[891] ), .A2(n8392), .B1(
        n11166), .B2(n11183), .ZN(n4383) );
  AOI22_X1 U14286 ( .A1(n11266), .A2(n11165), .B1(n8392), .B2(
        \DataPath/RF/bus_reg_dataout[892] ), .ZN(n4382) );
  AOI22_X1 U14287 ( .A1(\DataPath/RF/bus_reg_dataout[893] ), .A2(n11167), .B1(
        n11166), .B2(n11185), .ZN(n4381) );
  AOI22_X1 U14288 ( .A1(\DataPath/RF/bus_reg_dataout[894] ), .A2(n8392), .B1(
        n11166), .B2(n11219), .ZN(n4380) );
  AOI22_X1 U14289 ( .A1(\DataPath/RF/bus_reg_dataout[895] ), .A2(n8392), .B1(
        n11166), .B2(n11191), .ZN(n4377) );
  AOI22_X1 U14290 ( .A1(\DataPath/RF/bus_reg_dataout[832] ), .A2(n8393), .B1(
        n11169), .B2(n11174), .ZN(n4375) );
  AOI22_X1 U14291 ( .A1(\DataPath/RF/bus_reg_dataout[833] ), .A2(n8393), .B1(
        n11169), .B2(n11213), .ZN(n4374) );
  AOI22_X1 U14292 ( .A1(\DataPath/RF/bus_reg_dataout[834] ), .A2(n8393), .B1(
        n11169), .B2(n11203), .ZN(n4373) );
  AOI22_X1 U14293 ( .A1(\DataPath/RF/bus_reg_dataout[835] ), .A2(n11170), .B1(
        n11169), .B2(n11175), .ZN(n4372) );
  AOI22_X1 U14294 ( .A1(\DataPath/RF/bus_reg_dataout[836] ), .A2(n8393), .B1(
        n11169), .B2(n11189), .ZN(n4371) );
  AOI22_X1 U14295 ( .A1(\DataPath/RF/bus_reg_dataout[837] ), .A2(n11170), .B1(
        n11169), .B2(n11176), .ZN(n4370) );
  AOI22_X1 U14296 ( .A1(\DataPath/RF/bus_reg_dataout[838] ), .A2(n8393), .B1(
        n11169), .B2(n11227), .ZN(n4369) );
  AOI22_X1 U14297 ( .A1(\DataPath/RF/bus_reg_dataout[839] ), .A2(n11170), .B1(
        n11169), .B2(n11214), .ZN(n4368) );
  AOI22_X1 U14298 ( .A1(n11246), .A2(n11168), .B1(n8393), .B2(
        \DataPath/RF/bus_reg_dataout[840] ), .ZN(n4367) );
  AOI22_X1 U14299 ( .A1(\DataPath/RF/bus_reg_dataout[841] ), .A2(n8393), .B1(
        n11169), .B2(n11204), .ZN(n4366) );
  AOI22_X1 U14300 ( .A1(\DataPath/RF/bus_reg_dataout[842] ), .A2(n8393), .B1(
        n11169), .B2(n11228), .ZN(n4365) );
  AOI22_X1 U14301 ( .A1(\DataPath/RF/bus_reg_dataout[843] ), .A2(n8393), .B1(
        n11169), .B2(n11229), .ZN(n4364) );
  AOI22_X1 U14302 ( .A1(\DataPath/RF/bus_reg_dataout[844] ), .A2(n8393), .B1(
        n11169), .B2(n11178), .ZN(n4363) );
  AOI22_X1 U14303 ( .A1(\DataPath/RF/bus_reg_dataout[845] ), .A2(n8393), .B1(
        n11169), .B2(n11215), .ZN(n4362) );
  AOI22_X1 U14304 ( .A1(\DataPath/RF/bus_reg_dataout[846] ), .A2(n11170), .B1(
        n11169), .B2(n11216), .ZN(n4361) );
  AOI22_X1 U14305 ( .A1(\DataPath/RF/bus_reg_dataout[847] ), .A2(n11170), .B1(
        n11169), .B2(n11179), .ZN(n4360) );
  AOI22_X1 U14306 ( .A1(\DataPath/RF/bus_reg_dataout[848] ), .A2(n8393), .B1(
        n11169), .B2(n11205), .ZN(n4359) );
  AOI22_X1 U14307 ( .A1(\DataPath/RF/bus_reg_dataout[849] ), .A2(n11170), .B1(
        n11169), .B2(n11180), .ZN(n4358) );
  AOI22_X1 U14308 ( .A1(\DataPath/RF/bus_reg_dataout[850] ), .A2(n8393), .B1(
        n11169), .B2(n11230), .ZN(n4357) );
  AOI22_X1 U14309 ( .A1(\DataPath/RF/bus_reg_dataout[851] ), .A2(n11170), .B1(
        n11169), .B2(n11217), .ZN(n4356) );
  AOI22_X1 U14310 ( .A1(\DataPath/RF/bus_reg_dataout[852] ), .A2(n8393), .B1(
        n11169), .B2(n11231), .ZN(n4355) );
  AOI22_X1 U14311 ( .A1(\DataPath/RF/bus_reg_dataout[853] ), .A2(n8393), .B1(
        n11169), .B2(n11232), .ZN(n4354) );
  AOI22_X1 U14312 ( .A1(\DataPath/RF/bus_reg_dataout[854] ), .A2(n11170), .B1(
        n11169), .B2(n11218), .ZN(n4353) );
  AOI22_X1 U14313 ( .A1(\DataPath/RF/bus_reg_dataout[855] ), .A2(n8393), .B1(
        n11169), .B2(n11181), .ZN(n4352) );
  AOI22_X1 U14314 ( .A1(\DataPath/RF/bus_reg_dataout[856] ), .A2(n8393), .B1(
        n11169), .B2(n11206), .ZN(n4351) );
  AOI22_X1 U14315 ( .A1(\DataPath/RF/bus_reg_dataout[857] ), .A2(n8393), .B1(
        n11169), .B2(n11182), .ZN(n4350) );
  AOI22_X1 U14316 ( .A1(\DataPath/RF/bus_reg_dataout[858] ), .A2(n8393), .B1(
        n11169), .B2(n11207), .ZN(n4349) );
  AOI22_X1 U14317 ( .A1(n11265), .A2(n11168), .B1(n11170), .B2(
        \DataPath/RF/bus_reg_dataout[859] ), .ZN(n4348) );
  AOI22_X1 U14318 ( .A1(n11266), .A2(n11168), .B1(n8393), .B2(
        \DataPath/RF/bus_reg_dataout[860] ), .ZN(n4347) );
  AOI22_X1 U14319 ( .A1(\DataPath/RF/bus_reg_dataout[861] ), .A2(n8393), .B1(
        n11169), .B2(n11185), .ZN(n4346) );
  AOI22_X1 U14320 ( .A1(\DataPath/RF/bus_reg_dataout[862] ), .A2(n11170), .B1(
        n11169), .B2(n11219), .ZN(n4345) );
  AOI22_X1 U14321 ( .A1(\DataPath/RF/bus_reg_dataout[863] ), .A2(n8393), .B1(
        n11169), .B2(n11191), .ZN(n4342) );
  AOI22_X1 U14322 ( .A1(n11238), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[800] ), .ZN(n4340) );
  AOI22_X1 U14323 ( .A1(n11239), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[801] ), .ZN(n4339) );
  AOI22_X1 U14324 ( .A1(n11240), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[802] ), .ZN(n4338) );
  AOI22_X1 U14325 ( .A1(n11241), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[803] ), .ZN(n4337) );
  AOI22_X1 U14326 ( .A1(n11242), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[804] ), .ZN(n4336) );
  AOI22_X1 U14327 ( .A1(n11243), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[805] ), .ZN(n4335) );
  AOI22_X1 U14328 ( .A1(n11244), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[806] ), .ZN(n4334) );
  AOI22_X1 U14329 ( .A1(n11245), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[807] ), .ZN(n4333) );
  AOI22_X1 U14330 ( .A1(n11246), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[808] ), .ZN(n4332) );
  AOI22_X1 U14331 ( .A1(n11247), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[809] ), .ZN(n4331) );
  AOI22_X1 U14332 ( .A1(n11248), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[810] ), .ZN(n4330) );
  AOI22_X1 U14333 ( .A1(n11249), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[811] ), .ZN(n4329) );
  AOI22_X1 U14334 ( .A1(n11250), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[812] ), .ZN(n4328) );
  AOI22_X1 U14335 ( .A1(n11251), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[813] ), .ZN(n4327) );
  AOI22_X1 U14336 ( .A1(n11252), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[814] ), .ZN(n4326) );
  AOI22_X1 U14337 ( .A1(n11253), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[815] ), .ZN(n4325) );
  AOI22_X1 U14338 ( .A1(n11254), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[816] ), .ZN(n4324) );
  AOI22_X1 U14339 ( .A1(n11255), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[817] ), .ZN(n4323) );
  AOI22_X1 U14340 ( .A1(n11256), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[818] ), .ZN(n4322) );
  AOI22_X1 U14341 ( .A1(n11257), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[819] ), .ZN(n4321) );
  AOI22_X1 U14342 ( .A1(n11258), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[820] ), .ZN(n4320) );
  AOI22_X1 U14343 ( .A1(n11259), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[821] ), .ZN(n4319) );
  AOI22_X1 U14344 ( .A1(n11260), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[822] ), .ZN(n4318) );
  AOI22_X1 U14345 ( .A1(n11261), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[823] ), .ZN(n4317) );
  AOI22_X1 U14346 ( .A1(n11262), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[824] ), .ZN(n4316) );
  AOI22_X1 U14347 ( .A1(n11263), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[825] ), .ZN(n4315) );
  AOI22_X1 U14348 ( .A1(n11264), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[826] ), .ZN(n4314) );
  AOI22_X1 U14349 ( .A1(n11265), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[827] ), .ZN(n4313) );
  AOI22_X1 U14350 ( .A1(n11266), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[828] ), .ZN(n4312) );
  AOI22_X1 U14351 ( .A1(n11267), .A2(n11172), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[829] ), .ZN(n4311) );
  AOI22_X1 U14352 ( .A1(n11268), .A2(n8394), .B1(n8395), .B2(
        \DataPath/RF/bus_reg_dataout[830] ), .ZN(n4310) );
  AOI22_X1 U14353 ( .A1(n11270), .A2(n8394), .B1(n11171), .B2(
        \DataPath/RF/bus_reg_dataout[831] ), .ZN(n4307) );
  OAI22_X1 U14354 ( .A1(n11640), .A2(n11333), .B1(n11211), .B2(n11332), .ZN(
        n11173) );
  AOI22_X1 U14355 ( .A1(\DataPath/RF/bus_reg_dataout[768] ), .A2(n8396), .B1(
        n11186), .B2(n11174), .ZN(n4305) );
  AOI22_X1 U14356 ( .A1(\DataPath/RF/bus_reg_dataout[769] ), .A2(n8396), .B1(
        n11186), .B2(n11213), .ZN(n4304) );
  AOI22_X1 U14357 ( .A1(\DataPath/RF/bus_reg_dataout[770] ), .A2(n8396), .B1(
        n11186), .B2(n11203), .ZN(n4303) );
  AOI22_X1 U14358 ( .A1(\DataPath/RF/bus_reg_dataout[771] ), .A2(n11187), .B1(
        n11186), .B2(n11175), .ZN(n4302) );
  AOI22_X1 U14359 ( .A1(\DataPath/RF/bus_reg_dataout[772] ), .A2(n11187), .B1(
        n11186), .B2(n11189), .ZN(n4301) );
  AOI22_X1 U14360 ( .A1(\DataPath/RF/bus_reg_dataout[773] ), .A2(n11187), .B1(
        n11186), .B2(n11176), .ZN(n4300) );
  AOI22_X1 U14361 ( .A1(\DataPath/RF/bus_reg_dataout[774] ), .A2(n8396), .B1(
        n11186), .B2(n11227), .ZN(n4299) );
  AOI22_X1 U14362 ( .A1(\DataPath/RF/bus_reg_dataout[775] ), .A2(n11187), .B1(
        n11186), .B2(n11214), .ZN(n4298) );
  AOI22_X1 U14363 ( .A1(\DataPath/RF/bus_reg_dataout[776] ), .A2(n8396), .B1(
        n11186), .B2(n11177), .ZN(n4297) );
  AOI22_X1 U14364 ( .A1(\DataPath/RF/bus_reg_dataout[777] ), .A2(n8396), .B1(
        n11186), .B2(n11204), .ZN(n4296) );
  AOI22_X1 U14365 ( .A1(\DataPath/RF/bus_reg_dataout[778] ), .A2(n8396), .B1(
        n11186), .B2(n11228), .ZN(n4295) );
  AOI22_X1 U14366 ( .A1(\DataPath/RF/bus_reg_dataout[779] ), .A2(n8396), .B1(
        n11186), .B2(n11229), .ZN(n4294) );
  AOI22_X1 U14367 ( .A1(\DataPath/RF/bus_reg_dataout[780] ), .A2(n8396), .B1(
        n11186), .B2(n11178), .ZN(n4293) );
  AOI22_X1 U14368 ( .A1(\DataPath/RF/bus_reg_dataout[781] ), .A2(n11187), .B1(
        n11186), .B2(n11215), .ZN(n4292) );
  AOI22_X1 U14369 ( .A1(\DataPath/RF/bus_reg_dataout[782] ), .A2(n8396), .B1(
        n11186), .B2(n11216), .ZN(n4291) );
  AOI22_X1 U14370 ( .A1(\DataPath/RF/bus_reg_dataout[783] ), .A2(n8396), .B1(
        n11186), .B2(n11179), .ZN(n4290) );
  AOI22_X1 U14371 ( .A1(\DataPath/RF/bus_reg_dataout[784] ), .A2(n11187), .B1(
        n11186), .B2(n11205), .ZN(n4289) );
  AOI22_X1 U14372 ( .A1(\DataPath/RF/bus_reg_dataout[785] ), .A2(n8396), .B1(
        n11186), .B2(n11180), .ZN(n4288) );
  AOI22_X1 U14373 ( .A1(\DataPath/RF/bus_reg_dataout[786] ), .A2(n8396), .B1(
        n11186), .B2(n11230), .ZN(n4287) );
  AOI22_X1 U14374 ( .A1(\DataPath/RF/bus_reg_dataout[787] ), .A2(n8396), .B1(
        n11186), .B2(n11217), .ZN(n4286) );
  AOI22_X1 U14375 ( .A1(\DataPath/RF/bus_reg_dataout[788] ), .A2(n8396), .B1(
        n11186), .B2(n11231), .ZN(n4285) );
  AOI22_X1 U14376 ( .A1(\DataPath/RF/bus_reg_dataout[789] ), .A2(n8396), .B1(
        n11186), .B2(n11232), .ZN(n4284) );
  AOI22_X1 U14377 ( .A1(\DataPath/RF/bus_reg_dataout[790] ), .A2(n8396), .B1(
        n11186), .B2(n11218), .ZN(n4283) );
  AOI22_X1 U14378 ( .A1(\DataPath/RF/bus_reg_dataout[791] ), .A2(n11187), .B1(
        n11186), .B2(n11181), .ZN(n4282) );
  AOI22_X1 U14379 ( .A1(\DataPath/RF/bus_reg_dataout[792] ), .A2(n8396), .B1(
        n11186), .B2(n11206), .ZN(n4281) );
  AOI22_X1 U14380 ( .A1(\DataPath/RF/bus_reg_dataout[793] ), .A2(n11187), .B1(
        n11186), .B2(n11182), .ZN(n4280) );
  AOI22_X1 U14381 ( .A1(\DataPath/RF/bus_reg_dataout[794] ), .A2(n11187), .B1(
        n11186), .B2(n11207), .ZN(n4279) );
  AOI22_X1 U14382 ( .A1(\DataPath/RF/bus_reg_dataout[795] ), .A2(n8396), .B1(
        n11186), .B2(n11183), .ZN(n4278) );
  AOI22_X1 U14383 ( .A1(\DataPath/RF/bus_reg_dataout[796] ), .A2(n8396), .B1(
        n11186), .B2(n11184), .ZN(n4277) );
  AOI22_X1 U14384 ( .A1(\DataPath/RF/bus_reg_dataout[797] ), .A2(n8396), .B1(
        n11186), .B2(n11185), .ZN(n4276) );
  AOI22_X1 U14385 ( .A1(\DataPath/RF/bus_reg_dataout[798] ), .A2(n8396), .B1(
        n11186), .B2(n11219), .ZN(n4275) );
  AOI22_X1 U14386 ( .A1(\DataPath/RF/bus_reg_dataout[799] ), .A2(n11187), .B1(
        n11186), .B2(n11191), .ZN(n4272) );
  OAI22_X1 U14387 ( .A1(n11415), .A2(n11339), .B1(n11640), .B2(n11338), .ZN(
        n11188) );
  AOI22_X1 U14388 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[736] ), .B1(
        n11238), .B2(n11190), .ZN(n4270) );
  AOI22_X1 U14389 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[737] ), .B1(
        n11239), .B2(n11190), .ZN(n4269) );
  AOI22_X1 U14390 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[738] ), .B1(
        n11240), .B2(n11190), .ZN(n4268) );
  AOI22_X1 U14391 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[739] ), .B1(
        n11241), .B2(n11190), .ZN(n4267) );
  NOR2_X1 U14392 ( .A1(RST), .A2(n11193), .ZN(n11192) );
  AOI22_X1 U14393 ( .A1(\DataPath/RF/bus_reg_dataout[740] ), .A2(n11193), .B1(
        n11192), .B2(n11189), .ZN(n4266) );
  AOI22_X1 U14394 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[741] ), .B1(
        n11243), .B2(n11190), .ZN(n4265) );
  AOI22_X1 U14395 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[742] ), .B1(
        n11244), .B2(n11190), .ZN(n4264) );
  AOI22_X1 U14396 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[743] ), .B1(
        n11245), .B2(n11190), .ZN(n4263) );
  AOI22_X1 U14397 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[744] ), .B1(
        n11246), .B2(n11190), .ZN(n4262) );
  AOI22_X1 U14398 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[745] ), .B1(
        n11247), .B2(n11190), .ZN(n4261) );
  AOI22_X1 U14399 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[746] ), .B1(
        n11248), .B2(n11190), .ZN(n4260) );
  AOI22_X1 U14400 ( .A1(\DataPath/RF/bus_reg_dataout[747] ), .A2(n11193), .B1(
        n11192), .B2(n11229), .ZN(n4259) );
  AOI22_X1 U14401 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[748] ), .B1(
        n11250), .B2(n11190), .ZN(n4258) );
  AOI22_X1 U14402 ( .A1(\DataPath/RF/bus_reg_dataout[749] ), .A2(n11193), .B1(
        n11192), .B2(n11215), .ZN(n4257) );
  AOI22_X1 U14403 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[750] ), .B1(
        n11252), .B2(n11190), .ZN(n4256) );
  AOI22_X1 U14404 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[751] ), .B1(
        n11253), .B2(n11190), .ZN(n4255) );
  AOI22_X1 U14405 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[752] ), .B1(
        n11254), .B2(n11190), .ZN(n4254) );
  AOI22_X1 U14406 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[753] ), .B1(
        n11255), .B2(n11190), .ZN(n4253) );
  AOI22_X1 U14407 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[754] ), .B1(
        n11256), .B2(n11190), .ZN(n4252) );
  AOI22_X1 U14408 ( .A1(\DataPath/RF/bus_reg_dataout[755] ), .A2(n11193), .B1(
        n11192), .B2(n11217), .ZN(n4251) );
  AOI22_X1 U14409 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[756] ), .B1(
        n11258), .B2(n11190), .ZN(n4250) );
  AOI22_X1 U14410 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[757] ), .B1(
        n11259), .B2(n11190), .ZN(n4249) );
  AOI22_X1 U14411 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[758] ), .B1(
        n11260), .B2(n11190), .ZN(n4248) );
  AOI22_X1 U14412 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[759] ), .B1(
        n11261), .B2(n11190), .ZN(n4247) );
  AOI22_X1 U14413 ( .A1(\DataPath/RF/bus_reg_dataout[760] ), .A2(n11193), .B1(
        n11192), .B2(n11206), .ZN(n4246) );
  AOI22_X1 U14414 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[761] ), .B1(
        n11263), .B2(n11190), .ZN(n4245) );
  AOI22_X1 U14415 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[762] ), .B1(
        n11264), .B2(n11190), .ZN(n4244) );
  AOI22_X1 U14416 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[763] ), .B1(
        n11265), .B2(n11190), .ZN(n4243) );
  AOI22_X1 U14417 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[764] ), .B1(
        n11266), .B2(n11190), .ZN(n4242) );
  AOI22_X1 U14418 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[765] ), .B1(
        n11267), .B2(n11190), .ZN(n4241) );
  AOI22_X1 U14419 ( .A1(n11193), .A2(\DataPath/RF/bus_reg_dataout[766] ), .B1(
        n11268), .B2(n11190), .ZN(n4240) );
  AOI22_X1 U14420 ( .A1(\DataPath/RF/bus_reg_dataout[767] ), .A2(n11193), .B1(
        n11192), .B2(n11191), .ZN(n4237) );
  OAI22_X1 U14421 ( .A1(n11238), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[704] ), .B2(n11195), .ZN(n4235) );
  AOI22_X1 U14422 ( .A1(n11239), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[705] ), .ZN(n4234) );
  AOI22_X1 U14423 ( .A1(n11240), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[706] ), .ZN(n4233) );
  OAI22_X1 U14424 ( .A1(n11241), .A2(n11196), .B1(
        \DataPath/RF/bus_reg_dataout[707] ), .B2(n11195), .ZN(n4232) );
  AOI22_X1 U14425 ( .A1(n11242), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[708] ), .ZN(n4231) );
  AOI22_X1 U14426 ( .A1(n11243), .A2(n11195), .B1(n11196), .B2(
        \DataPath/RF/bus_reg_dataout[709] ), .ZN(n4230) );
  OAI22_X1 U14427 ( .A1(n11244), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[710] ), .B2(n11195), .ZN(n4229) );
  AOI22_X1 U14428 ( .A1(n11245), .A2(n11195), .B1(n11196), .B2(
        \DataPath/RF/bus_reg_dataout[711] ), .ZN(n4228) );
  OAI22_X1 U14429 ( .A1(n11246), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[712] ), .B2(n11195), .ZN(n4227) );
  AOI22_X1 U14430 ( .A1(n11247), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[713] ), .ZN(n4226) );
  OAI22_X1 U14431 ( .A1(n11248), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[714] ), .B2(n11195), .ZN(n4225) );
  OAI22_X1 U14432 ( .A1(n11249), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[715] ), .B2(n11195), .ZN(n4224) );
  OAI22_X1 U14433 ( .A1(n11250), .A2(n11196), .B1(
        \DataPath/RF/bus_reg_dataout[716] ), .B2(n11195), .ZN(n4223) );
  AOI22_X1 U14434 ( .A1(n11251), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[717] ), .ZN(n4222) );
  OAI22_X1 U14435 ( .A1(n11252), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[718] ), .B2(n11195), .ZN(n4221) );
  AOI22_X1 U14436 ( .A1(n11253), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[719] ), .ZN(n4220) );
  OAI22_X1 U14437 ( .A1(n11254), .A2(n11196), .B1(
        \DataPath/RF/bus_reg_dataout[720] ), .B2(n11195), .ZN(n4219) );
  OAI22_X1 U14438 ( .A1(n11255), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[721] ), .B2(n11195), .ZN(n4218) );
  OAI22_X1 U14439 ( .A1(n11256), .A2(n11196), .B1(
        \DataPath/RF/bus_reg_dataout[722] ), .B2(n11195), .ZN(n4217) );
  AOI22_X1 U14440 ( .A1(n11257), .A2(n11195), .B1(n11196), .B2(
        \DataPath/RF/bus_reg_dataout[723] ), .ZN(n4216) );
  AOI22_X1 U14441 ( .A1(n11258), .A2(n11195), .B1(n11196), .B2(
        \DataPath/RF/bus_reg_dataout[724] ), .ZN(n4215) );
  OAI22_X1 U14442 ( .A1(n11259), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[725] ), .B2(n11195), .ZN(n4214) );
  OAI22_X1 U14443 ( .A1(n11260), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[726] ), .B2(n11195), .ZN(n4213) );
  OAI22_X1 U14444 ( .A1(n11261), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[727] ), .B2(n11195), .ZN(n4212) );
  OAI22_X1 U14445 ( .A1(n11262), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[728] ), .B2(n11195), .ZN(n4211) );
  AOI22_X1 U14446 ( .A1(n11263), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[729] ), .ZN(n4210) );
  OAI22_X1 U14447 ( .A1(n11264), .A2(n11196), .B1(
        \DataPath/RF/bus_reg_dataout[730] ), .B2(n11195), .ZN(n4209) );
  AOI22_X1 U14448 ( .A1(n11265), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[731] ), .ZN(n4208) );
  AOI22_X1 U14449 ( .A1(n11266), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[732] ), .ZN(n4207) );
  AOI22_X1 U14450 ( .A1(n11267), .A2(n11195), .B1(n11196), .B2(
        \DataPath/RF/bus_reg_dataout[733] ), .ZN(n4206) );
  AOI22_X1 U14451 ( .A1(n11268), .A2(n11195), .B1(n8397), .B2(
        \DataPath/RF/bus_reg_dataout[734] ), .ZN(n4205) );
  OAI22_X1 U14452 ( .A1(n11270), .A2(n8397), .B1(
        \DataPath/RF/bus_reg_dataout[735] ), .B2(n11195), .ZN(n4202) );
  OAI22_X1 U14453 ( .A1(n11415), .A2(n11353), .B1(n11211), .B2(n11352), .ZN(
        n11197) );
  AOI22_X1 U14454 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[672] ), .B1(
        n11238), .B2(n11199), .ZN(n4200) );
  AOI22_X1 U14455 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[673] ), .B1(
        n11239), .B2(n11199), .ZN(n4199) );
  AOI22_X1 U14456 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[674] ), .B1(
        n11240), .B2(n11199), .ZN(n4198) );
  AOI22_X1 U14457 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[675] ), .B1(
        n11241), .B2(n11199), .ZN(n4197) );
  AOI22_X1 U14458 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[676] ), .B1(
        n11242), .B2(n11199), .ZN(n4196) );
  AOI22_X1 U14459 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[677] ), .B1(
        n11243), .B2(n11199), .ZN(n4195) );
  AOI22_X1 U14460 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[678] ), .B1(
        n11244), .B2(n11199), .ZN(n4194) );
  AOI22_X1 U14461 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[679] ), .B1(
        n11245), .B2(n11199), .ZN(n4193) );
  AOI22_X1 U14462 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[680] ), .B1(
        n11246), .B2(n11199), .ZN(n4192) );
  AOI22_X1 U14463 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[681] ), .B1(
        n11247), .B2(n11199), .ZN(n4191) );
  AOI22_X1 U14464 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[682] ), .B1(
        n11248), .B2(n11199), .ZN(n4190) );
  NOR2_X1 U14465 ( .A1(RST), .A2(n11200), .ZN(n11198) );
  AOI22_X1 U14466 ( .A1(\DataPath/RF/bus_reg_dataout[683] ), .A2(n11200), .B1(
        n11198), .B2(n11229), .ZN(n4189) );
  AOI22_X1 U14467 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[684] ), .B1(
        n11250), .B2(n11199), .ZN(n4188) );
  AOI22_X1 U14468 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[685] ), .B1(
        n11251), .B2(n11199), .ZN(n4187) );
  AOI22_X1 U14469 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[686] ), .B1(
        n11252), .B2(n11199), .ZN(n4186) );
  AOI22_X1 U14470 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[687] ), .B1(
        n11253), .B2(n11199), .ZN(n4185) );
  AOI22_X1 U14471 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[688] ), .B1(
        n11254), .B2(n11199), .ZN(n4184) );
  AOI22_X1 U14472 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[689] ), .B1(
        n11255), .B2(n11199), .ZN(n4183) );
  AOI22_X1 U14473 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[690] ), .B1(
        n11256), .B2(n11199), .ZN(n4182) );
  AOI22_X1 U14474 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[691] ), .B1(
        n11257), .B2(n11199), .ZN(n4181) );
  AOI22_X1 U14475 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[692] ), .B1(
        n11258), .B2(n11199), .ZN(n4180) );
  AOI22_X1 U14476 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[693] ), .B1(
        n11259), .B2(n11199), .ZN(n4179) );
  AOI22_X1 U14477 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[694] ), .B1(
        n11260), .B2(n11199), .ZN(n4178) );
  AOI22_X1 U14478 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[695] ), .B1(
        n11261), .B2(n11199), .ZN(n4177) );
  AOI22_X1 U14479 ( .A1(\DataPath/RF/bus_reg_dataout[696] ), .A2(n11200), .B1(
        n11198), .B2(n11206), .ZN(n4176) );
  AOI22_X1 U14480 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[697] ), .B1(
        n11263), .B2(n11199), .ZN(n4175) );
  AOI22_X1 U14481 ( .A1(\DataPath/RF/bus_reg_dataout[698] ), .A2(n11200), .B1(
        n11198), .B2(n11207), .ZN(n4174) );
  AOI22_X1 U14482 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[699] ), .B1(
        n11265), .B2(n11199), .ZN(n4173) );
  AOI22_X1 U14483 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[700] ), .B1(
        n11266), .B2(n11199), .ZN(n4172) );
  AOI22_X1 U14484 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[701] ), .B1(
        n11267), .B2(n11199), .ZN(n4171) );
  AOI22_X1 U14485 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[702] ), .B1(
        n11268), .B2(n11199), .ZN(n4170) );
  AOI22_X1 U14486 ( .A1(n11200), .A2(\DataPath/RF/bus_reg_dataout[703] ), .B1(
        n11270), .B2(n11199), .ZN(n4167) );
  OAI22_X1 U14487 ( .A1(n11415), .A2(n11360), .B1(n11211), .B2(n11361), .ZN(
        n11201) );
  AOI22_X1 U14488 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[640] ), .B1(
        n11238), .B2(n11209), .ZN(n4165) );
  AOI22_X1 U14489 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[641] ), .B1(
        n11239), .B2(n11209), .ZN(n4164) );
  AOI22_X1 U14490 ( .A1(\DataPath/RF/bus_reg_dataout[642] ), .A2(n11210), .B1(
        n11208), .B2(n11203), .ZN(n4163) );
  AOI22_X1 U14491 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[643] ), .B1(
        n11241), .B2(n11209), .ZN(n4162) );
  AOI22_X1 U14492 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[644] ), .B1(
        n11242), .B2(n11209), .ZN(n4161) );
  AOI22_X1 U14493 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[645] ), .B1(
        n11243), .B2(n11209), .ZN(n4160) );
  AOI22_X1 U14494 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[646] ), .B1(
        n11244), .B2(n11209), .ZN(n4159) );
  AOI22_X1 U14495 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[647] ), .B1(
        n11245), .B2(n11209), .ZN(n4158) );
  AOI22_X1 U14496 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[648] ), .B1(
        n11246), .B2(n11209), .ZN(n4157) );
  AOI22_X1 U14497 ( .A1(\DataPath/RF/bus_reg_dataout[649] ), .A2(n11210), .B1(
        n11208), .B2(n11204), .ZN(n4156) );
  AOI22_X1 U14498 ( .A1(\DataPath/RF/bus_reg_dataout[650] ), .A2(n11210), .B1(
        n11208), .B2(n11228), .ZN(n4155) );
  AOI22_X1 U14499 ( .A1(\DataPath/RF/bus_reg_dataout[651] ), .A2(n11210), .B1(
        n11208), .B2(n11229), .ZN(n4154) );
  AOI22_X1 U14500 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[652] ), .B1(
        n11250), .B2(n11209), .ZN(n4153) );
  AOI22_X1 U14501 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[653] ), .B1(
        n11251), .B2(n11209), .ZN(n4152) );
  AOI22_X1 U14502 ( .A1(\DataPath/RF/bus_reg_dataout[654] ), .A2(n11210), .B1(
        n11208), .B2(n11216), .ZN(n4151) );
  AOI22_X1 U14503 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[655] ), .B1(
        n11253), .B2(n11209), .ZN(n4150) );
  AOI22_X1 U14504 ( .A1(\DataPath/RF/bus_reg_dataout[656] ), .A2(n11210), .B1(
        n11208), .B2(n11205), .ZN(n4149) );
  AOI22_X1 U14505 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[657] ), .B1(
        n11255), .B2(n11209), .ZN(n4148) );
  AOI22_X1 U14506 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[658] ), .B1(
        n11256), .B2(n11209), .ZN(n4147) );
  AOI22_X1 U14507 ( .A1(\DataPath/RF/bus_reg_dataout[659] ), .A2(n11210), .B1(
        n11208), .B2(n11217), .ZN(n4146) );
  AOI22_X1 U14508 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[660] ), .B1(
        n11258), .B2(n11209), .ZN(n4145) );
  AOI22_X1 U14509 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[661] ), .B1(
        n11259), .B2(n11209), .ZN(n4144) );
  AOI22_X1 U14510 ( .A1(\DataPath/RF/bus_reg_dataout[662] ), .A2(n11210), .B1(
        n11208), .B2(n11218), .ZN(n4143) );
  AOI22_X1 U14511 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[663] ), .B1(
        n11261), .B2(n11209), .ZN(n4142) );
  AOI22_X1 U14512 ( .A1(\DataPath/RF/bus_reg_dataout[664] ), .A2(n11210), .B1(
        n11208), .B2(n11206), .ZN(n4141) );
  AOI22_X1 U14513 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[665] ), .B1(
        n11263), .B2(n11209), .ZN(n4140) );
  AOI22_X1 U14514 ( .A1(\DataPath/RF/bus_reg_dataout[666] ), .A2(n11210), .B1(
        n11208), .B2(n11207), .ZN(n4139) );
  AOI22_X1 U14515 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[667] ), .B1(
        n11265), .B2(n11209), .ZN(n4138) );
  AOI22_X1 U14516 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[668] ), .B1(
        n11266), .B2(n11209), .ZN(n4137) );
  AOI22_X1 U14517 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[669] ), .B1(
        n11267), .B2(n11209), .ZN(n4136) );
  AOI22_X1 U14518 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[670] ), .B1(
        n11268), .B2(n11209), .ZN(n4135) );
  AOI22_X1 U14519 ( .A1(n11210), .A2(\DataPath/RF/bus_reg_dataout[671] ), .B1(
        n11270), .B2(n11209), .ZN(n4132) );
  OAI22_X1 U14520 ( .A1(n11415), .A2(n11367), .B1(n11211), .B2(n11366), .ZN(
        n11212) );
  AOI22_X1 U14521 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[608] ), .B1(
        n11238), .B2(n11221), .ZN(n4130) );
  AOI22_X1 U14522 ( .A1(\DataPath/RF/bus_reg_dataout[609] ), .A2(n11222), .B1(
        n11220), .B2(n11213), .ZN(n4129) );
  AOI22_X1 U14523 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[610] ), .B1(
        n11240), .B2(n11221), .ZN(n4128) );
  AOI22_X1 U14524 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[611] ), .B1(
        n11241), .B2(n11221), .ZN(n4127) );
  AOI22_X1 U14525 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[612] ), .B1(
        n11242), .B2(n11221), .ZN(n4126) );
  AOI22_X1 U14526 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[613] ), .B1(
        n11243), .B2(n11221), .ZN(n4125) );
  AOI22_X1 U14527 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[614] ), .B1(
        n11244), .B2(n11221), .ZN(n4124) );
  AOI22_X1 U14528 ( .A1(\DataPath/RF/bus_reg_dataout[615] ), .A2(n11222), .B1(
        n11220), .B2(n11214), .ZN(n4123) );
  AOI22_X1 U14529 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[616] ), .B1(
        n11246), .B2(n11221), .ZN(n4122) );
  AOI22_X1 U14530 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[617] ), .B1(
        n11247), .B2(n11221), .ZN(n4121) );
  AOI22_X1 U14531 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[618] ), .B1(
        n11248), .B2(n11221), .ZN(n4120) );
  AOI22_X1 U14532 ( .A1(\DataPath/RF/bus_reg_dataout[619] ), .A2(n11222), .B1(
        n11220), .B2(n11229), .ZN(n4119) );
  AOI22_X1 U14533 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[620] ), .B1(
        n11250), .B2(n11221), .ZN(n4118) );
  AOI22_X1 U14534 ( .A1(\DataPath/RF/bus_reg_dataout[621] ), .A2(n11222), .B1(
        n11220), .B2(n11215), .ZN(n4117) );
  AOI22_X1 U14535 ( .A1(\DataPath/RF/bus_reg_dataout[622] ), .A2(n11222), .B1(
        n11220), .B2(n11216), .ZN(n4116) );
  AOI22_X1 U14536 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[623] ), .B1(
        n11253), .B2(n11221), .ZN(n4115) );
  AOI22_X1 U14537 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[624] ), .B1(
        n11254), .B2(n11221), .ZN(n4114) );
  AOI22_X1 U14538 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[625] ), .B1(
        n11255), .B2(n11221), .ZN(n4113) );
  AOI22_X1 U14539 ( .A1(\DataPath/RF/bus_reg_dataout[626] ), .A2(n11222), .B1(
        n11220), .B2(n11230), .ZN(n4112) );
  AOI22_X1 U14540 ( .A1(\DataPath/RF/bus_reg_dataout[627] ), .A2(n11222), .B1(
        n11220), .B2(n11217), .ZN(n4111) );
  AOI22_X1 U14541 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[628] ), .B1(
        n11258), .B2(n11221), .ZN(n4110) );
  AOI22_X1 U14542 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[629] ), .B1(
        n11259), .B2(n11221), .ZN(n4109) );
  AOI22_X1 U14543 ( .A1(\DataPath/RF/bus_reg_dataout[630] ), .A2(n11222), .B1(
        n11220), .B2(n11218), .ZN(n4108) );
  AOI22_X1 U14544 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[631] ), .B1(
        n11261), .B2(n11221), .ZN(n4107) );
  AOI22_X1 U14545 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[632] ), .B1(
        n11262), .B2(n11221), .ZN(n4106) );
  AOI22_X1 U14546 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[633] ), .B1(
        n11263), .B2(n11221), .ZN(n4105) );
  AOI22_X1 U14547 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[634] ), .B1(
        n11264), .B2(n11221), .ZN(n4104) );
  AOI22_X1 U14548 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[635] ), .B1(
        n11265), .B2(n11221), .ZN(n4103) );
  AOI22_X1 U14549 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[636] ), .B1(
        n11266), .B2(n11221), .ZN(n4102) );
  AOI22_X1 U14550 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[637] ), .B1(
        n11267), .B2(n11221), .ZN(n4101) );
  AOI22_X1 U14551 ( .A1(\DataPath/RF/bus_reg_dataout[638] ), .A2(n11222), .B1(
        n11220), .B2(n11219), .ZN(n4100) );
  AOI22_X1 U14552 ( .A1(n11222), .A2(\DataPath/RF/bus_reg_dataout[639] ), .B1(
        n11270), .B2(n11221), .ZN(n4097) );
  OAI22_X1 U14553 ( .A1(n11415), .A2(n11375), .B1(n11640), .B2(n11374), .ZN(
        n11223) );
  AOI22_X1 U14554 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[576] ), .B1(
        n11238), .B2(n11224), .ZN(n4095) );
  AOI22_X1 U14555 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[577] ), .B1(
        n11239), .B2(n11224), .ZN(n4094) );
  AOI22_X1 U14556 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[578] ), .B1(
        n11240), .B2(n11224), .ZN(n4093) );
  AOI22_X1 U14557 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[579] ), .B1(
        n11241), .B2(n11224), .ZN(n4092) );
  AOI22_X1 U14558 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[580] ), .B1(
        n11242), .B2(n11224), .ZN(n4091) );
  AOI22_X1 U14559 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[581] ), .B1(
        n11243), .B2(n11224), .ZN(n4090) );
  AOI22_X1 U14560 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[582] ), .B1(
        n11244), .B2(n11224), .ZN(n4089) );
  AOI22_X1 U14561 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[583] ), .B1(
        n11245), .B2(n11224), .ZN(n4088) );
  AOI22_X1 U14562 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[584] ), .B1(
        n11246), .B2(n11224), .ZN(n4087) );
  AOI22_X1 U14563 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[585] ), .B1(
        n11247), .B2(n11224), .ZN(n4086) );
  AOI22_X1 U14564 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[586] ), .B1(
        n11248), .B2(n11224), .ZN(n4085) );
  AOI22_X1 U14565 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[587] ), .B1(
        n11249), .B2(n11224), .ZN(n4084) );
  AOI22_X1 U14566 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[588] ), .B1(
        n11250), .B2(n11224), .ZN(n4083) );
  AOI22_X1 U14567 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[589] ), .B1(
        n11251), .B2(n11224), .ZN(n4082) );
  AOI22_X1 U14568 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[590] ), .B1(
        n11252), .B2(n11224), .ZN(n4081) );
  AOI22_X1 U14569 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[591] ), .B1(
        n11253), .B2(n11224), .ZN(n4080) );
  AOI22_X1 U14570 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[592] ), .B1(
        n11254), .B2(n11224), .ZN(n4079) );
  AOI22_X1 U14571 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[593] ), .B1(
        n11255), .B2(n11224), .ZN(n4078) );
  AOI22_X1 U14572 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[594] ), .B1(
        n11256), .B2(n11224), .ZN(n4077) );
  AOI22_X1 U14573 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[595] ), .B1(
        n11257), .B2(n11224), .ZN(n4076) );
  AOI22_X1 U14574 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[596] ), .B1(
        n11258), .B2(n11224), .ZN(n4075) );
  AOI22_X1 U14575 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[597] ), .B1(
        n11259), .B2(n11224), .ZN(n4074) );
  AOI22_X1 U14576 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[598] ), .B1(
        n11260), .B2(n11224), .ZN(n4073) );
  AOI22_X1 U14577 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[599] ), .B1(
        n11261), .B2(n11224), .ZN(n4072) );
  AOI22_X1 U14578 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[600] ), .B1(
        n11262), .B2(n11224), .ZN(n4071) );
  AOI22_X1 U14579 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[601] ), .B1(
        n11263), .B2(n11224), .ZN(n4070) );
  AOI22_X1 U14580 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[602] ), .B1(
        n11264), .B2(n11224), .ZN(n4069) );
  AOI22_X1 U14581 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[603] ), .B1(
        n11265), .B2(n11224), .ZN(n4068) );
  AOI22_X1 U14582 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[604] ), .B1(
        n11266), .B2(n11224), .ZN(n4067) );
  AOI22_X1 U14583 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[605] ), .B1(
        n11267), .B2(n11224), .ZN(n4066) );
  AOI22_X1 U14584 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[606] ), .B1(
        n11268), .B2(n11224), .ZN(n4065) );
  AOI22_X1 U14585 ( .A1(n11225), .A2(\DataPath/RF/bus_reg_dataout[607] ), .B1(
        n11270), .B2(n11224), .ZN(n4062) );
  OAI22_X1 U14586 ( .A1(n11415), .A2(n11407), .B1(n11640), .B2(n11406), .ZN(
        n11226) );
  AOI22_X1 U14587 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[544] ), .B1(
        n11238), .B2(n11234), .ZN(n4060) );
  AOI22_X1 U14588 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[545] ), .B1(
        n11239), .B2(n11234), .ZN(n4059) );
  AOI22_X1 U14589 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[546] ), .B1(
        n11240), .B2(n11234), .ZN(n4058) );
  AOI22_X1 U14590 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[547] ), .B1(
        n11241), .B2(n11234), .ZN(n4057) );
  AOI22_X1 U14591 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[548] ), .B1(
        n11242), .B2(n11234), .ZN(n4056) );
  AOI22_X1 U14592 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[549] ), .B1(
        n11243), .B2(n11234), .ZN(n4055) );
  NOR2_X1 U14593 ( .A1(RST), .A2(n11235), .ZN(n11233) );
  AOI22_X1 U14594 ( .A1(\DataPath/RF/bus_reg_dataout[550] ), .A2(n11235), .B1(
        n11233), .B2(n11227), .ZN(n4054) );
  AOI22_X1 U14595 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[551] ), .B1(
        n11245), .B2(n11234), .ZN(n4053) );
  AOI22_X1 U14596 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[552] ), .B1(
        n11246), .B2(n11234), .ZN(n4052) );
  AOI22_X1 U14597 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[553] ), .B1(
        n11247), .B2(n11234), .ZN(n4051) );
  AOI22_X1 U14598 ( .A1(\DataPath/RF/bus_reg_dataout[554] ), .A2(n11235), .B1(
        n11233), .B2(n11228), .ZN(n4050) );
  AOI22_X1 U14599 ( .A1(\DataPath/RF/bus_reg_dataout[555] ), .A2(n11235), .B1(
        n11233), .B2(n11229), .ZN(n4049) );
  AOI22_X1 U14600 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[556] ), .B1(
        n11250), .B2(n11234), .ZN(n4048) );
  AOI22_X1 U14601 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[557] ), .B1(
        n11251), .B2(n11234), .ZN(n4047) );
  AOI22_X1 U14602 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[558] ), .B1(
        n11252), .B2(n11234), .ZN(n4046) );
  AOI22_X1 U14603 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[559] ), .B1(
        n11253), .B2(n11234), .ZN(n4045) );
  AOI22_X1 U14604 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[560] ), .B1(
        n11254), .B2(n11234), .ZN(n4044) );
  AOI22_X1 U14605 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[561] ), .B1(
        n11255), .B2(n11234), .ZN(n4043) );
  AOI22_X1 U14606 ( .A1(\DataPath/RF/bus_reg_dataout[562] ), .A2(n11235), .B1(
        n11233), .B2(n11230), .ZN(n4042) );
  AOI22_X1 U14607 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[563] ), .B1(
        n11257), .B2(n11234), .ZN(n4041) );
  AOI22_X1 U14608 ( .A1(\DataPath/RF/bus_reg_dataout[564] ), .A2(n11235), .B1(
        n11233), .B2(n11231), .ZN(n4040) );
  AOI22_X1 U14609 ( .A1(\DataPath/RF/bus_reg_dataout[565] ), .A2(n11235), .B1(
        n11233), .B2(n11232), .ZN(n4039) );
  AOI22_X1 U14610 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[566] ), .B1(
        n11260), .B2(n11234), .ZN(n4038) );
  AOI22_X1 U14611 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[567] ), .B1(
        n11261), .B2(n11234), .ZN(n4037) );
  AOI22_X1 U14612 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[568] ), .B1(
        n11262), .B2(n11234), .ZN(n4036) );
  AOI22_X1 U14613 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[569] ), .B1(
        n11263), .B2(n11234), .ZN(n4035) );
  AOI22_X1 U14614 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[570] ), .B1(
        n11264), .B2(n11234), .ZN(n4034) );
  AOI22_X1 U14615 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[571] ), .B1(
        n11265), .B2(n11234), .ZN(n4033) );
  AOI22_X1 U14616 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[572] ), .B1(
        n11266), .B2(n11234), .ZN(n4032) );
  AOI22_X1 U14617 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[573] ), .B1(
        n11267), .B2(n11234), .ZN(n4031) );
  AOI22_X1 U14618 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[574] ), .B1(
        n11268), .B2(n11234), .ZN(n4030) );
  AOI22_X1 U14619 ( .A1(n11235), .A2(\DataPath/RF/bus_reg_dataout[575] ), .B1(
        n11270), .B2(n11234), .ZN(n4027) );
  OAI22_X1 U14620 ( .A1(n11415), .A2(n11416), .B1(n11640), .B2(n11414), .ZN(
        n11236) );
  AOI22_X1 U14621 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[512] ), .B1(
        n11238), .B2(n11269), .ZN(n4023) );
  AOI22_X1 U14622 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[513] ), .B1(
        n11239), .B2(n11269), .ZN(n4021) );
  AOI22_X1 U14623 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[514] ), .B1(
        n11240), .B2(n11269), .ZN(n4019) );
  AOI22_X1 U14624 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[515] ), .B1(
        n11241), .B2(n11269), .ZN(n4017) );
  AOI22_X1 U14625 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[516] ), .B1(
        n11242), .B2(n11269), .ZN(n4015) );
  AOI22_X1 U14626 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[517] ), .B1(
        n11243), .B2(n11269), .ZN(n4013) );
  AOI22_X1 U14627 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[518] ), .B1(
        n11244), .B2(n11269), .ZN(n4011) );
  AOI22_X1 U14628 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[519] ), .B1(
        n11245), .B2(n11269), .ZN(n4009) );
  AOI22_X1 U14629 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[520] ), .B1(
        n11246), .B2(n11269), .ZN(n4007) );
  AOI22_X1 U14630 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[521] ), .B1(
        n11247), .B2(n11269), .ZN(n4005) );
  AOI22_X1 U14631 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[522] ), .B1(
        n11248), .B2(n11269), .ZN(n4003) );
  AOI22_X1 U14632 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[523] ), .B1(
        n11249), .B2(n11269), .ZN(n4001) );
  AOI22_X1 U14633 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[524] ), .B1(
        n11250), .B2(n11269), .ZN(n3999) );
  AOI22_X1 U14634 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[525] ), .B1(
        n11251), .B2(n11269), .ZN(n3997) );
  AOI22_X1 U14635 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[526] ), .B1(
        n11252), .B2(n11269), .ZN(n3995) );
  AOI22_X1 U14636 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[527] ), .B1(
        n11253), .B2(n11269), .ZN(n3993) );
  AOI22_X1 U14637 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[528] ), .B1(
        n11254), .B2(n11269), .ZN(n3991) );
  AOI22_X1 U14638 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[529] ), .B1(
        n11255), .B2(n11269), .ZN(n3989) );
  AOI22_X1 U14639 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[530] ), .B1(
        n11256), .B2(n11269), .ZN(n3987) );
  AOI22_X1 U14640 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[531] ), .B1(
        n11257), .B2(n11269), .ZN(n3985) );
  AOI22_X1 U14641 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[532] ), .B1(
        n11258), .B2(n11269), .ZN(n3983) );
  AOI22_X1 U14642 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[533] ), .B1(
        n11259), .B2(n11269), .ZN(n3981) );
  AOI22_X1 U14643 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[534] ), .B1(
        n11260), .B2(n11269), .ZN(n3979) );
  AOI22_X1 U14644 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[535] ), .B1(
        n11261), .B2(n11269), .ZN(n3977) );
  AOI22_X1 U14645 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[536] ), .B1(
        n11262), .B2(n11269), .ZN(n3975) );
  AOI22_X1 U14646 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[537] ), .B1(
        n11263), .B2(n11269), .ZN(n3973) );
  AOI22_X1 U14647 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[538] ), .B1(
        n11264), .B2(n11269), .ZN(n3971) );
  AOI22_X1 U14648 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[539] ), .B1(
        n11265), .B2(n11269), .ZN(n3969) );
  AOI22_X1 U14649 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[540] ), .B1(
        n11266), .B2(n11269), .ZN(n3967) );
  AOI22_X1 U14650 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[541] ), .B1(
        n11267), .B2(n11269), .ZN(n3965) );
  AOI22_X1 U14651 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[542] ), .B1(
        n11268), .B2(n11269), .ZN(n3963) );
  AOI22_X1 U14652 ( .A1(n11271), .A2(\DataPath/RF/bus_reg_dataout[543] ), .B1(
        n11270), .B2(n11269), .ZN(n3959) );
  AOI22_X1 U14653 ( .A1(n11419), .A2(n11272), .B1(n11479), .B2(n7756), .ZN(
        n11378) );
  AOI22_X1 U14654 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[480] ), .B1(
        n11303), .B2(n11378), .ZN(n3955) );
  AOI22_X1 U14655 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[481] ), .B1(
        n11303), .B2(n11421), .ZN(n3953) );
  AOI22_X1 U14656 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[482] ), .B1(
        n11303), .B2(n11422), .ZN(n3951) );
  AOI22_X1 U14657 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[483] ), .B1(
        n11303), .B2(n11423), .ZN(n3949) );
  AOI22_X1 U14658 ( .A1(\DataPath/RF/bus_reg_dataout[484] ), .A2(n11306), .B1(
        n11424), .B2(n11305), .ZN(n3947) );
  AOI22_X1 U14659 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[485] ), .B1(
        n11303), .B2(n11380), .ZN(n3945) );
  AOI22_X1 U14660 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[486] ), .B1(
        n11303), .B2(n11426), .ZN(n3943) );
  AOI22_X1 U14661 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[487] ), .B1(
        n11303), .B2(n11381), .ZN(n3941) );
  AOI22_X1 U14662 ( .A1(n11419), .A2(n11280), .B1(n11487), .B2(n7756), .ZN(
        n11382) );
  AOI22_X1 U14663 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[488] ), .B1(
        n11303), .B2(n11382), .ZN(n3939) );
  AOI22_X1 U14664 ( .A1(n11419), .A2(n11281), .B1(n11488), .B2(n7756), .ZN(
        n11383) );
  AOI22_X1 U14665 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[489] ), .B1(
        n11303), .B2(n11383), .ZN(n3937) );
  AOI22_X1 U14666 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[490] ), .B1(
        n11303), .B2(n11384), .ZN(n3935) );
  AOI22_X1 U14667 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[491] ), .B1(
        n11303), .B2(n11385), .ZN(n3933) );
  AOI22_X1 U14668 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[492] ), .B1(
        n11303), .B2(n11386), .ZN(n3931) );
  AOI22_X1 U14669 ( .A1(n11419), .A2(n11285), .B1(n11492), .B2(n7756), .ZN(
        n11387) );
  AOI22_X1 U14670 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[493] ), .B1(
        n11303), .B2(n11387), .ZN(n3929) );
  AOI22_X1 U14671 ( .A1(n11419), .A2(n11286), .B1(n11493), .B2(n7756), .ZN(
        n11388) );
  AOI22_X1 U14672 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[494] ), .B1(
        n11303), .B2(n11388), .ZN(n3927) );
  AOI22_X1 U14673 ( .A1(n8410), .A2(n11287), .B1(n11494), .B2(n7756), .ZN(
        n11389) );
  AOI22_X1 U14674 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[495] ), .B1(
        n11303), .B2(n11389), .ZN(n3925) );
  AOI22_X1 U14675 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[496] ), .B1(
        n11303), .B2(n11390), .ZN(n3923) );
  OAI22_X1 U14676 ( .A1(n7756), .A2(n11289), .B1(n11496), .B2(n8410), .ZN(
        n11410) );
  AOI22_X1 U14677 ( .A1(\DataPath/RF/bus_reg_dataout[497] ), .A2(n8398), .B1(
        n11438), .B2(n11305), .ZN(n3921) );
  AOI22_X1 U14678 ( .A1(n8410), .A2(n11290), .B1(n11497), .B2(n7756), .ZN(
        n11391) );
  AOI22_X1 U14679 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[498] ), .B1(
        n11303), .B2(n11391), .ZN(n3919) );
  AOI22_X1 U14680 ( .A1(n8410), .A2(n11291), .B1(n11498), .B2(n7756), .ZN(
        n11392) );
  AOI22_X1 U14681 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[499] ), .B1(
        n11303), .B2(n11392), .ZN(n3917) );
  AOI22_X1 U14682 ( .A1(\DataPath/RF/bus_reg_dataout[500] ), .A2(n8398), .B1(
        n11305), .B2(n11441), .ZN(n3915) );
  OAI22_X1 U14683 ( .A1(n7756), .A2(n11293), .B1(n11500), .B2(n8410), .ZN(
        n11394) );
  AOI22_X1 U14684 ( .A1(\DataPath/RF/bus_reg_dataout[501] ), .A2(n8398), .B1(
        n11442), .B2(n11305), .ZN(n3913) );
  AOI22_X1 U14685 ( .A1(n11419), .A2(n11294), .B1(n11501), .B2(n7756), .ZN(
        n11395) );
  AOI22_X1 U14686 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[502] ), .B1(
        n11303), .B2(n11395), .ZN(n3911) );
  AOI22_X1 U14687 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[503] ), .B1(
        n11303), .B2(n11396), .ZN(n3909) );
  AOI22_X1 U14688 ( .A1(n8410), .A2(n11296), .B1(n11503), .B2(n7756), .ZN(
        n11397) );
  AOI22_X1 U14689 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[504] ), .B1(
        n11303), .B2(n11397), .ZN(n3907) );
  AOI22_X1 U14690 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[505] ), .B1(
        n11303), .B2(n11398), .ZN(n3905) );
  AOI22_X1 U14691 ( .A1(n11419), .A2(n11298), .B1(n11505), .B2(n7756), .ZN(
        n11399) );
  AOI22_X1 U14692 ( .A1(n11306), .A2(\DataPath/RF/bus_reg_dataout[506] ), .B1(
        n11303), .B2(n11399), .ZN(n3903) );
  OAI22_X1 U14693 ( .A1(n7756), .A2(n11299), .B1(n11506), .B2(n8410), .ZN(
        n11400) );
  AOI22_X1 U14694 ( .A1(\DataPath/RF/bus_reg_dataout[507] ), .A2(n8398), .B1(
        n11448), .B2(n11305), .ZN(n3901) );
  OAI22_X1 U14695 ( .A1(n7756), .A2(n11300), .B1(n11507), .B2(n8410), .ZN(
        n11401) );
  AOI22_X1 U14696 ( .A1(\DataPath/RF/bus_reg_dataout[508] ), .A2(n11306), .B1(
        n11449), .B2(n11305), .ZN(n3899) );
  AOI22_X1 U14697 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[509] ), .B1(
        n11303), .B2(n11402), .ZN(n3897) );
  AOI22_X1 U14698 ( .A1(n8398), .A2(\DataPath/RF/bus_reg_dataout[510] ), .B1(
        n11303), .B2(n11411), .ZN(n3895) );
  OAI22_X1 U14699 ( .A1(n7756), .A2(n11304), .B1(n11512), .B2(n8410), .ZN(
        n11403) );
  AOI22_X1 U14700 ( .A1(\DataPath/RF/bus_reg_dataout[511] ), .A2(n8398), .B1(
        n11597), .B2(n11305), .ZN(n3891) );
  AOI22_X1 U14701 ( .A1(\DataPath/RF/bus_reg_dataout[448] ), .A2(n8399), .B1(
        n11308), .B2(n11378), .ZN(n3889) );
  AOI22_X1 U14702 ( .A1(\DataPath/RF/bus_reg_dataout[449] ), .A2(n11309), .B1(
        n11308), .B2(n11421), .ZN(n3888) );
  AOI22_X1 U14703 ( .A1(\DataPath/RF/bus_reg_dataout[450] ), .A2(n8399), .B1(
        n11308), .B2(n11422), .ZN(n3887) );
  AOI22_X1 U14704 ( .A1(\DataPath/RF/bus_reg_dataout[451] ), .A2(n8399), .B1(
        n11308), .B2(n11423), .ZN(n3886) );
  AOI22_X1 U14705 ( .A1(\DataPath/RF/bus_reg_dataout[452] ), .A2(n11309), .B1(
        n11308), .B2(n11379), .ZN(n3885) );
  AOI22_X1 U14706 ( .A1(\DataPath/RF/bus_reg_dataout[453] ), .A2(n11309), .B1(
        n11308), .B2(n11380), .ZN(n3884) );
  AOI22_X1 U14707 ( .A1(\DataPath/RF/bus_reg_dataout[454] ), .A2(n8399), .B1(
        n11308), .B2(n11426), .ZN(n3883) );
  AOI22_X1 U14708 ( .A1(\DataPath/RF/bus_reg_dataout[455] ), .A2(n8399), .B1(
        n11308), .B2(n11381), .ZN(n3882) );
  AOI22_X1 U14709 ( .A1(\DataPath/RF/bus_reg_dataout[456] ), .A2(n11309), .B1(
        n11429), .B2(n11307), .ZN(n3881) );
  AOI22_X1 U14710 ( .A1(\DataPath/RF/bus_reg_dataout[457] ), .A2(n8399), .B1(
        n11430), .B2(n11307), .ZN(n3880) );
  AOI22_X1 U14711 ( .A1(\DataPath/RF/bus_reg_dataout[458] ), .A2(n11309), .B1(
        n11308), .B2(n11384), .ZN(n3879) );
  AOI22_X1 U14712 ( .A1(\DataPath/RF/bus_reg_dataout[459] ), .A2(n8399), .B1(
        n11308), .B2(n11385), .ZN(n3878) );
  AOI22_X1 U14713 ( .A1(\DataPath/RF/bus_reg_dataout[460] ), .A2(n8399), .B1(
        n11308), .B2(n11386), .ZN(n3877) );
  AOI22_X1 U14714 ( .A1(\DataPath/RF/bus_reg_dataout[461] ), .A2(n11309), .B1(
        n11308), .B2(n11387), .ZN(n3876) );
  AOI22_X1 U14715 ( .A1(\DataPath/RF/bus_reg_dataout[462] ), .A2(n8399), .B1(
        n11308), .B2(n11388), .ZN(n3875) );
  AOI22_X1 U14716 ( .A1(\DataPath/RF/bus_reg_dataout[463] ), .A2(n8399), .B1(
        n11308), .B2(n11389), .ZN(n3874) );
  AOI22_X1 U14717 ( .A1(\DataPath/RF/bus_reg_dataout[464] ), .A2(n8399), .B1(
        n11308), .B2(n11390), .ZN(n3873) );
  AOI22_X1 U14718 ( .A1(n11438), .A2(n11307), .B1(n8399), .B2(
        \DataPath/RF/bus_reg_dataout[465] ), .ZN(n3872) );
  AOI22_X1 U14719 ( .A1(\DataPath/RF/bus_reg_dataout[466] ), .A2(n8399), .B1(
        n11308), .B2(n11391), .ZN(n3871) );
  AOI22_X1 U14720 ( .A1(\DataPath/RF/bus_reg_dataout[467] ), .A2(n8399), .B1(
        n11308), .B2(n11392), .ZN(n3870) );
  OAI22_X1 U14721 ( .A1(n11309), .A2(n11441), .B1(
        \DataPath/RF/bus_reg_dataout[468] ), .B2(n11307), .ZN(n3869) );
  AOI22_X1 U14722 ( .A1(\DataPath/RF/bus_reg_dataout[469] ), .A2(n8399), .B1(
        n11308), .B2(n11394), .ZN(n3868) );
  AOI22_X1 U14723 ( .A1(\DataPath/RF/bus_reg_dataout[470] ), .A2(n8399), .B1(
        n11308), .B2(n11395), .ZN(n3867) );
  AOI22_X1 U14724 ( .A1(\DataPath/RF/bus_reg_dataout[471] ), .A2(n8399), .B1(
        n11308), .B2(n11396), .ZN(n3866) );
  AOI22_X1 U14725 ( .A1(\DataPath/RF/bus_reg_dataout[472] ), .A2(n11309), .B1(
        n11308), .B2(n11397), .ZN(n3865) );
  AOI22_X1 U14726 ( .A1(\DataPath/RF/bus_reg_dataout[473] ), .A2(n8399), .B1(
        n11308), .B2(n11398), .ZN(n3864) );
  AOI22_X1 U14727 ( .A1(\DataPath/RF/bus_reg_dataout[474] ), .A2(n8399), .B1(
        n11447), .B2(n11307), .ZN(n3863) );
  AOI22_X1 U14728 ( .A1(\DataPath/RF/bus_reg_dataout[475] ), .A2(n8399), .B1(
        n11308), .B2(n11400), .ZN(n3862) );
  AOI22_X1 U14729 ( .A1(\DataPath/RF/bus_reg_dataout[476] ), .A2(n11309), .B1(
        n11308), .B2(n11401), .ZN(n3861) );
  AOI22_X1 U14730 ( .A1(\DataPath/RF/bus_reg_dataout[477] ), .A2(n11309), .B1(
        n11308), .B2(n11402), .ZN(n3860) );
  AOI22_X1 U14731 ( .A1(\DataPath/RF/bus_reg_dataout[478] ), .A2(n8399), .B1(
        n11451), .B2(n11307), .ZN(n3859) );
  AOI22_X1 U14732 ( .A1(\DataPath/RF/bus_reg_dataout[479] ), .A2(n8399), .B1(
        n11308), .B2(n11403), .ZN(n3856) );
  AOI22_X1 U14733 ( .A1(\DataPath/RF/bus_reg_dataout[416] ), .A2(n8400), .B1(
        n11311), .B2(n11378), .ZN(n3854) );
  AOI22_X1 U14734 ( .A1(\DataPath/RF/bus_reg_dataout[417] ), .A2(n11312), .B1(
        n11311), .B2(n11421), .ZN(n3853) );
  AOI22_X1 U14735 ( .A1(\DataPath/RF/bus_reg_dataout[418] ), .A2(n11312), .B1(
        n11311), .B2(n11422), .ZN(n3852) );
  AOI22_X1 U14736 ( .A1(\DataPath/RF/bus_reg_dataout[419] ), .A2(n11312), .B1(
        n11311), .B2(n11423), .ZN(n3851) );
  AOI22_X1 U14737 ( .A1(\DataPath/RF/bus_reg_dataout[420] ), .A2(n8400), .B1(
        n11311), .B2(n11379), .ZN(n3850) );
  AOI22_X1 U14738 ( .A1(\DataPath/RF/bus_reg_dataout[421] ), .A2(n8400), .B1(
        n11311), .B2(n11380), .ZN(n3849) );
  AOI22_X1 U14739 ( .A1(\DataPath/RF/bus_reg_dataout[422] ), .A2(n8400), .B1(
        n11311), .B2(n11426), .ZN(n3848) );
  AOI22_X1 U14740 ( .A1(\DataPath/RF/bus_reg_dataout[423] ), .A2(n8400), .B1(
        n11311), .B2(n11381), .ZN(n3847) );
  AOI22_X1 U14741 ( .A1(n11429), .A2(n11310), .B1(n8400), .B2(
        \DataPath/RF/bus_reg_dataout[424] ), .ZN(n3846) );
  AOI22_X1 U14742 ( .A1(\DataPath/RF/bus_reg_dataout[425] ), .A2(n8400), .B1(
        n11311), .B2(n11383), .ZN(n3845) );
  AOI22_X1 U14743 ( .A1(\DataPath/RF/bus_reg_dataout[426] ), .A2(n8400), .B1(
        n11311), .B2(n11384), .ZN(n3844) );
  AOI22_X1 U14744 ( .A1(\DataPath/RF/bus_reg_dataout[427] ), .A2(n8400), .B1(
        n11311), .B2(n11385), .ZN(n3843) );
  AOI22_X1 U14745 ( .A1(\DataPath/RF/bus_reg_dataout[428] ), .A2(n8400), .B1(
        n11311), .B2(n11386), .ZN(n3842) );
  AOI22_X1 U14746 ( .A1(\DataPath/RF/bus_reg_dataout[429] ), .A2(n8400), .B1(
        n11434), .B2(n11310), .ZN(n3841) );
  AOI22_X1 U14747 ( .A1(\DataPath/RF/bus_reg_dataout[430] ), .A2(n11312), .B1(
        n11311), .B2(n11388), .ZN(n3840) );
  AOI22_X1 U14748 ( .A1(\DataPath/RF/bus_reg_dataout[431] ), .A2(n8400), .B1(
        n11436), .B2(n11310), .ZN(n3839) );
  AOI22_X1 U14749 ( .A1(\DataPath/RF/bus_reg_dataout[432] ), .A2(n11312), .B1(
        n11437), .B2(n11310), .ZN(n3838) );
  AOI22_X1 U14750 ( .A1(\DataPath/RF/bus_reg_dataout[433] ), .A2(n8400), .B1(
        n11311), .B2(n11410), .ZN(n3837) );
  AOI22_X1 U14751 ( .A1(\DataPath/RF/bus_reg_dataout[434] ), .A2(n8400), .B1(
        n11311), .B2(n11391), .ZN(n3836) );
  AOI22_X1 U14752 ( .A1(\DataPath/RF/bus_reg_dataout[435] ), .A2(n8400), .B1(
        n11311), .B2(n11392), .ZN(n3835) );
  AOI22_X1 U14753 ( .A1(\DataPath/RF/bus_reg_dataout[436] ), .A2(n8400), .B1(
        n11441), .B2(n11310), .ZN(n3834) );
  AOI22_X1 U14754 ( .A1(\DataPath/RF/bus_reg_dataout[437] ), .A2(n8400), .B1(
        n11311), .B2(n11394), .ZN(n3833) );
  AOI22_X1 U14755 ( .A1(\DataPath/RF/bus_reg_dataout[438] ), .A2(n8400), .B1(
        n11311), .B2(n11395), .ZN(n3832) );
  AOI22_X1 U14756 ( .A1(\DataPath/RF/bus_reg_dataout[439] ), .A2(n11312), .B1(
        n11311), .B2(n11396), .ZN(n3831) );
  AOI22_X1 U14757 ( .A1(\DataPath/RF/bus_reg_dataout[440] ), .A2(n11312), .B1(
        n11311), .B2(n11397), .ZN(n3830) );
  AOI22_X1 U14758 ( .A1(\DataPath/RF/bus_reg_dataout[441] ), .A2(n11312), .B1(
        n11311), .B2(n11398), .ZN(n3829) );
  AOI22_X1 U14759 ( .A1(n11447), .A2(n11310), .B1(n11312), .B2(
        \DataPath/RF/bus_reg_dataout[442] ), .ZN(n3828) );
  AOI22_X1 U14760 ( .A1(\DataPath/RF/bus_reg_dataout[443] ), .A2(n8400), .B1(
        n11311), .B2(n11400), .ZN(n3827) );
  AOI22_X1 U14761 ( .A1(n11449), .A2(n11310), .B1(n11312), .B2(
        \DataPath/RF/bus_reg_dataout[444] ), .ZN(n3826) );
  AOI22_X1 U14762 ( .A1(\DataPath/RF/bus_reg_dataout[445] ), .A2(n8400), .B1(
        n11311), .B2(n11402), .ZN(n3825) );
  AOI22_X1 U14763 ( .A1(n11451), .A2(n11310), .B1(n8400), .B2(
        \DataPath/RF/bus_reg_dataout[446] ), .ZN(n3824) );
  AOI22_X1 U14764 ( .A1(\DataPath/RF/bus_reg_dataout[447] ), .A2(n8400), .B1(
        n11311), .B2(n11403), .ZN(n3821) );
  AOI22_X1 U14765 ( .A1(\DataPath/RF/bus_reg_dataout[384] ), .A2(n8401), .B1(
        n11314), .B2(n11378), .ZN(n3819) );
  AOI22_X1 U14766 ( .A1(\DataPath/RF/bus_reg_dataout[385] ), .A2(n8401), .B1(
        n11314), .B2(n11421), .ZN(n3818) );
  AOI22_X1 U14767 ( .A1(\DataPath/RF/bus_reg_dataout[386] ), .A2(n8401), .B1(
        n11314), .B2(n11422), .ZN(n3817) );
  AOI22_X1 U14768 ( .A1(\DataPath/RF/bus_reg_dataout[387] ), .A2(n8401), .B1(
        n11314), .B2(n11423), .ZN(n3816) );
  AOI22_X1 U14769 ( .A1(\DataPath/RF/bus_reg_dataout[388] ), .A2(n8401), .B1(
        n11314), .B2(n11379), .ZN(n3815) );
  AOI22_X1 U14770 ( .A1(\DataPath/RF/bus_reg_dataout[389] ), .A2(n8401), .B1(
        n11314), .B2(n11380), .ZN(n3814) );
  AOI22_X1 U14771 ( .A1(\DataPath/RF/bus_reg_dataout[390] ), .A2(n8401), .B1(
        n11314), .B2(n11426), .ZN(n3813) );
  AOI22_X1 U14772 ( .A1(\DataPath/RF/bus_reg_dataout[391] ), .A2(n8401), .B1(
        n11314), .B2(n11381), .ZN(n3812) );
  AOI22_X1 U14773 ( .A1(n11429), .A2(n11316), .B1(n11315), .B2(
        \DataPath/RF/bus_reg_dataout[392] ), .ZN(n3811) );
  AOI22_X1 U14774 ( .A1(\DataPath/RF/bus_reg_dataout[393] ), .A2(n8401), .B1(
        n11314), .B2(n11383), .ZN(n3810) );
  AOI22_X1 U14775 ( .A1(\DataPath/RF/bus_reg_dataout[394] ), .A2(n8401), .B1(
        n11314), .B2(n11384), .ZN(n3809) );
  AOI22_X1 U14776 ( .A1(\DataPath/RF/bus_reg_dataout[395] ), .A2(n8401), .B1(
        n11432), .B2(n11316), .ZN(n3808) );
  AOI22_X1 U14777 ( .A1(\DataPath/RF/bus_reg_dataout[396] ), .A2(n8401), .B1(
        n11314), .B2(n11386), .ZN(n3807) );
  AOI22_X1 U14778 ( .A1(\DataPath/RF/bus_reg_dataout[397] ), .A2(n11315), .B1(
        n11314), .B2(n11387), .ZN(n3806) );
  AOI22_X1 U14779 ( .A1(\DataPath/RF/bus_reg_dataout[398] ), .A2(n11315), .B1(
        n11435), .B2(n11316), .ZN(n3805) );
  AOI22_X1 U14780 ( .A1(\DataPath/RF/bus_reg_dataout[399] ), .A2(n11315), .B1(
        n11314), .B2(n11389), .ZN(n3804) );
  AOI22_X1 U14781 ( .A1(\DataPath/RF/bus_reg_dataout[400] ), .A2(n8401), .B1(
        n11314), .B2(n11390), .ZN(n3803) );
  AOI22_X1 U14782 ( .A1(\DataPath/RF/bus_reg_dataout[401] ), .A2(n11315), .B1(
        n11314), .B2(n11410), .ZN(n3802) );
  AOI22_X1 U14783 ( .A1(\DataPath/RF/bus_reg_dataout[402] ), .A2(n8401), .B1(
        n11314), .B2(n11391), .ZN(n3801) );
  AOI22_X1 U14784 ( .A1(\DataPath/RF/bus_reg_dataout[403] ), .A2(n11315), .B1(
        n11440), .B2(n11316), .ZN(n3800) );
  INV_X1 U14785 ( .A(n11315), .ZN(n11313) );
  AOI22_X1 U14786 ( .A1(n8401), .A2(\DataPath/RF/bus_reg_dataout[404] ), .B1(
        n11441), .B2(n11313), .ZN(n3799) );
  AOI22_X1 U14787 ( .A1(n11442), .A2(n11316), .B1(n8401), .B2(
        \DataPath/RF/bus_reg_dataout[405] ), .ZN(n3798) );
  AOI22_X1 U14788 ( .A1(\DataPath/RF/bus_reg_dataout[406] ), .A2(n8401), .B1(
        n11443), .B2(n11316), .ZN(n3797) );
  AOI22_X1 U14789 ( .A1(\DataPath/RF/bus_reg_dataout[407] ), .A2(n8401), .B1(
        n11444), .B2(n11316), .ZN(n3796) );
  AOI22_X1 U14790 ( .A1(\DataPath/RF/bus_reg_dataout[408] ), .A2(n11315), .B1(
        n11314), .B2(n11397), .ZN(n3795) );
  AOI22_X1 U14791 ( .A1(\DataPath/RF/bus_reg_dataout[409] ), .A2(n8401), .B1(
        n11314), .B2(n11398), .ZN(n3794) );
  AOI22_X1 U14792 ( .A1(\DataPath/RF/bus_reg_dataout[410] ), .A2(n11315), .B1(
        n11314), .B2(n11399), .ZN(n3793) );
  AOI22_X1 U14793 ( .A1(n11448), .A2(n11316), .B1(n8401), .B2(
        \DataPath/RF/bus_reg_dataout[411] ), .ZN(n3792) );
  AOI22_X1 U14794 ( .A1(n11449), .A2(n11316), .B1(n8401), .B2(
        \DataPath/RF/bus_reg_dataout[412] ), .ZN(n3791) );
  AOI22_X1 U14795 ( .A1(\DataPath/RF/bus_reg_dataout[413] ), .A2(n8401), .B1(
        n11314), .B2(n11402), .ZN(n3790) );
  AOI22_X1 U14796 ( .A1(\DataPath/RF/bus_reg_dataout[414] ), .A2(n8401), .B1(
        n11314), .B2(n11411), .ZN(n3789) );
  AOI22_X1 U14797 ( .A1(n11597), .A2(n11316), .B1(n11315), .B2(
        \DataPath/RF/bus_reg_dataout[415] ), .ZN(n3786) );
  AOI22_X1 U14798 ( .A1(\DataPath/RF/bus_reg_dataout[352] ), .A2(n8402), .B1(
        n11420), .B2(n11318), .ZN(n3784) );
  AOI22_X1 U14799 ( .A1(\DataPath/RF/bus_reg_dataout[353] ), .A2(n8402), .B1(
        n11319), .B2(n11421), .ZN(n3783) );
  AOI22_X1 U14800 ( .A1(\DataPath/RF/bus_reg_dataout[354] ), .A2(n8402), .B1(
        n11319), .B2(n11422), .ZN(n3782) );
  AOI22_X1 U14801 ( .A1(\DataPath/RF/bus_reg_dataout[355] ), .A2(n8402), .B1(
        n11319), .B2(n11423), .ZN(n3781) );
  AOI22_X1 U14802 ( .A1(\DataPath/RF/bus_reg_dataout[356] ), .A2(n8402), .B1(
        n11319), .B2(n11379), .ZN(n3780) );
  AOI22_X1 U14803 ( .A1(\DataPath/RF/bus_reg_dataout[357] ), .A2(n8402), .B1(
        n11319), .B2(n11380), .ZN(n3779) );
  AOI22_X1 U14804 ( .A1(\DataPath/RF/bus_reg_dataout[358] ), .A2(n11320), .B1(
        n11319), .B2(n11426), .ZN(n3778) );
  AOI22_X1 U14805 ( .A1(\DataPath/RF/bus_reg_dataout[359] ), .A2(n11320), .B1(
        n11319), .B2(n11381), .ZN(n3777) );
  AOI22_X1 U14806 ( .A1(n11429), .A2(n11318), .B1(n8402), .B2(
        \DataPath/RF/bus_reg_dataout[360] ), .ZN(n3776) );
  AOI22_X1 U14807 ( .A1(\DataPath/RF/bus_reg_dataout[361] ), .A2(n8402), .B1(
        n11319), .B2(n11383), .ZN(n3775) );
  AOI22_X1 U14808 ( .A1(\DataPath/RF/bus_reg_dataout[362] ), .A2(n8402), .B1(
        n11319), .B2(n11384), .ZN(n3774) );
  AOI22_X1 U14809 ( .A1(n11432), .A2(n11318), .B1(n8402), .B2(
        \DataPath/RF/bus_reg_dataout[363] ), .ZN(n3773) );
  AOI22_X1 U14810 ( .A1(\DataPath/RF/bus_reg_dataout[364] ), .A2(n8402), .B1(
        n11319), .B2(n11386), .ZN(n3772) );
  AOI22_X1 U14811 ( .A1(\DataPath/RF/bus_reg_dataout[365] ), .A2(n8402), .B1(
        n11319), .B2(n11387), .ZN(n3771) );
  AOI22_X1 U14812 ( .A1(\DataPath/RF/bus_reg_dataout[366] ), .A2(n11320), .B1(
        n11319), .B2(n11388), .ZN(n3770) );
  AOI22_X1 U14813 ( .A1(\DataPath/RF/bus_reg_dataout[367] ), .A2(n8402), .B1(
        n11319), .B2(n11389), .ZN(n3769) );
  AOI22_X1 U14814 ( .A1(\DataPath/RF/bus_reg_dataout[368] ), .A2(n8402), .B1(
        n11319), .B2(n11390), .ZN(n3768) );
  AOI22_X1 U14815 ( .A1(n11438), .A2(n11318), .B1(n11320), .B2(
        \DataPath/RF/bus_reg_dataout[369] ), .ZN(n3767) );
  AOI22_X1 U14816 ( .A1(\DataPath/RF/bus_reg_dataout[370] ), .A2(n8402), .B1(
        n11319), .B2(n11391), .ZN(n3766) );
  AOI22_X1 U14817 ( .A1(\DataPath/RF/bus_reg_dataout[371] ), .A2(n11320), .B1(
        n11319), .B2(n11392), .ZN(n3765) );
  INV_X1 U14818 ( .A(n11320), .ZN(n11317) );
  AOI22_X1 U14819 ( .A1(n11320), .A2(\DataPath/RF/bus_reg_dataout[372] ), .B1(
        n11441), .B2(n11317), .ZN(n3764) );
  AOI22_X1 U14820 ( .A1(\DataPath/RF/bus_reg_dataout[373] ), .A2(n11320), .B1(
        n11319), .B2(n11394), .ZN(n3763) );
  AOI22_X1 U14821 ( .A1(n11443), .A2(n11318), .B1(n8402), .B2(
        \DataPath/RF/bus_reg_dataout[374] ), .ZN(n3762) );
  AOI22_X1 U14822 ( .A1(\DataPath/RF/bus_reg_dataout[375] ), .A2(n8402), .B1(
        n11319), .B2(n11396), .ZN(n3761) );
  AOI22_X1 U14823 ( .A1(\DataPath/RF/bus_reg_dataout[376] ), .A2(n8402), .B1(
        n11445), .B2(n11318), .ZN(n3760) );
  AOI22_X1 U14824 ( .A1(\DataPath/RF/bus_reg_dataout[377] ), .A2(n8402), .B1(
        n11446), .B2(n11318), .ZN(n3759) );
  AOI22_X1 U14825 ( .A1(n11447), .A2(n11318), .B1(n11320), .B2(
        \DataPath/RF/bus_reg_dataout[378] ), .ZN(n3758) );
  AOI22_X1 U14826 ( .A1(n11448), .A2(n11318), .B1(n8402), .B2(
        \DataPath/RF/bus_reg_dataout[379] ), .ZN(n3757) );
  AOI22_X1 U14827 ( .A1(n11449), .A2(n11318), .B1(n11320), .B2(
        \DataPath/RF/bus_reg_dataout[380] ), .ZN(n3756) );
  AOI22_X1 U14828 ( .A1(\DataPath/RF/bus_reg_dataout[381] ), .A2(n8402), .B1(
        n11319), .B2(n11402), .ZN(n3755) );
  AOI22_X1 U14829 ( .A1(\DataPath/RF/bus_reg_dataout[382] ), .A2(n8402), .B1(
        n11319), .B2(n11411), .ZN(n3754) );
  AOI22_X1 U14830 ( .A1(\DataPath/RF/bus_reg_dataout[383] ), .A2(n8402), .B1(
        n11319), .B2(n11403), .ZN(n3751) );
  AOI22_X1 U14831 ( .A1(n11420), .A2(n11323), .B1(n8403), .B2(
        \DataPath/RF/bus_reg_dataout[320] ), .ZN(n3747) );
  AOI22_X1 U14832 ( .A1(\DataPath/RF/bus_reg_dataout[321] ), .A2(n11325), .B1(
        n11324), .B2(n11421), .ZN(n3746) );
  AOI22_X1 U14833 ( .A1(\DataPath/RF/bus_reg_dataout[322] ), .A2(n8403), .B1(
        n11324), .B2(n11422), .ZN(n3745) );
  AOI22_X1 U14834 ( .A1(\DataPath/RF/bus_reg_dataout[323] ), .A2(n11325), .B1(
        n11324), .B2(n11423), .ZN(n3744) );
  AOI22_X1 U14835 ( .A1(\DataPath/RF/bus_reg_dataout[324] ), .A2(n8403), .B1(
        n11324), .B2(n11379), .ZN(n3743) );
  AOI22_X1 U14836 ( .A1(\DataPath/RF/bus_reg_dataout[325] ), .A2(n8403), .B1(
        n11324), .B2(n11380), .ZN(n3742) );
  AOI22_X1 U14837 ( .A1(\DataPath/RF/bus_reg_dataout[326] ), .A2(n8403), .B1(
        n11324), .B2(n11426), .ZN(n3741) );
  AOI22_X1 U14838 ( .A1(\DataPath/RF/bus_reg_dataout[327] ), .A2(n8403), .B1(
        n11428), .B2(n11323), .ZN(n3740) );
  AOI22_X1 U14839 ( .A1(\DataPath/RF/bus_reg_dataout[328] ), .A2(n8403), .B1(
        n11324), .B2(n11382), .ZN(n3739) );
  AOI22_X1 U14840 ( .A1(\DataPath/RF/bus_reg_dataout[329] ), .A2(n11325), .B1(
        n11324), .B2(n11383), .ZN(n3738) );
  AOI22_X1 U14841 ( .A1(\DataPath/RF/bus_reg_dataout[330] ), .A2(n8403), .B1(
        n11324), .B2(n11384), .ZN(n3737) );
  AOI22_X1 U14842 ( .A1(\DataPath/RF/bus_reg_dataout[331] ), .A2(n8403), .B1(
        n11324), .B2(n11385), .ZN(n3736) );
  AOI22_X1 U14843 ( .A1(\DataPath/RF/bus_reg_dataout[332] ), .A2(n8403), .B1(
        n11324), .B2(n11386), .ZN(n3735) );
  AOI22_X1 U14844 ( .A1(n11434), .A2(n11323), .B1(n8403), .B2(
        \DataPath/RF/bus_reg_dataout[333] ), .ZN(n3734) );
  AOI22_X1 U14845 ( .A1(n11435), .A2(n11323), .B1(n11325), .B2(
        \DataPath/RF/bus_reg_dataout[334] ), .ZN(n3733) );
  AOI22_X1 U14846 ( .A1(\DataPath/RF/bus_reg_dataout[335] ), .A2(n8403), .B1(
        n11324), .B2(n11389), .ZN(n3732) );
  AOI22_X1 U14847 ( .A1(\DataPath/RF/bus_reg_dataout[336] ), .A2(n8403), .B1(
        n11324), .B2(n11390), .ZN(n3731) );
  AOI22_X1 U14848 ( .A1(n11438), .A2(n11323), .B1(n8403), .B2(
        \DataPath/RF/bus_reg_dataout[337] ), .ZN(n3730) );
  AOI22_X1 U14849 ( .A1(\DataPath/RF/bus_reg_dataout[338] ), .A2(n8403), .B1(
        n11439), .B2(n11323), .ZN(n3729) );
  AOI22_X1 U14850 ( .A1(\DataPath/RF/bus_reg_dataout[339] ), .A2(n11325), .B1(
        n11324), .B2(n11392), .ZN(n3728) );
  AOI22_X1 U14851 ( .A1(\DataPath/RF/bus_reg_dataout[340] ), .A2(n8403), .B1(
        n11441), .B2(n11323), .ZN(n3727) );
  AOI22_X1 U14852 ( .A1(\DataPath/RF/bus_reg_dataout[341] ), .A2(n11325), .B1(
        n11324), .B2(n11394), .ZN(n3726) );
  AOI22_X1 U14853 ( .A1(n11443), .A2(n11323), .B1(n11325), .B2(
        \DataPath/RF/bus_reg_dataout[342] ), .ZN(n3725) );
  AOI22_X1 U14854 ( .A1(\DataPath/RF/bus_reg_dataout[343] ), .A2(n8403), .B1(
        n11324), .B2(n11396), .ZN(n3724) );
  AOI22_X1 U14855 ( .A1(n11445), .A2(n11323), .B1(n8403), .B2(
        \DataPath/RF/bus_reg_dataout[344] ), .ZN(n3723) );
  AOI22_X1 U14856 ( .A1(\DataPath/RF/bus_reg_dataout[345] ), .A2(n8403), .B1(
        n11324), .B2(n11398), .ZN(n3722) );
  AOI22_X1 U14857 ( .A1(\DataPath/RF/bus_reg_dataout[346] ), .A2(n8403), .B1(
        n11324), .B2(n11399), .ZN(n3721) );
  AOI22_X1 U14858 ( .A1(\DataPath/RF/bus_reg_dataout[347] ), .A2(n8403), .B1(
        n11324), .B2(n11400), .ZN(n3720) );
  AOI22_X1 U14859 ( .A1(\DataPath/RF/bus_reg_dataout[348] ), .A2(n11325), .B1(
        n11324), .B2(n11401), .ZN(n3719) );
  AOI22_X1 U14860 ( .A1(\DataPath/RF/bus_reg_dataout[349] ), .A2(n8403), .B1(
        n11450), .B2(n11323), .ZN(n3718) );
  AOI22_X1 U14861 ( .A1(n11451), .A2(n11323), .B1(n11325), .B2(
        \DataPath/RF/bus_reg_dataout[350] ), .ZN(n3717) );
  AOI22_X1 U14862 ( .A1(\DataPath/RF/bus_reg_dataout[351] ), .A2(n11325), .B1(
        n11324), .B2(n11403), .ZN(n3714) );
  AOI22_X1 U14863 ( .A1(\DataPath/RF/bus_reg_dataout[288] ), .A2(n8404), .B1(
        n11330), .B2(n11378), .ZN(n3710) );
  AOI22_X1 U14864 ( .A1(\DataPath/RF/bus_reg_dataout[289] ), .A2(n8404), .B1(
        n11330), .B2(n11421), .ZN(n3709) );
  AOI22_X1 U14865 ( .A1(\DataPath/RF/bus_reg_dataout[290] ), .A2(n8404), .B1(
        n11330), .B2(n11422), .ZN(n3708) );
  AOI22_X1 U14866 ( .A1(\DataPath/RF/bus_reg_dataout[291] ), .A2(n8404), .B1(
        n11330), .B2(n11423), .ZN(n3707) );
  AOI22_X1 U14867 ( .A1(\DataPath/RF/bus_reg_dataout[292] ), .A2(n8404), .B1(
        n11330), .B2(n11379), .ZN(n3706) );
  AOI22_X1 U14868 ( .A1(\DataPath/RF/bus_reg_dataout[293] ), .A2(n8404), .B1(
        n11330), .B2(n11380), .ZN(n3705) );
  AOI22_X1 U14869 ( .A1(\DataPath/RF/bus_reg_dataout[294] ), .A2(n11331), .B1(
        n11330), .B2(n11426), .ZN(n3704) );
  AOI22_X1 U14870 ( .A1(\DataPath/RF/bus_reg_dataout[295] ), .A2(n8404), .B1(
        n11330), .B2(n11381), .ZN(n3703) );
  AOI22_X1 U14871 ( .A1(\DataPath/RF/bus_reg_dataout[296] ), .A2(n11331), .B1(
        n11330), .B2(n11382), .ZN(n3702) );
  AOI22_X1 U14872 ( .A1(\DataPath/RF/bus_reg_dataout[297] ), .A2(n8404), .B1(
        n11330), .B2(n11383), .ZN(n3701) );
  AOI22_X1 U14873 ( .A1(\DataPath/RF/bus_reg_dataout[298] ), .A2(n8404), .B1(
        n11330), .B2(n11384), .ZN(n3700) );
  AOI22_X1 U14874 ( .A1(n11432), .A2(n11329), .B1(n11331), .B2(
        \DataPath/RF/bus_reg_dataout[299] ), .ZN(n3699) );
  AOI22_X1 U14875 ( .A1(\DataPath/RF/bus_reg_dataout[300] ), .A2(n8404), .B1(
        n11330), .B2(n11386), .ZN(n3698) );
  AOI22_X1 U14876 ( .A1(\DataPath/RF/bus_reg_dataout[301] ), .A2(n11331), .B1(
        n11330), .B2(n11387), .ZN(n3697) );
  AOI22_X1 U14877 ( .A1(n11435), .A2(n11329), .B1(n8404), .B2(
        \DataPath/RF/bus_reg_dataout[302] ), .ZN(n3696) );
  AOI22_X1 U14878 ( .A1(\DataPath/RF/bus_reg_dataout[303] ), .A2(n11331), .B1(
        n11330), .B2(n11389), .ZN(n3695) );
  AOI22_X1 U14879 ( .A1(\DataPath/RF/bus_reg_dataout[304] ), .A2(n8404), .B1(
        n11330), .B2(n11390), .ZN(n3694) );
  AOI22_X1 U14880 ( .A1(\DataPath/RF/bus_reg_dataout[305] ), .A2(n8404), .B1(
        n11330), .B2(n11410), .ZN(n3693) );
  AOI22_X1 U14881 ( .A1(\DataPath/RF/bus_reg_dataout[306] ), .A2(n8404), .B1(
        n11330), .B2(n11391), .ZN(n3692) );
  AOI22_X1 U14882 ( .A1(\DataPath/RF/bus_reg_dataout[307] ), .A2(n11331), .B1(
        n11330), .B2(n11392), .ZN(n3691) );
  INV_X1 U14883 ( .A(n11331), .ZN(n11328) );
  AOI22_X1 U14884 ( .A1(n8404), .A2(\DataPath/RF/bus_reg_dataout[308] ), .B1(
        n11441), .B2(n11328), .ZN(n3690) );
  AOI22_X1 U14885 ( .A1(\DataPath/RF/bus_reg_dataout[309] ), .A2(n8404), .B1(
        n11330), .B2(n11394), .ZN(n3689) );
  AOI22_X1 U14886 ( .A1(n11443), .A2(n11329), .B1(n11331), .B2(
        \DataPath/RF/bus_reg_dataout[310] ), .ZN(n3688) );
  AOI22_X1 U14887 ( .A1(\DataPath/RF/bus_reg_dataout[311] ), .A2(n8404), .B1(
        n11330), .B2(n11396), .ZN(n3687) );
  AOI22_X1 U14888 ( .A1(\DataPath/RF/bus_reg_dataout[312] ), .A2(n8404), .B1(
        n11330), .B2(n11397), .ZN(n3686) );
  AOI22_X1 U14889 ( .A1(\DataPath/RF/bus_reg_dataout[313] ), .A2(n8404), .B1(
        n11330), .B2(n11398), .ZN(n3685) );
  AOI22_X1 U14890 ( .A1(\DataPath/RF/bus_reg_dataout[314] ), .A2(n11331), .B1(
        n11330), .B2(n11399), .ZN(n3684) );
  AOI22_X1 U14891 ( .A1(\DataPath/RF/bus_reg_dataout[315] ), .A2(n8404), .B1(
        n11330), .B2(n11400), .ZN(n3683) );
  AOI22_X1 U14892 ( .A1(\DataPath/RF/bus_reg_dataout[316] ), .A2(n8404), .B1(
        n11330), .B2(n11401), .ZN(n3682) );
  AOI22_X1 U14893 ( .A1(\DataPath/RF/bus_reg_dataout[317] ), .A2(n8404), .B1(
        n11330), .B2(n11402), .ZN(n3681) );
  AOI22_X1 U14894 ( .A1(\DataPath/RF/bus_reg_dataout[318] ), .A2(n11331), .B1(
        n11330), .B2(n11411), .ZN(n3680) );
  AOI22_X1 U14895 ( .A1(\DataPath/RF/bus_reg_dataout[319] ), .A2(n8404), .B1(
        n11330), .B2(n11403), .ZN(n3677) );
  AOI22_X1 U14896 ( .A1(\DataPath/RF/bus_reg_dataout[256] ), .A2(n8405), .B1(
        n11336), .B2(n11378), .ZN(n3673) );
  AOI22_X1 U14897 ( .A1(\DataPath/RF/bus_reg_dataout[257] ), .A2(n8405), .B1(
        n11336), .B2(n11421), .ZN(n3672) );
  AOI22_X1 U14898 ( .A1(\DataPath/RF/bus_reg_dataout[258] ), .A2(n8405), .B1(
        n11336), .B2(n11422), .ZN(n3671) );
  AOI22_X1 U14899 ( .A1(\DataPath/RF/bus_reg_dataout[259] ), .A2(n8405), .B1(
        n11336), .B2(n11423), .ZN(n3670) );
  AOI22_X1 U14900 ( .A1(\DataPath/RF/bus_reg_dataout[260] ), .A2(n8405), .B1(
        n11336), .B2(n11379), .ZN(n3669) );
  AOI22_X1 U14901 ( .A1(\DataPath/RF/bus_reg_dataout[261] ), .A2(n8405), .B1(
        n11336), .B2(n11380), .ZN(n3668) );
  AOI22_X1 U14902 ( .A1(\DataPath/RF/bus_reg_dataout[262] ), .A2(n11337), .B1(
        n11336), .B2(n11426), .ZN(n3667) );
  AOI22_X1 U14903 ( .A1(\DataPath/RF/bus_reg_dataout[263] ), .A2(n8405), .B1(
        n11336), .B2(n11381), .ZN(n3666) );
  AOI22_X1 U14904 ( .A1(\DataPath/RF/bus_reg_dataout[264] ), .A2(n11337), .B1(
        n11336), .B2(n11382), .ZN(n3665) );
  AOI22_X1 U14905 ( .A1(\DataPath/RF/bus_reg_dataout[265] ), .A2(n8405), .B1(
        n11336), .B2(n11383), .ZN(n3664) );
  AOI22_X1 U14906 ( .A1(\DataPath/RF/bus_reg_dataout[266] ), .A2(n8405), .B1(
        n11336), .B2(n11384), .ZN(n3663) );
  AOI22_X1 U14907 ( .A1(\DataPath/RF/bus_reg_dataout[267] ), .A2(n8405), .B1(
        n11336), .B2(n11385), .ZN(n3662) );
  AOI22_X1 U14908 ( .A1(\DataPath/RF/bus_reg_dataout[268] ), .A2(n8405), .B1(
        n11336), .B2(n11386), .ZN(n3661) );
  AOI22_X1 U14909 ( .A1(\DataPath/RF/bus_reg_dataout[269] ), .A2(n11337), .B1(
        n11336), .B2(n11387), .ZN(n3660) );
  AOI22_X1 U14910 ( .A1(\DataPath/RF/bus_reg_dataout[270] ), .A2(n8405), .B1(
        n11336), .B2(n11388), .ZN(n3659) );
  AOI22_X1 U14911 ( .A1(\DataPath/RF/bus_reg_dataout[271] ), .A2(n8405), .B1(
        n11336), .B2(n11389), .ZN(n3658) );
  AOI22_X1 U14912 ( .A1(\DataPath/RF/bus_reg_dataout[272] ), .A2(n8405), .B1(
        n11336), .B2(n11390), .ZN(n3657) );
  AOI22_X1 U14913 ( .A1(\DataPath/RF/bus_reg_dataout[273] ), .A2(n11337), .B1(
        n11336), .B2(n11410), .ZN(n3656) );
  AOI22_X1 U14914 ( .A1(\DataPath/RF/bus_reg_dataout[274] ), .A2(n8405), .B1(
        n11336), .B2(n11391), .ZN(n3655) );
  AOI22_X1 U14915 ( .A1(\DataPath/RF/bus_reg_dataout[275] ), .A2(n8405), .B1(
        n11336), .B2(n11392), .ZN(n3654) );
  INV_X1 U14916 ( .A(n11337), .ZN(n11334) );
  AOI22_X1 U14917 ( .A1(n8405), .A2(\DataPath/RF/bus_reg_dataout[276] ), .B1(
        n11441), .B2(n11334), .ZN(n3653) );
  AOI22_X1 U14918 ( .A1(\DataPath/RF/bus_reg_dataout[277] ), .A2(n8405), .B1(
        n11336), .B2(n11394), .ZN(n3652) );
  AOI22_X1 U14919 ( .A1(\DataPath/RF/bus_reg_dataout[278] ), .A2(n11337), .B1(
        n11336), .B2(n11395), .ZN(n3651) );
  AOI22_X1 U14920 ( .A1(\DataPath/RF/bus_reg_dataout[279] ), .A2(n11337), .B1(
        n11336), .B2(n11396), .ZN(n3650) );
  AOI22_X1 U14921 ( .A1(n11445), .A2(n11335), .B1(n11337), .B2(
        \DataPath/RF/bus_reg_dataout[280] ), .ZN(n3649) );
  AOI22_X1 U14922 ( .A1(n11446), .A2(n11335), .B1(n8405), .B2(
        \DataPath/RF/bus_reg_dataout[281] ), .ZN(n3648) );
  AOI22_X1 U14923 ( .A1(\DataPath/RF/bus_reg_dataout[282] ), .A2(n8405), .B1(
        n11336), .B2(n11399), .ZN(n3647) );
  AOI22_X1 U14924 ( .A1(n11448), .A2(n11335), .B1(n11337), .B2(
        \DataPath/RF/bus_reg_dataout[283] ), .ZN(n3646) );
  AOI22_X1 U14925 ( .A1(\DataPath/RF/bus_reg_dataout[284] ), .A2(n8405), .B1(
        n11336), .B2(n11401), .ZN(n3645) );
  AOI22_X1 U14926 ( .A1(\DataPath/RF/bus_reg_dataout[285] ), .A2(n8405), .B1(
        n11336), .B2(n11402), .ZN(n3644) );
  AOI22_X1 U14927 ( .A1(\DataPath/RF/bus_reg_dataout[286] ), .A2(n11337), .B1(
        n11336), .B2(n11411), .ZN(n3643) );
  AOI22_X1 U14928 ( .A1(\DataPath/RF/bus_reg_dataout[287] ), .A2(n8405), .B1(
        n11336), .B2(n11403), .ZN(n3640) );
  OAI22_X1 U14929 ( .A1(n8450), .A2(n11339), .B1(n11415), .B2(n11338), .ZN(
        n11340) );
  AOI22_X1 U14930 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[224] ), .B1(
        n11420), .B2(n11343), .ZN(n3635) );
  NOR2_X1 U14931 ( .A1(RST), .A2(n11344), .ZN(n11342) );
  AOI22_X1 U14932 ( .A1(\DataPath/RF/bus_reg_dataout[225] ), .A2(n11344), .B1(
        n11342), .B2(n11421), .ZN(n3634) );
  AOI22_X1 U14933 ( .A1(\DataPath/RF/bus_reg_dataout[226] ), .A2(n11344), .B1(
        n11342), .B2(n11422), .ZN(n3633) );
  AOI22_X1 U14934 ( .A1(\DataPath/RF/bus_reg_dataout[227] ), .A2(n11344), .B1(
        n11342), .B2(n11423), .ZN(n3632) );
  AOI22_X1 U14935 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[228] ), .B1(
        n11424), .B2(n11343), .ZN(n3631) );
  AOI22_X1 U14936 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[229] ), .B1(
        n11425), .B2(n11343), .ZN(n3630) );
  AOI22_X1 U14937 ( .A1(\DataPath/RF/bus_reg_dataout[230] ), .A2(n11344), .B1(
        n11342), .B2(n11426), .ZN(n3629) );
  AOI22_X1 U14938 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[231] ), .B1(
        n11428), .B2(n11343), .ZN(n3628) );
  AOI22_X1 U14939 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[232] ), .B1(
        n11429), .B2(n11343), .ZN(n3627) );
  AOI22_X1 U14940 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[233] ), .B1(
        n11430), .B2(n11343), .ZN(n3626) );
  AOI22_X1 U14941 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[234] ), .B1(
        n11431), .B2(n11343), .ZN(n3625) );
  AOI22_X1 U14942 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[235] ), .B1(
        n11432), .B2(n11343), .ZN(n3624) );
  AOI22_X1 U14943 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[236] ), .B1(
        n11433), .B2(n11343), .ZN(n3623) );
  AOI22_X1 U14944 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[237] ), .B1(
        n11434), .B2(n11343), .ZN(n3622) );
  AOI22_X1 U14945 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[238] ), .B1(
        n11435), .B2(n11343), .ZN(n3621) );
  AOI22_X1 U14946 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[239] ), .B1(
        n11436), .B2(n11343), .ZN(n3620) );
  AOI22_X1 U14947 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[240] ), .B1(
        n11437), .B2(n11343), .ZN(n3619) );
  AOI22_X1 U14948 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[241] ), .B1(
        n11438), .B2(n11343), .ZN(n3618) );
  AOI22_X1 U14949 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[242] ), .B1(
        n11439), .B2(n11343), .ZN(n3617) );
  AOI22_X1 U14950 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[243] ), .B1(
        n11440), .B2(n11343), .ZN(n3616) );
  AOI22_X1 U14951 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[244] ), .B1(
        n11441), .B2(n11343), .ZN(n3615) );
  AOI22_X1 U14952 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[245] ), .B1(
        n11442), .B2(n11343), .ZN(n3614) );
  AOI22_X1 U14953 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[246] ), .B1(
        n11443), .B2(n11343), .ZN(n3613) );
  AOI22_X1 U14954 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[247] ), .B1(
        n11444), .B2(n11343), .ZN(n3612) );
  AOI22_X1 U14955 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[248] ), .B1(
        n11445), .B2(n11343), .ZN(n3611) );
  AOI22_X1 U14956 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[249] ), .B1(
        n11446), .B2(n11343), .ZN(n3610) );
  AOI22_X1 U14957 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[250] ), .B1(
        n11447), .B2(n11343), .ZN(n3609) );
  AOI22_X1 U14958 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[251] ), .B1(
        n11448), .B2(n11343), .ZN(n3608) );
  AOI22_X1 U14959 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[252] ), .B1(
        n11449), .B2(n11343), .ZN(n3607) );
  AOI22_X1 U14960 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[253] ), .B1(
        n11450), .B2(n11343), .ZN(n3606) );
  AOI22_X1 U14961 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[254] ), .B1(
        n11451), .B2(n11343), .ZN(n3605) );
  AOI22_X1 U14962 ( .A1(n11344), .A2(\DataPath/RF/bus_reg_dataout[255] ), .B1(
        n11597), .B2(n11343), .ZN(n3602) );
  OAI22_X1 U14963 ( .A1(n8450), .A2(n11346), .B1(n7756), .B2(n11345), .ZN(
        n11347) );
  AOI22_X1 U14964 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[192] ), .B1(
        n11420), .B2(n11350), .ZN(n3597) );
  NOR2_X1 U14965 ( .A1(RST), .A2(n11351), .ZN(n11349) );
  AOI22_X1 U14966 ( .A1(\DataPath/RF/bus_reg_dataout[193] ), .A2(n11351), .B1(
        n11349), .B2(n11421), .ZN(n3596) );
  AOI22_X1 U14967 ( .A1(\DataPath/RF/bus_reg_dataout[194] ), .A2(n11351), .B1(
        n11349), .B2(n11422), .ZN(n3595) );
  AOI22_X1 U14968 ( .A1(\DataPath/RF/bus_reg_dataout[195] ), .A2(n11351), .B1(
        n11349), .B2(n11423), .ZN(n3594) );
  AOI22_X1 U14969 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[196] ), .B1(
        n11424), .B2(n11350), .ZN(n3593) );
  AOI22_X1 U14970 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[197] ), .B1(
        n11425), .B2(n11350), .ZN(n3592) );
  AOI22_X1 U14971 ( .A1(\DataPath/RF/bus_reg_dataout[198] ), .A2(n11351), .B1(
        n11349), .B2(n11426), .ZN(n3591) );
  AOI22_X1 U14972 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[199] ), .B1(
        n11428), .B2(n11350), .ZN(n3590) );
  AOI22_X1 U14973 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[200] ), .B1(
        n11429), .B2(n11350), .ZN(n3589) );
  AOI22_X1 U14974 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[201] ), .B1(
        n11430), .B2(n11350), .ZN(n3588) );
  AOI22_X1 U14975 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[202] ), .B1(
        n11431), .B2(n11350), .ZN(n3587) );
  AOI22_X1 U14976 ( .A1(\DataPath/RF/bus_reg_dataout[203] ), .A2(n11351), .B1(
        n11349), .B2(n11385), .ZN(n3586) );
  AOI22_X1 U14977 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[204] ), .B1(
        n11433), .B2(n11350), .ZN(n3585) );
  AOI22_X1 U14978 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[205] ), .B1(
        n11434), .B2(n11350), .ZN(n3584) );
  AOI22_X1 U14979 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[206] ), .B1(
        n11435), .B2(n11350), .ZN(n3583) );
  AOI22_X1 U14980 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[207] ), .B1(
        n11436), .B2(n11350), .ZN(n3582) );
  AOI22_X1 U14981 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[208] ), .B1(
        n11437), .B2(n11350), .ZN(n3581) );
  AOI22_X1 U14982 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[209] ), .B1(
        n11438), .B2(n11350), .ZN(n3580) );
  AOI22_X1 U14983 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[210] ), .B1(
        n11439), .B2(n11350), .ZN(n3579) );
  AOI22_X1 U14984 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[211] ), .B1(
        n11440), .B2(n11350), .ZN(n3578) );
  AOI22_X1 U14985 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[212] ), .B1(
        n11441), .B2(n11350), .ZN(n3577) );
  AOI22_X1 U14986 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[213] ), .B1(
        n11442), .B2(n11350), .ZN(n3576) );
  AOI22_X1 U14987 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[214] ), .B1(
        n11443), .B2(n11350), .ZN(n3575) );
  AOI22_X1 U14988 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[215] ), .B1(
        n11444), .B2(n11350), .ZN(n3574) );
  AOI22_X1 U14989 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[216] ), .B1(
        n11445), .B2(n11350), .ZN(n3573) );
  AOI22_X1 U14990 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[217] ), .B1(
        n11446), .B2(n11350), .ZN(n3572) );
  AOI22_X1 U14991 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[218] ), .B1(
        n11447), .B2(n11350), .ZN(n3571) );
  AOI22_X1 U14992 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[219] ), .B1(
        n11448), .B2(n11350), .ZN(n3570) );
  AOI22_X1 U14993 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[220] ), .B1(
        n11449), .B2(n11350), .ZN(n3569) );
  AOI22_X1 U14994 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[221] ), .B1(
        n11450), .B2(n11350), .ZN(n3568) );
  AOI22_X1 U14995 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[222] ), .B1(
        n11451), .B2(n11350), .ZN(n3567) );
  AOI22_X1 U14996 ( .A1(n11351), .A2(\DataPath/RF/bus_reg_dataout[223] ), .B1(
        n11597), .B2(n11350), .ZN(n3564) );
  OAI22_X1 U14997 ( .A1(n8450), .A2(n11353), .B1(n7756), .B2(n11352), .ZN(
        n11354) );
  AOI22_X1 U14998 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[160] ), .B1(
        n11420), .B2(n11357), .ZN(n3559) );
  AOI22_X1 U14999 ( .A1(\DataPath/RF/bus_reg_dataout[161] ), .A2(n11358), .B1(
        n11356), .B2(n11421), .ZN(n3558) );
  AOI22_X1 U15000 ( .A1(\DataPath/RF/bus_reg_dataout[162] ), .A2(n11358), .B1(
        n11356), .B2(n11422), .ZN(n3557) );
  AOI22_X1 U15001 ( .A1(\DataPath/RF/bus_reg_dataout[163] ), .A2(n11358), .B1(
        n11356), .B2(n11423), .ZN(n3556) );
  AOI22_X1 U15002 ( .A1(\DataPath/RF/bus_reg_dataout[164] ), .A2(n11358), .B1(
        n11356), .B2(n11379), .ZN(n3555) );
  AOI22_X1 U15003 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[165] ), .B1(
        n11425), .B2(n11357), .ZN(n3554) );
  AOI22_X1 U15004 ( .A1(\DataPath/RF/bus_reg_dataout[166] ), .A2(n11358), .B1(
        n11356), .B2(n11426), .ZN(n3553) );
  AOI22_X1 U15005 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[167] ), .B1(
        n11428), .B2(n11357), .ZN(n3552) );
  AOI22_X1 U15006 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[168] ), .B1(
        n11429), .B2(n11357), .ZN(n3551) );
  AOI22_X1 U15007 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[169] ), .B1(
        n11430), .B2(n11357), .ZN(n3550) );
  AOI22_X1 U15008 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[170] ), .B1(
        n11431), .B2(n11357), .ZN(n3549) );
  AOI22_X1 U15009 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[171] ), .B1(
        n11432), .B2(n11357), .ZN(n3548) );
  AOI22_X1 U15010 ( .A1(\DataPath/RF/bus_reg_dataout[172] ), .A2(n11358), .B1(
        n11356), .B2(n11386), .ZN(n3547) );
  AOI22_X1 U15011 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[173] ), .B1(
        n11434), .B2(n11357), .ZN(n3546) );
  AOI22_X1 U15012 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[174] ), .B1(
        n11435), .B2(n11357), .ZN(n3545) );
  AOI22_X1 U15013 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[175] ), .B1(
        n11436), .B2(n11357), .ZN(n3544) );
  AOI22_X1 U15014 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[176] ), .B1(
        n11437), .B2(n11357), .ZN(n3543) );
  AOI22_X1 U15015 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[177] ), .B1(
        n11438), .B2(n11357), .ZN(n3542) );
  AOI22_X1 U15016 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[178] ), .B1(
        n11439), .B2(n11357), .ZN(n3541) );
  AOI22_X1 U15017 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[179] ), .B1(
        n11440), .B2(n11357), .ZN(n3540) );
  AOI22_X1 U15018 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[180] ), .B1(
        n11441), .B2(n11357), .ZN(n3539) );
  AOI22_X1 U15019 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[181] ), .B1(
        n11442), .B2(n11357), .ZN(n3538) );
  AOI22_X1 U15020 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[182] ), .B1(
        n11443), .B2(n11357), .ZN(n3537) );
  AOI22_X1 U15021 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[183] ), .B1(
        n11444), .B2(n11357), .ZN(n3536) );
  AOI22_X1 U15022 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[184] ), .B1(
        n11445), .B2(n11357), .ZN(n3535) );
  AOI22_X1 U15023 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[185] ), .B1(
        n11446), .B2(n11357), .ZN(n3534) );
  AOI22_X1 U15024 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[186] ), .B1(
        n11447), .B2(n11357), .ZN(n3533) );
  AOI22_X1 U15025 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[187] ), .B1(
        n11448), .B2(n11357), .ZN(n3532) );
  AOI22_X1 U15026 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[188] ), .B1(
        n11449), .B2(n11357), .ZN(n3531) );
  AOI22_X1 U15027 ( .A1(\DataPath/RF/bus_reg_dataout[189] ), .A2(n11358), .B1(
        n11356), .B2(n11402), .ZN(n3530) );
  AOI22_X1 U15028 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[190] ), .B1(
        n11451), .B2(n11357), .ZN(n3529) );
  AOI22_X1 U15029 ( .A1(n11358), .A2(\DataPath/RF/bus_reg_dataout[191] ), .B1(
        n11597), .B2(n11357), .ZN(n3526) );
  OAI222_X1 U15030 ( .A1(n11361), .A2(n7756), .B1(n11360), .B2(n8173), .C1(
        n11359), .C2(n11415), .ZN(n11362) );
  AOI22_X1 U15031 ( .A1(\DataPath/RF/bus_reg_dataout[128] ), .A2(n8406), .B1(
        n11364), .B2(n11378), .ZN(n3521) );
  AOI22_X1 U15032 ( .A1(\DataPath/RF/bus_reg_dataout[129] ), .A2(n8406), .B1(
        n11364), .B2(n11421), .ZN(n3520) );
  AOI22_X1 U15033 ( .A1(\DataPath/RF/bus_reg_dataout[130] ), .A2(n8406), .B1(
        n11364), .B2(n11422), .ZN(n3519) );
  AOI22_X1 U15034 ( .A1(\DataPath/RF/bus_reg_dataout[131] ), .A2(n8406), .B1(
        n11364), .B2(n11423), .ZN(n3518) );
  AOI22_X1 U15035 ( .A1(\DataPath/RF/bus_reg_dataout[132] ), .A2(n8406), .B1(
        n11364), .B2(n11379), .ZN(n3517) );
  AOI22_X1 U15036 ( .A1(\DataPath/RF/bus_reg_dataout[133] ), .A2(n8406), .B1(
        n11364), .B2(n11380), .ZN(n3516) );
  AOI22_X1 U15037 ( .A1(\DataPath/RF/bus_reg_dataout[134] ), .A2(n8406), .B1(
        n11364), .B2(n11426), .ZN(n3515) );
  AOI22_X1 U15038 ( .A1(\DataPath/RF/bus_reg_dataout[135] ), .A2(n11365), .B1(
        n11364), .B2(n11381), .ZN(n3514) );
  AOI22_X1 U15039 ( .A1(\DataPath/RF/bus_reg_dataout[136] ), .A2(n8406), .B1(
        n11364), .B2(n11382), .ZN(n3513) );
  AOI22_X1 U15040 ( .A1(\DataPath/RF/bus_reg_dataout[137] ), .A2(n8406), .B1(
        n11364), .B2(n11383), .ZN(n3512) );
  AOI22_X1 U15041 ( .A1(\DataPath/RF/bus_reg_dataout[138] ), .A2(n8406), .B1(
        n11364), .B2(n11384), .ZN(n3511) );
  AOI22_X1 U15042 ( .A1(\DataPath/RF/bus_reg_dataout[139] ), .A2(n11365), .B1(
        n11364), .B2(n11385), .ZN(n3510) );
  AOI22_X1 U15043 ( .A1(\DataPath/RF/bus_reg_dataout[140] ), .A2(n8406), .B1(
        n11364), .B2(n11386), .ZN(n3509) );
  AOI22_X1 U15044 ( .A1(\DataPath/RF/bus_reg_dataout[141] ), .A2(n8406), .B1(
        n11364), .B2(n11387), .ZN(n3508) );
  AOI22_X1 U15045 ( .A1(\DataPath/RF/bus_reg_dataout[142] ), .A2(n11365), .B1(
        n11364), .B2(n11388), .ZN(n3507) );
  AOI22_X1 U15046 ( .A1(\DataPath/RF/bus_reg_dataout[143] ), .A2(n11365), .B1(
        n11364), .B2(n11389), .ZN(n3506) );
  AOI22_X1 U15047 ( .A1(\DataPath/RF/bus_reg_dataout[144] ), .A2(n8406), .B1(
        n11364), .B2(n11390), .ZN(n3505) );
  AOI22_X1 U15048 ( .A1(\DataPath/RF/bus_reg_dataout[145] ), .A2(n8406), .B1(
        n11364), .B2(n11410), .ZN(n3504) );
  AOI22_X1 U15049 ( .A1(\DataPath/RF/bus_reg_dataout[146] ), .A2(n11365), .B1(
        n11364), .B2(n11391), .ZN(n3503) );
  AOI22_X1 U15050 ( .A1(\DataPath/RF/bus_reg_dataout[147] ), .A2(n8406), .B1(
        n11364), .B2(n11392), .ZN(n3502) );
  INV_X1 U15051 ( .A(n11365), .ZN(n11363) );
  AOI22_X1 U15052 ( .A1(n11365), .A2(\DataPath/RF/bus_reg_dataout[148] ), .B1(
        n11441), .B2(n11363), .ZN(n3501) );
  AOI22_X1 U15053 ( .A1(\DataPath/RF/bus_reg_dataout[149] ), .A2(n8406), .B1(
        n11364), .B2(n11394), .ZN(n3500) );
  AOI22_X1 U15054 ( .A1(\DataPath/RF/bus_reg_dataout[150] ), .A2(n8406), .B1(
        n11364), .B2(n11395), .ZN(n3499) );
  AOI22_X1 U15055 ( .A1(\DataPath/RF/bus_reg_dataout[151] ), .A2(n8406), .B1(
        n11364), .B2(n11396), .ZN(n3498) );
  AOI22_X1 U15056 ( .A1(\DataPath/RF/bus_reg_dataout[152] ), .A2(n8406), .B1(
        n11364), .B2(n11397), .ZN(n3497) );
  AOI22_X1 U15057 ( .A1(\DataPath/RF/bus_reg_dataout[153] ), .A2(n8406), .B1(
        n11364), .B2(n11398), .ZN(n3496) );
  AOI22_X1 U15058 ( .A1(\DataPath/RF/bus_reg_dataout[154] ), .A2(n8406), .B1(
        n11364), .B2(n11399), .ZN(n3495) );
  AOI22_X1 U15059 ( .A1(\DataPath/RF/bus_reg_dataout[155] ), .A2(n11365), .B1(
        n11364), .B2(n11400), .ZN(n3494) );
  AOI22_X1 U15060 ( .A1(\DataPath/RF/bus_reg_dataout[156] ), .A2(n8406), .B1(
        n11364), .B2(n11401), .ZN(n3493) );
  AOI22_X1 U15061 ( .A1(\DataPath/RF/bus_reg_dataout[157] ), .A2(n8406), .B1(
        n11364), .B2(n11402), .ZN(n3492) );
  AOI22_X1 U15062 ( .A1(\DataPath/RF/bus_reg_dataout[158] ), .A2(n8406), .B1(
        n11364), .B2(n11411), .ZN(n3491) );
  AOI22_X1 U15063 ( .A1(\DataPath/RF/bus_reg_dataout[159] ), .A2(n8406), .B1(
        n11364), .B2(n11403), .ZN(n3488) );
  OAI22_X1 U15064 ( .A1(n8450), .A2(n11367), .B1(n7756), .B2(n11366), .ZN(
        n11368) );
  AOI22_X1 U15065 ( .A1(\DataPath/RF/bus_reg_dataout[96] ), .A2(n11372), .B1(
        n11370), .B2(n11378), .ZN(n3483) );
  AOI22_X1 U15066 ( .A1(\DataPath/RF/bus_reg_dataout[97] ), .A2(n11372), .B1(
        n11370), .B2(n11421), .ZN(n3482) );
  AOI22_X1 U15067 ( .A1(\DataPath/RF/bus_reg_dataout[98] ), .A2(n11372), .B1(
        n11370), .B2(n11422), .ZN(n3481) );
  AOI22_X1 U15068 ( .A1(\DataPath/RF/bus_reg_dataout[99] ), .A2(n11372), .B1(
        n11370), .B2(n11423), .ZN(n3480) );
  AOI22_X1 U15069 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[100] ), .B1(
        n11424), .B2(n11371), .ZN(n3479) );
  AOI22_X1 U15070 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[101] ), .B1(
        n11425), .B2(n11371), .ZN(n3478) );
  AOI22_X1 U15071 ( .A1(\DataPath/RF/bus_reg_dataout[102] ), .A2(n11372), .B1(
        n11370), .B2(n11426), .ZN(n3477) );
  AOI22_X1 U15072 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[103] ), .B1(
        n11428), .B2(n11371), .ZN(n3476) );
  AOI22_X1 U15073 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[104] ), .B1(
        n11429), .B2(n11371), .ZN(n3475) );
  AOI22_X1 U15074 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[105] ), .B1(
        n11430), .B2(n11371), .ZN(n3474) );
  AOI22_X1 U15075 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[106] ), .B1(
        n11431), .B2(n11371), .ZN(n3473) );
  AOI22_X1 U15076 ( .A1(\DataPath/RF/bus_reg_dataout[107] ), .A2(n11372), .B1(
        n11370), .B2(n11385), .ZN(n3472) );
  AOI22_X1 U15077 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[108] ), .B1(
        n11433), .B2(n11371), .ZN(n3471) );
  AOI22_X1 U15078 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[109] ), .B1(
        n11434), .B2(n11371), .ZN(n3470) );
  AOI22_X1 U15079 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[110] ), .B1(
        n11435), .B2(n11371), .ZN(n3469) );
  AOI22_X1 U15080 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[111] ), .B1(
        n11436), .B2(n11371), .ZN(n3468) );
  AOI22_X1 U15081 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[112] ), .B1(
        n11437), .B2(n11371), .ZN(n3467) );
  AOI22_X1 U15082 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[113] ), .B1(
        n11438), .B2(n11371), .ZN(n3466) );
  AOI22_X1 U15083 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[114] ), .B1(
        n11439), .B2(n11371), .ZN(n3465) );
  AOI22_X1 U15084 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[115] ), .B1(
        n11440), .B2(n11371), .ZN(n3464) );
  AOI22_X1 U15085 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[116] ), .B1(
        n11441), .B2(n11371), .ZN(n3463) );
  AOI22_X1 U15086 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[117] ), .B1(
        n11442), .B2(n11371), .ZN(n3462) );
  AOI22_X1 U15087 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[118] ), .B1(
        n11443), .B2(n11371), .ZN(n3461) );
  AOI22_X1 U15088 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[119] ), .B1(
        n11444), .B2(n11371), .ZN(n3460) );
  AOI22_X1 U15089 ( .A1(\DataPath/RF/bus_reg_dataout[120] ), .A2(n11372), .B1(
        n11370), .B2(n11397), .ZN(n3459) );
  AOI22_X1 U15090 ( .A1(\DataPath/RF/bus_reg_dataout[121] ), .A2(n11372), .B1(
        n11370), .B2(n11398), .ZN(n3458) );
  AOI22_X1 U15091 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[122] ), .B1(
        n11447), .B2(n11371), .ZN(n3457) );
  AOI22_X1 U15092 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[123] ), .B1(
        n11448), .B2(n11371), .ZN(n3456) );
  AOI22_X1 U15093 ( .A1(\DataPath/RF/bus_reg_dataout[124] ), .A2(n11372), .B1(
        n11370), .B2(n11401), .ZN(n3455) );
  AOI22_X1 U15094 ( .A1(\DataPath/RF/bus_reg_dataout[125] ), .A2(n11372), .B1(
        n11370), .B2(n11402), .ZN(n3454) );
  AOI22_X1 U15095 ( .A1(\DataPath/RF/bus_reg_dataout[126] ), .A2(n11372), .B1(
        n11370), .B2(n11411), .ZN(n3453) );
  AOI22_X1 U15096 ( .A1(n11372), .A2(\DataPath/RF/bus_reg_dataout[127] ), .B1(
        n11597), .B2(n11371), .ZN(n3450) );
  INV_X1 U15097 ( .A(n11373), .ZN(n11376) );
  OAI222_X1 U15098 ( .A1(n11376), .A2(n7756), .B1(n11375), .B2(n8173), .C1(
        n11415), .C2(n11374), .ZN(n11377) );
  AOI22_X1 U15099 ( .A1(\DataPath/RF/bus_reg_dataout[64] ), .A2(n8407), .B1(
        n11404), .B2(n11378), .ZN(n3445) );
  AOI22_X1 U15100 ( .A1(\DataPath/RF/bus_reg_dataout[65] ), .A2(n8407), .B1(
        n11404), .B2(n11421), .ZN(n3444) );
  AOI22_X1 U15101 ( .A1(\DataPath/RF/bus_reg_dataout[66] ), .A2(n8407), .B1(
        n11404), .B2(n11422), .ZN(n3443) );
  AOI22_X1 U15102 ( .A1(\DataPath/RF/bus_reg_dataout[67] ), .A2(n8407), .B1(
        n11404), .B2(n11423), .ZN(n3442) );
  AOI22_X1 U15103 ( .A1(\DataPath/RF/bus_reg_dataout[68] ), .A2(n8407), .B1(
        n11404), .B2(n11379), .ZN(n3441) );
  AOI22_X1 U15104 ( .A1(\DataPath/RF/bus_reg_dataout[69] ), .A2(n8407), .B1(
        n11404), .B2(n11380), .ZN(n3440) );
  AOI22_X1 U15105 ( .A1(\DataPath/RF/bus_reg_dataout[70] ), .A2(n8407), .B1(
        n11404), .B2(n11426), .ZN(n3439) );
  AOI22_X1 U15106 ( .A1(\DataPath/RF/bus_reg_dataout[71] ), .A2(n11405), .B1(
        n11404), .B2(n11381), .ZN(n3438) );
  AOI22_X1 U15107 ( .A1(\DataPath/RF/bus_reg_dataout[72] ), .A2(n8407), .B1(
        n11404), .B2(n11382), .ZN(n3437) );
  AOI22_X1 U15108 ( .A1(\DataPath/RF/bus_reg_dataout[73] ), .A2(n8407), .B1(
        n11404), .B2(n11383), .ZN(n3436) );
  AOI22_X1 U15109 ( .A1(\DataPath/RF/bus_reg_dataout[74] ), .A2(n8407), .B1(
        n11404), .B2(n11384), .ZN(n3435) );
  AOI22_X1 U15110 ( .A1(\DataPath/RF/bus_reg_dataout[75] ), .A2(n11405), .B1(
        n11404), .B2(n11385), .ZN(n3434) );
  AOI22_X1 U15111 ( .A1(\DataPath/RF/bus_reg_dataout[76] ), .A2(n8407), .B1(
        n11404), .B2(n11386), .ZN(n3433) );
  AOI22_X1 U15112 ( .A1(\DataPath/RF/bus_reg_dataout[77] ), .A2(n8407), .B1(
        n11404), .B2(n11387), .ZN(n3432) );
  AOI22_X1 U15113 ( .A1(\DataPath/RF/bus_reg_dataout[78] ), .A2(n11405), .B1(
        n11404), .B2(n11388), .ZN(n3431) );
  AOI22_X1 U15114 ( .A1(\DataPath/RF/bus_reg_dataout[79] ), .A2(n8407), .B1(
        n11404), .B2(n11389), .ZN(n3430) );
  AOI22_X1 U15115 ( .A1(\DataPath/RF/bus_reg_dataout[80] ), .A2(n8407), .B1(
        n11404), .B2(n11390), .ZN(n3429) );
  AOI22_X1 U15116 ( .A1(\DataPath/RF/bus_reg_dataout[81] ), .A2(n8407), .B1(
        n11404), .B2(n11410), .ZN(n3428) );
  AOI22_X1 U15117 ( .A1(\DataPath/RF/bus_reg_dataout[82] ), .A2(n11405), .B1(
        n11404), .B2(n11391), .ZN(n3427) );
  AOI22_X1 U15118 ( .A1(\DataPath/RF/bus_reg_dataout[83] ), .A2(n8407), .B1(
        n11404), .B2(n11392), .ZN(n3426) );
  INV_X1 U15119 ( .A(n11405), .ZN(n11393) );
  AOI22_X1 U15120 ( .A1(n11405), .A2(\DataPath/RF/bus_reg_dataout[84] ), .B1(
        n11441), .B2(n11393), .ZN(n3425) );
  AOI22_X1 U15121 ( .A1(\DataPath/RF/bus_reg_dataout[85] ), .A2(n8407), .B1(
        n11404), .B2(n11394), .ZN(n3424) );
  AOI22_X1 U15122 ( .A1(\DataPath/RF/bus_reg_dataout[86] ), .A2(n8407), .B1(
        n11404), .B2(n11395), .ZN(n3423) );
  AOI22_X1 U15123 ( .A1(\DataPath/RF/bus_reg_dataout[87] ), .A2(n8407), .B1(
        n11404), .B2(n11396), .ZN(n3422) );
  AOI22_X1 U15124 ( .A1(\DataPath/RF/bus_reg_dataout[88] ), .A2(n11405), .B1(
        n11404), .B2(n11397), .ZN(n3421) );
  AOI22_X1 U15125 ( .A1(\DataPath/RF/bus_reg_dataout[89] ), .A2(n8407), .B1(
        n11404), .B2(n11398), .ZN(n3420) );
  AOI22_X1 U15126 ( .A1(\DataPath/RF/bus_reg_dataout[90] ), .A2(n8407), .B1(
        n11404), .B2(n11399), .ZN(n3419) );
  AOI22_X1 U15127 ( .A1(\DataPath/RF/bus_reg_dataout[91] ), .A2(n11405), .B1(
        n11404), .B2(n11400), .ZN(n3418) );
  AOI22_X1 U15128 ( .A1(\DataPath/RF/bus_reg_dataout[92] ), .A2(n8407), .B1(
        n11404), .B2(n11401), .ZN(n3417) );
  AOI22_X1 U15129 ( .A1(\DataPath/RF/bus_reg_dataout[93] ), .A2(n8407), .B1(
        n11404), .B2(n11402), .ZN(n3416) );
  AOI22_X1 U15130 ( .A1(\DataPath/RF/bus_reg_dataout[94] ), .A2(n8407), .B1(
        n11404), .B2(n11411), .ZN(n3415) );
  AOI22_X1 U15131 ( .A1(\DataPath/RF/bus_reg_dataout[95] ), .A2(n8407), .B1(
        n11404), .B2(n11403), .ZN(n3412) );
  OAI22_X1 U15132 ( .A1(n8450), .A2(n11407), .B1(n11415), .B2(n11406), .ZN(
        n11408) );
  AOI22_X1 U15133 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[32] ), .B1(
        n11420), .B2(n8409), .ZN(n3407) );
  AOI22_X1 U15134 ( .A1(\DataPath/RF/bus_reg_dataout[33] ), .A2(n8408), .B1(
        n11412), .B2(n11421), .ZN(n3406) );
  AOI22_X1 U15135 ( .A1(\DataPath/RF/bus_reg_dataout[34] ), .A2(n8408), .B1(
        n11412), .B2(n11422), .ZN(n3405) );
  AOI22_X1 U15136 ( .A1(\DataPath/RF/bus_reg_dataout[35] ), .A2(n8408), .B1(
        n11412), .B2(n11423), .ZN(n3404) );
  AOI22_X1 U15137 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[36] ), .B1(
        n11424), .B2(n8409), .ZN(n3403) );
  AOI22_X1 U15138 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[37] ), .B1(
        n11425), .B2(n8409), .ZN(n3402) );
  AOI22_X1 U15139 ( .A1(\DataPath/RF/bus_reg_dataout[38] ), .A2(n8408), .B1(
        n11412), .B2(n11426), .ZN(n3401) );
  AOI22_X1 U15140 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[39] ), .B1(
        n11428), .B2(n8409), .ZN(n3400) );
  AOI22_X1 U15141 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[40] ), .B1(
        n11429), .B2(n8409), .ZN(n3399) );
  AOI22_X1 U15142 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[41] ), .B1(
        n11430), .B2(n8409), .ZN(n3398) );
  AOI22_X1 U15143 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[42] ), .B1(
        n11431), .B2(n8409), .ZN(n3397) );
  AOI22_X1 U15144 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[43] ), .B1(
        n11432), .B2(n8409), .ZN(n3396) );
  AOI22_X1 U15145 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[44] ), .B1(
        n11433), .B2(n8409), .ZN(n3395) );
  AOI22_X1 U15146 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[45] ), .B1(
        n11434), .B2(n8409), .ZN(n3394) );
  AOI22_X1 U15147 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[46] ), .B1(
        n11435), .B2(n8409), .ZN(n3393) );
  AOI22_X1 U15148 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[47] ), .B1(
        n11436), .B2(n8409), .ZN(n3392) );
  AOI22_X1 U15149 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[48] ), .B1(
        n11437), .B2(n8409), .ZN(n3391) );
  AOI22_X1 U15150 ( .A1(\DataPath/RF/bus_reg_dataout[49] ), .A2(n8408), .B1(
        n11412), .B2(n11410), .ZN(n3390) );
  AOI22_X1 U15151 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[50] ), .B1(
        n11439), .B2(n8409), .ZN(n3389) );
  AOI22_X1 U15152 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[51] ), .B1(
        n11440), .B2(n8409), .ZN(n3388) );
  AOI22_X1 U15153 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[52] ), .B1(
        n11441), .B2(n8409), .ZN(n3387) );
  AOI22_X1 U15154 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[53] ), .B1(
        n11442), .B2(n8409), .ZN(n3386) );
  AOI22_X1 U15155 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[54] ), .B1(
        n11443), .B2(n8409), .ZN(n3385) );
  AOI22_X1 U15156 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[55] ), .B1(
        n11444), .B2(n8409), .ZN(n3384) );
  AOI22_X1 U15157 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[56] ), .B1(
        n11445), .B2(n8409), .ZN(n3383) );
  AOI22_X1 U15158 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[57] ), .B1(
        n11446), .B2(n8409), .ZN(n3382) );
  AOI22_X1 U15159 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[58] ), .B1(
        n11447), .B2(n8409), .ZN(n3381) );
  AOI22_X1 U15160 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[59] ), .B1(
        n11448), .B2(n8409), .ZN(n3380) );
  AOI22_X1 U15161 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[60] ), .B1(
        n11449), .B2(n8409), .ZN(n3379) );
  AOI22_X1 U15162 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[61] ), .B1(
        n11450), .B2(n8409), .ZN(n3378) );
  AOI22_X1 U15163 ( .A1(\DataPath/RF/bus_reg_dataout[62] ), .A2(n8408), .B1(
        n11412), .B2(n11411), .ZN(n3377) );
  AOI22_X1 U15164 ( .A1(n8408), .A2(\DataPath/RF/bus_reg_dataout[63] ), .B1(
        n11597), .B2(n8409), .ZN(n3374) );
  OAI22_X1 U15165 ( .A1(n8450), .A2(n11416), .B1(n11415), .B2(n11414), .ZN(
        n11417) );
  AOI22_X1 U15166 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[0] ), .B1(
        n11420), .B2(n8420), .ZN(n3367) );
  NOR2_X1 U15167 ( .A1(RST), .A2(n8419), .ZN(n11427) );
  AOI22_X1 U15168 ( .A1(\DataPath/RF/bus_reg_dataout[1] ), .A2(n8418), .B1(
        n11427), .B2(n11421), .ZN(n3365) );
  AOI22_X1 U15169 ( .A1(\DataPath/RF/bus_reg_dataout[2] ), .A2(n8418), .B1(
        n11427), .B2(n11422), .ZN(n3363) );
  AOI22_X1 U15170 ( .A1(\DataPath/RF/bus_reg_dataout[3] ), .A2(n8418), .B1(
        n11427), .B2(n11423), .ZN(n3361) );
  AOI22_X1 U15171 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[4] ), .B1(
        n11424), .B2(n8420), .ZN(n3359) );
  AOI22_X1 U15172 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[5] ), .B1(
        n11425), .B2(n8420), .ZN(n3357) );
  AOI22_X1 U15173 ( .A1(\DataPath/RF/bus_reg_dataout[6] ), .A2(n8418), .B1(
        n11427), .B2(n11426), .ZN(n3355) );
  AOI22_X1 U15174 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[7] ), .B1(
        n11428), .B2(n8420), .ZN(n3353) );
  AOI22_X1 U15175 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[8] ), .B1(
        n11429), .B2(n8420), .ZN(n3351) );
  AOI22_X1 U15176 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[9] ), .B1(
        n11430), .B2(n8420), .ZN(n3349) );
  AOI22_X1 U15177 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[10] ), .B1(
        n11431), .B2(n8420), .ZN(n3347) );
  AOI22_X1 U15178 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[11] ), .B1(
        n11432), .B2(n8420), .ZN(n3345) );
  AOI22_X1 U15179 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[12] ), .B1(
        n11433), .B2(n8420), .ZN(n3343) );
  AOI22_X1 U15180 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[13] ), .B1(
        n11434), .B2(n8420), .ZN(n3341) );
  AOI22_X1 U15181 ( .A1(n8419), .A2(\DataPath/RF/bus_reg_dataout[14] ), .B1(
        n11435), .B2(n8420), .ZN(n3339) );
  AOI22_X1 U15182 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[15] ), .B1(
        n11436), .B2(n8420), .ZN(n3337) );
  AOI22_X1 U15183 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[16] ), .B1(
        n11437), .B2(n8420), .ZN(n3335) );
  AOI22_X1 U15184 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[17] ), .B1(
        n11438), .B2(n8420), .ZN(n3333) );
  AOI22_X1 U15185 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[18] ), .B1(
        n11439), .B2(n8420), .ZN(n3331) );
  AOI22_X1 U15186 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[19] ), .B1(
        n11440), .B2(n8420), .ZN(n3329) );
  AOI22_X1 U15187 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[20] ), .B1(
        n11441), .B2(n8420), .ZN(n3327) );
  AOI22_X1 U15188 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[21] ), .B1(
        n11442), .B2(n8420), .ZN(n3325) );
  AOI22_X1 U15189 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[22] ), .B1(
        n11443), .B2(n8420), .ZN(n3323) );
  AOI22_X1 U15190 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[23] ), .B1(
        n11444), .B2(n8420), .ZN(n3321) );
  AOI22_X1 U15191 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[24] ), .B1(
        n11445), .B2(n8420), .ZN(n3319) );
  AOI22_X1 U15192 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[25] ), .B1(
        n11446), .B2(n8420), .ZN(n3317) );
  AOI22_X1 U15193 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[26] ), .B1(
        n11447), .B2(n8420), .ZN(n3315) );
  AOI22_X1 U15194 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[27] ), .B1(
        n11448), .B2(n8420), .ZN(n3313) );
  AOI22_X1 U15195 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[28] ), .B1(
        n11449), .B2(n8420), .ZN(n3311) );
  AOI22_X1 U15196 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[29] ), .B1(
        n11450), .B2(n8420), .ZN(n3309) );
  AOI22_X1 U15197 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[30] ), .B1(
        n11451), .B2(n8420), .ZN(n3307) );
  NAND2_X1 U15198 ( .A1(n11452), .A2(n11476), .ZN(n11453) );
  OAI22_X1 U15199 ( .A1(n11479), .A2(n11455), .B1(n802), .B2(n11454), .ZN(
        n6984) );
  OAI22_X1 U15200 ( .A1(n11480), .A2(n11455), .B1(n803), .B2(n11454), .ZN(
        n6983) );
  OAI22_X1 U15201 ( .A1(n11481), .A2(n11455), .B1(n804), .B2(n11454), .ZN(
        n6982) );
  OAI22_X1 U15202 ( .A1(n11482), .A2(n11455), .B1(n805), .B2(n11454), .ZN(
        n6981) );
  OAI22_X1 U15203 ( .A1(n11483), .A2(n11455), .B1(n806), .B2(n11454), .ZN(
        n6980) );
  OAI22_X1 U15204 ( .A1(n11484), .A2(n11455), .B1(n807), .B2(n11454), .ZN(
        n6979) );
  OAI22_X1 U15205 ( .A1(n11485), .A2(n11455), .B1(n808), .B2(n11454), .ZN(
        n6978) );
  OAI22_X1 U15206 ( .A1(n11486), .A2(n11455), .B1(n809), .B2(n11454), .ZN(
        n6977) );
  OAI22_X1 U15207 ( .A1(n11487), .A2(n11455), .B1(n810), .B2(n11454), .ZN(
        n6976) );
  OAI22_X1 U15208 ( .A1(n11488), .A2(n11455), .B1(n811), .B2(n11454), .ZN(
        n6975) );
  OAI22_X1 U15209 ( .A1(n11489), .A2(n8411), .B1(n812), .B2(n11454), .ZN(n6974) );
  OAI22_X1 U15210 ( .A1(n11490), .A2(n8411), .B1(n813), .B2(n11454), .ZN(n6973) );
  OAI22_X1 U15211 ( .A1(n11491), .A2(n8411), .B1(n814), .B2(n11454), .ZN(n6972) );
  OAI22_X1 U15212 ( .A1(n11492), .A2(n8411), .B1(n815), .B2(n11454), .ZN(n6971) );
  OAI22_X1 U15213 ( .A1(n11493), .A2(n8411), .B1(n816), .B2(n11454), .ZN(n6970) );
  OAI22_X1 U15214 ( .A1(n11494), .A2(n8411), .B1(n817), .B2(n11454), .ZN(n6969) );
  OAI22_X1 U15215 ( .A1(n11495), .A2(n8411), .B1(n818), .B2(n11454), .ZN(n6968) );
  OAI22_X1 U15216 ( .A1(n11496), .A2(n8411), .B1(n819), .B2(n11454), .ZN(n6967) );
  OAI22_X1 U15217 ( .A1(n11497), .A2(n8411), .B1(n820), .B2(n11454), .ZN(n6966) );
  OAI22_X1 U15218 ( .A1(n11498), .A2(n8411), .B1(n821), .B2(n11454), .ZN(n6965) );
  OAI22_X1 U15219 ( .A1(n11499), .A2(n8411), .B1(n822), .B2(n11454), .ZN(n6964) );
  OAI22_X1 U15220 ( .A1(n11500), .A2(n8411), .B1(n823), .B2(n11454), .ZN(n6963) );
  OAI22_X1 U15221 ( .A1(n11501), .A2(n11455), .B1(n824), .B2(n11454), .ZN(
        n6962) );
  OAI22_X1 U15222 ( .A1(n11502), .A2(n11455), .B1(n825), .B2(n11454), .ZN(
        n6961) );
  OAI22_X1 U15223 ( .A1(n11503), .A2(n11455), .B1(n826), .B2(n11454), .ZN(
        n6960) );
  OAI22_X1 U15224 ( .A1(n11504), .A2(n11455), .B1(n827), .B2(n11454), .ZN(
        n6959) );
  OAI22_X1 U15225 ( .A1(n11505), .A2(n8411), .B1(n828), .B2(n11454), .ZN(n6958) );
  OAI22_X1 U15226 ( .A1(n11506), .A2(n11455), .B1(n829), .B2(n11454), .ZN(
        n6957) );
  OAI22_X1 U15227 ( .A1(n11507), .A2(n8411), .B1(n830), .B2(n11454), .ZN(n6956) );
  OAI22_X1 U15228 ( .A1(n11508), .A2(n8411), .B1(n831), .B2(n11454), .ZN(n6955) );
  OAI22_X1 U15229 ( .A1(n11509), .A2(n8411), .B1(n832), .B2(n11454), .ZN(n6954) );
  OAI22_X1 U15230 ( .A1(n11512), .A2(n8411), .B1(n833), .B2(n11454), .ZN(n6953) );
  AOI21_X1 U15231 ( .B1(n11456), .B2(n11476), .A(RST), .ZN(n11457) );
  OAI22_X1 U15232 ( .A1(n11479), .A2(n11459), .B1(n770), .B2(n11458), .ZN(
        n6952) );
  OAI22_X1 U15233 ( .A1(n11480), .A2(n11459), .B1(n771), .B2(n11458), .ZN(
        n6951) );
  OAI22_X1 U15234 ( .A1(n11481), .A2(n11459), .B1(n772), .B2(n11458), .ZN(
        n6950) );
  OAI22_X1 U15235 ( .A1(n11482), .A2(n11459), .B1(n773), .B2(n11458), .ZN(
        n6949) );
  OAI22_X1 U15236 ( .A1(n11483), .A2(n11459), .B1(n774), .B2(n11458), .ZN(
        n6948) );
  OAI22_X1 U15237 ( .A1(n11484), .A2(n11459), .B1(n775), .B2(n11458), .ZN(
        n6947) );
  OAI22_X1 U15238 ( .A1(n11485), .A2(n11459), .B1(n776), .B2(n11458), .ZN(
        n6946) );
  OAI22_X1 U15239 ( .A1(n11486), .A2(n11459), .B1(n777), .B2(n11458), .ZN(
        n6945) );
  OAI22_X1 U15240 ( .A1(n11487), .A2(n11459), .B1(n778), .B2(n11458), .ZN(
        n6944) );
  OAI22_X1 U15241 ( .A1(n11488), .A2(n11459), .B1(n779), .B2(n11458), .ZN(
        n6943) );
  OAI22_X1 U15242 ( .A1(n11489), .A2(n8412), .B1(n780), .B2(n11458), .ZN(n6942) );
  OAI22_X1 U15243 ( .A1(n11490), .A2(n8412), .B1(n781), .B2(n11458), .ZN(n6941) );
  OAI22_X1 U15244 ( .A1(n11491), .A2(n8412), .B1(n782), .B2(n11458), .ZN(n6940) );
  OAI22_X1 U15245 ( .A1(n11492), .A2(n8412), .B1(n783), .B2(n11458), .ZN(n6939) );
  OAI22_X1 U15246 ( .A1(n11493), .A2(n8412), .B1(n784), .B2(n11458), .ZN(n6938) );
  OAI22_X1 U15247 ( .A1(n11494), .A2(n8412), .B1(n785), .B2(n11458), .ZN(n6937) );
  OAI22_X1 U15248 ( .A1(n11495), .A2(n8412), .B1(n786), .B2(n11458), .ZN(n6936) );
  OAI22_X1 U15249 ( .A1(n11496), .A2(n8412), .B1(n787), .B2(n11458), .ZN(n6935) );
  OAI22_X1 U15250 ( .A1(n11497), .A2(n8412), .B1(n788), .B2(n11458), .ZN(n6934) );
  OAI22_X1 U15251 ( .A1(n11498), .A2(n8412), .B1(n789), .B2(n11458), .ZN(n6933) );
  OAI22_X1 U15252 ( .A1(n11499), .A2(n8412), .B1(n790), .B2(n11458), .ZN(n6932) );
  OAI22_X1 U15253 ( .A1(n11500), .A2(n8412), .B1(n791), .B2(n11458), .ZN(n6931) );
  OAI22_X1 U15254 ( .A1(n11501), .A2(n11459), .B1(n792), .B2(n11458), .ZN(
        n6930) );
  OAI22_X1 U15255 ( .A1(n11502), .A2(n11459), .B1(n793), .B2(n11458), .ZN(
        n6929) );
  OAI22_X1 U15256 ( .A1(n11503), .A2(n11459), .B1(n794), .B2(n11458), .ZN(
        n6928) );
  OAI22_X1 U15257 ( .A1(n11504), .A2(n11459), .B1(n795), .B2(n11458), .ZN(
        n6927) );
  OAI22_X1 U15258 ( .A1(n11505), .A2(n8412), .B1(n796), .B2(n11458), .ZN(n6926) );
  OAI22_X1 U15259 ( .A1(n11506), .A2(n11459), .B1(n797), .B2(n11458), .ZN(
        n6925) );
  OAI22_X1 U15260 ( .A1(n11507), .A2(n8412), .B1(n798), .B2(n11458), .ZN(n6924) );
  OAI22_X1 U15261 ( .A1(n11508), .A2(n8412), .B1(n799), .B2(n11458), .ZN(n6923) );
  OAI22_X1 U15262 ( .A1(n11509), .A2(n8412), .B1(n800), .B2(n11458), .ZN(n6922) );
  OAI22_X1 U15263 ( .A1(n11512), .A2(n8412), .B1(n801), .B2(n11458), .ZN(n6921) );
  AOI21_X1 U15264 ( .B1(n11460), .B2(n11476), .A(RST), .ZN(n11461) );
  OAI22_X1 U15265 ( .A1(n11479), .A2(n11463), .B1(n738), .B2(n11462), .ZN(
        n6920) );
  OAI22_X1 U15266 ( .A1(n11480), .A2(n11463), .B1(n739), .B2(n11462), .ZN(
        n6919) );
  OAI22_X1 U15267 ( .A1(n11481), .A2(n11463), .B1(n740), .B2(n11462), .ZN(
        n6918) );
  OAI22_X1 U15268 ( .A1(n11482), .A2(n11463), .B1(n741), .B2(n11462), .ZN(
        n6917) );
  OAI22_X1 U15269 ( .A1(n11483), .A2(n11463), .B1(n742), .B2(n11462), .ZN(
        n6916) );
  OAI22_X1 U15270 ( .A1(n11484), .A2(n11463), .B1(n743), .B2(n11462), .ZN(
        n6915) );
  OAI22_X1 U15271 ( .A1(n11485), .A2(n11463), .B1(n744), .B2(n11462), .ZN(
        n6914) );
  OAI22_X1 U15272 ( .A1(n11486), .A2(n11463), .B1(n745), .B2(n11462), .ZN(
        n6913) );
  OAI22_X1 U15273 ( .A1(n11487), .A2(n11463), .B1(n746), .B2(n11462), .ZN(
        n6912) );
  OAI22_X1 U15274 ( .A1(n11488), .A2(n11463), .B1(n747), .B2(n11462), .ZN(
        n6911) );
  OAI22_X1 U15275 ( .A1(n11489), .A2(n11463), .B1(n748), .B2(n11462), .ZN(
        n6910) );
  OAI22_X1 U15276 ( .A1(n11490), .A2(n8413), .B1(n749), .B2(n11462), .ZN(n6909) );
  OAI22_X1 U15277 ( .A1(n11491), .A2(n8413), .B1(n750), .B2(n11462), .ZN(n6908) );
  OAI22_X1 U15278 ( .A1(n11492), .A2(n8413), .B1(n751), .B2(n11462), .ZN(n6907) );
  OAI22_X1 U15279 ( .A1(n11493), .A2(n8413), .B1(n752), .B2(n11462), .ZN(n6906) );
  OAI22_X1 U15280 ( .A1(n11494), .A2(n8413), .B1(n753), .B2(n11462), .ZN(n6905) );
  OAI22_X1 U15281 ( .A1(n11495), .A2(n8413), .B1(n754), .B2(n11462), .ZN(n6904) );
  OAI22_X1 U15282 ( .A1(n11496), .A2(n8413), .B1(n755), .B2(n11462), .ZN(n6903) );
  OAI22_X1 U15283 ( .A1(n11497), .A2(n8413), .B1(n756), .B2(n11462), .ZN(n6902) );
  OAI22_X1 U15284 ( .A1(n11498), .A2(n8413), .B1(n757), .B2(n11462), .ZN(n6901) );
  OAI22_X1 U15285 ( .A1(n11499), .A2(n8413), .B1(n758), .B2(n11462), .ZN(n6900) );
  OAI22_X1 U15286 ( .A1(n11500), .A2(n8413), .B1(n759), .B2(n11462), .ZN(n6899) );
  OAI22_X1 U15287 ( .A1(n11501), .A2(n11463), .B1(n760), .B2(n11462), .ZN(
        n6898) );
  OAI22_X1 U15288 ( .A1(n11502), .A2(n11463), .B1(n761), .B2(n11462), .ZN(
        n6897) );
  OAI22_X1 U15289 ( .A1(n11503), .A2(n11463), .B1(n762), .B2(n11462), .ZN(
        n6896) );
  OAI22_X1 U15290 ( .A1(n11504), .A2(n11463), .B1(n763), .B2(n11462), .ZN(
        n6895) );
  OAI22_X1 U15291 ( .A1(n11505), .A2(n8413), .B1(n764), .B2(n11462), .ZN(n6894) );
  OAI22_X1 U15292 ( .A1(n11506), .A2(n11463), .B1(n765), .B2(n11462), .ZN(
        n6893) );
  OAI22_X1 U15293 ( .A1(n11507), .A2(n8413), .B1(n766), .B2(n11462), .ZN(n6892) );
  OAI22_X1 U15294 ( .A1(n11508), .A2(n8413), .B1(n767), .B2(n11462), .ZN(n6891) );
  OAI22_X1 U15295 ( .A1(n11509), .A2(n8413), .B1(n768), .B2(n11462), .ZN(n6890) );
  OAI22_X1 U15296 ( .A1(n11512), .A2(n8413), .B1(n769), .B2(n11462), .ZN(n6889) );
  AOI21_X1 U15297 ( .B1(n11464), .B2(n11476), .A(RST), .ZN(n11465) );
  OAI22_X1 U15298 ( .A1(n11479), .A2(n11467), .B1(n706), .B2(n11466), .ZN(
        n6888) );
  OAI22_X1 U15299 ( .A1(n11480), .A2(n11467), .B1(n707), .B2(n11466), .ZN(
        n6887) );
  OAI22_X1 U15300 ( .A1(n11481), .A2(n11467), .B1(n708), .B2(n11466), .ZN(
        n6886) );
  OAI22_X1 U15301 ( .A1(n11482), .A2(n11467), .B1(n709), .B2(n11466), .ZN(
        n6885) );
  OAI22_X1 U15302 ( .A1(n11483), .A2(n11467), .B1(n710), .B2(n11466), .ZN(
        n6884) );
  OAI22_X1 U15303 ( .A1(n11484), .A2(n11467), .B1(n711), .B2(n11466), .ZN(
        n6883) );
  OAI22_X1 U15304 ( .A1(n11485), .A2(n11467), .B1(n712), .B2(n11466), .ZN(
        n6882) );
  OAI22_X1 U15305 ( .A1(n11486), .A2(n11467), .B1(n713), .B2(n11466), .ZN(
        n6881) );
  OAI22_X1 U15306 ( .A1(n11487), .A2(n11467), .B1(n714), .B2(n11466), .ZN(
        n6880) );
  OAI22_X1 U15307 ( .A1(n11488), .A2(n11467), .B1(n715), .B2(n11466), .ZN(
        n6879) );
  OAI22_X1 U15308 ( .A1(n11489), .A2(n11467), .B1(n716), .B2(n11466), .ZN(
        n6878) );
  OAI22_X1 U15309 ( .A1(n11490), .A2(n8414), .B1(n717), .B2(n11466), .ZN(n6877) );
  OAI22_X1 U15310 ( .A1(n11491), .A2(n8414), .B1(n718), .B2(n11466), .ZN(n6876) );
  OAI22_X1 U15311 ( .A1(n11492), .A2(n8414), .B1(n719), .B2(n11466), .ZN(n6875) );
  OAI22_X1 U15312 ( .A1(n11493), .A2(n8414), .B1(n720), .B2(n11466), .ZN(n6874) );
  OAI22_X1 U15313 ( .A1(n11494), .A2(n8414), .B1(n721), .B2(n11466), .ZN(n6873) );
  OAI22_X1 U15314 ( .A1(n11495), .A2(n8414), .B1(n722), .B2(n11466), .ZN(n6872) );
  OAI22_X1 U15315 ( .A1(n11496), .A2(n8414), .B1(n723), .B2(n11466), .ZN(n6871) );
  OAI22_X1 U15316 ( .A1(n11497), .A2(n8414), .B1(n724), .B2(n11466), .ZN(n6870) );
  OAI22_X1 U15317 ( .A1(n11498), .A2(n8414), .B1(n725), .B2(n11466), .ZN(n6869) );
  OAI22_X1 U15318 ( .A1(n11499), .A2(n8414), .B1(n726), .B2(n11466), .ZN(n6868) );
  OAI22_X1 U15319 ( .A1(n11500), .A2(n8414), .B1(n727), .B2(n11466), .ZN(n6867) );
  OAI22_X1 U15320 ( .A1(n11501), .A2(n11467), .B1(n728), .B2(n11466), .ZN(
        n6866) );
  OAI22_X1 U15321 ( .A1(n11502), .A2(n11467), .B1(n729), .B2(n11466), .ZN(
        n6865) );
  OAI22_X1 U15322 ( .A1(n11503), .A2(n11467), .B1(n730), .B2(n11466), .ZN(
        n6864) );
  OAI22_X1 U15323 ( .A1(n11504), .A2(n11467), .B1(n731), .B2(n11466), .ZN(
        n6863) );
  OAI22_X1 U15324 ( .A1(n11505), .A2(n8414), .B1(n732), .B2(n11466), .ZN(n6862) );
  OAI22_X1 U15325 ( .A1(n11506), .A2(n11467), .B1(n733), .B2(n11466), .ZN(
        n6861) );
  OAI22_X1 U15326 ( .A1(n11507), .A2(n8414), .B1(n734), .B2(n11466), .ZN(n6860) );
  OAI22_X1 U15327 ( .A1(n11508), .A2(n8414), .B1(n735), .B2(n11466), .ZN(n6859) );
  OAI22_X1 U15328 ( .A1(n11509), .A2(n8414), .B1(n736), .B2(n11466), .ZN(n6858) );
  OAI22_X1 U15329 ( .A1(n11512), .A2(n8414), .B1(n737), .B2(n11466), .ZN(n6857) );
  AOI21_X1 U15330 ( .B1(n11468), .B2(n11476), .A(RST), .ZN(n11469) );
  OAI22_X1 U15331 ( .A1(n11479), .A2(n11471), .B1(n674), .B2(n11470), .ZN(
        n6856) );
  OAI22_X1 U15332 ( .A1(n11480), .A2(n11471), .B1(n675), .B2(n11470), .ZN(
        n6855) );
  OAI22_X1 U15333 ( .A1(n11481), .A2(n11471), .B1(n676), .B2(n11470), .ZN(
        n6854) );
  OAI22_X1 U15334 ( .A1(n11482), .A2(n11471), .B1(n677), .B2(n11470), .ZN(
        n6853) );
  OAI22_X1 U15335 ( .A1(n11483), .A2(n11471), .B1(n678), .B2(n11470), .ZN(
        n6852) );
  OAI22_X1 U15336 ( .A1(n11484), .A2(n11471), .B1(n679), .B2(n11470), .ZN(
        n6851) );
  OAI22_X1 U15337 ( .A1(n11485), .A2(n11471), .B1(n680), .B2(n11470), .ZN(
        n6850) );
  OAI22_X1 U15338 ( .A1(n11486), .A2(n11471), .B1(n681), .B2(n11470), .ZN(
        n6849) );
  OAI22_X1 U15339 ( .A1(n11487), .A2(n11471), .B1(n682), .B2(n11470), .ZN(
        n6848) );
  OAI22_X1 U15340 ( .A1(n11488), .A2(n11471), .B1(n683), .B2(n11470), .ZN(
        n6847) );
  OAI22_X1 U15341 ( .A1(n11489), .A2(n8415), .B1(n684), .B2(n11470), .ZN(n6846) );
  OAI22_X1 U15342 ( .A1(n11490), .A2(n8415), .B1(n685), .B2(n11470), .ZN(n6845) );
  OAI22_X1 U15343 ( .A1(n11491), .A2(n8415), .B1(n686), .B2(n11470), .ZN(n6844) );
  OAI22_X1 U15344 ( .A1(n11492), .A2(n8415), .B1(n687), .B2(n11470), .ZN(n6843) );
  OAI22_X1 U15345 ( .A1(n11493), .A2(n8415), .B1(n688), .B2(n11470), .ZN(n6842) );
  OAI22_X1 U15346 ( .A1(n11494), .A2(n8415), .B1(n689), .B2(n11470), .ZN(n6841) );
  OAI22_X1 U15347 ( .A1(n11495), .A2(n8415), .B1(n690), .B2(n11470), .ZN(n6840) );
  OAI22_X1 U15348 ( .A1(n11496), .A2(n8415), .B1(n691), .B2(n11470), .ZN(n6839) );
  OAI22_X1 U15349 ( .A1(n11497), .A2(n8415), .B1(n692), .B2(n11470), .ZN(n6838) );
  OAI22_X1 U15350 ( .A1(n11498), .A2(n8415), .B1(n693), .B2(n11470), .ZN(n6837) );
  OAI22_X1 U15351 ( .A1(n11499), .A2(n8415), .B1(n694), .B2(n11470), .ZN(n6836) );
  OAI22_X1 U15352 ( .A1(n11500), .A2(n8415), .B1(n695), .B2(n11470), .ZN(n6835) );
  OAI22_X1 U15353 ( .A1(n11501), .A2(n11471), .B1(n696), .B2(n11470), .ZN(
        n6834) );
  OAI22_X1 U15354 ( .A1(n11502), .A2(n11471), .B1(n697), .B2(n11470), .ZN(
        n6833) );
  OAI22_X1 U15355 ( .A1(n11503), .A2(n11471), .B1(n698), .B2(n11470), .ZN(
        n6832) );
  OAI22_X1 U15356 ( .A1(n11504), .A2(n11471), .B1(n699), .B2(n11470), .ZN(
        n6831) );
  OAI22_X1 U15357 ( .A1(n11505), .A2(n8415), .B1(n700), .B2(n11470), .ZN(n6830) );
  OAI22_X1 U15358 ( .A1(n11506), .A2(n11471), .B1(n701), .B2(n11470), .ZN(
        n6829) );
  OAI22_X1 U15359 ( .A1(n11507), .A2(n8415), .B1(n702), .B2(n11470), .ZN(n6828) );
  OAI22_X1 U15360 ( .A1(n11508), .A2(n8415), .B1(n703), .B2(n11470), .ZN(n6827) );
  OAI22_X1 U15361 ( .A1(n11509), .A2(n8415), .B1(n704), .B2(n11470), .ZN(n6826) );
  OAI22_X1 U15362 ( .A1(n11512), .A2(n8415), .B1(n705), .B2(n11470), .ZN(n6825) );
  NAND2_X1 U15363 ( .A1(n11472), .A2(n11476), .ZN(n11473) );
  OAI22_X1 U15364 ( .A1(n11479), .A2(n11475), .B1(n642), .B2(n11474), .ZN(
        n6824) );
  OAI22_X1 U15365 ( .A1(n11480), .A2(n11475), .B1(n643), .B2(n11474), .ZN(
        n6823) );
  OAI22_X1 U15366 ( .A1(n11481), .A2(n11475), .B1(n644), .B2(n11474), .ZN(
        n6822) );
  OAI22_X1 U15367 ( .A1(n11482), .A2(n11475), .B1(n645), .B2(n11474), .ZN(
        n6821) );
  OAI22_X1 U15368 ( .A1(n11483), .A2(n11475), .B1(n646), .B2(n11474), .ZN(
        n6820) );
  OAI22_X1 U15369 ( .A1(n11484), .A2(n11475), .B1(n647), .B2(n11474), .ZN(
        n6819) );
  OAI22_X1 U15370 ( .A1(n11485), .A2(n11475), .B1(n648), .B2(n11474), .ZN(
        n6818) );
  OAI22_X1 U15371 ( .A1(n11486), .A2(n11475), .B1(n649), .B2(n11474), .ZN(
        n6817) );
  OAI22_X1 U15372 ( .A1(n11487), .A2(n11475), .B1(n650), .B2(n11474), .ZN(
        n6816) );
  OAI22_X1 U15373 ( .A1(n11488), .A2(n11475), .B1(n651), .B2(n11474), .ZN(
        n6815) );
  OAI22_X1 U15374 ( .A1(n11489), .A2(n8416), .B1(n652), .B2(n11474), .ZN(n6814) );
  OAI22_X1 U15375 ( .A1(n11490), .A2(n8416), .B1(n653), .B2(n11474), .ZN(n6813) );
  OAI22_X1 U15376 ( .A1(n11491), .A2(n8416), .B1(n654), .B2(n11474), .ZN(n6812) );
  OAI22_X1 U15377 ( .A1(n11492), .A2(n8416), .B1(n655), .B2(n11474), .ZN(n6811) );
  OAI22_X1 U15378 ( .A1(n11493), .A2(n8416), .B1(n656), .B2(n11474), .ZN(n6810) );
  OAI22_X1 U15379 ( .A1(n11494), .A2(n8416), .B1(n657), .B2(n11474), .ZN(n6809) );
  OAI22_X1 U15380 ( .A1(n11495), .A2(n8416), .B1(n658), .B2(n11474), .ZN(n6808) );
  OAI22_X1 U15381 ( .A1(n11496), .A2(n8416), .B1(n659), .B2(n11474), .ZN(n6807) );
  OAI22_X1 U15382 ( .A1(n11497), .A2(n8416), .B1(n660), .B2(n11474), .ZN(n6806) );
  OAI22_X1 U15383 ( .A1(n11498), .A2(n8416), .B1(n661), .B2(n11474), .ZN(n6805) );
  OAI22_X1 U15384 ( .A1(n11499), .A2(n8416), .B1(n662), .B2(n11474), .ZN(n6804) );
  OAI22_X1 U15385 ( .A1(n11500), .A2(n8416), .B1(n663), .B2(n11474), .ZN(n6803) );
  OAI22_X1 U15386 ( .A1(n11501), .A2(n11475), .B1(n664), .B2(n11474), .ZN(
        n6802) );
  OAI22_X1 U15387 ( .A1(n11502), .A2(n11475), .B1(n665), .B2(n11474), .ZN(
        n6801) );
  OAI22_X1 U15388 ( .A1(n11503), .A2(n11475), .B1(n666), .B2(n11474), .ZN(
        n6800) );
  OAI22_X1 U15389 ( .A1(n11504), .A2(n11475), .B1(n667), .B2(n11474), .ZN(
        n6799) );
  OAI22_X1 U15390 ( .A1(n11505), .A2(n8416), .B1(n668), .B2(n11474), .ZN(n6798) );
  OAI22_X1 U15391 ( .A1(n11506), .A2(n11475), .B1(n669), .B2(n11474), .ZN(
        n6797) );
  OAI22_X1 U15392 ( .A1(n11507), .A2(n8416), .B1(n670), .B2(n11474), .ZN(n6796) );
  OAI22_X1 U15393 ( .A1(n11508), .A2(n8416), .B1(n671), .B2(n11474), .ZN(n6795) );
  OAI22_X1 U15394 ( .A1(n11509), .A2(n8416), .B1(n672), .B2(n11474), .ZN(n6794) );
  OAI22_X1 U15395 ( .A1(n11512), .A2(n8416), .B1(n673), .B2(n11474), .ZN(n6793) );
  NAND2_X1 U15396 ( .A1(n11477), .A2(n11476), .ZN(n11478) );
  OAI22_X1 U15397 ( .A1(n11479), .A2(n11511), .B1(n610), .B2(n11510), .ZN(
        n6792) );
  OAI22_X1 U15398 ( .A1(n11480), .A2(n11511), .B1(n611), .B2(n11510), .ZN(
        n6791) );
  OAI22_X1 U15399 ( .A1(n11481), .A2(n11511), .B1(n612), .B2(n11510), .ZN(
        n6790) );
  OAI22_X1 U15400 ( .A1(n11482), .A2(n11511), .B1(n613), .B2(n11510), .ZN(
        n6789) );
  OAI22_X1 U15401 ( .A1(n11483), .A2(n11511), .B1(n614), .B2(n11510), .ZN(
        n6788) );
  OAI22_X1 U15402 ( .A1(n11484), .A2(n11511), .B1(n615), .B2(n11510), .ZN(
        n6787) );
  OAI22_X1 U15403 ( .A1(n11485), .A2(n11511), .B1(n616), .B2(n11510), .ZN(
        n6786) );
  OAI22_X1 U15404 ( .A1(n11486), .A2(n11511), .B1(n617), .B2(n11510), .ZN(
        n6785) );
  OAI22_X1 U15405 ( .A1(n11487), .A2(n11511), .B1(n618), .B2(n11510), .ZN(
        n6784) );
  OAI22_X1 U15406 ( .A1(n11488), .A2(n11511), .B1(n619), .B2(n11510), .ZN(
        n6783) );
  OAI22_X1 U15407 ( .A1(n11489), .A2(n11511), .B1(n620), .B2(n11510), .ZN(
        n6782) );
  OAI22_X1 U15408 ( .A1(n11490), .A2(n8417), .B1(n621), .B2(n11510), .ZN(n6781) );
  OAI22_X1 U15409 ( .A1(n11491), .A2(n8417), .B1(n622), .B2(n11510), .ZN(n6780) );
  OAI22_X1 U15410 ( .A1(n11492), .A2(n8417), .B1(n623), .B2(n11510), .ZN(n6779) );
  OAI22_X1 U15411 ( .A1(n11493), .A2(n8417), .B1(n624), .B2(n11510), .ZN(n6778) );
  OAI22_X1 U15412 ( .A1(n11494), .A2(n8417), .B1(n625), .B2(n11510), .ZN(n6777) );
  OAI22_X1 U15413 ( .A1(n11495), .A2(n8417), .B1(n626), .B2(n11510), .ZN(n6776) );
  OAI22_X1 U15414 ( .A1(n11496), .A2(n8417), .B1(n627), .B2(n11510), .ZN(n6775) );
  OAI22_X1 U15415 ( .A1(n11497), .A2(n8417), .B1(n628), .B2(n11510), .ZN(n6774) );
  OAI22_X1 U15416 ( .A1(n11498), .A2(n8417), .B1(n629), .B2(n11510), .ZN(n6773) );
  OAI22_X1 U15417 ( .A1(n11499), .A2(n8417), .B1(n630), .B2(n11510), .ZN(n6772) );
  OAI22_X1 U15418 ( .A1(n11500), .A2(n8417), .B1(n631), .B2(n11510), .ZN(n6771) );
  OAI22_X1 U15419 ( .A1(n11501), .A2(n11511), .B1(n632), .B2(n11510), .ZN(
        n6770) );
  OAI22_X1 U15420 ( .A1(n11502), .A2(n11511), .B1(n633), .B2(n11510), .ZN(
        n6769) );
  OAI22_X1 U15421 ( .A1(n11503), .A2(n11511), .B1(n634), .B2(n11510), .ZN(
        n6768) );
  OAI22_X1 U15422 ( .A1(n11504), .A2(n11511), .B1(n635), .B2(n11510), .ZN(
        n6767) );
  OAI22_X1 U15423 ( .A1(n11505), .A2(n8417), .B1(n636), .B2(n11510), .ZN(n6766) );
  OAI22_X1 U15424 ( .A1(n11506), .A2(n11511), .B1(n637), .B2(n11510), .ZN(
        n6765) );
  OAI22_X1 U15425 ( .A1(n11507), .A2(n8417), .B1(n638), .B2(n11510), .ZN(n6764) );
  OAI22_X1 U15426 ( .A1(n11508), .A2(n8417), .B1(n639), .B2(n11510), .ZN(n6763) );
  OAI22_X1 U15427 ( .A1(n11509), .A2(n8417), .B1(n640), .B2(n11510), .ZN(n6762) );
  OAI22_X1 U15428 ( .A1(n11512), .A2(n8417), .B1(n641), .B2(n11510), .ZN(n6761) );
  AOI22_X1 U15429 ( .A1(i_RD1[0]), .A2(n8423), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_A[0] ), .ZN(n3256) );
  AOI22_X1 U15430 ( .A1(i_RD1[1]), .A2(n7753), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[1] ), .ZN(n11514) );
  INV_X1 U15431 ( .A(n11514), .ZN(n6728) );
  AOI22_X1 U15432 ( .A1(i_RD1[2]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_A[2] ), .ZN(n3255) );
  AOI22_X1 U15433 ( .A1(i_RD1[3]), .A2(n8424), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_A[3] ), .ZN(n11515) );
  INV_X1 U15434 ( .A(n11515), .ZN(n6727) );
  AOI22_X1 U15435 ( .A1(i_RD1[4]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[4] ), .ZN(n3254) );
  AOI22_X1 U15436 ( .A1(i_RD1[5]), .A2(n8424), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_A[5] ), .ZN(n3253) );
  AOI22_X1 U15437 ( .A1(i_RD1[6]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[6] ), .ZN(n3252) );
  AOI22_X1 U15438 ( .A1(i_RD1[7]), .A2(n8424), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_A[7] ), .ZN(n3251) );
  AOI22_X1 U15439 ( .A1(i_RD1[8]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[8] ), .ZN(n11516) );
  INV_X1 U15440 ( .A(n11516), .ZN(n6726) );
  AOI22_X1 U15441 ( .A1(i_RD1[9]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[9] ), .ZN(n3250) );
  AOI22_X1 U15442 ( .A1(i_RD1[10]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[10] ), .ZN(n3249) );
  AOI22_X1 U15443 ( .A1(i_RD1[11]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[11] ), .ZN(n3248) );
  AOI22_X1 U15444 ( .A1(i_RD1[12]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[12] ), .ZN(n3247) );
  AOI22_X1 U15445 ( .A1(i_RD1[13]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[13] ), .ZN(n11517) );
  INV_X1 U15446 ( .A(n11517), .ZN(n6725) );
  AOI22_X1 U15447 ( .A1(i_RD1[14]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[14] ), .ZN(n11518) );
  INV_X1 U15448 ( .A(n11518), .ZN(n6724) );
  AOI22_X1 U15449 ( .A1(i_RD1[15]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[15] ), .ZN(n3246) );
  AOI22_X1 U15450 ( .A1(i_RD1[16]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[16] ), .ZN(n3245) );
  AOI22_X1 U15451 ( .A1(i_RD1[17]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[17] ), .ZN(n3244) );
  AOI22_X1 U15452 ( .A1(i_RD1[18]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[18] ), .ZN(n3243) );
  AOI22_X1 U15453 ( .A1(i_RD1[19]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[19] ), .ZN(n3242) );
  AOI22_X1 U15454 ( .A1(i_RD1[20]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[20] ), .ZN(n11519) );
  INV_X1 U15455 ( .A(n11519), .ZN(n6723) );
  AOI22_X1 U15456 ( .A1(i_RD1[21]), .A2(n8424), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[21] ), .ZN(n3241) );
  AOI22_X1 U15457 ( .A1(i_RD1[22]), .A2(n8423), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[22] ), .ZN(n3240) );
  AOI22_X1 U15458 ( .A1(i_RD1[23]), .A2(n8423), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[23] ), .ZN(n3239) );
  AOI22_X1 U15459 ( .A1(i_RD1[24]), .A2(n8423), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[24] ), .ZN(n3238) );
  AOI22_X1 U15460 ( .A1(i_RD1[25]), .A2(n8423), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[25] ), .ZN(n3237) );
  AOI22_X1 U15461 ( .A1(i_RD1[26]), .A2(n8423), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[26] ), .ZN(n3236) );
  AOI22_X1 U15462 ( .A1(i_RD1[27]), .A2(n8423), .B1(n8427), .B2(
        \DataPath/i_PIPLIN_A[27] ), .ZN(n3235) );
  AOI22_X1 U15463 ( .A1(i_RD1[28]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_A[28] ), .ZN(n3234) );
  AOI22_X1 U15464 ( .A1(i_RD1[29]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_A[29] ), .ZN(n3233) );
  AOI22_X1 U15465 ( .A1(i_RD1[30]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_A[30] ), .ZN(n3232) );
  AOI22_X1 U15466 ( .A1(i_RD1[31]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_A[31] ), .ZN(n3231) );
  NAND2_X1 U15467 ( .A1(n8460), .A2(n11520), .ZN(n3230) );
  NAND2_X1 U15468 ( .A1(n8459), .A2(n11521), .ZN(n3229) );
  NAND2_X1 U15469 ( .A1(n8460), .A2(n11522), .ZN(n3228) );
  NAND2_X1 U15470 ( .A1(n8460), .A2(n11523), .ZN(n3227) );
  NAND2_X1 U15471 ( .A1(n8459), .A2(n11524), .ZN(n3226) );
  NAND2_X1 U15472 ( .A1(n8459), .A2(n11525), .ZN(n3225) );
  NAND2_X1 U15473 ( .A1(n8459), .A2(n11526), .ZN(n3224) );
  NAND2_X1 U15474 ( .A1(n8459), .A2(n11527), .ZN(n3223) );
  NAND2_X1 U15475 ( .A1(n8460), .A2(n11528), .ZN(n3222) );
  NAND2_X1 U15476 ( .A1(n8459), .A2(n11529), .ZN(n3221) );
  NAND2_X1 U15477 ( .A1(n8459), .A2(n11530), .ZN(n3220) );
  NAND2_X1 U15478 ( .A1(n8459), .A2(n11531), .ZN(n3219) );
  NAND2_X1 U15479 ( .A1(n8459), .A2(n11532), .ZN(n3218) );
  NAND2_X1 U15480 ( .A1(n8459), .A2(n11533), .ZN(n3217) );
  NAND2_X1 U15481 ( .A1(n8457), .A2(n11534), .ZN(n3216) );
  NAND2_X1 U15482 ( .A1(n8458), .A2(n11535), .ZN(n3215) );
  NAND2_X1 U15483 ( .A1(n8458), .A2(n11536), .ZN(n3214) );
  NAND2_X1 U15484 ( .A1(n8458), .A2(n11537), .ZN(n3213) );
  NAND2_X1 U15485 ( .A1(n8460), .A2(n11538), .ZN(n3212) );
  NAND2_X1 U15486 ( .A1(n8458), .A2(n11539), .ZN(n3211) );
  NAND2_X1 U15487 ( .A1(n8458), .A2(n11540), .ZN(n3210) );
  NAND2_X1 U15488 ( .A1(n8458), .A2(n11541), .ZN(n3209) );
  NAND2_X1 U15489 ( .A1(n8458), .A2(n11542), .ZN(n3208) );
  NAND2_X1 U15490 ( .A1(n8459), .A2(n11543), .ZN(n3207) );
  NAND2_X1 U15491 ( .A1(n8458), .A2(n11544), .ZN(n3206) );
  NAND2_X1 U15492 ( .A1(n8458), .A2(n11545), .ZN(n3205) );
  NAND2_X1 U15493 ( .A1(n8458), .A2(n11546), .ZN(n3204) );
  NAND2_X1 U15494 ( .A1(n8458), .A2(n11547), .ZN(n3203) );
  NAND2_X1 U15495 ( .A1(n8459), .A2(n11548), .ZN(n3202) );
  NAND2_X1 U15496 ( .A1(n8457), .A2(n11549), .ZN(n3201) );
  NAND2_X1 U15497 ( .A1(n8458), .A2(n11550), .ZN(n3200) );
  NAND2_X1 U15498 ( .A1(n8457), .A2(n11551), .ZN(n3197) );
  NOR2_X1 U15499 ( .A1(n555), .A2(n556), .ZN(n11553) );
  NAND2_X1 U15500 ( .A1(\DECODEhw/i_tickcounter[2] ), .A2(n11553), .ZN(n11555)
         );
  NAND2_X1 U15501 ( .A1(\DECODEhw/i_tickcounter[4] ), .A2(n11556), .ZN(n11558)
         );
  NAND2_X1 U15502 ( .A1(\DECODEhw/i_tickcounter[6] ), .A2(n11559), .ZN(n11561)
         );
  NAND2_X1 U15503 ( .A1(\DECODEhw/i_tickcounter[8] ), .A2(n11562), .ZN(n11564)
         );
  NAND2_X1 U15504 ( .A1(\DECODEhw/i_tickcounter[10] ), .A2(n11565), .ZN(n11567) );
  NAND2_X1 U15505 ( .A1(\DECODEhw/i_tickcounter[12] ), .A2(n11568), .ZN(n11570) );
  NAND2_X1 U15506 ( .A1(\DECODEhw/i_tickcounter[14] ), .A2(n11571), .ZN(n11573) );
  NAND2_X1 U15507 ( .A1(\DECODEhw/i_tickcounter[16] ), .A2(n11574), .ZN(n11576) );
  NAND2_X1 U15508 ( .A1(\DECODEhw/i_tickcounter[18] ), .A2(n11577), .ZN(n11579) );
  NAND2_X1 U15509 ( .A1(\DECODEhw/i_tickcounter[20] ), .A2(n11580), .ZN(n11582) );
  NAND2_X1 U15510 ( .A1(\DECODEhw/i_tickcounter[22] ), .A2(n11583), .ZN(n11585) );
  NAND2_X1 U15511 ( .A1(\DECODEhw/i_tickcounter[24] ), .A2(n11586), .ZN(n11588) );
  NOR2_X1 U15512 ( .A1(n580), .A2(n11588), .ZN(n11589) );
  NAND2_X1 U15513 ( .A1(\DECODEhw/i_tickcounter[26] ), .A2(n11589), .ZN(n11592) );
  NOR2_X1 U15514 ( .A1(n582), .A2(n11592), .ZN(n11591) );
  INV_X1 U15515 ( .A(n11591), .ZN(n11593) );
  NOR2_X1 U15516 ( .A1(n583), .A2(n11593), .ZN(n11594) );
  NAND2_X1 U15517 ( .A1(\DECODEhw/i_tickcounter[29] ), .A2(n11594), .ZN(n11596) );
  NOR2_X1 U15518 ( .A1(n584), .A2(n11596), .ZN(n11595) );
  OAI21_X1 U15519 ( .B1(\DECODEhw/i_tickcounter[31] ), .B2(n11595), .A(n8458), 
        .ZN(n11552) );
  AOI21_X1 U15520 ( .B1(\DECODEhw/i_tickcounter[31] ), .B2(n11595), .A(n11552), 
        .ZN(n7170) );
  AND2_X1 U15521 ( .A1(n8462), .A2(n555), .ZN(n7169) );
  AOI211_X1 U15522 ( .C1(n556), .C2(n555), .A(RST), .B(n11553), .ZN(n7168) );
  OAI211_X1 U15523 ( .C1(\DECODEhw/i_tickcounter[2] ), .C2(n11553), .A(n11555), 
        .B(n8461), .ZN(n11554) );
  AOI211_X1 U15524 ( .C1(n558), .C2(n11555), .A(RST), .B(n11556), .ZN(n7166)
         );
  OAI211_X1 U15525 ( .C1(\DECODEhw/i_tickcounter[4] ), .C2(n11556), .A(n11558), 
        .B(n8458), .ZN(n11557) );
  AOI211_X1 U15526 ( .C1(n560), .C2(n11558), .A(RST), .B(n11559), .ZN(n7164)
         );
  OAI211_X1 U15527 ( .C1(\DECODEhw/i_tickcounter[6] ), .C2(n11559), .A(n11561), 
        .B(n8463), .ZN(n11560) );
  INV_X1 U15528 ( .A(n11560), .ZN(n7163) );
  AOI211_X1 U15529 ( .C1(n562), .C2(n11561), .A(RST), .B(n11562), .ZN(n7162)
         );
  OAI211_X1 U15530 ( .C1(\DECODEhw/i_tickcounter[8] ), .C2(n11562), .A(n11564), 
        .B(n8466), .ZN(n11563) );
  INV_X1 U15531 ( .A(n11563), .ZN(n7161) );
  AOI211_X1 U15532 ( .C1(n564), .C2(n11564), .A(RST), .B(n11565), .ZN(n7160)
         );
  OAI211_X1 U15533 ( .C1(\DECODEhw/i_tickcounter[10] ), .C2(n11565), .A(n11567), .B(n8457), .ZN(n11566) );
  INV_X1 U15534 ( .A(n11566), .ZN(n7159) );
  AOI211_X1 U15535 ( .C1(n566), .C2(n11567), .A(RST), .B(n11568), .ZN(n7158)
         );
  OAI211_X1 U15536 ( .C1(\DECODEhw/i_tickcounter[12] ), .C2(n11568), .A(n11570), .B(n8463), .ZN(n11569) );
  INV_X1 U15537 ( .A(n11569), .ZN(n7157) );
  AOI211_X1 U15538 ( .C1(n568), .C2(n11570), .A(RST), .B(n11571), .ZN(n7156)
         );
  OAI211_X1 U15539 ( .C1(\DECODEhw/i_tickcounter[14] ), .C2(n11571), .A(n11573), .B(n8462), .ZN(n11572) );
  INV_X1 U15540 ( .A(n11572), .ZN(n7155) );
  AOI211_X1 U15541 ( .C1(n570), .C2(n11573), .A(RST), .B(n11574), .ZN(n7154)
         );
  OAI211_X1 U15542 ( .C1(\DECODEhw/i_tickcounter[16] ), .C2(n11574), .A(n11576), .B(n8457), .ZN(n11575) );
  INV_X1 U15543 ( .A(n11575), .ZN(n7153) );
  AOI211_X1 U15544 ( .C1(n572), .C2(n11576), .A(RST), .B(n11577), .ZN(n7152)
         );
  OAI211_X1 U15545 ( .C1(\DECODEhw/i_tickcounter[18] ), .C2(n11577), .A(n11579), .B(n8467), .ZN(n11578) );
  INV_X1 U15546 ( .A(n11578), .ZN(n7151) );
  AOI211_X1 U15547 ( .C1(n574), .C2(n11579), .A(RST), .B(n11580), .ZN(n7150)
         );
  OAI211_X1 U15548 ( .C1(\DECODEhw/i_tickcounter[20] ), .C2(n11580), .A(n11582), .B(n8468), .ZN(n11581) );
  INV_X1 U15549 ( .A(n11581), .ZN(n7149) );
  AOI211_X1 U15550 ( .C1(n576), .C2(n11582), .A(RST), .B(n11583), .ZN(n7148)
         );
  OAI211_X1 U15551 ( .C1(\DECODEhw/i_tickcounter[22] ), .C2(n11583), .A(n11585), .B(n8463), .ZN(n11584) );
  INV_X1 U15552 ( .A(n11584), .ZN(n7147) );
  AOI211_X1 U15553 ( .C1(n578), .C2(n11585), .A(RST), .B(n11586), .ZN(n7146)
         );
  OAI211_X1 U15554 ( .C1(\DECODEhw/i_tickcounter[24] ), .C2(n11586), .A(n11588), .B(n8467), .ZN(n11587) );
  INV_X1 U15555 ( .A(n11587), .ZN(n7145) );
  AOI211_X1 U15556 ( .C1(n580), .C2(n11588), .A(RST), .B(n11589), .ZN(n7144)
         );
  OAI211_X1 U15557 ( .C1(\DECODEhw/i_tickcounter[26] ), .C2(n11589), .A(n11592), .B(n8464), .ZN(n11590) );
  INV_X1 U15558 ( .A(n11590), .ZN(n7143) );
  AOI211_X1 U15559 ( .C1(n582), .C2(n11592), .A(RST), .B(n11591), .ZN(n7142)
         );
  AOI211_X1 U15560 ( .C1(n583), .C2(n11593), .A(RST), .B(n11594), .ZN(n7141)
         );
  OAI211_X1 U15561 ( .C1(\DECODEhw/i_tickcounter[29] ), .C2(n11594), .A(n11596), .B(n8466), .ZN(n3153) );
  AOI211_X1 U15562 ( .C1(n584), .C2(n11596), .A(RST), .B(n11595), .ZN(n7140)
         );
  AOI22_X1 U15563 ( .A1(n8418), .A2(\DataPath/RF/bus_reg_dataout[31] ), .B1(
        n11597), .B2(n8420), .ZN(n3147) );
  OR2_X1 U15564 ( .A1(IR[9]), .A2(IR[10]), .ZN(n11599) );
  NOR4_X1 U15565 ( .A1(IR[8]), .A2(IR[7]), .A3(IR[6]), .A4(n11599), .ZN(n11617) );
  NAND3_X1 U15566 ( .A1(IR[5]), .A2(IR[3]), .A3(n11617), .ZN(n11618) );
  AOI21_X1 U15567 ( .B1(IR[2]), .B2(IR[1]), .A(n11618), .ZN(n11623) );
  OAI21_X1 U15568 ( .B1(n8101), .B2(n8294), .A(n11600), .ZN(n7139) );
  OAI21_X1 U15569 ( .B1(n8294), .B2(n184), .A(n11601), .ZN(n7138) );
  OAI21_X1 U15570 ( .B1(n8294), .B2(n183), .A(n11602), .ZN(n7137) );
  OAI21_X1 U15571 ( .B1(n8294), .B2(n182), .A(n11603), .ZN(n7136) );
  OAI21_X1 U15572 ( .B1(n8294), .B2(n181), .A(n11604), .ZN(n7135) );
  OAI21_X1 U15573 ( .B1(n8294), .B2(n180), .A(n11605), .ZN(n7134) );
  OAI21_X1 U15574 ( .B1(n8294), .B2(n179), .A(n11606), .ZN(n7133) );
  OAI21_X1 U15575 ( .B1(n8294), .B2(n178), .A(n11607), .ZN(n7132) );
  OAI21_X1 U15576 ( .B1(n8294), .B2(n177), .A(n11608), .ZN(n7131) );
  OAI21_X1 U15577 ( .B1(n8294), .B2(n176), .A(n11609), .ZN(n7130) );
  OAI21_X1 U15578 ( .B1(n8294), .B2(n175), .A(n11610), .ZN(n7129) );
  OAI21_X1 U15579 ( .B1(n8294), .B2(n174), .A(n11611), .ZN(n7128) );
  OAI21_X1 U15580 ( .B1(n8294), .B2(n173), .A(n11612), .ZN(n7127) );
  INV_X1 U15581 ( .A(IRAM_DATA[26]), .ZN(n11613) );
  INV_X1 U15582 ( .A(IRAM_DATA[28]), .ZN(n11614) );
  INV_X1 U15583 ( .A(IRAM_DATA[30]), .ZN(n11615) );
  OAI22_X1 U15584 ( .A1(DRAM_READNOTWRITE), .A2(n11828), .B1(n11830), .B2(
        n8203), .ZN(n7121) );
  AOI22_X1 U15585 ( .A1(n10300), .A2(\CU_I/CW_ID[WB_EN] ), .B1(n11626), .B2(
        \CU_I/CW_EX[WB_EN] ), .ZN(n2853) );
  AOI22_X1 U15586 ( .A1(n10300), .A2(\CU_I/CW_ID[WB_MUX_SEL] ), .B1(n11626), 
        .B2(\CU_I/CW_EX[WB_MUX_SEL] ), .ZN(n2852) );
  AOI22_X1 U15587 ( .A1(n10300), .A2(\CU_I/CW_EX[WB_EN] ), .B1(n11626), .B2(
        \CU_I/CW_MEM[WB_EN] ), .ZN(n2847) );
  AOI22_X1 U15588 ( .A1(n10300), .A2(\CU_I/CW_EX[WB_MUX_SEL] ), .B1(n11626), 
        .B2(\CU_I/CW_MEM[WB_MUX_SEL] ), .ZN(n2846) );
  AOI21_X1 U15589 ( .B1(n8246), .B2(n8199), .A(RST), .ZN(n7094) );
  OAI22_X1 U15590 ( .A1(n380), .A2(n11828), .B1(n11830), .B2(n8202), .ZN(n7093) );
  OAI22_X1 U15591 ( .A1(n381), .A2(n11828), .B1(n11830), .B2(n8201), .ZN(n7092) );
  OAI22_X1 U15592 ( .A1(n11616), .A2(n11828), .B1(n11830), .B2(n8200), .ZN(
        n7091) );
  NOR2_X1 U15593 ( .A1(IR[2]), .A2(IR[1]), .ZN(n11622) );
  OAI222_X1 U15594 ( .A1(n11621), .A2(n11620), .B1(n11828), .B2(n223), .C1(
        n11619), .C2(n172), .ZN(n7083) );
  INV_X1 U15595 ( .A(\CU_I/CW_ID[MUXB_SEL] ), .ZN(n11624) );
  NAND2_X1 U15596 ( .A1(n10300), .A2(\CU_I/CW_ID[MUXA_SEL] ), .ZN(n11625) );
  OAI21_X1 U15597 ( .B1(n11828), .B2(n7732), .A(n11625), .ZN(n7080) );
  AOI22_X1 U15598 ( .A1(n10300), .A2(\CU_I/CW_ID[EX_EN] ), .B1(
        \CU_I/CW_EX[EX_EN] ), .B2(n11626), .ZN(n2780) );
  AOI22_X1 U15599 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_WRB1[0] ), .B1(n7764), 
        .B2(\DataPath/i_PIPLIN_WRB2[0] ), .ZN(n2779) );
  AOI22_X1 U15600 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_WRB1[1] ), .B1(n7764), 
        .B2(\DataPath/i_PIPLIN_WRB2[1] ), .ZN(n2778) );
  AOI22_X1 U15601 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_WRB1[2] ), .B1(n7764), 
        .B2(\DataPath/i_PIPLIN_WRB2[2] ), .ZN(n2777) );
  AOI22_X1 U15602 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_WRB1[3] ), .B1(n7764), 
        .B2(\DataPath/i_PIPLIN_WRB2[3] ), .ZN(n2776) );
  AOI22_X1 U15603 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_WRB1[4] ), .B1(n7764), 
        .B2(\DataPath/i_PIPLIN_WRB2[4] ), .ZN(n2775) );
  OAI22_X1 U15604 ( .A1(n218), .A2(n11828), .B1(n10298), .B2(n11830), .ZN(
        n7079) );
  OAI22_X1 U15605 ( .A1(n217), .A2(n11828), .B1(n218), .B2(n11830), .ZN(n7078)
         );
  AOI22_X1 U15606 ( .A1(i_RD2[0]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[0] ), .ZN(n11627) );
  INV_X1 U15607 ( .A(n11627), .ZN(n7077) );
  AOI22_X1 U15608 ( .A1(i_RD2[1]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[1] ), .ZN(n2767) );
  AOI22_X1 U15609 ( .A1(i_RD2[2]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[2] ), .ZN(n2766) );
  AOI22_X1 U15610 ( .A1(i_RD2[3]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[3] ), .ZN(n11628) );
  INV_X1 U15611 ( .A(n11628), .ZN(n7076) );
  AOI22_X1 U15612 ( .A1(i_RD2[5]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[5] ), .ZN(n2765) );
  OAI22_X1 U15613 ( .A1(n481), .A2(n11838), .B1(n11629), .B2(n11839), .ZN(
        n7074) );
  AOI22_X1 U15614 ( .A1(i_RD2[7]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[7] ), .ZN(n2764) );
  AOI22_X1 U15615 ( .A1(i_RD2[8]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[8] ), .ZN(n11630) );
  INV_X1 U15616 ( .A(n11630), .ZN(n7073) );
  AOI22_X1 U15617 ( .A1(i_RD2[9]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[9] ), .ZN(n2763) );
  AOI22_X1 U15618 ( .A1(i_RD2[10]), .A2(n8422), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[10] ), .ZN(n2762) );
  AOI22_X1 U15619 ( .A1(i_RD2[11]), .A2(n8422), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[11] ), .ZN(n2761) );
  AOI22_X1 U15620 ( .A1(i_RD2[12]), .A2(n8422), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[12] ), .ZN(n2760) );
  AOI22_X1 U15621 ( .A1(i_RD2[13]), .A2(n8422), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[13] ), .ZN(n11631) );
  INV_X1 U15622 ( .A(n11631), .ZN(n7072) );
  AOI22_X1 U15623 ( .A1(i_RD2[14]), .A2(n8422), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[14] ), .ZN(n11632) );
  INV_X1 U15624 ( .A(n11632), .ZN(n7071) );
  AOI22_X1 U15625 ( .A1(i_RD2[15]), .A2(n8422), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[15] ), .ZN(n2759) );
  AOI22_X1 U15626 ( .A1(i_RD2[16]), .A2(n8422), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[16] ), .ZN(n2758) );
  AOI22_X1 U15627 ( .A1(i_RD2[17]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[17] ), .ZN(n2757) );
  AOI22_X1 U15628 ( .A1(i_RD2[18]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[18] ), .ZN(n2756) );
  AOI22_X1 U15629 ( .A1(i_RD2[19]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[19] ), .ZN(n2755) );
  AOI22_X1 U15630 ( .A1(i_RD2[20]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[20] ), .ZN(n2754) );
  AOI22_X1 U15631 ( .A1(i_RD2[21]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[21] ), .ZN(n2753) );
  AOI22_X1 U15632 ( .A1(i_RD2[22]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[22] ), .ZN(n2752) );
  AOI22_X1 U15633 ( .A1(i_RD2[23]), .A2(n8422), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_B[23] ), .ZN(n2751) );
  AOI22_X1 U15634 ( .A1(i_RD2[24]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[24] ), .ZN(n2750) );
  AOI22_X1 U15635 ( .A1(i_RD2[25]), .A2(n8422), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_B[25] ), .ZN(n2749) );
  AOI22_X1 U15636 ( .A1(i_RD2[26]), .A2(n8422), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_B[26] ), .ZN(n2748) );
  AOI22_X1 U15637 ( .A1(i_RD2[27]), .A2(n8422), .B1(n11679), .B2(
        \DataPath/i_PIPLIN_B[27] ), .ZN(n2747) );
  AOI22_X1 U15638 ( .A1(i_RD2[28]), .A2(n8422), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_B[28] ), .ZN(n2746) );
  AOI22_X1 U15639 ( .A1(i_RD2[29]), .A2(n8424), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_B[29] ), .ZN(n2745) );
  AOI22_X1 U15640 ( .A1(i_RD2[30]), .A2(n7753), .B1(n8425), .B2(
        \DataPath/i_PIPLIN_B[30] ), .ZN(n2744) );
  AOI22_X1 U15641 ( .A1(i_RD2[31]), .A2(n8423), .B1(n8426), .B2(
        \DataPath/i_PIPLIN_B[31] ), .ZN(n2743) );
  AOI22_X1 U15642 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[0] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[0] ), .ZN(n2742) );
  AOI22_X1 U15643 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[1] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[1] ), .ZN(n2741) );
  AOI22_X1 U15644 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[2] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[2] ), .ZN(n2740) );
  AOI22_X1 U15645 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[3] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[3] ), .ZN(n2739) );
  AOI22_X1 U15646 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[4] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[4] ), .ZN(n2738) );
  AOI22_X1 U15647 ( .A1(n10290), .A2(\DataPath/i_PIPLIN_B[5] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[5] ), .ZN(n2737) );
  OAI22_X1 U15648 ( .A1(n481), .A2(n11694), .B1(n11734), .B2(n8223), .ZN(n7070) );
  AOI22_X1 U15649 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[7] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[7] ), .ZN(n2736) );
  AOI22_X1 U15650 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[8] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[8] ), .ZN(n2735) );
  AOI22_X1 U15651 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[9] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[9] ), .ZN(n2734) );
  AOI22_X1 U15652 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[10] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[10] ), .ZN(n2733) );
  AOI22_X1 U15653 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[11] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[11] ), .ZN(n2732) );
  AOI22_X1 U15654 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[12] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[12] ), .ZN(n2731) );
  AOI22_X1 U15655 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[13] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[13] ), .ZN(n2730) );
  AOI22_X1 U15656 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[14] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[14] ), .ZN(n2729) );
  AOI22_X1 U15657 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[15] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[15] ), .ZN(n2728) );
  AOI22_X1 U15658 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[16] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[16] ), .ZN(n2727) );
  AOI22_X1 U15659 ( .A1(n10290), .A2(\DataPath/i_PIPLIN_B[17] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[17] ), .ZN(n2726) );
  AOI22_X1 U15660 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[18] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[18] ), .ZN(n2725) );
  AOI22_X1 U15661 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[19] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[19] ), .ZN(n2724) );
  AOI22_X1 U15662 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[20] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[20] ), .ZN(n2723) );
  AOI22_X1 U15663 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[21] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[21] ), .ZN(n2722) );
  AOI22_X1 U15664 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[22] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[22] ), .ZN(n2721) );
  AOI22_X1 U15665 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[23] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[23] ), .ZN(n2720) );
  AOI22_X1 U15666 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[24] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[24] ), .ZN(n2719) );
  AOI22_X1 U15667 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[25] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[25] ), .ZN(n2718) );
  AOI22_X1 U15668 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[26] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[26] ), .ZN(n2717) );
  AOI22_X1 U15669 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[27] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[27] ), .ZN(n2716) );
  AOI22_X1 U15670 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[28] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[28] ), .ZN(n2715) );
  AOI22_X1 U15671 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[29] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[29] ), .ZN(n2714) );
  AOI22_X1 U15672 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[30] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[30] ), .ZN(n2713) );
  AOI22_X1 U15673 ( .A1(n7769), .A2(\DataPath/i_PIPLIN_B[31] ), .B1(n7764), 
        .B2(\DataPath/i_REG_ME_DATA_DATAMEM[31] ), .ZN(n2712) );
  INV_X1 U15674 ( .A(n11633), .ZN(n11635) );
  OAI21_X1 U15675 ( .B1(n11635), .B2(n11634), .A(n11649), .ZN(n11636) );
  NAND2_X1 U15676 ( .A1(n11637), .A2(n11636), .ZN(n11639) );
  NOR2_X1 U15677 ( .A1(n11637), .A2(n11636), .ZN(n11645) );
  INV_X1 U15678 ( .A(n11639), .ZN(n11644) );
  NOR2_X1 U15679 ( .A1(n11645), .A2(n11644), .ZN(n11643) );
  AOI22_X1 U15680 ( .A1(n7648), .A2(n11645), .B1(\DataPath/RF/c_win[0] ), .B2(
        n11643), .ZN(n11638) );
  OAI211_X1 U15681 ( .C1(n11640), .C2(n11639), .A(n11638), .B(n8463), .ZN(
        n7069) );
  AOI222_X1 U15682 ( .A1(\DataPath/RF/c_win[2] ), .A2(n11644), .B1(n8275), 
        .B2(n11643), .C1(\DataPath/RF/c_win[0] ), .C2(n11645), .ZN(n11641) );
  NOR2_X1 U15683 ( .A1(RST), .A2(n11641), .ZN(n7068) );
  AOI222_X1 U15684 ( .A1(\DataPath/RF/c_win[2] ), .A2(n11645), .B1(n11644), 
        .B2(n7648), .C1(\DataPath/RF/c_win[3] ), .C2(n11643), .ZN(n11642) );
  NOR2_X1 U15685 ( .A1(RST), .A2(n11642), .ZN(n7066) );
  NOR2_X1 U15686 ( .A1(n11846), .A2(n11646), .ZN(n11648) );
  NAND2_X1 U15687 ( .A1(\DataPath/RF/PUSH_ADDRGEN/curr_state[0] ), .A2(n11647), 
        .ZN(n11847) );
  AOI21_X1 U15688 ( .B1(n11648), .B2(n11847), .A(RST), .ZN(n7064) );
  NOR2_X1 U15689 ( .A1(n11649), .A2(n11846), .ZN(n11656) );
  INV_X1 U15690 ( .A(n11656), .ZN(n11652) );
  NOR2_X1 U15691 ( .A1(n11650), .A2(n9270), .ZN(n11658) );
  NOR2_X1 U15692 ( .A1(n11658), .A2(n11656), .ZN(n11657) );
  AOI22_X1 U15693 ( .A1(\DataPath/RF/c_swin[0] ), .A2(n11657), .B1(n8281), 
        .B2(n11658), .ZN(n11651) );
  OAI211_X1 U15694 ( .C1(n835), .C2(n11652), .A(n11651), .B(n8460), .ZN(n7063)
         );
  AOI222_X1 U15695 ( .A1(\DataPath/RF/c_swin[1] ), .A2(n11657), .B1(n11658), 
        .B2(\DataPath/RF/c_swin[0] ), .C1(\DataPath/RF/c_swin[2] ), .C2(n11656), .ZN(n11653) );
  NOR2_X1 U15696 ( .A1(RST), .A2(n11653), .ZN(n7062) );
  AOI222_X1 U15697 ( .A1(\DataPath/RF/c_swin[3] ), .A2(n11656), .B1(
        \DataPath/RF/c_swin[1] ), .B2(n11658), .C1(\DataPath/RF/c_swin[2] ), 
        .C2(n11657), .ZN(n11654) );
  NOR2_X1 U15698 ( .A1(RST), .A2(n11654), .ZN(n7061) );
  NOR2_X1 U15699 ( .A1(RST), .A2(n11655), .ZN(n7060) );
  AOI222_X1 U15700 ( .A1(\DataPath/RF/c_swin[3] ), .A2(n11658), .B1(n8281), 
        .B2(n11657), .C1(\DataPath/RF/c_swin[0] ), .C2(n11656), .ZN(n11659) );
  NOR2_X1 U15701 ( .A1(RST), .A2(n11659), .ZN(n7059) );
  NAND2_X1 U15702 ( .A1(n11662), .A2(n11661), .ZN(n11663) );
  OAI21_X1 U15703 ( .B1(n11663), .B2(n11666), .A(n8459), .ZN(n11664) );
  AOI21_X1 U15704 ( .B1(n877), .B2(n11666), .A(n11664), .ZN(n7058) );
  AOI211_X1 U15705 ( .C1(n8207), .C2(n11666), .A(RST), .B(n11665), .ZN(n7057)
         );
  INV_X1 U15706 ( .A(i_RD1[1]), .ZN(n11668) );
  OAI21_X1 U15707 ( .B1(n11670), .B2(n11678), .A(n11669), .ZN(n7047) );
  INV_X1 U15708 ( .A(i_RD1[12]), .ZN(n11671) );
  AND2_X1 U15709 ( .A1(n11672), .A2(IRAM_ADDRESS[17]), .ZN(n11673) );
  OAI21_X1 U15710 ( .B1(n11678), .B2(n11675), .A(n11674), .ZN(n7038) );
  OAI21_X1 U15711 ( .B1(n11677), .B2(n11678), .A(n11676), .ZN(n7037) );
  NOR2_X1 U15712 ( .A1(n8095), .A2(n8085), .ZN(n11681) );
  INV_X1 U15713 ( .A(n11681), .ZN(n11716) );
  NOR2_X1 U15714 ( .A1(i_ALU_OP[2]), .A2(n11731), .ZN(n11680) );
  NOR2_X1 U15715 ( .A1(n8084), .A2(n8085), .ZN(n11682) );
  INV_X1 U15716 ( .A(n11682), .ZN(n11683) );
  NAND2_X1 U15717 ( .A1(n11716), .A2(n11683), .ZN(n11718) );
  NAND3_X1 U15718 ( .A1(n8084), .A2(n8095), .A3(i_ALU_OP[4]), .ZN(n11725) );
  INV_X1 U15719 ( .A(n11725), .ZN(n11720) );
  NOR2_X1 U15720 ( .A1(n8095), .A2(n11732), .ZN(n11685) );
  INV_X1 U15721 ( .A(n11680), .ZN(n11684) );
  NAND2_X1 U15722 ( .A1(n8084), .A2(n8085), .ZN(n11722) );
  OAI21_X1 U15723 ( .B1(n506), .B2(n223), .A(\DataPath/i_LGET[0] ), .ZN(n11686) );
  OAI21_X1 U15724 ( .B1(\DataPath/i_LGET[0] ), .B2(n222), .A(n11686), .ZN(
        n11689) );
  AOI22_X1 U15725 ( .A1(\i_SEL_LGET[1] ), .A2(n8106), .B1(n222), .B2(n8198), 
        .ZN(n11687) );
  OAI221_X1 U15726 ( .B1(\DataPath/i_LGET[0] ), .B2(n222), .C1(n8197), .C2(
        n11687), .A(n223), .ZN(n11688) );
  OAI211_X1 U15727 ( .C1(\i_SEL_LGET[1] ), .C2(n11689), .A(i_SEL_ALU_SETCMP), 
        .B(n11688), .ZN(n11690) );
  OAI211_X1 U15728 ( .C1(n11692), .C2(n11691), .A(n7769), .B(n11690), .ZN(
        n11693) );
  OAI21_X1 U15729 ( .B1(n507), .B2(n11734), .A(n11693), .ZN(n7013) );
  AOI22_X1 U15730 ( .A1(n11835), .A2(DRAM_DATA_OUT[0]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[0] ), .ZN(n2223) );
  AOI22_X1 U15731 ( .A1(n11835), .A2(DRAM_DATA_OUT[1]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[1] ), .ZN(n2222) );
  AOI22_X1 U15732 ( .A1(n11835), .A2(DRAM_DATA_OUT[2]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[2] ), .ZN(n2221) );
  AOI22_X1 U15733 ( .A1(n11835), .A2(DRAM_DATA_OUT[3]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[3] ), .ZN(n2220) );
  AOI22_X1 U15734 ( .A1(n11835), .A2(DRAM_DATA_OUT[4]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[4] ), .ZN(n2219) );
  AOI22_X1 U15735 ( .A1(n11835), .A2(DRAM_DATA_OUT[5]), .B1(n8441), .B2(
        \DataPath/i_REG_LDSTR_OUT[5] ), .ZN(n2218) );
  AOI22_X1 U15736 ( .A1(n11835), .A2(DRAM_DATA_OUT[6]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[6] ), .ZN(n2217) );
  AOI22_X1 U15737 ( .A1(n11835), .A2(DRAM_DATA_OUT[7]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[7] ), .ZN(n2216) );
  AOI22_X1 U15738 ( .A1(n11835), .A2(DRAM_DATA_OUT[8]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[8] ), .ZN(n2215) );
  AOI22_X1 U15739 ( .A1(n11835), .A2(DRAM_DATA_OUT[9]), .B1(n8441), .B2(
        \DataPath/i_REG_LDSTR_OUT[9] ), .ZN(n2214) );
  AOI22_X1 U15740 ( .A1(n11835), .A2(DRAM_DATA_OUT[10]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[10] ), .ZN(n2213) );
  AOI22_X1 U15741 ( .A1(n11835), .A2(DRAM_DATA_OUT[11]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[11] ), .ZN(n2212) );
  AOI22_X1 U15742 ( .A1(n11835), .A2(DRAM_DATA_OUT[12]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[12] ), .ZN(n2211) );
  AOI22_X1 U15743 ( .A1(n11835), .A2(DRAM_DATA_OUT[13]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[13] ), .ZN(n2210) );
  AOI22_X1 U15744 ( .A1(n11835), .A2(DRAM_DATA_OUT[14]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[14] ), .ZN(n2209) );
  AOI22_X1 U15745 ( .A1(n11835), .A2(DRAM_DATA_OUT[15]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[15] ), .ZN(n2208) );
  AOI22_X1 U15746 ( .A1(n11835), .A2(DRAM_DATA_OUT[16]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[16] ), .ZN(n2207) );
  AOI22_X1 U15747 ( .A1(n11835), .A2(DRAM_DATA_OUT[17]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[17] ), .ZN(n2206) );
  AOI22_X1 U15748 ( .A1(n11835), .A2(DRAM_DATA_OUT[18]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[18] ), .ZN(n2205) );
  AOI22_X1 U15749 ( .A1(n11835), .A2(DRAM_DATA_OUT[19]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[19] ), .ZN(n2204) );
  AOI22_X1 U15750 ( .A1(n11835), .A2(DRAM_DATA_OUT[20]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[20] ), .ZN(n2203) );
  AOI22_X1 U15751 ( .A1(n11835), .A2(DRAM_DATA_OUT[21]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[21] ), .ZN(n2202) );
  AOI22_X1 U15752 ( .A1(n11835), .A2(DRAM_DATA_OUT[22]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[22] ), .ZN(n2201) );
  AOI22_X1 U15753 ( .A1(n11835), .A2(DRAM_DATA_OUT[23]), .B1(n11836), .B2(
        \DataPath/i_REG_LDSTR_OUT[23] ), .ZN(n2200) );
  AOI22_X1 U15754 ( .A1(n11835), .A2(DRAM_DATA_OUT[24]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[24] ), .ZN(n2199) );
  AOI22_X1 U15755 ( .A1(n11835), .A2(DRAM_DATA_OUT[25]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[25] ), .ZN(n2198) );
  AOI22_X1 U15756 ( .A1(n11835), .A2(DRAM_DATA_OUT[26]), .B1(n8441), .B2(
        \DataPath/i_REG_LDSTR_OUT[26] ), .ZN(n2197) );
  AOI22_X1 U15757 ( .A1(n11835), .A2(DRAM_DATA_OUT[27]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[27] ), .ZN(n2196) );
  AOI22_X1 U15758 ( .A1(n11835), .A2(DRAM_DATA_OUT[28]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[28] ), .ZN(n2195) );
  AOI22_X1 U15759 ( .A1(n11835), .A2(DRAM_DATA_OUT[29]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[29] ), .ZN(n2194) );
  AOI22_X1 U15760 ( .A1(n11835), .A2(DRAM_DATA_OUT[30]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[30] ), .ZN(n2193) );
  AOI22_X1 U15761 ( .A1(n11835), .A2(DRAM_DATA_OUT[31]), .B1(n7757), .B2(
        \DataPath/i_REG_LDSTR_OUT[31] ), .ZN(n2192) );
  NOR2_X1 U15762 ( .A1(n10282), .A2(n11695), .ZN(n11697) );
  NAND4_X1 U15763 ( .A1(n11702), .A2(n11701), .A3(n11700), .A4(n11699), .ZN(
        n11703) );
  NAND4_X1 U15764 ( .A1(n11707), .A2(n11706), .A3(n11705), .A4(n11704), .ZN(
        n11711) );
  OAI21_X1 U15765 ( .B1(n10277), .B2(n11713), .A(n10278), .ZN(n11708) );
  AOI21_X1 U15766 ( .B1(n10277), .B2(n11713), .A(n11708), .ZN(n11710) );
  AOI211_X1 U15767 ( .C1(n10287), .C2(n11711), .A(n11710), .B(n11709), .ZN(
        n11712) );
  OAI22_X1 U15768 ( .A1(n510), .A2(n11734), .B1(n11712), .B2(n11735), .ZN(
        n7009) );
  NAND2_X1 U15769 ( .A1(i_ALU_OP[3]), .A2(n10299), .ZN(n11726) );
  OAI22_X1 U15770 ( .A1(n511), .A2(n11734), .B1(n11714), .B2(n11735), .ZN(
        n7008) );
  OAI22_X1 U15771 ( .A1(n512), .A2(n11734), .B1(n11715), .B2(n11735), .ZN(
        n7006) );
  NAND2_X1 U15772 ( .A1(n10285), .A2(n11716), .ZN(n11717) );
  NOR2_X1 U15773 ( .A1(n11724), .A2(n8428), .ZN(n11727) );
  AOI22_X1 U15774 ( .A1(\DataPath/i_REG_MEM_ALUOUT[0] ), .A2(n7757), .B1(
        n11835), .B2(n8208), .ZN(n1163) );
  AOI22_X1 U15775 ( .A1(\DataPath/i_REG_MEM_ALUOUT[1] ), .A2(n7757), .B1(
        n11835), .B2(n8168), .ZN(n1162) );
  AOI22_X1 U15776 ( .A1(n11835), .A2(DRAM_ADDRESS[2]), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[2] ), .ZN(n1161) );
  AOI22_X1 U15777 ( .A1(DRAM_ADDRESS[3]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[3] ), .ZN(n1160) );
  AOI22_X1 U15778 ( .A1(\DataPath/i_REG_MEM_ALUOUT[4] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[4]), .ZN(n1159) );
  AOI22_X1 U15779 ( .A1(n11835), .A2(DRAM_ADDRESS[5]), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[5] ), .ZN(n1158) );
  AOI22_X1 U15780 ( .A1(\DataPath/i_REG_MEM_ALUOUT[6] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[6]), .ZN(n1157) );
  AOI22_X1 U15781 ( .A1(DRAM_ADDRESS[7]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[7] ), .ZN(n1156) );
  AOI22_X1 U15782 ( .A1(\DataPath/i_REG_MEM_ALUOUT[8] ), .A2(n7757), .B1(
        n11835), .B2(DRAM_ADDRESS[8]), .ZN(n1155) );
  AOI22_X1 U15783 ( .A1(DRAM_ADDRESS[9]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[9] ), .ZN(n1154) );
  AOI22_X1 U15784 ( .A1(\DataPath/i_REG_MEM_ALUOUT[10] ), .A2(n7757), .B1(
        n11835), .B2(DRAM_ADDRESS[10]), .ZN(n1153) );
  AOI22_X1 U15785 ( .A1(\DataPath/i_REG_MEM_ALUOUT[11] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[11]), .ZN(n1152) );
  AOI22_X1 U15786 ( .A1(\DataPath/i_REG_MEM_ALUOUT[12] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[12]), .ZN(n1151) );
  AOI22_X1 U15787 ( .A1(DRAM_ADDRESS[13]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[13] ), .ZN(n1150) );
  AOI22_X1 U15788 ( .A1(\DataPath/i_REG_MEM_ALUOUT[14] ), .A2(n7757), .B1(
        n11835), .B2(DRAM_ADDRESS[14]), .ZN(n1149) );
  AOI22_X1 U15789 ( .A1(\DataPath/i_REG_MEM_ALUOUT[15] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[15]), .ZN(n1148) );
  AOI22_X1 U15790 ( .A1(\DataPath/i_REG_MEM_ALUOUT[16] ), .A2(n11836), .B1(
        n11835), .B2(DRAM_ADDRESS[16]), .ZN(n1147) );
  AOI22_X1 U15791 ( .A1(DRAM_ADDRESS[17]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[17] ), .ZN(n1146) );
  AOI22_X1 U15792 ( .A1(\DataPath/i_REG_MEM_ALUOUT[18] ), .A2(n7757), .B1(
        n11835), .B2(DRAM_ADDRESS[18]), .ZN(n1145) );
  AOI22_X1 U15793 ( .A1(\DataPath/i_REG_MEM_ALUOUT[19] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[19]), .ZN(n1144) );
  AOI22_X1 U15794 ( .A1(\DataPath/i_REG_MEM_ALUOUT[20] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[20]), .ZN(n1143) );
  AOI22_X1 U15795 ( .A1(DRAM_ADDRESS[21]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[21] ), .ZN(n1142) );
  AOI22_X1 U15796 ( .A1(\DataPath/i_REG_MEM_ALUOUT[22] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[22]), .ZN(n1141) );
  AOI22_X1 U15797 ( .A1(\DataPath/i_REG_MEM_ALUOUT[23] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[23]), .ZN(n1140) );
  AOI22_X1 U15798 ( .A1(\DataPath/i_REG_MEM_ALUOUT[24] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[24]), .ZN(n1139) );
  AOI22_X1 U15799 ( .A1(DRAM_ADDRESS[25]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[25] ), .ZN(n1138) );
  AOI22_X1 U15800 ( .A1(\DataPath/i_REG_MEM_ALUOUT[26] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[26]), .ZN(n1137) );
  AOI22_X1 U15801 ( .A1(\DataPath/i_REG_MEM_ALUOUT[27] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[27]), .ZN(n1136) );
  AOI22_X1 U15802 ( .A1(\DataPath/i_REG_MEM_ALUOUT[28] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[28]), .ZN(n1135) );
  AOI22_X1 U15803 ( .A1(DRAM_ADDRESS[29]), .A2(n11835), .B1(n7757), .B2(
        \DataPath/i_REG_MEM_ALUOUT[29] ), .ZN(n1134) );
  AOI22_X1 U15804 ( .A1(\DataPath/i_REG_MEM_ALUOUT[30] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[30]), .ZN(n1133) );
  AOI22_X1 U15805 ( .A1(\DataPath/i_REG_MEM_ALUOUT[31] ), .A2(n8441), .B1(
        n11835), .B2(DRAM_ADDRESS[31]), .ZN(n1130) );
  AOI22_X1 U15806 ( .A1(n11804), .A2(n8429), .B1(n8430), .B2(
        \DataPath/RF/bus_reg_dataout[2528] ), .ZN(n1126) );
  AOI22_X1 U15807 ( .A1(\DataPath/RF/bus_reg_dataout[2529] ), .A2(n8430), .B1(
        n11805), .B2(n8429), .ZN(n1125) );
  AOI22_X1 U15808 ( .A1(\DataPath/RF/bus_reg_dataout[2530] ), .A2(n8430), .B1(
        n11806), .B2(n8429), .ZN(n1124) );
  AOI22_X1 U15809 ( .A1(\DataPath/RF/bus_reg_dataout[2531] ), .A2(n8430), .B1(
        n11807), .B2(n8429), .ZN(n1123) );
  AOI22_X1 U15810 ( .A1(\DataPath/RF/bus_reg_dataout[2532] ), .A2(n8430), .B1(
        n11808), .B2(n8429), .ZN(n1122) );
  AOI22_X1 U15811 ( .A1(\DataPath/RF/bus_reg_dataout[2533] ), .A2(n8430), .B1(
        n11809), .B2(n8429), .ZN(n1121) );
  AOI22_X1 U15812 ( .A1(\DataPath/RF/bus_reg_dataout[2534] ), .A2(n8430), .B1(
        n11810), .B2(n11738), .ZN(n1120) );
  AOI22_X1 U15813 ( .A1(\DataPath/RF/bus_reg_dataout[2535] ), .A2(n8430), .B1(
        n11811), .B2(n11738), .ZN(n1119) );
  AOI22_X1 U15814 ( .A1(\DataPath/RF/bus_reg_dataout[2536] ), .A2(n8430), .B1(
        n11812), .B2(n11738), .ZN(n1118) );
  AOI22_X1 U15815 ( .A1(\DataPath/RF/bus_reg_dataout[2537] ), .A2(n8430), .B1(
        n11813), .B2(n11738), .ZN(n1117) );
  AOI22_X1 U15816 ( .A1(\DataPath/RF/bus_reg_dataout[2538] ), .A2(n8430), .B1(
        n11814), .B2(n11738), .ZN(n1116) );
  AOI22_X1 U15817 ( .A1(\DataPath/RF/bus_reg_dataout[2539] ), .A2(n8430), .B1(
        n11815), .B2(n11738), .ZN(n1115) );
  AOI22_X1 U15818 ( .A1(\DataPath/RF/bus_reg_dataout[2540] ), .A2(n8430), .B1(
        n11816), .B2(n11738), .ZN(n1114) );
  AOI22_X1 U15819 ( .A1(\DataPath/RF/bus_reg_dataout[2541] ), .A2(n8430), .B1(
        n11817), .B2(n11738), .ZN(n1113) );
  AOI22_X1 U15820 ( .A1(\DataPath/RF/bus_reg_dataout[2542] ), .A2(n8430), .B1(
        n11818), .B2(n11738), .ZN(n1112) );
  AOI22_X1 U15821 ( .A1(\DataPath/RF/bus_reg_dataout[2543] ), .A2(n8430), .B1(
        n11819), .B2(n8429), .ZN(n1111) );
  AOI22_X1 U15822 ( .A1(\DataPath/RF/bus_reg_dataout[2544] ), .A2(n8430), .B1(
        n11820), .B2(n8429), .ZN(n1110) );
  AOI22_X1 U15823 ( .A1(\DataPath/RF/bus_reg_dataout[2545] ), .A2(n8430), .B1(
        n11823), .B2(n8429), .ZN(n1109) );
  AOI22_X1 U15824 ( .A1(\DataPath/RF/bus_reg_dataout[2546] ), .A2(n8430), .B1(
        n11746), .B2(n8429), .ZN(n1108) );
  AOI22_X1 U15825 ( .A1(\DataPath/RF/bus_reg_dataout[2547] ), .A2(n8430), .B1(
        n11747), .B2(n8429), .ZN(n1107) );
  AOI22_X1 U15826 ( .A1(\DataPath/RF/bus_reg_dataout[2548] ), .A2(n8430), .B1(
        n11748), .B2(n8429), .ZN(n1106) );
  AOI22_X1 U15827 ( .A1(\DataPath/RF/bus_reg_dataout[2549] ), .A2(n11739), 
        .B1(n11749), .B2(n8429), .ZN(n1105) );
  AOI22_X1 U15828 ( .A1(\DataPath/RF/bus_reg_dataout[2550] ), .A2(n11739), 
        .B1(n11791), .B2(n8429), .ZN(n1104) );
  AOI22_X1 U15829 ( .A1(\DataPath/RF/bus_reg_dataout[2551] ), .A2(n11739), 
        .B1(n11750), .B2(n8429), .ZN(n1103) );
  AOI22_X1 U15830 ( .A1(\DataPath/RF/bus_reg_dataout[2552] ), .A2(n11739), 
        .B1(n11793), .B2(n8429), .ZN(n1102) );
  AOI22_X1 U15831 ( .A1(\DataPath/RF/bus_reg_dataout[2553] ), .A2(n11739), 
        .B1(n11794), .B2(n8429), .ZN(n1101) );
  AOI22_X1 U15832 ( .A1(\DataPath/RF/bus_reg_dataout[2554] ), .A2(n11739), 
        .B1(n11751), .B2(n8429), .ZN(n1100) );
  AOI22_X1 U15833 ( .A1(\DataPath/RF/bus_reg_dataout[2555] ), .A2(n11739), 
        .B1(n11796), .B2(n8429), .ZN(n1099) );
  AOI22_X1 U15834 ( .A1(\DataPath/RF/bus_reg_dataout[2556] ), .A2(n11739), 
        .B1(n11752), .B2(n8429), .ZN(n1098) );
  AOI22_X1 U15835 ( .A1(\DataPath/RF/bus_reg_dataout[2557] ), .A2(n11739), 
        .B1(n11753), .B2(n8429), .ZN(n1097) );
  AOI22_X1 U15836 ( .A1(\DataPath/RF/bus_reg_dataout[2558] ), .A2(n11739), 
        .B1(n11754), .B2(n8429), .ZN(n1096) );
  AOI22_X1 U15837 ( .A1(\DataPath/RF/bus_reg_dataout[2559] ), .A2(n8430), .B1(
        n11803), .B2(n8429), .ZN(n1093) );
  AOI22_X1 U15838 ( .A1(n11804), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2496] ), .ZN(n1089) );
  AOI22_X1 U15839 ( .A1(n11805), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2497] ), .ZN(n1088) );
  AOI22_X1 U15840 ( .A1(n11806), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2498] ), .ZN(n1087) );
  AOI22_X1 U15841 ( .A1(n11807), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2499] ), .ZN(n1086) );
  AOI22_X1 U15842 ( .A1(n11808), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2500] ), .ZN(n1085) );
  AOI22_X1 U15843 ( .A1(n11809), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2501] ), .ZN(n1084) );
  AOI22_X1 U15844 ( .A1(n11810), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2502] ), .ZN(n1083) );
  AOI22_X1 U15845 ( .A1(n11811), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2503] ), .ZN(n1082) );
  AOI22_X1 U15846 ( .A1(n11812), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2504] ), .ZN(n1081) );
  AOI22_X1 U15847 ( .A1(n11813), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2505] ), .ZN(n1080) );
  AOI22_X1 U15848 ( .A1(n11814), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2506] ), .ZN(n1079) );
  AOI22_X1 U15849 ( .A1(n11815), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2507] ), .ZN(n1078) );
  AOI22_X1 U15850 ( .A1(n11816), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2508] ), .ZN(n1077) );
  AOI22_X1 U15851 ( .A1(n11817), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2509] ), .ZN(n1076) );
  AOI22_X1 U15852 ( .A1(n11818), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2510] ), .ZN(n1075) );
  AOI22_X1 U15853 ( .A1(n11819), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2511] ), .ZN(n1074) );
  AOI22_X1 U15854 ( .A1(n11820), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2512] ), .ZN(n1073) );
  AOI22_X1 U15855 ( .A1(n11823), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2513] ), .ZN(n1072) );
  AOI22_X1 U15856 ( .A1(n11746), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2514] ), .ZN(n1071) );
  AOI22_X1 U15857 ( .A1(n11747), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2515] ), .ZN(n1070) );
  AOI22_X1 U15858 ( .A1(n11748), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2516] ), .ZN(n1069) );
  AOI22_X1 U15859 ( .A1(n11749), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2517] ), .ZN(n1068) );
  AOI22_X1 U15860 ( .A1(n11791), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2518] ), .ZN(n1067) );
  AOI22_X1 U15861 ( .A1(n11750), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2519] ), .ZN(n1066) );
  AOI22_X1 U15862 ( .A1(n11793), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2520] ), .ZN(n1065) );
  AOI22_X1 U15863 ( .A1(n11794), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2521] ), .ZN(n1064) );
  AOI22_X1 U15864 ( .A1(n11751), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2522] ), .ZN(n1063) );
  AOI22_X1 U15865 ( .A1(n11796), .A2(n8432), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2523] ), .ZN(n1062) );
  AOI22_X1 U15866 ( .A1(n11752), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2524] ), .ZN(n1061) );
  AOI22_X1 U15867 ( .A1(n11753), .A2(n8432), .B1(n11742), .B2(
        \DataPath/RF/bus_reg_dataout[2525] ), .ZN(n1060) );
  AOI22_X1 U15868 ( .A1(n11754), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2526] ), .ZN(n1059) );
  AOI22_X1 U15869 ( .A1(n11803), .A2(n11743), .B1(n8431), .B2(
        \DataPath/RF/bus_reg_dataout[2527] ), .ZN(n1056) );
  AOI22_X1 U15870 ( .A1(n11804), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2464] ), .ZN(n1052) );
  AOI22_X1 U15871 ( .A1(n11805), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2465] ), .ZN(n1051) );
  AOI22_X1 U15872 ( .A1(n11806), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2466] ), .ZN(n1050) );
  AOI22_X1 U15873 ( .A1(n11807), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2467] ), .ZN(n1049) );
  AOI22_X1 U15874 ( .A1(n11808), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2468] ), .ZN(n1048) );
  AOI22_X1 U15875 ( .A1(n11809), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2469] ), .ZN(n1047) );
  AOI22_X1 U15876 ( .A1(n11810), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2470] ), .ZN(n1046) );
  AOI22_X1 U15877 ( .A1(n11811), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2471] ), .ZN(n1045) );
  AOI22_X1 U15878 ( .A1(n11812), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2472] ), .ZN(n1044) );
  AOI22_X1 U15879 ( .A1(n11813), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2473] ), .ZN(n1043) );
  AOI22_X1 U15880 ( .A1(n11814), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2474] ), .ZN(n1042) );
  AOI22_X1 U15881 ( .A1(n11815), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2475] ), .ZN(n1041) );
  AOI22_X1 U15882 ( .A1(n11816), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2476] ), .ZN(n1040) );
  AOI22_X1 U15883 ( .A1(n11817), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2477] ), .ZN(n1039) );
  AOI22_X1 U15884 ( .A1(n11818), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2478] ), .ZN(n1038) );
  AOI22_X1 U15885 ( .A1(n11819), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2479] ), .ZN(n1037) );
  AOI22_X1 U15886 ( .A1(n11820), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2480] ), .ZN(n1036) );
  AOI22_X1 U15887 ( .A1(n11823), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2481] ), .ZN(n1035) );
  AOI22_X1 U15888 ( .A1(n11746), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2482] ), .ZN(n1034) );
  AOI22_X1 U15889 ( .A1(n11747), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2483] ), .ZN(n1033) );
  AOI22_X1 U15890 ( .A1(n11748), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2484] ), .ZN(n1032) );
  AOI22_X1 U15891 ( .A1(n11749), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2485] ), .ZN(n1031) );
  AOI22_X1 U15892 ( .A1(n11791), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2486] ), .ZN(n1030) );
  AOI22_X1 U15893 ( .A1(n11750), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2487] ), .ZN(n1029) );
  AOI22_X1 U15894 ( .A1(n11793), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2488] ), .ZN(n1028) );
  AOI22_X1 U15895 ( .A1(n11794), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2489] ), .ZN(n1027) );
  AOI22_X1 U15896 ( .A1(n11751), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2490] ), .ZN(n1026) );
  AOI22_X1 U15897 ( .A1(n11796), .A2(n8434), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2491] ), .ZN(n1025) );
  AOI22_X1 U15898 ( .A1(n11752), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2492] ), .ZN(n1024) );
  AOI22_X1 U15899 ( .A1(n11753), .A2(n8434), .B1(n11755), .B2(
        \DataPath/RF/bus_reg_dataout[2493] ), .ZN(n1023) );
  AOI22_X1 U15900 ( .A1(n11754), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2494] ), .ZN(n1022) );
  AOI22_X1 U15901 ( .A1(n11803), .A2(n11756), .B1(n8433), .B2(
        \DataPath/RF/bus_reg_dataout[2495] ), .ZN(n1019) );
  OAI22_X1 U15902 ( .A1(n8173), .A2(n11758), .B1(n8437), .B2(n11757), .ZN(
        n11759) );
  AOI22_X1 U15903 ( .A1(\DataPath/RF/bus_reg_dataout[2432] ), .A2(n8435), .B1(
        n11770), .B2(n11774), .ZN(n1015) );
  AOI22_X1 U15904 ( .A1(\DataPath/RF/bus_reg_dataout[2433] ), .A2(n11771), 
        .B1(n11770), .B2(n11775), .ZN(n1014) );
  AOI22_X1 U15905 ( .A1(\DataPath/RF/bus_reg_dataout[2434] ), .A2(n8435), .B1(
        n11770), .B2(n11776), .ZN(n1013) );
  AOI22_X1 U15906 ( .A1(\DataPath/RF/bus_reg_dataout[2435] ), .A2(n11771), 
        .B1(n11770), .B2(n11777), .ZN(n1012) );
  AOI22_X1 U15907 ( .A1(\DataPath/RF/bus_reg_dataout[2436] ), .A2(n11771), 
        .B1(n11770), .B2(n11778), .ZN(n1011) );
  AOI22_X1 U15908 ( .A1(\DataPath/RF/bus_reg_dataout[2437] ), .A2(n11771), 
        .B1(n11770), .B2(n11779), .ZN(n1010) );
  AOI22_X1 U15909 ( .A1(\DataPath/RF/bus_reg_dataout[2438] ), .A2(n11771), 
        .B1(n11770), .B2(n11780), .ZN(n1009) );
  AOI22_X1 U15910 ( .A1(\DataPath/RF/bus_reg_dataout[2439] ), .A2(n8435), .B1(
        n11770), .B2(n11781), .ZN(n1008) );
  OAI22_X1 U15911 ( .A1(n11812), .A2(n11771), .B1(
        \DataPath/RF/bus_reg_dataout[2440] ), .B2(n11759), .ZN(n1007) );
  AOI22_X1 U15912 ( .A1(\DataPath/RF/bus_reg_dataout[2441] ), .A2(n8435), .B1(
        n11770), .B2(n11760), .ZN(n1006) );
  AOI22_X1 U15913 ( .A1(\DataPath/RF/bus_reg_dataout[2442] ), .A2(n8435), .B1(
        n11770), .B2(n11783), .ZN(n1005) );
  AOI22_X1 U15914 ( .A1(\DataPath/RF/bus_reg_dataout[2443] ), .A2(n8435), .B1(
        n11770), .B2(n11784), .ZN(n1004) );
  AOI22_X1 U15915 ( .A1(\DataPath/RF/bus_reg_dataout[2444] ), .A2(n8435), .B1(
        n11770), .B2(n11761), .ZN(n1003) );
  AOI22_X1 U15916 ( .A1(\DataPath/RF/bus_reg_dataout[2445] ), .A2(n8435), .B1(
        n11770), .B2(n11785), .ZN(n1002) );
  AOI22_X1 U15917 ( .A1(\DataPath/RF/bus_reg_dataout[2446] ), .A2(n8435), .B1(
        n11770), .B2(n11786), .ZN(n1001) );
  AOI22_X1 U15918 ( .A1(\DataPath/RF/bus_reg_dataout[2447] ), .A2(n8435), .B1(
        n11770), .B2(n11762), .ZN(n1000) );
  AOI22_X1 U15919 ( .A1(\DataPath/RF/bus_reg_dataout[2448] ), .A2(n8435), .B1(
        n11770), .B2(n11763), .ZN(n999) );
  AOI22_X1 U15920 ( .A1(\DataPath/RF/bus_reg_dataout[2449] ), .A2(n8435), .B1(
        n11770), .B2(n11764), .ZN(n998) );
  AOI22_X1 U15921 ( .A1(\DataPath/RF/bus_reg_dataout[2450] ), .A2(n8435), .B1(
        n11770), .B2(n11787), .ZN(n997) );
  AOI22_X1 U15922 ( .A1(\DataPath/RF/bus_reg_dataout[2451] ), .A2(n8435), .B1(
        n11770), .B2(n11788), .ZN(n996) );
  AOI22_X1 U15923 ( .A1(\DataPath/RF/bus_reg_dataout[2452] ), .A2(n8435), .B1(
        n11770), .B2(n11789), .ZN(n995) );
  AOI22_X1 U15924 ( .A1(\DataPath/RF/bus_reg_dataout[2453] ), .A2(n11771), 
        .B1(n11770), .B2(n11790), .ZN(n994) );
  AOI22_X1 U15925 ( .A1(\DataPath/RF/bus_reg_dataout[2454] ), .A2(n11771), 
        .B1(n11770), .B2(n11765), .ZN(n993) );
  AOI22_X1 U15926 ( .A1(\DataPath/RF/bus_reg_dataout[2455] ), .A2(n11771), 
        .B1(n11770), .B2(n11792), .ZN(n992) );
  AOI22_X1 U15927 ( .A1(\DataPath/RF/bus_reg_dataout[2456] ), .A2(n8435), .B1(
        n11770), .B2(n11766), .ZN(n991) );
  AOI22_X1 U15928 ( .A1(\DataPath/RF/bus_reg_dataout[2457] ), .A2(n8435), .B1(
        n11770), .B2(n11767), .ZN(n990) );
  AOI22_X1 U15929 ( .A1(\DataPath/RF/bus_reg_dataout[2458] ), .A2(n11771), 
        .B1(n11770), .B2(n11795), .ZN(n989) );
  AOI22_X1 U15930 ( .A1(\DataPath/RF/bus_reg_dataout[2459] ), .A2(n8435), .B1(
        n11770), .B2(n11768), .ZN(n988) );
  AOI22_X1 U15931 ( .A1(\DataPath/RF/bus_reg_dataout[2460] ), .A2(n8435), .B1(
        n11770), .B2(n11797), .ZN(n987) );
  AOI22_X1 U15932 ( .A1(\DataPath/RF/bus_reg_dataout[2461] ), .A2(n8435), .B1(
        n11770), .B2(n11798), .ZN(n986) );
  AOI22_X1 U15933 ( .A1(\DataPath/RF/bus_reg_dataout[2462] ), .A2(n8435), .B1(
        n11770), .B2(n11799), .ZN(n985) );
  AOI22_X1 U15934 ( .A1(\DataPath/RF/bus_reg_dataout[2463] ), .A2(n8435), .B1(
        n11770), .B2(n11769), .ZN(n982) );
  AOI22_X1 U15935 ( .A1(\DataPath/RF/bus_reg_dataout[2400] ), .A2(n8438), .B1(
        n11800), .B2(n11774), .ZN(n977) );
  AOI22_X1 U15936 ( .A1(\DataPath/RF/bus_reg_dataout[2401] ), .A2(n8438), .B1(
        n11800), .B2(n11775), .ZN(n976) );
  AOI22_X1 U15937 ( .A1(\DataPath/RF/bus_reg_dataout[2402] ), .A2(n8438), .B1(
        n11800), .B2(n11776), .ZN(n975) );
  AOI22_X1 U15938 ( .A1(\DataPath/RF/bus_reg_dataout[2403] ), .A2(n8438), .B1(
        n11800), .B2(n11777), .ZN(n974) );
  AOI22_X1 U15939 ( .A1(\DataPath/RF/bus_reg_dataout[2404] ), .A2(n8438), .B1(
        n11800), .B2(n11778), .ZN(n973) );
  AOI22_X1 U15940 ( .A1(\DataPath/RF/bus_reg_dataout[2405] ), .A2(n8438), .B1(
        n11800), .B2(n11779), .ZN(n972) );
  AOI22_X1 U15941 ( .A1(\DataPath/RF/bus_reg_dataout[2406] ), .A2(n8438), .B1(
        n11800), .B2(n11780), .ZN(n971) );
  AOI22_X1 U15942 ( .A1(\DataPath/RF/bus_reg_dataout[2407] ), .A2(n8438), .B1(
        n11800), .B2(n11781), .ZN(n970) );
  AOI22_X1 U15943 ( .A1(\DataPath/RF/bus_reg_dataout[2408] ), .A2(n8438), .B1(
        n11800), .B2(n11782), .ZN(n969) );
  AOI22_X1 U15944 ( .A1(n11813), .A2(n11802), .B1(n11801), .B2(
        \DataPath/RF/bus_reg_dataout[2409] ), .ZN(n968) );
  AOI22_X1 U15945 ( .A1(\DataPath/RF/bus_reg_dataout[2410] ), .A2(n8438), .B1(
        n11800), .B2(n11783), .ZN(n967) );
  AOI22_X1 U15946 ( .A1(\DataPath/RF/bus_reg_dataout[2411] ), .A2(n8438), .B1(
        n11800), .B2(n11784), .ZN(n966) );
  AOI22_X1 U15947 ( .A1(n11816), .A2(n11802), .B1(n11801), .B2(
        \DataPath/RF/bus_reg_dataout[2412] ), .ZN(n965) );
  AOI22_X1 U15948 ( .A1(\DataPath/RF/bus_reg_dataout[2413] ), .A2(n8438), .B1(
        n11800), .B2(n11785), .ZN(n964) );
  AOI22_X1 U15949 ( .A1(\DataPath/RF/bus_reg_dataout[2414] ), .A2(n11801), 
        .B1(n11800), .B2(n11786), .ZN(n963) );
  AOI22_X1 U15950 ( .A1(n11819), .A2(n11802), .B1(n11801), .B2(
        \DataPath/RF/bus_reg_dataout[2415] ), .ZN(n962) );
  AOI22_X1 U15951 ( .A1(n11820), .A2(n11802), .B1(n11801), .B2(
        \DataPath/RF/bus_reg_dataout[2416] ), .ZN(n961) );
  AOI22_X1 U15952 ( .A1(n11823), .A2(n11802), .B1(n11801), .B2(
        \DataPath/RF/bus_reg_dataout[2417] ), .ZN(n960) );
  AOI22_X1 U15953 ( .A1(\DataPath/RF/bus_reg_dataout[2418] ), .A2(n11801), 
        .B1(n11800), .B2(n11787), .ZN(n958) );
  AOI22_X1 U15954 ( .A1(\DataPath/RF/bus_reg_dataout[2419] ), .A2(n8438), .B1(
        n11800), .B2(n11788), .ZN(n956) );
  AOI22_X1 U15955 ( .A1(\DataPath/RF/bus_reg_dataout[2420] ), .A2(n8438), .B1(
        n11800), .B2(n11789), .ZN(n954) );
  AOI22_X1 U15956 ( .A1(\DataPath/RF/bus_reg_dataout[2421] ), .A2(n11801), 
        .B1(n11800), .B2(n11790), .ZN(n952) );
  AOI22_X1 U15957 ( .A1(n11791), .A2(n11802), .B1(n11801), .B2(
        \DataPath/RF/bus_reg_dataout[2422] ), .ZN(n950) );
  AOI22_X1 U15958 ( .A1(\DataPath/RF/bus_reg_dataout[2423] ), .A2(n8438), .B1(
        n11800), .B2(n11792), .ZN(n948) );
  AOI22_X1 U15959 ( .A1(n11793), .A2(n11802), .B1(n8438), .B2(
        \DataPath/RF/bus_reg_dataout[2424] ), .ZN(n946) );
  AOI22_X1 U15960 ( .A1(n11794), .A2(n11802), .B1(n8438), .B2(
        \DataPath/RF/bus_reg_dataout[2425] ), .ZN(n944) );
  AOI22_X1 U15961 ( .A1(\DataPath/RF/bus_reg_dataout[2426] ), .A2(n11801), 
        .B1(n11800), .B2(n11795), .ZN(n942) );
  AOI22_X1 U15962 ( .A1(n11796), .A2(n11802), .B1(n8438), .B2(
        \DataPath/RF/bus_reg_dataout[2427] ), .ZN(n940) );
  AOI22_X1 U15963 ( .A1(\DataPath/RF/bus_reg_dataout[2428] ), .A2(n8438), .B1(
        n11800), .B2(n11797), .ZN(n938) );
  AOI22_X1 U15964 ( .A1(\DataPath/RF/bus_reg_dataout[2429] ), .A2(n8438), .B1(
        n11800), .B2(n11798), .ZN(n936) );
  AOI22_X1 U15965 ( .A1(\DataPath/RF/bus_reg_dataout[2430] ), .A2(n8438), .B1(
        n11800), .B2(n11799), .ZN(n934) );
  AOI22_X1 U15966 ( .A1(n11803), .A2(n11802), .B1(n8438), .B2(
        \DataPath/RF/bus_reg_dataout[2431] ), .ZN(n930) );
  AOI22_X1 U15967 ( .A1(n11804), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2368] ), .ZN(n928) );
  AOI22_X1 U15968 ( .A1(n11805), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2369] ), .ZN(n926) );
  AOI22_X1 U15969 ( .A1(n11806), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2370] ), .ZN(n924) );
  AOI22_X1 U15970 ( .A1(n11807), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2371] ), .ZN(n922) );
  AOI22_X1 U15971 ( .A1(n11808), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2372] ), .ZN(n920) );
  AOI22_X1 U15972 ( .A1(n11809), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2373] ), .ZN(n918) );
  AOI22_X1 U15973 ( .A1(n11810), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2374] ), .ZN(n916) );
  AOI22_X1 U15974 ( .A1(n11811), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2375] ), .ZN(n914) );
  AOI22_X1 U15975 ( .A1(n11812), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2376] ), .ZN(n912) );
  AOI22_X1 U15976 ( .A1(n11813), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2377] ), .ZN(n910) );
  AOI22_X1 U15977 ( .A1(n11814), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2378] ), .ZN(n908) );
  AOI22_X1 U15978 ( .A1(n11815), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2379] ), .ZN(n906) );
  AOI22_X1 U15979 ( .A1(n11816), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2380] ), .ZN(n904) );
  AOI22_X1 U15980 ( .A1(n11817), .A2(n8440), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2381] ), .ZN(n902) );
  AOI22_X1 U15981 ( .A1(n11818), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2382] ), .ZN(n900) );
  AOI22_X1 U15982 ( .A1(n11819), .A2(n8440), .B1(n11821), .B2(
        \DataPath/RF/bus_reg_dataout[2383] ), .ZN(n898) );
  AOI22_X1 U15983 ( .A1(n11820), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2384] ), .ZN(n896) );
  AOI22_X1 U15984 ( .A1(n11823), .A2(n11822), .B1(n8439), .B2(
        \DataPath/RF/bus_reg_dataout[2385] ), .ZN(n892) );
  INV_X1 U15985 ( .A(\CU_I/CW_ID[DRAM_RE] ), .ZN(n11824) );
  OAI22_X1 U15986 ( .A1(n11830), .A2(n11824), .B1(n11828), .B2(n8200), .ZN(
        n370) );
  INV_X1 U15987 ( .A(\CU_I/CW_ID[DATA_SIZE][1] ), .ZN(n11825) );
  OAI22_X1 U15988 ( .A1(n11830), .A2(n11825), .B1(n11828), .B2(n8201), .ZN(
        n369) );
  INV_X1 U15989 ( .A(\CU_I/CW_ID[DATA_SIZE][0] ), .ZN(n11826) );
  OAI22_X1 U15990 ( .A1(n11830), .A2(n11826), .B1(n11828), .B2(n8202), .ZN(
        n368) );
  INV_X1 U15991 ( .A(\CU_I/CW_ID[MEM_EN] ), .ZN(n11827) );
  OAI22_X1 U15992 ( .A1(n11830), .A2(n11827), .B1(n11828), .B2(n8199), .ZN(
        n367) );
  INV_X1 U15993 ( .A(\CU_I/CW_ID[DRAM_WE] ), .ZN(n11829) );
  OAI22_X1 U15994 ( .A1(n11830), .A2(n11829), .B1(n11828), .B2(n8203), .ZN(
        n366) );
  AOI22_X1 U15995 ( .A1(n11835), .A2(\DataPath/i_PIPLIN_WRB2[4] ), .B1(n7757), 
        .B2(i_ADD_WB[4]), .ZN(n11831) );
  INV_X1 U15996 ( .A(n11831), .ZN(n363) );
  AOI22_X1 U15997 ( .A1(n11835), .A2(\DataPath/i_PIPLIN_WRB2[3] ), .B1(n7757), 
        .B2(i_ADD_WB[3]), .ZN(n11832) );
  INV_X1 U15998 ( .A(n11832), .ZN(n362) );
  AOI22_X1 U15999 ( .A1(i_ADD_WB[2]), .A2(n8441), .B1(n11835), .B2(
        \DataPath/i_PIPLIN_WRB2[2] ), .ZN(n11833) );
  INV_X1 U16000 ( .A(n11833), .ZN(n361) );
  AOI22_X1 U16001 ( .A1(n11835), .A2(\DataPath/i_PIPLIN_WRB2[1] ), .B1(n7757), 
        .B2(i_ADD_WB[1]), .ZN(n11834) );
  INV_X1 U16002 ( .A(n11834), .ZN(n360) );
  AOI22_X1 U16003 ( .A1(i_ADD_WB[0]), .A2(n8441), .B1(n11835), .B2(
        \DataPath/i_PIPLIN_WRB2[0] ), .ZN(n11837) );
  INV_X1 U16004 ( .A(n11837), .ZN(n359) );
  AOI22_X1 U16005 ( .A1(n470), .A2(n11841), .B1(n471), .B2(n11840), .ZN(n11844) );
  NAND2_X1 U16006 ( .A1(n10293), .A2(n9270), .ZN(n11842) );
  OAI21_X1 U16007 ( .B1(n10295), .B2(n470), .A(n11842), .ZN(n11843) );
  AOI21_X1 U16008 ( .B1(n11844), .B2(n11843), .A(RST), .ZN(n99) );
  OAI21_X1 U16009 ( .B1(n10295), .B2(n11846), .A(n11845), .ZN(DRAMRF_ISSUE) );
  AND2_X1 U16010 ( .A1(n11848), .A2(n11847), .ZN(n90) );
  OAI21_X1 U16011 ( .B1(n8294), .B2(n185), .A(n11849), .ZN(n43) );
  OAI21_X1 U16012 ( .B1(n8294), .B2(n186), .A(n11850), .ZN(n42) );
  OAI21_X1 U16013 ( .B1(n8107), .B2(n8294), .A(n11851), .ZN(n40) );
  OAI21_X1 U16014 ( .B1(n8196), .B2(n8294), .A(n11852), .ZN(n36) );
endmodule

