package CONSTANTS is
   constant IVDELAY : time := 0.1 ns;
   constant NDDELAY : time := 0.2 ns;
   constant NRDELAY : time := 0.2 ns;
end CONSTANTS;
