library ieee;
use ieee.std_logic_1164.all;
use work.myTypes.all;
 
package record_CU is

	-- Control word bits
	type control_word is record
		fetch_en            : std_logic; -- F
		fecth_stall         : std_logic; -- S
		pc_en               : std_logic; -- P
		jump_en             : std_logic; -- J
		call                : std_logic; -- L
		ret                 : std_logic; -- E
		rf_rd1_en           : std_logic; -- 1
		rf_rd2_en           : std_logic; -- 2
		sel_cmpb            : std_logic; -- P
		unsigned_id         : std_logic; -- U
		npc_sel             : std_logic; -- N
		hazard_table_wr1    : std_logic; -- H
		id_en               : std_logic; -- D
		ex_en               : std_logic; -- X
		muxa_sel            : std_logic; -- A
		muxb_sel            : std_logic; -- B
		alu_opcode          : alu_op_sig_t; -- -----
		set_cmp             : set_op_sig_t; -- +++
		sel_alu             : std_logic; -- T
		dram_we             : std_logic; -- W
		dram_re             : std_logic; -- R
		data_size           : std_logic_vector(1 downto 0); -- 10
		mem_en              : std_logic; -- M
		wb_mux_sel          : std_logic; -- C
		wb_en               : std_logic; -- K
	end record control_word;

	constant R_TYPE_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        => ALU_ADD,
		set_cmp           => SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant VOID_RECORD: control_word := (
		fetch_en          => '0', 
		fecth_stall       => '0',
		pc_en             => '0',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        => ALU_ADD,
		set_cmp           => SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant J_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant JAL_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant BEQZ_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant BNEZ_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant ADDI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant ADDUI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SUBI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SUB,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SUBUI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SUB,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant ANDI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_AND,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant ORI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_OR,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant XORI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_XOR,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant LHI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '1',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SLL,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant JR_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '1',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant JALR_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '1',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SLLI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SLL,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant NOP_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant SRLI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SRL,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SRAI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SRA,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SEQI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SNEI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SNE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SLTI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SGTI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SLEI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SGEI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant CALL_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RET_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '1',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '1',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant LB_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "10",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant LH_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "01",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant LW_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant LBU_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "10",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant LHU_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "01",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant SB_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '1',
		dram_re           => '0',
		data_size         => "10",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant SH_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '1',
		dram_re           => '0',
		data_size         => "01",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant SW_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '1',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant BGT_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant BGE_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant BLT_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant BLE_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant TICKTMR_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SLTUI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SGTUI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SLEUI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant SGEUI_RECORD: control_word := (
		fetch_en          => '1', 
		fecth_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

end package record_CU;