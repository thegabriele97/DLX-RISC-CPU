
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_registerfile_generic_NBIT_DATA32_NBIT_ADD5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_registerfile_generic_NBIT_DATA32_NBIT_ADD5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_registerfile_generic_NBIT_DATA32_NBIT_ADD5.all;

entity registerfile_generic_NBIT_DATA32_NBIT_ADD5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end registerfile_generic_NBIT_DATA32_NBIT_ADD5;

architecture SYN_behavioural of registerfile_generic_NBIT_DATA32_NBIT_ADD5 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, 
      N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, 
      N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, 
      N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, 
      N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, 
      N467, N468, N469, N470, N471, n1180, n1181, n1182, n1183, n1184, n1185, 
      n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, 
      n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, 
      n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, 
      n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, 
      n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
      n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, 
      n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, 
      n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, 
      n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
      n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, 
      n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, 
      n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, 
      n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, 
      n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, 
      n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
      n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, 
      n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
      n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, 
      n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, 
      n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
      n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, 
      n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
      n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, 
      n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, 
      n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, 
      n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, 
      n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, 
      n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, 
      n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, 
      n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, 
      n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, 
      n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, 
      n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, 
      n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, 
      n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, 
      n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, 
      n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, 
      n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, 
      n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, 
      n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, 
      n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, 
      n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, 
      n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, 
      n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, 
      n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, 
      n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
      n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
      n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, 
      n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, 
      n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, 
      n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, 
      n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, 
      n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, 
      n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, 
      n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, 
      n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
      n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, 
      n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, 
      n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, 
      n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n6682, n6683, 
      n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
      n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, 
      n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n7741, 
      n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, 
      n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, 
      n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, 
      n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, 
      n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, 
      n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, 
      n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, 
      n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, 
      n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, 
      n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, 
      n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, 
      n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, 
      n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, 
      n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, 
      n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, 
      n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, 
      n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, 
      n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, 
      n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, 
      n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, 
      n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, 
      n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, 
      n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, 
      n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, 
      n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, 
      n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, 
      n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, 
      n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, 
      n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, 
      n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, 
      n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, 
      n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, 
      n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, 
      n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, 
      n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, 
      n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, 
      n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, 
      n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, 
      n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, 
      n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, 
      n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, 
      n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, 
      n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, 
      n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, 
      n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, 
      n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, 
      n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, 
      n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, 
      n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, 
      n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, 
      n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, 
      n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, 
      n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, 
      n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, 
      n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, 
      n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, 
      n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, 
      n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, 
      n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, 
      n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, 
      n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, 
      n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, 
      n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, 
      n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, 
      n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, 
      n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, 
      n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, 
      n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, 
      n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, 
      n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, 
      n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, 
      n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, 
      n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, 
      n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, 
      n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, 
      n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, 
      n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, 
      n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, 
      n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, 
      n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, 
      n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, 
      n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, 
      n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, 
      n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, 
      n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, 
      n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, 
      n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, 
      n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, 
      n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, 
      n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, 
      n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, 
      n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, 
      n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, 
      n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, 
      n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, 
      n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, 
      n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, 
      n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, 
      n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, 
      n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, 
      n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, 
      n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, 
      n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, 
      n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, 
      n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, 
      n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, 
      n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, 
      n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, 
      n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, 
      n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, 
      n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, 
      n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, 
      n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, 
      n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, 
      n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, 
      n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, 
      n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, 
      n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, 
      n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, 
      n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, 
      n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, 
      n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, 
      n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, 
      n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, 
      n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, 
      n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, 
      n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, 
      n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, 
      n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, 
      n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, 
      n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, 
      n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, 
      n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, 
      n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, 
      n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, 
      n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, 
      n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, 
      n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, 
      n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, 
      n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, 
      n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, 
      n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, 
      n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, 
      n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, 
      n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, 
      n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, 
      n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, 
      n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, 
      n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, 
      n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, 
      n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, 
      n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, 
      n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, 
      n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, 
      n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, 
      n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, 
      n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, 
      n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, 
      n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, 
      n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, 
      n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, 
      n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, 
      n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, 
      n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, 
      n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, 
      n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, 
      n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, 
      n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, 
      n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, 
      n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, 
      n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, 
      n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, 
      n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, 
      n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, 
      n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, 
      n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, 
      n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, 
      n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, 
      n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, 
      n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, 
      n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, 
      n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, 
      n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, 
      n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, 
      n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, 
      n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, 
      n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, 
      n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, 
      n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, 
      n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, 
      n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, 
      n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, 
      n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, 
      n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, 
      n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, 
      n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, 
      n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, 
      n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, 
      n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, 
      n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, 
      n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, 
      n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, 
      n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, 
      n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, 
      n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, 
      n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, 
      n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, 
      n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, 
      n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, 
      n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, 
      n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, 
      n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, 
      n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, 
      n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, 
      n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, 
      n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, 
      n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, 
      n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, 
      n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, 
      n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, 
      n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, 
      n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, 
      n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, 
      n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, 
      n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, 
      n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, 
      n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, 
      n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, 
      n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, 
      n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, 
      n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, 
      n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, 
      n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, 
      n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, 
      n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, 
      n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, 
      n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, 
      n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, 
      n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, 
      n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, 
      n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, 
      n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, 
      n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, 
      n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, 
      n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, 
      n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, 
      n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, 
      n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, 
      n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, 
      n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, 
      n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, 
      n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, 
      n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, 
      n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, 
      n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, 
      n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, 
      n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, 
      n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, 
      n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, 
      n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, 
      n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, 
      n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, 
      n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, 
      n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, 
      n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, 
      n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, 
      n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, 
      n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, 
      n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, 
      n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, 
      n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, 
      n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, 
      n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, 
      n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, 
      n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, 
      n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, 
      n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, 
      n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, 
      n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, 
      n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, 
      n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, 
      n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, 
      n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, 
      n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, 
      n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, 
      n10533, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, 
      n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, 
      n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, 
      n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, 
      n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, 
      n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, 
      n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, 
      n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, 
      n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, 
      n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, 
      n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, 
      n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, 
      n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, 
      n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, 
      n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, 
      n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, 
      n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, 
      n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, 
      n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, 
      n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, 
      n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, 
      n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, 
      n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, 
      n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, 
      n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, 
      n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, 
      n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, 
      n_1575 : std_logic;

begin
   
   OUT1_reg_17_inst : DFF_X1 port map( D => N457, CK => CLK, Q => OUT1(17), QN 
                           => n_1000);
   OUT1_reg_16_inst : DFF_X1 port map( D => N456, CK => CLK, Q => OUT1(16), QN 
                           => n_1001);
   OUT1_reg_15_inst : DFF_X1 port map( D => N455, CK => CLK, Q => OUT1(15), QN 
                           => n_1002);
   OUT1_reg_14_inst : DFF_X1 port map( D => N454, CK => CLK, Q => OUT1(14), QN 
                           => n_1003);
   OUT1_reg_13_inst : DFF_X1 port map( D => N453, CK => CLK, Q => OUT1(13), QN 
                           => n_1004);
   OUT1_reg_12_inst : DFF_X1 port map( D => N452, CK => CLK, Q => OUT1(12), QN 
                           => n_1005);
   OUT1_reg_11_inst : DFF_X1 port map( D => N451, CK => CLK, Q => OUT1(11), QN 
                           => n_1006);
   OUT1_reg_10_inst : DFF_X1 port map( D => N450, CK => CLK, Q => OUT1(10), QN 
                           => n_1007);
   OUT1_reg_9_inst : DFF_X1 port map( D => N449, CK => CLK, Q => OUT1(9), QN =>
                           n_1008);
   OUT1_reg_8_inst : DFF_X1 port map( D => N448, CK => CLK, Q => OUT1(8), QN =>
                           n_1009);
   OUT1_reg_7_inst : DFF_X1 port map( D => N447, CK => CLK, Q => OUT1(7), QN =>
                           n_1010);
   OUT1_reg_6_inst : DFF_X1 port map( D => N446, CK => CLK, Q => OUT1(6), QN =>
                           n_1011);
   OUT1_reg_5_inst : DFF_X1 port map( D => N445, CK => CLK, Q => OUT1(5), QN =>
                           n_1012);
   OUT1_reg_4_inst : DFF_X1 port map( D => N444, CK => CLK, Q => OUT1(4), QN =>
                           n_1013);
   OUT1_reg_3_inst : DFF_X1 port map( D => N443, CK => CLK, Q => OUT1(3), QN =>
                           n_1014);
   OUT1_reg_2_inst : DFF_X1 port map( D => N442, CK => CLK, Q => OUT1(2), QN =>
                           n_1015);
   OUT1_reg_1_inst : DFF_X1 port map( D => N441, CK => CLK, Q => OUT1(1), QN =>
                           n_1016);
   OUT1_reg_0_inst : DFF_X1 port map( D => N440, CK => CLK, Q => OUT1(0), QN =>
                           n_1017);
   OUT2_reg_13_inst : DFF_X1 port map( D => N421, CK => CLK, Q => OUT2(13), QN 
                           => n_1018);
   OUT2_reg_12_inst : DFF_X1 port map( D => N420, CK => CLK, Q => OUT2(12), QN 
                           => n_1019);
   OUT2_reg_11_inst : DFF_X1 port map( D => N419, CK => CLK, Q => OUT2(11), QN 
                           => n_1020);
   OUT2_reg_10_inst : DFF_X1 port map( D => N418, CK => CLK, Q => OUT2(10), QN 
                           => n_1021);
   OUT2_reg_9_inst : DFF_X1 port map( D => N417, CK => CLK, Q => OUT2(9), QN =>
                           n_1022);
   OUT2_reg_8_inst : DFF_X1 port map( D => N416, CK => CLK, Q => OUT2(8), QN =>
                           n_1023);
   OUT2_reg_7_inst : DFF_X1 port map( D => N415, CK => CLK, Q => OUT2(7), QN =>
                           n_1024);
   OUT2_reg_6_inst : DFF_X1 port map( D => N414, CK => CLK, Q => OUT2(6), QN =>
                           n_1025);
   OUT2_reg_5_inst : DFF_X1 port map( D => N413, CK => CLK, Q => OUT2(5), QN =>
                           n_1026);
   OUT2_reg_4_inst : DFF_X1 port map( D => N412, CK => CLK, Q => OUT2(4), QN =>
                           n_1027);
   OUT2_reg_3_inst : DFF_X1 port map( D => N411, CK => CLK, Q => OUT2(3), QN =>
                           n_1028);
   OUT2_reg_2_inst : DFF_X1 port map( D => N410, CK => CLK, Q => OUT2(2), QN =>
                           n_1029);
   OUT2_reg_1_inst : DFF_X1 port map( D => N409, CK => CLK, Q => OUT2(1), QN =>
                           n_1030);
   OUT2_reg_0_inst : DFF_X1 port map( D => N408, CK => CLK, Q => OUT2(0), QN =>
                           n_1031);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n1211, CK => CLK, Q => 
                           n_1032, QN => n6682);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n1210, CK => CLK, Q => 
                           n_1033, QN => n6683);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n1209, CK => CLK, Q => 
                           n_1034, QN => n6684);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n1208, CK => CLK, Q => 
                           n_1035, QN => n6685);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n1207, CK => CLK, Q => 
                           n_1036, QN => n6686);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n1206, CK => CLK, Q => 
                           n_1037, QN => n6687);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n1205, CK => CLK, Q => 
                           n_1038, QN => n6688);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n1204, CK => CLK, Q => 
                           n_1039, QN => n6689);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n1203, CK => CLK, Q => 
                           n_1040, QN => n6690);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n1202, CK => CLK, Q => 
                           n_1041, QN => n6691);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n1201, CK => CLK, Q => 
                           n_1042, QN => n6692);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n1200, CK => CLK, Q => 
                           n_1043, QN => n6693);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n1199, CK => CLK, Q => 
                           n_1044, QN => n6694);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n1198, CK => CLK, Q => 
                           n_1045, QN => n6695);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n1197, CK => CLK, Q => 
                           n_1046, QN => n6696);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n1196, CK => CLK, Q => 
                           n_1047, QN => n6697);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n1195, CK => CLK, Q => 
                           n_1048, QN => n6698);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n1194, CK => CLK, Q => 
                           n_1049, QN => n6699);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n1193, CK => CLK, Q => 
                           n_1050, QN => n6700);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n1192, CK => CLK, Q => 
                           n_1051, QN => n6701);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n1191, CK => CLK, Q => 
                           n_1052, QN => n6702);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n1190, CK => CLK, Q => 
                           n_1053, QN => n6703);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n1189, CK => CLK, Q => 
                           n_1054, QN => n6704);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n1188, CK => CLK, Q => 
                           n_1055, QN => n6705);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n1187, CK => CLK, Q => 
                           n_1056, QN => n6706);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n1186, CK => CLK, Q => 
                           n_1057, QN => n6707);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n1185, CK => CLK, Q => 
                           n_1058, QN => n6708);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n1184, CK => CLK, Q => 
                           n_1059, QN => n6709);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n1183, CK => CLK, Q => 
                           n_1060, QN => n6710);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n1182, CK => CLK, Q => 
                           n_1061, QN => n6711);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n1181, CK => CLK, Q => 
                           n_1062, QN => n6712);
   U7554 : NAND3_X1 port map( A1 => n7744, A2 => n7743, A3 => n8785, ZN => 
                           n8777);
   U7555 : NAND3_X1 port map( A1 => n8785, A2 => n7743, A3 => ADD_WR(2), ZN => 
                           n8787);
   U7556 : NAND3_X1 port map( A1 => n8785, A2 => n7744, A3 => ADD_WR(3), ZN => 
                           n8792);
   U7557 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n8785, A3 => ADD_WR(3), ZN
                           => n8797);
   U7558 : NAND3_X1 port map( A1 => n7744, A2 => n7743, A3 => n8806, ZN => 
                           n8802);
   U7559 : NAND3_X1 port map( A1 => ADD_WR(2), A2 => n7743, A3 => n8806, ZN => 
                           n8808);
   U7560 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n7744, A3 => n8806, ZN => 
                           n8813);
   U7561 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), A3 => n8806, ZN
                           => n8818);
   U7562 : NAND3_X1 port map( A1 => ENABLE, A2 => n10533, A3 => RD1, ZN => 
                           n8823);
   U7563 : NAND3_X1 port map( A1 => ENABLE, A2 => n10533, A3 => RD2, ZN => 
                           n8855);
   U7564 : NAND3_X1 port map( A1 => ADD_RD1(4), A2 => n7747, A3 => ADD_RD1(2), 
                           ZN => n8864);
   U7565 : NAND3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), A3 => 
                           ADD_RD1(2), ZN => n8863);
   U7566 : NAND3_X1 port map( A1 => n7748, A2 => n7747, A3 => ADD_RD1(4), ZN =>
                           n8869);
   U7567 : NAND3_X1 port map( A1 => ADD_RD1(3), A2 => n7748, A3 => ADD_RD1(4), 
                           ZN => n8868);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n1180, CK => CLK, Q => 
                           n_1063, QN => n8709);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => 
                           n_1064, QN => n8453);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => 
                           n_1065, QN => n8454);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => 
                           n_1066, QN => n8455);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => 
                           n_1067, QN => n8456);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => 
                           n_1068, QN => n8457);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => 
                           n_1069, QN => n8458);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => 
                           n_1070, QN => n8459);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => 
                           n_1071, QN => n8460);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => 
                           n_1072, QN => n8421);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => 
                           n_1073, QN => n8422);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => 
                           n_1074, QN => n8423);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => 
                           n_1075, QN => n8424);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => 
                           n_1076, QN => n8425);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => 
                           n_1077, QN => n8426);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => 
                           n_1078, QN => n8427);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => 
                           n_1079, QN => n8428);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => 
                           n_1080, QN => n8389);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => 
                           n_1081, QN => n8390);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => 
                           n_1082, QN => n8391);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => 
                           n_1083, QN => n8392);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => 
                           n_1084, QN => n8393);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => 
                           n_1085, QN => n8394);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => 
                           n_1086, QN => n8395);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => 
                           n_1087, QN => n8396);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => 
                           n_1088, QN => n8357);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => 
                           n_1089, QN => n8358);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => 
                           n_1090, QN => n8359);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => 
                           n_1091, QN => n8360);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => 
                           n_1092, QN => n8361);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => 
                           n_1093, QN => n8362);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => 
                           n_1094, QN => n8363);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => 
                           n_1095, QN => n8364);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => 
                           n_1096, QN => n8325);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => 
                           n_1097, QN => n8326);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => 
                           n_1098, QN => n8327);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => 
                           n_1099, QN => n8328);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => 
                           n_1100, QN => n8329);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => 
                           n_1101, QN => n8330);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => 
                           n_1102, QN => n8331);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => 
                           n_1103, QN => n8332);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => 
                           n_1104, QN => n8293);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => 
                           n_1105, QN => n8294);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => 
                           n_1106, QN => n8295);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => 
                           n_1107, QN => n8296);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => 
                           n_1108, QN => n8297);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => 
                           n_1109, QN => n8298);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => 
                           n_1110, QN => n8299);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => 
                           n_1111, QN => n8300);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => 
                           n_1112, QN => n8261);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => 
                           n_1113, QN => n8262);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => 
                           n_1114, QN => n8263);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => 
                           n_1115, QN => n8264);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => 
                           n_1116, QN => n8265);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => 
                           n_1117, QN => n8266);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => 
                           n_1118, QN => n8267);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => 
                           n_1119, QN => n8268);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => 
                           n_1120, QN => n8229);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => 
                           n_1121, QN => n8230);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => 
                           n_1122, QN => n8231);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => 
                           n_1123, QN => n8232);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => 
                           n_1124, QN => n8233);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => 
                           n_1125, QN => n8234);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => 
                           n_1126, QN => n8235);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => 
                           n_1127, QN => n8236);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n1243, CK => CLK, Q => 
                           n_1128, QN => n8677);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n1242, CK => CLK, Q => 
                           n_1129, QN => n8678);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n1241, CK => CLK, Q => 
                           n_1130, QN => n8679);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n1240, CK => CLK, Q => 
                           n_1131, QN => n8680);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n1239, CK => CLK, Q => 
                           n_1132, QN => n8681);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n1238, CK => CLK, Q => 
                           n_1133, QN => n8682);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n1237, CK => CLK, Q => 
                           n_1134, QN => n8683);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n1236, CK => CLK, Q => 
                           n_1135, QN => n8684);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n1275, CK => CLK, Q => 
                           n_1136, QN => n8645);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n1274, CK => CLK, Q => 
                           n_1137, QN => n8646);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n1273, CK => CLK, Q => 
                           n_1138, QN => n8647);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n1272, CK => CLK, Q => 
                           n_1139, QN => n8648);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n1271, CK => CLK, Q => 
                           n_1140, QN => n8649);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n1270, CK => CLK, Q => 
                           n_1141, QN => n8650);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n1269, CK => CLK, Q => 
                           n_1142, QN => n8651);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n1268, CK => CLK, Q => 
                           n_1143, QN => n8652);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n1307, CK => CLK, Q => 
                           n_1144, QN => n8613);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n1306, CK => CLK, Q => 
                           n_1145, QN => n8614);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n1305, CK => CLK, Q => 
                           n_1146, QN => n8615);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n1304, CK => CLK, Q => 
                           n_1147, QN => n8616);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n1303, CK => CLK, Q => 
                           n_1148, QN => n8617);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n1302, CK => CLK, Q => 
                           n_1149, QN => n8618);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n1301, CK => CLK, Q => 
                           n_1150, QN => n8619);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n1300, CK => CLK, Q => 
                           n_1151, QN => n8620);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => 
                           n_1152, QN => n8581);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => 
                           n_1153, QN => n8582);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => 
                           n_1154, QN => n8583);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => 
                           n_1155, QN => n8584);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => 
                           n_1156, QN => n8585);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => 
                           n_1157, QN => n8586);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => 
                           n_1158, QN => n8587);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => 
                           n_1159, QN => n8588);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => 
                           n_1160, QN => n8549);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => 
                           n_1161, QN => n8550);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => 
                           n_1162, QN => n8551);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => 
                           n_1163, QN => n8552);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => 
                           n_1164, QN => n8553);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => 
                           n_1165, QN => n8554);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => 
                           n_1166, QN => n8555);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => 
                           n_1167, QN => n8556);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => 
                           n_1168, QN => n8517);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => 
                           n_1169, QN => n8518);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => 
                           n_1170, QN => n8519);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => 
                           n_1171, QN => n8520);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => 
                           n_1172, QN => n8521);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => 
                           n_1173, QN => n8522);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => 
                           n_1174, QN => n8523);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => 
                           n_1175, QN => n8524);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => 
                           n_1176, QN => n8485);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => 
                           n_1177, QN => n8486);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => 
                           n_1178, QN => n8487);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => 
                           n_1179, QN => n8488);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => 
                           n_1180, QN => n8489);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => 
                           n_1181, QN => n8490);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => 
                           n_1182, QN => n8491);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => 
                           n_1183, QN => n8492);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => 
                           n_1184, QN => n8461);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => 
                           n_1185, QN => n8462);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => 
                           n_1186, QN => n8463);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => 
                           n_1187, QN => n8464);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => 
                           n_1188, QN => n8465);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => 
                           n_1189, QN => n8466);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => 
                           n_1190, QN => n8467);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => 
                           n_1191, QN => n8468);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => 
                           n_1192, QN => n8469);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => 
                           n_1193, QN => n8470);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => 
                           n_1194, QN => n8471);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => 
                           n_1195, QN => n8472);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => 
                           n_1196, QN => n8473);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => 
                           n_1197, QN => n8474);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => 
                           n_1198, QN => n8475);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => 
                           n_1199, QN => n8476);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => 
                           n_1200, QN => n8477);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => 
                           n_1201, QN => n8478);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => 
                           n_1202, QN => n8479);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => 
                           n_1203, QN => n8480);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => 
                           n_1204, QN => n8481);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => 
                           n_1205, QN => n8482);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => 
                           n_1206, QN => n8483);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => 
                           n_1207, QN => n8484);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => 
                           n_1208, QN => n8429);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => 
                           n_1209, QN => n8430);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => 
                           n_1210, QN => n8431);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => 
                           n_1211, QN => n8432);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => 
                           n_1212, QN => n8433);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => 
                           n_1213, QN => n8434);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => 
                           n_1214, QN => n8435);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => 
                           n_1215, QN => n8436);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => 
                           n_1216, QN => n8437);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => 
                           n_1217, QN => n8438);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => 
                           n_1218, QN => n8439);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => 
                           n_1219, QN => n8440);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => 
                           n_1220, QN => n8441);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => 
                           n_1221, QN => n8442);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => 
                           n_1222, QN => n8443);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => 
                           n_1223, QN => n8444);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => 
                           n_1224, QN => n8445);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => 
                           n_1225, QN => n8446);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => 
                           n_1226, QN => n8447);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => 
                           n_1227, QN => n8448);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => 
                           n_1228, QN => n8449);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => 
                           n_1229, QN => n8450);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => 
                           n_1230, QN => n8451);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => 
                           n_1231, QN => n8452);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => 
                           n_1232, QN => n8397);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => 
                           n_1233, QN => n8398);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => 
                           n_1234, QN => n8399);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => 
                           n_1235, QN => n8400);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => 
                           n_1236, QN => n8401);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => 
                           n_1237, QN => n8402);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => 
                           n_1238, QN => n8403);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => 
                           n_1239, QN => n8404);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => 
                           n_1240, QN => n8405);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => 
                           n_1241, QN => n8406);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => 
                           n_1242, QN => n8407);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => 
                           n_1243, QN => n8408);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => 
                           n_1244, QN => n8409);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => 
                           n_1245, QN => n8410);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => 
                           n_1246, QN => n8411);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => 
                           n_1247, QN => n8412);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => 
                           n_1248, QN => n8413);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => 
                           n_1249, QN => n8414);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => 
                           n_1250, QN => n8415);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => 
                           n_1251, QN => n8416);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => 
                           n_1252, QN => n8417);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => 
                           n_1253, QN => n8418);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => 
                           n_1254, QN => n8419);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => 
                           n_1255, QN => n8420);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => 
                           n_1256, QN => n8365);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => 
                           n_1257, QN => n8366);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => 
                           n_1258, QN => n8367);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => 
                           n_1259, QN => n8368);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => 
                           n_1260, QN => n8369);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => 
                           n_1261, QN => n8370);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => 
                           n_1262, QN => n8371);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => 
                           n_1263, QN => n8372);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => 
                           n_1264, QN => n8373);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => 
                           n_1265, QN => n8374);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => 
                           n_1266, QN => n8375);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => 
                           n_1267, QN => n8376);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => 
                           n_1268, QN => n8377);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => 
                           n_1269, QN => n8378);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => 
                           n_1270, QN => n8379);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => 
                           n_1271, QN => n8380);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => 
                           n_1272, QN => n8381);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => 
                           n_1273, QN => n8382);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => 
                           n_1274, QN => n8383);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => 
                           n_1275, QN => n8384);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => 
                           n_1276, QN => n8385);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => 
                           n_1277, QN => n8386);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => 
                           n_1278, QN => n8387);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => 
                           n_1279, QN => n8388);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => 
                           n_1280, QN => n8333);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => 
                           n_1281, QN => n8334);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => 
                           n_1282, QN => n8335);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => 
                           n_1283, QN => n8336);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => 
                           n_1284, QN => n8337);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => 
                           n_1285, QN => n8338);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => 
                           n_1286, QN => n8339);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => 
                           n_1287, QN => n8340);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => 
                           n_1288, QN => n8341);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => 
                           n_1289, QN => n8342);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => 
                           n_1290, QN => n8343);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => 
                           n_1291, QN => n8344);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => 
                           n_1292, QN => n8345);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => 
                           n_1293, QN => n8346);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => 
                           n_1294, QN => n8347);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => 
                           n_1295, QN => n8348);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => 
                           n_1296, QN => n8349);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => 
                           n_1297, QN => n8350);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => 
                           n_1298, QN => n8351);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => 
                           n_1299, QN => n8352);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => 
                           n_1300, QN => n8353);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => 
                           n_1301, QN => n8354);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => 
                           n_1302, QN => n8355);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => 
                           n_1303, QN => n8356);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => 
                           n_1304, QN => n8301);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => 
                           n_1305, QN => n8302);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => 
                           n_1306, QN => n8303);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => 
                           n_1307, QN => n8304);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => 
                           n_1308, QN => n8305);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => 
                           n_1309, QN => n8306);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => 
                           n_1310, QN => n8307);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => 
                           n_1311, QN => n8308);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => 
                           n_1312, QN => n8309);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => 
                           n_1313, QN => n8310);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => 
                           n_1314, QN => n8311);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => 
                           n_1315, QN => n8312);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => 
                           n_1316, QN => n8313);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => 
                           n_1317, QN => n8314);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => 
                           n_1318, QN => n8315);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => 
                           n_1319, QN => n8316);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => 
                           n_1320, QN => n8317);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => 
                           n_1321, QN => n8318);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => 
                           n_1322, QN => n8319);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => 
                           n_1323, QN => n8320);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => 
                           n_1324, QN => n8321);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => 
                           n_1325, QN => n8322);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => 
                           n_1326, QN => n8323);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => 
                           n_1327, QN => n8324);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => 
                           n_1328, QN => n8269);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => 
                           n_1329, QN => n8270);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => 
                           n_1330, QN => n8271);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => 
                           n_1331, QN => n8272);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => 
                           n_1332, QN => n8273);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => 
                           n_1333, QN => n8274);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => 
                           n_1334, QN => n8275);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => 
                           n_1335, QN => n8276);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => 
                           n_1336, QN => n8277);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => 
                           n_1337, QN => n8278);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => 
                           n_1338, QN => n8279);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => 
                           n_1339, QN => n8280);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => 
                           n_1340, QN => n8281);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => 
                           n_1341, QN => n8282);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => 
                           n_1342, QN => n8283);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => 
                           n_1343, QN => n8284);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => 
                           n_1344, QN => n8285);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => 
                           n_1345, QN => n8286);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => 
                           n_1346, QN => n8287);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => 
                           n_1347, QN => n8288);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => 
                           n_1348, QN => n8289);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => 
                           n_1349, QN => n8290);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => 
                           n_1350, QN => n8291);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => 
                           n_1351, QN => n8292);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => 
                           n_1352, QN => n8237);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => 
                           n_1353, QN => n8238);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => 
                           n_1354, QN => n8239);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => 
                           n_1355, QN => n8240);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => 
                           n_1356, QN => n8241);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => 
                           n_1357, QN => n8242);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => 
                           n_1358, QN => n8243);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => 
                           n_1359, QN => n8244);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => 
                           n_1360, QN => n8245);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => 
                           n_1361, QN => n8246);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => 
                           n_1362, QN => n8247);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => 
                           n_1363, QN => n8248);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => 
                           n_1364, QN => n8249);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => 
                           n_1365, QN => n8250);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => 
                           n_1366, QN => n8251);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => 
                           n_1367, QN => n8252);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => 
                           n_1368, QN => n8253);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => 
                           n_1369, QN => n8254);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => 
                           n_1370, QN => n8255);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => 
                           n_1371, QN => n8256);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => 
                           n_1372, QN => n8257);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => 
                           n_1373, QN => n8258);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => 
                           n_1374, QN => n8259);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => 
                           n_1375, QN => n8260);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n1235, CK => CLK, Q => 
                           n_1376, QN => n8685);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n1234, CK => CLK, Q => 
                           n_1377, QN => n8686);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n1233, CK => CLK, Q => 
                           n_1378, QN => n8687);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n1232, CK => CLK, Q => 
                           n_1379, QN => n8688);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n1231, CK => CLK, Q => 
                           n_1380, QN => n8689);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n1230, CK => CLK, Q => 
                           n_1381, QN => n8690);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n1229, CK => CLK, Q => 
                           n_1382, QN => n8691);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n1228, CK => CLK, Q => 
                           n_1383, QN => n8692);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n1227, CK => CLK, Q => 
                           n_1384, QN => n8693);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n1226, CK => CLK, Q => 
                           n_1385, QN => n8694);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n1225, CK => CLK, Q => 
                           n_1386, QN => n8695);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n1224, CK => CLK, Q => 
                           n_1387, QN => n8696);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n1223, CK => CLK, Q => 
                           n_1388, QN => n8697);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n1222, CK => CLK, Q => 
                           n_1389, QN => n8698);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n1221, CK => CLK, Q => 
                           n_1390, QN => n8699);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n1220, CK => CLK, Q => 
                           n_1391, QN => n8700);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n1219, CK => CLK, Q => 
                           n_1392, QN => n8701);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n1218, CK => CLK, Q => 
                           n_1393, QN => n8702);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n1217, CK => CLK, Q => 
                           n_1394, QN => n8703);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n1216, CK => CLK, Q => 
                           n_1395, QN => n8704);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n1215, CK => CLK, Q => 
                           n_1396, QN => n8705);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n1214, CK => CLK, Q => 
                           n_1397, QN => n8706);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n1213, CK => CLK, Q => 
                           n_1398, QN => n8707);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n1212, CK => CLK, Q => 
                           n_1399, QN => n8708);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n1267, CK => CLK, Q => 
                           n_1400, QN => n8653);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n1266, CK => CLK, Q => 
                           n_1401, QN => n8654);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n1265, CK => CLK, Q => 
                           n_1402, QN => n8655);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n1264, CK => CLK, Q => 
                           n_1403, QN => n8656);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n1263, CK => CLK, Q => 
                           n_1404, QN => n8657);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n1262, CK => CLK, Q => 
                           n_1405, QN => n8658);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n1261, CK => CLK, Q => 
                           n_1406, QN => n8659);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n1260, CK => CLK, Q => 
                           n_1407, QN => n8660);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n1259, CK => CLK, Q => 
                           n_1408, QN => n8661);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n1258, CK => CLK, Q => 
                           n_1409, QN => n8662);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n1257, CK => CLK, Q => 
                           n_1410, QN => n8663);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n1256, CK => CLK, Q => 
                           n_1411, QN => n8664);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n1255, CK => CLK, Q => 
                           n_1412, QN => n8665);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n1254, CK => CLK, Q => 
                           n_1413, QN => n8666);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n1253, CK => CLK, Q => 
                           n_1414, QN => n8667);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n1252, CK => CLK, Q => 
                           n_1415, QN => n8668);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n1251, CK => CLK, Q => 
                           n_1416, QN => n8669);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n1250, CK => CLK, Q => 
                           n_1417, QN => n8670);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n1249, CK => CLK, Q => 
                           n_1418, QN => n8671);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n1248, CK => CLK, Q => 
                           n_1419, QN => n8672);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n1247, CK => CLK, Q => 
                           n_1420, QN => n8673);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n1246, CK => CLK, Q => 
                           n_1421, QN => n8674);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n1245, CK => CLK, Q => 
                           n_1422, QN => n8675);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n1244, CK => CLK, Q => 
                           n_1423, QN => n8676);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n1299, CK => CLK, Q => 
                           n_1424, QN => n8621);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n1298, CK => CLK, Q => 
                           n_1425, QN => n8622);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n1297, CK => CLK, Q => 
                           n_1426, QN => n8623);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n1296, CK => CLK, Q => 
                           n_1427, QN => n8624);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n1295, CK => CLK, Q => 
                           n_1428, QN => n8625);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n1294, CK => CLK, Q => 
                           n_1429, QN => n8626);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n1293, CK => CLK, Q => 
                           n_1430, QN => n8627);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n1292, CK => CLK, Q => 
                           n_1431, QN => n8628);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n1291, CK => CLK, Q => 
                           n_1432, QN => n8629);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n1290, CK => CLK, Q => 
                           n_1433, QN => n8630);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n1289, CK => CLK, Q => 
                           n_1434, QN => n8631);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n1288, CK => CLK, Q => 
                           n_1435, QN => n8632);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n1287, CK => CLK, Q => 
                           n_1436, QN => n8633);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n1286, CK => CLK, Q => 
                           n_1437, QN => n8634);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n1285, CK => CLK, Q => 
                           n_1438, QN => n8635);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n1284, CK => CLK, Q => 
                           n_1439, QN => n8636);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n1283, CK => CLK, Q => 
                           n_1440, QN => n8637);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n1282, CK => CLK, Q => 
                           n_1441, QN => n8638);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n1281, CK => CLK, Q => 
                           n_1442, QN => n8639);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n1280, CK => CLK, Q => 
                           n_1443, QN => n8640);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n1279, CK => CLK, Q => 
                           n_1444, QN => n8641);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n1278, CK => CLK, Q => 
                           n_1445, QN => n8642);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n1277, CK => CLK, Q => 
                           n_1446, QN => n8643);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n1276, CK => CLK, Q => 
                           n_1447, QN => n8644);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => 
                           n_1448, QN => n8589);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => 
                           n_1449, QN => n8590);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => 
                           n_1450, QN => n8591);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => 
                           n_1451, QN => n8592);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => 
                           n_1452, QN => n8593);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => 
                           n_1453, QN => n8594);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => 
                           n_1454, QN => n8595);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => 
                           n_1455, QN => n8596);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => 
                           n_1456, QN => n8597);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => 
                           n_1457, QN => n8598);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => 
                           n_1458, QN => n8599);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => 
                           n_1459, QN => n8600);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => 
                           n_1460, QN => n8601);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => 
                           n_1461, QN => n8602);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => 
                           n_1462, QN => n8603);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => 
                           n_1463, QN => n8604);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => 
                           n_1464, QN => n8605);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => 
                           n_1465, QN => n8606);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => 
                           n_1466, QN => n8607);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => 
                           n_1467, QN => n8608);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => 
                           n_1468, QN => n8609);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => 
                           n_1469, QN => n8610);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n1309, CK => CLK, Q => 
                           n_1470, QN => n8611);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n1308, CK => CLK, Q => 
                           n_1471, QN => n8612);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => 
                           n_1472, QN => n8557);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => 
                           n_1473, QN => n8558);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => 
                           n_1474, QN => n8559);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => 
                           n_1475, QN => n8560);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => 
                           n_1476, QN => n8561);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => 
                           n_1477, QN => n8562);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => 
                           n_1478, QN => n8563);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => 
                           n_1479, QN => n8564);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => 
                           n_1480, QN => n8565);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => 
                           n_1481, QN => n8566);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => 
                           n_1482, QN => n8567);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => 
                           n_1483, QN => n8568);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => 
                           n_1484, QN => n8569);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => 
                           n_1485, QN => n8570);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => 
                           n_1486, QN => n8571);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => 
                           n_1487, QN => n8572);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => 
                           n_1488, QN => n8573);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => 
                           n_1489, QN => n8574);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => 
                           n_1490, QN => n8575);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => 
                           n_1491, QN => n8576);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => 
                           n_1492, QN => n8577);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => 
                           n_1493, QN => n8578);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => 
                           n_1494, QN => n8579);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => 
                           n_1495, QN => n8580);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => 
                           n_1496, QN => n8525);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => 
                           n_1497, QN => n8526);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => 
                           n_1498, QN => n8527);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => 
                           n_1499, QN => n8528);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => 
                           n_1500, QN => n8529);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => 
                           n_1501, QN => n8530);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => 
                           n_1502, QN => n8531);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => 
                           n_1503, QN => n8532);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => 
                           n_1504, QN => n8533);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => 
                           n_1505, QN => n8534);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => 
                           n_1506, QN => n8535);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => 
                           n_1507, QN => n8536);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => 
                           n_1508, QN => n8537);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => 
                           n_1509, QN => n8538);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => 
                           n_1510, QN => n8539);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => 
                           n_1511, QN => n8540);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => 
                           n_1512, QN => n8541);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => 
                           n_1513, QN => n8542);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => 
                           n_1514, QN => n8543);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => 
                           n_1515, QN => n8544);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => 
                           n_1516, QN => n8545);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => 
                           n_1517, QN => n8546);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => 
                           n_1518, QN => n8547);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => 
                           n_1519, QN => n8548);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => 
                           n_1520, QN => n8493);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => 
                           n_1521, QN => n8494);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => 
                           n_1522, QN => n8495);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => 
                           n_1523, QN => n8496);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => 
                           n_1524, QN => n8497);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => 
                           n_1525, QN => n8498);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => 
                           n_1526, QN => n8499);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => 
                           n_1527, QN => n8500);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => 
                           n_1528, QN => n8501);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => 
                           n_1529, QN => n8502);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => 
                           n_1530, QN => n8503);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => 
                           n_1531, QN => n8504);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => 
                           n_1532, QN => n8505);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => 
                           n_1533, QN => n8506);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => 
                           n_1534, QN => n8507);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => 
                           n_1535, QN => n8508);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => 
                           n_1536, QN => n8509);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => 
                           n_1537, QN => n8510);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => 
                           n_1538, QN => n8511);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => 
                           n_1539, QN => n8512);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => 
                           n_1540, QN => n8513);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => 
                           n_1541, QN => n8514);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => 
                           n_1542, QN => n8515);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => 
                           n_1543, QN => n8516);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n1979, CK => CLK, Q => n9567
                           , QN => n7975);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n1978, CK => CLK, Q => n9566
                           , QN => n7976);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n1977, CK => CLK, Q => n9565
                           , QN => n7977);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n1976, CK => CLK, Q => n9564
                           , QN => n7978);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n1975, CK => CLK, Q => n9563
                           , QN => n7979);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n1974, CK => CLK, Q => n9562
                           , QN => n7980);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n1973, CK => CLK, Q => n9561
                           , QN => n7981);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n1972, CK => CLK, Q => n9560
                           , QN => n7982);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n2011, CK => CLK, Q => n9575
                           , QN => n7943);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n2010, CK => CLK, Q => n9574
                           , QN => n7944);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n2009, CK => CLK, Q => n9573
                           , QN => n7945);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n2008, CK => CLK, Q => n9572
                           , QN => n7946);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n2007, CK => CLK, Q => n9571
                           , QN => n7947);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n2006, CK => CLK, Q => n9570
                           , QN => n7948);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n2005, CK => CLK, Q => n9569
                           , QN => n7949);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n2004, CK => CLK, Q => n9568
                           , QN => n7950);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n2043, CK => CLK, Q => n9583
                           , QN => n7911);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n2042, CK => CLK, Q => n9582
                           , QN => n7912);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n2041, CK => CLK, Q => n9581
                           , QN => n7913);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n2040, CK => CLK, Q => n9580
                           , QN => n7914);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n2039, CK => CLK, Q => n9579
                           , QN => n7915);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n2038, CK => CLK, Q => n9578
                           , QN => n7916);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n2037, CK => CLK, Q => n9577
                           , QN => n7917);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n2036, CK => CLK, Q => n9576
                           , QN => n7918);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n2075, CK => CLK, Q => n9585
                           , QN => n7879);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n2074, CK => CLK, Q => n9584
                           , QN => n7880);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n2073, CK => CLK, Q => 
                           n10019, QN => n7881);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n2072, CK => CLK, Q => 
                           n10015, QN => n7882);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n2071, CK => CLK, Q => 
                           n10011, QN => n7883);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n2070, CK => CLK, Q => 
                           n10007, QN => n7884);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n2069, CK => CLK, Q => 
                           n10003, QN => n7885);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n2068, CK => CLK, Q => n9999
                           , QN => n7886);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n2107, CK => CLK, Q => n9593
                           , QN => n7847);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n2106, CK => CLK, Q => n9592
                           , QN => n7848);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n2105, CK => CLK, Q => n9591
                           , QN => n7849);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n2104, CK => CLK, Q => n9590
                           , QN => n7850);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n2103, CK => CLK, Q => n9589
                           , QN => n7851);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n2102, CK => CLK, Q => n9588
                           , QN => n7852);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n2101, CK => CLK, Q => n9587
                           , QN => n7853);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n2100, CK => CLK, Q => n9586
                           , QN => n7854);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n2139, CK => CLK, Q => n9601
                           , QN => n7815);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n2138, CK => CLK, Q => n9600
                           , QN => n7816);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n2137, CK => CLK, Q => n9599
                           , QN => n7817);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n2136, CK => CLK, Q => n9598
                           , QN => n7818);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n2135, CK => CLK, Q => n9597
                           , QN => n7819);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n2134, CK => CLK, Q => n9596
                           , QN => n7820);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n2133, CK => CLK, Q => n9595
                           , QN => n7821);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n2132, CK => CLK, Q => n9594
                           , QN => n7822);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n2171, CK => CLK, Q => n9609
                           , QN => n7783);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n2170, CK => CLK, Q => n9608
                           , QN => n7784);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n2169, CK => CLK, Q => n9607
                           , QN => n7785);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n2168, CK => CLK, Q => n9606
                           , QN => n7786);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n2167, CK => CLK, Q => n9605
                           , QN => n7787);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n2166, CK => CLK, Q => n9604
                           , QN => n7788);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n2165, CK => CLK, Q => n9603
                           , QN => n7789);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n2164, CK => CLK, Q => n9602
                           , QN => n7790);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n2203, CK => CLK, Q => n9611
                           , QN => n7751);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n2202, CK => CLK, Q => n9610
                           , QN => n7752);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n2201, CK => CLK, Q => 
                           n10017, QN => n7753);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n2200, CK => CLK, Q => 
                           n10013, QN => n7754);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n2199, CK => CLK, Q => 
                           n10009, QN => n7755);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n2198, CK => CLK, Q => 
                           n10005, QN => n7756);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n2197, CK => CLK, Q => 
                           n10001, QN => n7757);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n2196, CK => CLK, Q => n9997
                           , QN => n7758);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n1723, CK => CLK, Q => 
                           n9515, QN => n8710);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n1722, CK => CLK, Q => 
                           n9514, QN => n8711);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n1721, CK => CLK, Q => 
                           n9513, QN => n8712);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n1720, CK => CLK, Q => 
                           n9512, QN => n8713);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n1719, CK => CLK, Q => 
                           n9511, QN => n8714);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n1718, CK => CLK, Q => 
                           n9510, QN => n8715);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n1717, CK => CLK, Q => 
                           n9509, QN => n8716);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n1716, CK => CLK, Q => 
                           n9508, QN => n8717);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n1755, CK => CLK, Q => 
                           n9523, QN => n8718);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n1754, CK => CLK, Q => 
                           n9522, QN => n8719);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n1753, CK => CLK, Q => 
                           n9521, QN => n8720);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n1752, CK => CLK, Q => 
                           n9520, QN => n8721);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n1751, CK => CLK, Q => 
                           n9519, QN => n8722);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n1750, CK => CLK, Q => 
                           n9518, QN => n8723);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n1749, CK => CLK, Q => 
                           n9517, QN => n8724);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n1748, CK => CLK, Q => 
                           n9516, QN => n8725);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n1787, CK => CLK, Q => 
                           n9531, QN => n8726);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n1786, CK => CLK, Q => 
                           n9530, QN => n8727);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n1785, CK => CLK, Q => 
                           n9529, QN => n8728);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n1784, CK => CLK, Q => 
                           n9528, QN => n8729);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n1783, CK => CLK, Q => 
                           n9527, QN => n8730);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n1782, CK => CLK, Q => 
                           n9526, QN => n8731);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n1781, CK => CLK, Q => 
                           n9525, QN => n8732);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n1780, CK => CLK, Q => 
                           n9524, QN => n8733);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n1819, CK => CLK, Q => 
                           n9533, QN => n8734);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n1818, CK => CLK, Q => 
                           n9532, QN => n8735);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n1817, CK => CLK, Q => 
                           n10018, QN => n8736);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n1816, CK => CLK, Q => 
                           n10014, QN => n8737);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n1815, CK => CLK, Q => 
                           n10010, QN => n8738);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n1814, CK => CLK, Q => 
                           n10006, QN => n8739);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n1813, CK => CLK, Q => 
                           n10002, QN => n8740);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n1812, CK => CLK, Q => 
                           n9998, QN => n8741);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n1851, CK => CLK, Q => 
                           n9541, QN => n8742);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n1850, CK => CLK, Q => 
                           n9540, QN => n8743);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n1849, CK => CLK, Q => 
                           n9539, QN => n8103);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n1848, CK => CLK, Q => 
                           n9538, QN => n8104);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n1847, CK => CLK, Q => 
                           n9537, QN => n8105);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n1846, CK => CLK, Q => 
                           n9536, QN => n8106);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n1845, CK => CLK, Q => 
                           n9535, QN => n8107);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n1844, CK => CLK, Q => 
                           n9534, QN => n8108);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n1883, CK => CLK, Q => 
                           n9549, QN => n8071);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n1882, CK => CLK, Q => 
                           n9548, QN => n8072);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n1881, CK => CLK, Q => 
                           n9547, QN => n8073);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n1880, CK => CLK, Q => 
                           n9546, QN => n8074);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n1879, CK => CLK, Q => 
                           n9545, QN => n8075);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n1878, CK => CLK, Q => 
                           n9544, QN => n8076);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n1877, CK => CLK, Q => 
                           n9543, QN => n8077);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n1876, CK => CLK, Q => 
                           n9542, QN => n8078);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n1915, CK => CLK, Q => n9557
                           , QN => n8039);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n1914, CK => CLK, Q => n9556
                           , QN => n8040);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n1913, CK => CLK, Q => n9555
                           , QN => n8041);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n1912, CK => CLK, Q => n9554
                           , QN => n8042);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n1911, CK => CLK, Q => n9553
                           , QN => n8043);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n1910, CK => CLK, Q => n9552
                           , QN => n8044);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n1909, CK => CLK, Q => n9551
                           , QN => n8045);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n1908, CK => CLK, Q => n9550
                           , QN => n8046);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n1947, CK => CLK, Q => n9559
                           , QN => n8007);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n1946, CK => CLK, Q => n9558
                           , QN => n8008);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n1945, CK => CLK, Q => 
                           n10016, QN => n8009);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n1944, CK => CLK, Q => 
                           n10012, QN => n8010);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n1943, CK => CLK, Q => 
                           n10008, QN => n8011);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n1942, CK => CLK, Q => 
                           n10004, QN => n8012);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n1941, CK => CLK, Q => 
                           n10000, QN => n8013);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n1940, CK => CLK, Q => n9996
                           , QN => n8014);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n1971, CK => CLK, Q => n9779
                           , QN => n7983);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n1970, CK => CLK, Q => n9778
                           , QN => n7984);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n1969, CK => CLK, Q => n9777
                           , QN => n7985);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n1968, CK => CLK, Q => n9776
                           , QN => n7986);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n1967, CK => CLK, Q => n9775
                           , QN => n7987);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n1966, CK => CLK, Q => n9774
                           , QN => n7988);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n1965, CK => CLK, Q => n9773
                           , QN => n7989);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n1964, CK => CLK, Q => n9772
                           , QN => n7990);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n1963, CK => CLK, Q => n9771
                           , QN => n7991);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n1962, CK => CLK, Q => n9770
                           , QN => n7992);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n1961, CK => CLK, Q => n9769
                           , QN => n7993);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n1960, CK => CLK, Q => n9768
                           , QN => n7994);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n1959, CK => CLK, Q => n9767
                           , QN => n7995);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n1958, CK => CLK, Q => n9766
                           , QN => n7996);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n1957, CK => CLK, Q => n9765,
                           QN => n7997);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n1956, CK => CLK, Q => n9764,
                           QN => n7998);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n1955, CK => CLK, Q => n9763,
                           QN => n7999);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n1954, CK => CLK, Q => n9762,
                           QN => n8000);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n1953, CK => CLK, Q => n9761,
                           QN => n8001);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n1952, CK => CLK, Q => n9760,
                           QN => n8002);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n1951, CK => CLK, Q => n9759,
                           QN => n8003);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n1950, CK => CLK, Q => n9758,
                           QN => n8004);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n1949, CK => CLK, Q => n9757,
                           QN => n8005);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n1948, CK => CLK, Q => n9756,
                           QN => n8006);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n2003, CK => CLK, Q => n9803
                           , QN => n7951);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n2002, CK => CLK, Q => n9802
                           , QN => n7952);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n2001, CK => CLK, Q => n9801
                           , QN => n7953);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n2000, CK => CLK, Q => n9800
                           , QN => n7954);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n1999, CK => CLK, Q => n9799
                           , QN => n7955);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n1998, CK => CLK, Q => n9798
                           , QN => n7956);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n1997, CK => CLK, Q => n9797
                           , QN => n7957);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n1996, CK => CLK, Q => n9796
                           , QN => n7958);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n1995, CK => CLK, Q => n9795
                           , QN => n7959);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n1994, CK => CLK, Q => n9794
                           , QN => n7960);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n1993, CK => CLK, Q => n9793
                           , QN => n7961);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n1992, CK => CLK, Q => n9792
                           , QN => n7962);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n1991, CK => CLK, Q => n9791
                           , QN => n7963);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n1990, CK => CLK, Q => n9790
                           , QN => n7964);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n1989, CK => CLK, Q => n9789,
                           QN => n7965);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n1988, CK => CLK, Q => n9788,
                           QN => n7966);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n1987, CK => CLK, Q => n9787,
                           QN => n7967);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n1986, CK => CLK, Q => n9786,
                           QN => n7968);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n1985, CK => CLK, Q => n9785,
                           QN => n7969);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n1984, CK => CLK, Q => n9784,
                           QN => n7970);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n1983, CK => CLK, Q => n9783,
                           QN => n7971);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n1982, CK => CLK, Q => n9782,
                           QN => n7972);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n1981, CK => CLK, Q => n9781,
                           QN => n7973);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n1980, CK => CLK, Q => n9780,
                           QN => n7974);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n2035, CK => CLK, Q => n9827
                           , QN => n7919);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n2034, CK => CLK, Q => n9826
                           , QN => n7920);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n2033, CK => CLK, Q => n9825
                           , QN => n7921);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n2032, CK => CLK, Q => n9824
                           , QN => n7922);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n2031, CK => CLK, Q => n9823
                           , QN => n7923);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n2030, CK => CLK, Q => n9822
                           , QN => n7924);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n2029, CK => CLK, Q => n9821
                           , QN => n7925);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n2028, CK => CLK, Q => n9820
                           , QN => n7926);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n2027, CK => CLK, Q => n9819
                           , QN => n7927);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n2026, CK => CLK, Q => n9818
                           , QN => n7928);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n2025, CK => CLK, Q => n9817
                           , QN => n7929);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n2024, CK => CLK, Q => n9816
                           , QN => n7930);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n2023, CK => CLK, Q => n9815
                           , QN => n7931);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n2022, CK => CLK, Q => n9814
                           , QN => n7932);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n2021, CK => CLK, Q => n9813,
                           QN => n7933);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n2020, CK => CLK, Q => n9812,
                           QN => n7934);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n2019, CK => CLK, Q => n9811,
                           QN => n7935);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n2018, CK => CLK, Q => n9810,
                           QN => n7936);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n2017, CK => CLK, Q => n9809,
                           QN => n7937);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n2016, CK => CLK, Q => n9808,
                           QN => n7938);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n2015, CK => CLK, Q => n9807,
                           QN => n7939);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n2014, CK => CLK, Q => n9806,
                           QN => n7940);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n2013, CK => CLK, Q => n9805,
                           QN => n7941);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n2012, CK => CLK, Q => n9804,
                           QN => n7942);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n2067, CK => CLK, Q => n9995
                           , QN => n7887);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n2066, CK => CLK, Q => n9991
                           , QN => n7888);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n2065, CK => CLK, Q => n9987
                           , QN => n7889);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n2064, CK => CLK, Q => n9983
                           , QN => n7890);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n2063, CK => CLK, Q => n9979
                           , QN => n7891);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n2062, CK => CLK, Q => n9975
                           , QN => n7892);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n2061, CK => CLK, Q => n9971
                           , QN => n7893);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n2060, CK => CLK, Q => n9967
                           , QN => n7894);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n2059, CK => CLK, Q => n9963
                           , QN => n7895);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n2058, CK => CLK, Q => n9959
                           , QN => n7896);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n2057, CK => CLK, Q => n9955
                           , QN => n7897);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n2056, CK => CLK, Q => n9951
                           , QN => n7898);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n2055, CK => CLK, Q => n9947
                           , QN => n7899);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n2054, CK => CLK, Q => n9943
                           , QN => n7900);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n2053, CK => CLK, Q => n9939,
                           QN => n7901);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n2052, CK => CLK, Q => n9935,
                           QN => n7902);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n2051, CK => CLK, Q => n9931,
                           QN => n7903);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n2050, CK => CLK, Q => n9927,
                           QN => n7904);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n2049, CK => CLK, Q => n9923,
                           QN => n7905);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n2048, CK => CLK, Q => n9919,
                           QN => n7906);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n2047, CK => CLK, Q => n9915,
                           QN => n7907);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n2046, CK => CLK, Q => n9911,
                           QN => n7908);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n2045, CK => CLK, Q => n9907,
                           QN => n7909);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n2044, CK => CLK, Q => n9903,
                           QN => n7910);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n2099, CK => CLK, Q => n9851
                           , QN => n7855);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n2098, CK => CLK, Q => n9850
                           , QN => n7856);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n2097, CK => CLK, Q => n9849
                           , QN => n7857);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n2096, CK => CLK, Q => n9848
                           , QN => n7858);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n2095, CK => CLK, Q => n9847
                           , QN => n7859);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n2094, CK => CLK, Q => n9846
                           , QN => n7860);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n2093, CK => CLK, Q => n9845
                           , QN => n7861);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n2092, CK => CLK, Q => n9844
                           , QN => n7862);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n2091, CK => CLK, Q => n9843
                           , QN => n7863);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n2090, CK => CLK, Q => n9842
                           , QN => n7864);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n2089, CK => CLK, Q => n9841
                           , QN => n7865);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n2088, CK => CLK, Q => n9840
                           , QN => n7866);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n2087, CK => CLK, Q => n9839
                           , QN => n7867);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n2086, CK => CLK, Q => n9838
                           , QN => n7868);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n2085, CK => CLK, Q => n9837,
                           QN => n7869);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n2084, CK => CLK, Q => n9836,
                           QN => n7870);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n2083, CK => CLK, Q => n9835,
                           QN => n7871);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n2082, CK => CLK, Q => n9834,
                           QN => n7872);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n2081, CK => CLK, Q => n9833,
                           QN => n7873);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n2080, CK => CLK, Q => n9832,
                           QN => n7874);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n2079, CK => CLK, Q => n9831,
                           QN => n7875);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n2078, CK => CLK, Q => n9830,
                           QN => n7876);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n2077, CK => CLK, Q => n9829,
                           QN => n7877);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n2076, CK => CLK, Q => n9828,
                           QN => n7878);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n2131, CK => CLK, Q => n9875
                           , QN => n7823);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n2130, CK => CLK, Q => n9874
                           , QN => n7824);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n2129, CK => CLK, Q => n9873
                           , QN => n7825);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n2128, CK => CLK, Q => n9872
                           , QN => n7826);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n2127, CK => CLK, Q => n9871
                           , QN => n7827);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n2126, CK => CLK, Q => n9870
                           , QN => n7828);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n2125, CK => CLK, Q => n9869
                           , QN => n7829);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n2124, CK => CLK, Q => n9868
                           , QN => n7830);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n2123, CK => CLK, Q => n9867
                           , QN => n7831);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n2122, CK => CLK, Q => n9866
                           , QN => n7832);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n2121, CK => CLK, Q => n9865
                           , QN => n7833);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n2120, CK => CLK, Q => n9864
                           , QN => n7834);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n2119, CK => CLK, Q => n9863
                           , QN => n7835);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n2118, CK => CLK, Q => n9862
                           , QN => n7836);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n2117, CK => CLK, Q => n9861,
                           QN => n7837);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n2116, CK => CLK, Q => n9860,
                           QN => n7838);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n2115, CK => CLK, Q => n9859,
                           QN => n7839);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n2114, CK => CLK, Q => n9858,
                           QN => n7840);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n2113, CK => CLK, Q => n9857,
                           QN => n7841);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n2112, CK => CLK, Q => n9856,
                           QN => n7842);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n2111, CK => CLK, Q => n9855,
                           QN => n7843);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n2110, CK => CLK, Q => n9854,
                           QN => n7844);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n2109, CK => CLK, Q => n9853,
                           QN => n7845);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n2108, CK => CLK, Q => n9852,
                           QN => n7846);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n2163, CK => CLK, Q => n9899
                           , QN => n7791);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n2162, CK => CLK, Q => n9898
                           , QN => n7792);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n2161, CK => CLK, Q => n9897
                           , QN => n7793);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n2160, CK => CLK, Q => n9896
                           , QN => n7794);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n2159, CK => CLK, Q => n9895
                           , QN => n7795);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n2158, CK => CLK, Q => n9894
                           , QN => n7796);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n2157, CK => CLK, Q => n9893
                           , QN => n7797);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n2156, CK => CLK, Q => n9892
                           , QN => n7798);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n2155, CK => CLK, Q => n9891
                           , QN => n7799);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n2154, CK => CLK, Q => n9890
                           , QN => n7800);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n2153, CK => CLK, Q => n9889
                           , QN => n7801);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n2152, CK => CLK, Q => n9888
                           , QN => n7802);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n2151, CK => CLK, Q => n9887
                           , QN => n7803);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n2150, CK => CLK, Q => n9886
                           , QN => n7804);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n2149, CK => CLK, Q => n9885,
                           QN => n7805);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n2148, CK => CLK, Q => n9884,
                           QN => n7806);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n2147, CK => CLK, Q => n9883,
                           QN => n7807);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n2146, CK => CLK, Q => n9882,
                           QN => n7808);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n2145, CK => CLK, Q => n9881,
                           QN => n7809);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n2144, CK => CLK, Q => n9880,
                           QN => n7810);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n2143, CK => CLK, Q => n9879,
                           QN => n7811);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n2142, CK => CLK, Q => n9878,
                           QN => n7812);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n2141, CK => CLK, Q => n9877,
                           QN => n7813);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n2140, CK => CLK, Q => n9876,
                           QN => n7814);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n2195, CK => CLK, Q => n9993
                           , QN => n7759);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n2194, CK => CLK, Q => n9989
                           , QN => n7760);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n2193, CK => CLK, Q => n9985
                           , QN => n7761);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n2192, CK => CLK, Q => n9981
                           , QN => n7762);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n2191, CK => CLK, Q => n9977
                           , QN => n7763);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n2190, CK => CLK, Q => n9973
                           , QN => n7764);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n2189, CK => CLK, Q => n9969
                           , QN => n7765);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n2188, CK => CLK, Q => n9965
                           , QN => n7766);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n2187, CK => CLK, Q => n9961
                           , QN => n7767);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n2186, CK => CLK, Q => n9957
                           , QN => n7768);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n2185, CK => CLK, Q => n9953
                           , QN => n7769);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n2184, CK => CLK, Q => n9949
                           , QN => n7770);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n2183, CK => CLK, Q => n9945
                           , QN => n7771);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n2182, CK => CLK, Q => n9941
                           , QN => n7772);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n2181, CK => CLK, Q => n9937,
                           QN => n7773);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n2180, CK => CLK, Q => n9933,
                           QN => n7774);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n2179, CK => CLK, Q => n9929,
                           QN => n7775);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n2178, CK => CLK, Q => n9925,
                           QN => n7776);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n2177, CK => CLK, Q => n9921,
                           QN => n7777);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n2176, CK => CLK, Q => n9917,
                           QN => n7778);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n2175, CK => CLK, Q => n9913,
                           QN => n7779);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n2174, CK => CLK, Q => n9909,
                           QN => n7780);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n2173, CK => CLK, Q => n9905,
                           QN => n7781);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n2172, CK => CLK, Q => n9901,
                           QN => n7782);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n1715, CK => CLK, Q => 
                           n9635, QN => n8205);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n1714, CK => CLK, Q => 
                           n9634, QN => n8206);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n1713, CK => CLK, Q => 
                           n9633, QN => n8207);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n1712, CK => CLK, Q => 
                           n9632, QN => n8208);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n1711, CK => CLK, Q => 
                           n9631, QN => n8209);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n1710, CK => CLK, Q => 
                           n9630, QN => n8210);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n1709, CK => CLK, Q => 
                           n9629, QN => n8211);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n1708, CK => CLK, Q => 
                           n9628, QN => n8212);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n1707, CK => CLK, Q => 
                           n9627, QN => n8213);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n1706, CK => CLK, Q => 
                           n9626, QN => n8214);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n1705, CK => CLK, Q => 
                           n9625, QN => n8215);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n1704, CK => CLK, Q => 
                           n9624, QN => n8216);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n1703, CK => CLK, Q => 
                           n9623, QN => n8217);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n1702, CK => CLK, Q => 
                           n9622, QN => n8218);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n1701, CK => CLK, Q => n9621
                           , QN => n8219);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n1700, CK => CLK, Q => n9620
                           , QN => n8220);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n1699, CK => CLK, Q => n9619
                           , QN => n8221);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n1698, CK => CLK, Q => n9618
                           , QN => n8222);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n1697, CK => CLK, Q => n9617
                           , QN => n8223);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n1696, CK => CLK, Q => n9616
                           , QN => n8224);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n1695, CK => CLK, Q => n9615
                           , QN => n8225);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n1694, CK => CLK, Q => n9614
                           , QN => n8226);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => n9613
                           , QN => n8227);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => n9612
                           , QN => n8228);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n1747, CK => CLK, Q => 
                           n9659, QN => n8181);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n1746, CK => CLK, Q => 
                           n9658, QN => n8182);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n1745, CK => CLK, Q => 
                           n9657, QN => n8183);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n1744, CK => CLK, Q => 
                           n9656, QN => n8184);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n1743, CK => CLK, Q => 
                           n9655, QN => n8185);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n1742, CK => CLK, Q => 
                           n9654, QN => n8186);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n1741, CK => CLK, Q => 
                           n9653, QN => n8187);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n1740, CK => CLK, Q => 
                           n9652, QN => n8188);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n1739, CK => CLK, Q => 
                           n9651, QN => n8189);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n1738, CK => CLK, Q => 
                           n9650, QN => n8190);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n1737, CK => CLK, Q => 
                           n9649, QN => n8191);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n1736, CK => CLK, Q => 
                           n9648, QN => n8192);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n1735, CK => CLK, Q => 
                           n9647, QN => n8193);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n1734, CK => CLK, Q => 
                           n9646, QN => n8194);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n1733, CK => CLK, Q => n9645
                           , QN => n8195);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n1732, CK => CLK, Q => n9644
                           , QN => n8196);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n1731, CK => CLK, Q => n9643
                           , QN => n8197);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n1730, CK => CLK, Q => n9642
                           , QN => n8198);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n1729, CK => CLK, Q => n9641
                           , QN => n8199);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n1728, CK => CLK, Q => n9640
                           , QN => n8200);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n1727, CK => CLK, Q => n9639
                           , QN => n8201);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n1726, CK => CLK, Q => n9638
                           , QN => n8202);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n1725, CK => CLK, Q => n9637
                           , QN => n8203);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n1724, CK => CLK, Q => n9636
                           , QN => n8204);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n1779, CK => CLK, Q => 
                           n9683, QN => n8157);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n1778, CK => CLK, Q => 
                           n9682, QN => n8158);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n1777, CK => CLK, Q => 
                           n9681, QN => n8159);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n1776, CK => CLK, Q => 
                           n9680, QN => n8160);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n1775, CK => CLK, Q => 
                           n9679, QN => n8161);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n1774, CK => CLK, Q => 
                           n9678, QN => n8162);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n1773, CK => CLK, Q => 
                           n9677, QN => n8163);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n1772, CK => CLK, Q => 
                           n9676, QN => n8164);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n1771, CK => CLK, Q => 
                           n9675, QN => n8165);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n1770, CK => CLK, Q => 
                           n9674, QN => n8166);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n1769, CK => CLK, Q => 
                           n9673, QN => n8167);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n1768, CK => CLK, Q => 
                           n9672, QN => n8168);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n1767, CK => CLK, Q => 
                           n9671, QN => n8169);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n1766, CK => CLK, Q => 
                           n9670, QN => n8170);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n1765, CK => CLK, Q => n9669
                           , QN => n8171);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n1764, CK => CLK, Q => n9668
                           , QN => n8172);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n1763, CK => CLK, Q => n9667
                           , QN => n8173);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n1762, CK => CLK, Q => n9666
                           , QN => n8174);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n1761, CK => CLK, Q => n9665
                           , QN => n8175);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n1760, CK => CLK, Q => n9664
                           , QN => n8176);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n1759, CK => CLK, Q => n9663
                           , QN => n8177);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n1758, CK => CLK, Q => n9662
                           , QN => n8178);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n1757, CK => CLK, Q => n9661
                           , QN => n8179);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n1756, CK => CLK, Q => n9660
                           , QN => n8180);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n1811, CK => CLK, Q => 
                           n9994, QN => n8133);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n1810, CK => CLK, Q => 
                           n9990, QN => n8134);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n1809, CK => CLK, Q => 
                           n9986, QN => n8135);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n1808, CK => CLK, Q => 
                           n9982, QN => n8136);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n1807, CK => CLK, Q => 
                           n9978, QN => n8137);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n1806, CK => CLK, Q => 
                           n9974, QN => n8138);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n1805, CK => CLK, Q => 
                           n9970, QN => n8139);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n1804, CK => CLK, Q => 
                           n9966, QN => n8140);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n1803, CK => CLK, Q => 
                           n9962, QN => n8141);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n1802, CK => CLK, Q => 
                           n9958, QN => n8142);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n1801, CK => CLK, Q => 
                           n9954, QN => n8143);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n1800, CK => CLK, Q => 
                           n9950, QN => n8144);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n1799, CK => CLK, Q => 
                           n9946, QN => n8145);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n1798, CK => CLK, Q => 
                           n9942, QN => n8146);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n1797, CK => CLK, Q => n9938
                           , QN => n8147);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n1796, CK => CLK, Q => n9934
                           , QN => n8148);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n1795, CK => CLK, Q => n9930
                           , QN => n8149);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n1794, CK => CLK, Q => n9926
                           , QN => n8150);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n1793, CK => CLK, Q => n9922
                           , QN => n8151);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n1792, CK => CLK, Q => n9918
                           , QN => n8152);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n1791, CK => CLK, Q => n9914
                           , QN => n8153);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n1790, CK => CLK, Q => n9910
                           , QN => n8154);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n1789, CK => CLK, Q => n9906
                           , QN => n8155);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n1788, CK => CLK, Q => n9902
                           , QN => n8156);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n1843, CK => CLK, Q => 
                           n9707, QN => n8109);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n1842, CK => CLK, Q => 
                           n9706, QN => n8110);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n1841, CK => CLK, Q => 
                           n9705, QN => n8111);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n1840, CK => CLK, Q => 
                           n9704, QN => n8112);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n1839, CK => CLK, Q => 
                           n9703, QN => n8113);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n1838, CK => CLK, Q => 
                           n9702, QN => n8114);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n1837, CK => CLK, Q => 
                           n9701, QN => n8115);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n1836, CK => CLK, Q => 
                           n9700, QN => n8116);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n1835, CK => CLK, Q => 
                           n9699, QN => n8117);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n1834, CK => CLK, Q => 
                           n9698, QN => n8118);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n1833, CK => CLK, Q => 
                           n9697, QN => n8119);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n1832, CK => CLK, Q => 
                           n9696, QN => n8120);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n1831, CK => CLK, Q => 
                           n9695, QN => n8121);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n1830, CK => CLK, Q => 
                           n9694, QN => n8122);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n1829, CK => CLK, Q => n9693
                           , QN => n8123);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n1828, CK => CLK, Q => n9692
                           , QN => n8124);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n1827, CK => CLK, Q => n9691
                           , QN => n8125);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n1826, CK => CLK, Q => n9690
                           , QN => n8126);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n1825, CK => CLK, Q => n9689
                           , QN => n8127);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n1824, CK => CLK, Q => n9688
                           , QN => n8128);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n1823, CK => CLK, Q => n9687
                           , QN => n8129);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n1822, CK => CLK, Q => n9686
                           , QN => n8130);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n1821, CK => CLK, Q => n9685
                           , QN => n8131);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n1820, CK => CLK, Q => n9684
                           , QN => n8132);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n1875, CK => CLK, Q => 
                           n9731, QN => n8079);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n1874, CK => CLK, Q => 
                           n9730, QN => n8080);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n1873, CK => CLK, Q => 
                           n9729, QN => n8081);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n1872, CK => CLK, Q => 
                           n9728, QN => n8082);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n1871, CK => CLK, Q => 
                           n9727, QN => n8083);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n1870, CK => CLK, Q => 
                           n9726, QN => n8084);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n1869, CK => CLK, Q => 
                           n9725, QN => n8085);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n1868, CK => CLK, Q => 
                           n9724, QN => n8086);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n1867, CK => CLK, Q => 
                           n9723, QN => n8087);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n1866, CK => CLK, Q => 
                           n9722, QN => n8088);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n1865, CK => CLK, Q => 
                           n9721, QN => n8089);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n1864, CK => CLK, Q => 
                           n9720, QN => n8090);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n1863, CK => CLK, Q => 
                           n9719, QN => n8091);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n1862, CK => CLK, Q => 
                           n9718, QN => n8092);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n1861, CK => CLK, Q => n9717
                           , QN => n8093);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n1860, CK => CLK, Q => n9716
                           , QN => n8094);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n1859, CK => CLK, Q => n9715
                           , QN => n8095);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n1858, CK => CLK, Q => n9714
                           , QN => n8096);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n1857, CK => CLK, Q => n9713
                           , QN => n8097);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n1856, CK => CLK, Q => n9712
                           , QN => n8098);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n1855, CK => CLK, Q => n9711
                           , QN => n8099);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n1854, CK => CLK, Q => n9710
                           , QN => n8100);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n1853, CK => CLK, Q => n9709
                           , QN => n8101);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n1852, CK => CLK, Q => n9708
                           , QN => n8102);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n1907, CK => CLK, Q => n9755
                           , QN => n8047);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n1906, CK => CLK, Q => n9754
                           , QN => n8048);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n1905, CK => CLK, Q => n9753
                           , QN => n8049);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n1904, CK => CLK, Q => n9752
                           , QN => n8050);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n1903, CK => CLK, Q => n9751
                           , QN => n8051);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n1902, CK => CLK, Q => n9750
                           , QN => n8052);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n1901, CK => CLK, Q => n9749
                           , QN => n8053);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n1900, CK => CLK, Q => n9748
                           , QN => n8054);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n1899, CK => CLK, Q => n9747
                           , QN => n8055);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n1898, CK => CLK, Q => n9746
                           , QN => n8056);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n1897, CK => CLK, Q => n9745
                           , QN => n8057);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n1896, CK => CLK, Q => n9744
                           , QN => n8058);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n1895, CK => CLK, Q => n9743
                           , QN => n8059);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n1894, CK => CLK, Q => n9742
                           , QN => n8060);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n1893, CK => CLK, Q => n9741,
                           QN => n8061);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n1892, CK => CLK, Q => n9740,
                           QN => n8062);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n1891, CK => CLK, Q => n9739,
                           QN => n8063);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n1890, CK => CLK, Q => n9738,
                           QN => n8064);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n1889, CK => CLK, Q => n9737,
                           QN => n8065);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n1888, CK => CLK, Q => n9736,
                           QN => n8066);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n1887, CK => CLK, Q => n9735,
                           QN => n8067);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n1886, CK => CLK, Q => n9734,
                           QN => n8068);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n1885, CK => CLK, Q => n9733,
                           QN => n8069);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n1884, CK => CLK, Q => n9732,
                           QN => n8070);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n1939, CK => CLK, Q => n9992
                           , QN => n8015);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n1938, CK => CLK, Q => n9988
                           , QN => n8016);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n1937, CK => CLK, Q => n9984
                           , QN => n8017);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n1936, CK => CLK, Q => n9980
                           , QN => n8018);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n1935, CK => CLK, Q => n9976
                           , QN => n8019);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n1934, CK => CLK, Q => n9972
                           , QN => n8020);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n1933, CK => CLK, Q => n9968
                           , QN => n8021);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n1932, CK => CLK, Q => n9964
                           , QN => n8022);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n1931, CK => CLK, Q => n9960
                           , QN => n8023);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n1930, CK => CLK, Q => n9956
                           , QN => n8024);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n1929, CK => CLK, Q => n9952
                           , QN => n8025);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n1928, CK => CLK, Q => n9948
                           , QN => n8026);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n1927, CK => CLK, Q => n9944
                           , QN => n8027);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n1926, CK => CLK, Q => n9940
                           , QN => n8028);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n1925, CK => CLK, Q => n9936,
                           QN => n8029);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n1924, CK => CLK, Q => n9932,
                           QN => n8030);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n1923, CK => CLK, Q => n9928,
                           QN => n8031);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n1922, CK => CLK, Q => n9924,
                           QN => n8032);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n1921, CK => CLK, Q => n9920,
                           QN => n8033);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n1920, CK => CLK, Q => n9916,
                           QN => n8034);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n1919, CK => CLK, Q => n9912,
                           QN => n8035);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n1918, CK => CLK, Q => n9908,
                           QN => n8036);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n1917, CK => CLK, Q => n9904,
                           QN => n8037);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n1916, CK => CLK, Q => n9900,
                           QN => n8038);
   OUT2_reg_31_inst : DFF_X1 port map( D => N439, CK => CLK, Q => OUT2(31), QN 
                           => n_1544);
   OUT2_reg_30_inst : DFF_X1 port map( D => N438, CK => CLK, Q => OUT2(30), QN 
                           => n_1545);
   OUT1_reg_31_inst : DFF_X1 port map( D => N471, CK => CLK, Q => OUT1(31), QN 
                           => n_1546);
   OUT1_reg_30_inst : DFF_X1 port map( D => N470, CK => CLK, Q => OUT1(30), QN 
                           => n_1547);
   OUT2_reg_29_inst : DFF_X1 port map( D => N437, CK => CLK, Q => OUT2(29), QN 
                           => n_1548);
   OUT2_reg_28_inst : DFF_X1 port map( D => N436, CK => CLK, Q => OUT2(28), QN 
                           => n_1549);
   OUT2_reg_27_inst : DFF_X1 port map( D => N435, CK => CLK, Q => OUT2(27), QN 
                           => n_1550);
   OUT2_reg_26_inst : DFF_X1 port map( D => N434, CK => CLK, Q => OUT2(26), QN 
                           => n_1551);
   OUT2_reg_25_inst : DFF_X1 port map( D => N433, CK => CLK, Q => OUT2(25), QN 
                           => n_1552);
   OUT2_reg_24_inst : DFF_X1 port map( D => N432, CK => CLK, Q => OUT2(24), QN 
                           => n_1553);
   OUT1_reg_29_inst : DFF_X1 port map( D => N469, CK => CLK, Q => OUT1(29), QN 
                           => n_1554);
   OUT1_reg_28_inst : DFF_X1 port map( D => N468, CK => CLK, Q => OUT1(28), QN 
                           => n_1555);
   OUT1_reg_27_inst : DFF_X1 port map( D => N467, CK => CLK, Q => OUT1(27), QN 
                           => n_1556);
   OUT1_reg_26_inst : DFF_X1 port map( D => N466, CK => CLK, Q => OUT1(26), QN 
                           => n_1557);
   OUT1_reg_25_inst : DFF_X1 port map( D => N465, CK => CLK, Q => OUT1(25), QN 
                           => n_1558);
   OUT1_reg_24_inst : DFF_X1 port map( D => N464, CK => CLK, Q => OUT1(24), QN 
                           => n_1559);
   OUT2_reg_23_inst : DFF_X1 port map( D => N431, CK => CLK, Q => OUT2(23), QN 
                           => n_1560);
   OUT2_reg_22_inst : DFF_X1 port map( D => N430, CK => CLK, Q => OUT2(22), QN 
                           => n_1561);
   OUT2_reg_21_inst : DFF_X1 port map( D => N429, CK => CLK, Q => OUT2(21), QN 
                           => n_1562);
   OUT2_reg_20_inst : DFF_X1 port map( D => N428, CK => CLK, Q => OUT2(20), QN 
                           => n_1563);
   OUT2_reg_19_inst : DFF_X1 port map( D => N427, CK => CLK, Q => OUT2(19), QN 
                           => n_1564);
   OUT2_reg_18_inst : DFF_X1 port map( D => N426, CK => CLK, Q => OUT2(18), QN 
                           => n_1565);
   OUT1_reg_23_inst : DFF_X1 port map( D => N463, CK => CLK, Q => OUT1(23), QN 
                           => n_1566);
   OUT1_reg_22_inst : DFF_X1 port map( D => N462, CK => CLK, Q => OUT1(22), QN 
                           => n_1567);
   OUT1_reg_21_inst : DFF_X1 port map( D => N461, CK => CLK, Q => OUT1(21), QN 
                           => n_1568);
   OUT1_reg_20_inst : DFF_X1 port map( D => N460, CK => CLK, Q => OUT1(20), QN 
                           => n_1569);
   OUT1_reg_19_inst : DFF_X1 port map( D => N459, CK => CLK, Q => OUT1(19), QN 
                           => n_1570);
   OUT1_reg_18_inst : DFF_X1 port map( D => N458, CK => CLK, Q => OUT1(18), QN 
                           => n_1571);
   OUT2_reg_17_inst : DFF_X1 port map( D => N425, CK => CLK, Q => OUT2(17), QN 
                           => n_1572);
   OUT2_reg_16_inst : DFF_X1 port map( D => N424, CK => CLK, Q => OUT2(16), QN 
                           => n_1573);
   OUT2_reg_15_inst : DFF_X1 port map( D => N423, CK => CLK, Q => OUT2(15), QN 
                           => n_1574);
   OUT2_reg_14_inst : DFF_X1 port map( D => N422, CK => CLK, Q => OUT2(14), QN 
                           => n_1575);
   U7568 : INV_X1 port map( A => n10286, ZN => n10279);
   U7569 : INV_X1 port map( A => n10523, ZN => n10516);
   U7570 : INV_X1 port map( A => n10160, ZN => n10153);
   U7571 : INV_X1 port map( A => n10169, ZN => n10162);
   U7572 : INV_X1 port map( A => n10178, ZN => n10171);
   U7573 : INV_X1 port map( A => n10187, ZN => n10180);
   U7574 : INV_X1 port map( A => n10196, ZN => n10189);
   U7575 : INV_X1 port map( A => n10205, ZN => n10198);
   U7576 : INV_X1 port map( A => n10214, ZN => n10207);
   U7577 : INV_X1 port map( A => n10223, ZN => n10216);
   U7578 : INV_X1 port map( A => n10232, ZN => n10225);
   U7579 : INV_X1 port map( A => n10241, ZN => n10234);
   U7580 : INV_X1 port map( A => n10250, ZN => n10243);
   U7581 : INV_X1 port map( A => n10259, ZN => n10252);
   U7582 : INV_X1 port map( A => n10268, ZN => n10261);
   U7583 : INV_X1 port map( A => n10277, ZN => n10270);
   U7584 : INV_X1 port map( A => n10295, ZN => n10288);
   U7585 : INV_X1 port map( A => n10304, ZN => n10297);
   U7586 : INV_X1 port map( A => n10313, ZN => n10306);
   U7587 : INV_X1 port map( A => n10322, ZN => n10315);
   U7588 : INV_X1 port map( A => n10331, ZN => n10324);
   U7589 : INV_X1 port map( A => n10340, ZN => n10333);
   U7590 : INV_X1 port map( A => n10349, ZN => n10342);
   U7591 : INV_X1 port map( A => n10358, ZN => n10351);
   U7592 : INV_X1 port map( A => n10367, ZN => n10360);
   U7593 : INV_X1 port map( A => n10376, ZN => n10369);
   U7594 : INV_X1 port map( A => n10385, ZN => n10378);
   U7595 : INV_X1 port map( A => n10394, ZN => n10387);
   U7596 : INV_X1 port map( A => n10403, ZN => n10396);
   U7597 : INV_X1 port map( A => n10412, ZN => n10405);
   U7598 : INV_X1 port map( A => n10421, ZN => n10414);
   U7599 : BUF_X1 port map( A => n10287, Z => n10280);
   U7600 : BUF_X1 port map( A => n10287, Z => n10281);
   U7601 : BUF_X1 port map( A => n10287, Z => n10282);
   U7602 : BUF_X1 port map( A => n10287, Z => n10283);
   U7603 : BUF_X1 port map( A => n10287, Z => n10284);
   U7604 : BUF_X1 port map( A => n10287, Z => n10285);
   U7605 : BUF_X1 port map( A => n10524, Z => n10517);
   U7606 : BUF_X1 port map( A => n10524, Z => n10518);
   U7607 : BUF_X1 port map( A => n10524, Z => n10519);
   U7608 : BUF_X1 port map( A => n10524, Z => n10520);
   U7609 : BUF_X1 port map( A => n10524, Z => n10521);
   U7610 : BUF_X1 port map( A => n10524, Z => n10522);
   U7611 : BUF_X1 port map( A => n10287, Z => n10286);
   U7612 : BUF_X1 port map( A => n10524, Z => n10523);
   U7613 : BUF_X1 port map( A => n10152, Z => n10151);
   U7614 : BUF_X1 port map( A => n10152, Z => n10144);
   U7615 : BUF_X1 port map( A => n10151, Z => n10145);
   U7616 : BUF_X1 port map( A => n10152, Z => n10146);
   U7617 : BUF_X1 port map( A => n10151, Z => n10147);
   U7618 : BUF_X1 port map( A => n10152, Z => n10148);
   U7619 : BUF_X1 port map( A => n10152, Z => n10149);
   U7620 : BUF_X1 port map( A => n10152, Z => n10150);
   U7621 : BUF_X1 port map( A => n10146, Z => n10143);
   U7622 : NOR2_X1 port map( A1 => n8830, A2 => n10138, ZN => N432);
   U7623 : NOR2_X1 port map( A1 => n8829, A2 => n10138, ZN => N433);
   U7624 : NOR2_X1 port map( A1 => n8828, A2 => n10138, ZN => N434);
   U7625 : NOR2_X1 port map( A1 => n8827, A2 => n10138, ZN => N435);
   U7626 : NOR2_X1 port map( A1 => n8826, A2 => n10138, ZN => N436);
   U7627 : NOR2_X1 port map( A1 => n8825, A2 => n10138, ZN => N437);
   U7628 : NOR2_X1 port map( A1 => n8824, A2 => n10138, ZN => N438);
   U7629 : NOR2_X1 port map( A1 => n8822, A2 => n10138, ZN => N439);
   U7630 : NOR2_X1 port map( A1 => n8830, A2 => n10141, ZN => N464);
   U7631 : NOR2_X1 port map( A1 => n8829, A2 => n10141, ZN => N465);
   U7632 : NOR2_X1 port map( A1 => n8828, A2 => n10141, ZN => N466);
   U7633 : NOR2_X1 port map( A1 => n8827, A2 => n10141, ZN => N467);
   U7634 : NOR2_X1 port map( A1 => n8826, A2 => n10141, ZN => N468);
   U7635 : NOR2_X1 port map( A1 => n8825, A2 => n10141, ZN => N469);
   U7636 : NOR2_X1 port map( A1 => n8824, A2 => n10141, ZN => N470);
   U7637 : NOR2_X1 port map( A1 => n8822, A2 => n10141, ZN => N471);
   U7638 : NOR2_X1 port map( A1 => n8854, A2 => n10136, ZN => N408);
   U7639 : NOR2_X1 port map( A1 => n8853, A2 => n10136, ZN => N409);
   U7640 : NOR2_X1 port map( A1 => n8852, A2 => n10136, ZN => N410);
   U7641 : NOR2_X1 port map( A1 => n8851, A2 => n10136, ZN => N411);
   U7642 : NOR2_X1 port map( A1 => n8850, A2 => n10136, ZN => N412);
   U7643 : NOR2_X1 port map( A1 => n8849, A2 => n10136, ZN => N413);
   U7644 : NOR2_X1 port map( A1 => n8848, A2 => n10136, ZN => N414);
   U7645 : NOR2_X1 port map( A1 => n8847, A2 => n10136, ZN => N415);
   U7646 : NOR2_X1 port map( A1 => n8846, A2 => n10136, ZN => N416);
   U7647 : NOR2_X1 port map( A1 => n8845, A2 => n10136, ZN => N417);
   U7648 : NOR2_X1 port map( A1 => n8844, A2 => n10136, ZN => N418);
   U7649 : NOR2_X1 port map( A1 => n8843, A2 => n10136, ZN => N419);
   U7650 : NOR2_X1 port map( A1 => n8842, A2 => n10137, ZN => N420);
   U7651 : NOR2_X1 port map( A1 => n8841, A2 => n10137, ZN => N421);
   U7652 : NOR2_X1 port map( A1 => n8840, A2 => n10137, ZN => N422);
   U7653 : NOR2_X1 port map( A1 => n8839, A2 => n10137, ZN => N423);
   U7654 : NOR2_X1 port map( A1 => n8838, A2 => n10137, ZN => N424);
   U7655 : NOR2_X1 port map( A1 => n8837, A2 => n10137, ZN => N425);
   U7656 : NOR2_X1 port map( A1 => n8836, A2 => n10137, ZN => N426);
   U7657 : NOR2_X1 port map( A1 => n8835, A2 => n10137, ZN => N427);
   U7658 : NOR2_X1 port map( A1 => n8834, A2 => n10137, ZN => N428);
   U7659 : NOR2_X1 port map( A1 => n8833, A2 => n10137, ZN => N429);
   U7660 : NOR2_X1 port map( A1 => n8832, A2 => n10137, ZN => N430);
   U7661 : NOR2_X1 port map( A1 => n8831, A2 => n10137, ZN => N431);
   U7662 : NOR2_X1 port map( A1 => n8854, A2 => n10139, ZN => N440);
   U7663 : NOR2_X1 port map( A1 => n8853, A2 => n10139, ZN => N441);
   U7664 : NOR2_X1 port map( A1 => n8852, A2 => n10139, ZN => N442);
   U7665 : NOR2_X1 port map( A1 => n8851, A2 => n10139, ZN => N443);
   U7666 : NOR2_X1 port map( A1 => n8850, A2 => n10139, ZN => N444);
   U7667 : NOR2_X1 port map( A1 => n8849, A2 => n10139, ZN => N445);
   U7668 : NOR2_X1 port map( A1 => n8848, A2 => n10139, ZN => N446);
   U7669 : NOR2_X1 port map( A1 => n8847, A2 => n10139, ZN => N447);
   U7670 : NOR2_X1 port map( A1 => n8846, A2 => n10139, ZN => N448);
   U7671 : NOR2_X1 port map( A1 => n8845, A2 => n10139, ZN => N449);
   U7672 : NOR2_X1 port map( A1 => n8844, A2 => n10139, ZN => N450);
   U7673 : NOR2_X1 port map( A1 => n8843, A2 => n10139, ZN => N451);
   U7674 : NOR2_X1 port map( A1 => n8842, A2 => n10140, ZN => N452);
   U7675 : NOR2_X1 port map( A1 => n8841, A2 => n10140, ZN => N453);
   U7676 : NOR2_X1 port map( A1 => n8840, A2 => n10140, ZN => N454);
   U7677 : NOR2_X1 port map( A1 => n8839, A2 => n10140, ZN => N455);
   U7678 : NOR2_X1 port map( A1 => n8838, A2 => n10140, ZN => N456);
   U7679 : NOR2_X1 port map( A1 => n8837, A2 => n10140, ZN => N457);
   U7680 : NOR2_X1 port map( A1 => n8836, A2 => n10140, ZN => N458);
   U7681 : NOR2_X1 port map( A1 => n8835, A2 => n10140, ZN => N459);
   U7682 : NOR2_X1 port map( A1 => n8834, A2 => n10140, ZN => N460);
   U7683 : NOR2_X1 port map( A1 => n8833, A2 => n10140, ZN => N461);
   U7684 : NOR2_X1 port map( A1 => n8832, A2 => n10140, ZN => N462);
   U7685 : NOR2_X1 port map( A1 => n8831, A2 => n10140, ZN => N463);
   U7686 : BUF_X1 port map( A => n8885, Z => n10020);
   U7687 : BUF_X1 port map( A => n8885, Z => n10021);
   U7688 : BUF_X1 port map( A => n10107, Z => n10109);
   U7689 : BUF_X1 port map( A => n10055, Z => n10057);
   U7690 : BUF_X1 port map( A => n10107, Z => n10110);
   U7691 : BUF_X1 port map( A => n10055, Z => n10058);
   U7692 : BUF_X1 port map( A => n10107, Z => n10111);
   U7693 : BUF_X1 port map( A => n10055, Z => n10059);
   U7694 : BUF_X1 port map( A => n10107, Z => n10112);
   U7695 : BUF_X1 port map( A => n10055, Z => n10060);
   U7696 : BUF_X1 port map( A => n10107, Z => n10113);
   U7697 : BUF_X1 port map( A => n10055, Z => n10061);
   U7698 : BUF_X1 port map( A => n10107, Z => n10114);
   U7699 : BUF_X1 port map( A => n10055, Z => n10062);
   U7700 : BUF_X1 port map( A => n10108, Z => n10115);
   U7701 : BUF_X1 port map( A => n10056, Z => n10063);
   U7702 : BUF_X1 port map( A => n10108, Z => n10116);
   U7703 : BUF_X1 port map( A => n10056, Z => n10064);
   U7704 : BUF_X1 port map( A => n10108, Z => n10117);
   U7705 : BUF_X1 port map( A => n10056, Z => n10065);
   U7706 : BUF_X1 port map( A => n10108, Z => n10118);
   U7707 : BUF_X1 port map( A => n10056, Z => n10066);
   U7708 : BUF_X1 port map( A => n10094, Z => n10096);
   U7709 : BUF_X1 port map( A => n10042, Z => n10044);
   U7710 : BUF_X1 port map( A => n10094, Z => n10097);
   U7711 : BUF_X1 port map( A => n10042, Z => n10045);
   U7712 : BUF_X1 port map( A => n10094, Z => n10098);
   U7713 : BUF_X1 port map( A => n10042, Z => n10046);
   U7714 : BUF_X1 port map( A => n10094, Z => n10099);
   U7715 : BUF_X1 port map( A => n10042, Z => n10047);
   U7716 : BUF_X1 port map( A => n10094, Z => n10100);
   U7717 : BUF_X1 port map( A => n10042, Z => n10048);
   U7718 : BUF_X1 port map( A => n10094, Z => n10101);
   U7719 : BUF_X1 port map( A => n10042, Z => n10049);
   U7720 : BUF_X1 port map( A => n10095, Z => n10102);
   U7721 : BUF_X1 port map( A => n10043, Z => n10050);
   U7722 : BUF_X1 port map( A => n10095, Z => n10103);
   U7723 : BUF_X1 port map( A => n10043, Z => n10051);
   U7724 : BUF_X1 port map( A => n10095, Z => n10104);
   U7725 : BUF_X1 port map( A => n10043, Z => n10052);
   U7726 : BUF_X1 port map( A => n10095, Z => n10105);
   U7727 : BUF_X1 port map( A => n10043, Z => n10053);
   U7728 : BUF_X1 port map( A => n10120, Z => n10122);
   U7729 : BUF_X1 port map( A => n10068, Z => n10070);
   U7730 : BUF_X1 port map( A => n10120, Z => n10123);
   U7731 : BUF_X1 port map( A => n10068, Z => n10071);
   U7732 : BUF_X1 port map( A => n10120, Z => n10124);
   U7733 : BUF_X1 port map( A => n10068, Z => n10072);
   U7734 : BUF_X1 port map( A => n10120, Z => n10125);
   U7735 : BUF_X1 port map( A => n10068, Z => n10073);
   U7736 : BUF_X1 port map( A => n10120, Z => n10126);
   U7737 : BUF_X1 port map( A => n10068, Z => n10074);
   U7738 : BUF_X1 port map( A => n10120, Z => n10127);
   U7739 : BUF_X1 port map( A => n10068, Z => n10075);
   U7740 : BUF_X1 port map( A => n10121, Z => n10128);
   U7741 : BUF_X1 port map( A => n10069, Z => n10076);
   U7742 : BUF_X1 port map( A => n10121, Z => n10129);
   U7743 : BUF_X1 port map( A => n10069, Z => n10077);
   U7744 : BUF_X1 port map( A => n10121, Z => n10130);
   U7745 : BUF_X1 port map( A => n10069, Z => n10078);
   U7746 : BUF_X1 port map( A => n10121, Z => n10131);
   U7747 : BUF_X1 port map( A => n10069, Z => n10079);
   U7748 : BUF_X1 port map( A => n10081, Z => n10083);
   U7749 : BUF_X1 port map( A => n10029, Z => n10031);
   U7750 : BUF_X1 port map( A => n10081, Z => n10084);
   U7751 : BUF_X1 port map( A => n10029, Z => n10032);
   U7752 : BUF_X1 port map( A => n10081, Z => n10085);
   U7753 : BUF_X1 port map( A => n10029, Z => n10033);
   U7754 : BUF_X1 port map( A => n10081, Z => n10086);
   U7755 : BUF_X1 port map( A => n10029, Z => n10034);
   U7756 : BUF_X1 port map( A => n10081, Z => n10087);
   U7757 : BUF_X1 port map( A => n10029, Z => n10035);
   U7758 : BUF_X1 port map( A => n10081, Z => n10088);
   U7759 : BUF_X1 port map( A => n10029, Z => n10036);
   U7760 : BUF_X1 port map( A => n10082, Z => n10089);
   U7761 : BUF_X1 port map( A => n10030, Z => n10037);
   U7762 : BUF_X1 port map( A => n10082, Z => n10090);
   U7763 : BUF_X1 port map( A => n10030, Z => n10038);
   U7764 : BUF_X1 port map( A => n10082, Z => n10091);
   U7765 : BUF_X1 port map( A => n10030, Z => n10039);
   U7766 : BUF_X1 port map( A => n10082, Z => n10092);
   U7767 : BUF_X1 port map( A => n10030, Z => n10040);
   U7768 : BUF_X1 port map( A => n8885, Z => n10022);
   U7769 : BUF_X1 port map( A => n10323, Z => n10321);
   U7770 : BUF_X1 port map( A => n10314, Z => n10312);
   U7771 : BUF_X1 port map( A => n10305, Z => n10303);
   U7772 : BUF_X1 port map( A => n10296, Z => n10294);
   U7773 : BUF_X1 port map( A => n10161, Z => n10154);
   U7774 : BUF_X1 port map( A => n10161, Z => n10155);
   U7775 : BUF_X1 port map( A => n10161, Z => n10156);
   U7776 : BUF_X1 port map( A => n10161, Z => n10157);
   U7777 : BUF_X1 port map( A => n10161, Z => n10158);
   U7778 : BUF_X1 port map( A => n10161, Z => n10159);
   U7779 : BUF_X1 port map( A => n10170, Z => n10163);
   U7780 : BUF_X1 port map( A => n10170, Z => n10164);
   U7781 : BUF_X1 port map( A => n10170, Z => n10165);
   U7782 : BUF_X1 port map( A => n10170, Z => n10166);
   U7783 : BUF_X1 port map( A => n10170, Z => n10167);
   U7784 : BUF_X1 port map( A => n10170, Z => n10168);
   U7785 : BUF_X1 port map( A => n10179, Z => n10172);
   U7786 : BUF_X1 port map( A => n10179, Z => n10173);
   U7787 : BUF_X1 port map( A => n10179, Z => n10174);
   U7788 : BUF_X1 port map( A => n10179, Z => n10175);
   U7789 : BUF_X1 port map( A => n10179, Z => n10176);
   U7790 : BUF_X1 port map( A => n10179, Z => n10177);
   U7791 : BUF_X1 port map( A => n10188, Z => n10181);
   U7792 : BUF_X1 port map( A => n10188, Z => n10182);
   U7793 : BUF_X1 port map( A => n10188, Z => n10183);
   U7794 : BUF_X1 port map( A => n10188, Z => n10184);
   U7795 : BUF_X1 port map( A => n10188, Z => n10185);
   U7796 : BUF_X1 port map( A => n10188, Z => n10186);
   U7797 : BUF_X1 port map( A => n10197, Z => n10190);
   U7798 : BUF_X1 port map( A => n10197, Z => n10191);
   U7799 : BUF_X1 port map( A => n10197, Z => n10192);
   U7800 : BUF_X1 port map( A => n10197, Z => n10193);
   U7801 : BUF_X1 port map( A => n10197, Z => n10194);
   U7802 : BUF_X1 port map( A => n10197, Z => n10195);
   U7803 : BUF_X1 port map( A => n10206, Z => n10199);
   U7804 : BUF_X1 port map( A => n10206, Z => n10200);
   U7805 : BUF_X1 port map( A => n10206, Z => n10201);
   U7806 : BUF_X1 port map( A => n10206, Z => n10202);
   U7807 : BUF_X1 port map( A => n10206, Z => n10203);
   U7808 : BUF_X1 port map( A => n10206, Z => n10204);
   U7809 : BUF_X1 port map( A => n10215, Z => n10208);
   U7810 : BUF_X1 port map( A => n10215, Z => n10209);
   U7811 : BUF_X1 port map( A => n10215, Z => n10210);
   U7812 : BUF_X1 port map( A => n10215, Z => n10211);
   U7813 : BUF_X1 port map( A => n10215, Z => n10212);
   U7814 : BUF_X1 port map( A => n10215, Z => n10213);
   U7815 : BUF_X1 port map( A => n10224, Z => n10217);
   U7816 : BUF_X1 port map( A => n10224, Z => n10218);
   U7817 : BUF_X1 port map( A => n10224, Z => n10219);
   U7818 : BUF_X1 port map( A => n10224, Z => n10220);
   U7819 : BUF_X1 port map( A => n10224, Z => n10221);
   U7820 : BUF_X1 port map( A => n10224, Z => n10222);
   U7821 : BUF_X1 port map( A => n10233, Z => n10226);
   U7822 : BUF_X1 port map( A => n10233, Z => n10227);
   U7823 : BUF_X1 port map( A => n10233, Z => n10228);
   U7824 : BUF_X1 port map( A => n10233, Z => n10229);
   U7825 : BUF_X1 port map( A => n10233, Z => n10230);
   U7826 : BUF_X1 port map( A => n10233, Z => n10231);
   U7827 : BUF_X1 port map( A => n10242, Z => n10235);
   U7828 : BUF_X1 port map( A => n10242, Z => n10236);
   U7829 : BUF_X1 port map( A => n10242, Z => n10237);
   U7830 : BUF_X1 port map( A => n10242, Z => n10238);
   U7831 : BUF_X1 port map( A => n10242, Z => n10239);
   U7832 : BUF_X1 port map( A => n10242, Z => n10240);
   U7833 : BUF_X1 port map( A => n10251, Z => n10244);
   U7834 : BUF_X1 port map( A => n10251, Z => n10245);
   U7835 : BUF_X1 port map( A => n10251, Z => n10246);
   U7836 : BUF_X1 port map( A => n10251, Z => n10247);
   U7837 : BUF_X1 port map( A => n10251, Z => n10248);
   U7838 : BUF_X1 port map( A => n10251, Z => n10249);
   U7839 : BUF_X1 port map( A => n10260, Z => n10253);
   U7840 : BUF_X1 port map( A => n10260, Z => n10254);
   U7841 : BUF_X1 port map( A => n10260, Z => n10255);
   U7842 : BUF_X1 port map( A => n10260, Z => n10256);
   U7843 : BUF_X1 port map( A => n10260, Z => n10257);
   U7844 : BUF_X1 port map( A => n10260, Z => n10258);
   U7845 : BUF_X1 port map( A => n10269, Z => n10262);
   U7846 : BUF_X1 port map( A => n10269, Z => n10263);
   U7847 : BUF_X1 port map( A => n10269, Z => n10264);
   U7848 : BUF_X1 port map( A => n10269, Z => n10265);
   U7849 : BUF_X1 port map( A => n10269, Z => n10266);
   U7850 : BUF_X1 port map( A => n10269, Z => n10267);
   U7851 : BUF_X1 port map( A => n10278, Z => n10271);
   U7852 : BUF_X1 port map( A => n10278, Z => n10272);
   U7853 : BUF_X1 port map( A => n10278, Z => n10273);
   U7854 : BUF_X1 port map( A => n10278, Z => n10274);
   U7855 : BUF_X1 port map( A => n10278, Z => n10275);
   U7856 : BUF_X1 port map( A => n10278, Z => n10276);
   U7857 : BUF_X1 port map( A => n10296, Z => n10289);
   U7858 : BUF_X1 port map( A => n10296, Z => n10290);
   U7859 : BUF_X1 port map( A => n10296, Z => n10291);
   U7860 : BUF_X1 port map( A => n10296, Z => n10292);
   U7861 : BUF_X1 port map( A => n10296, Z => n10293);
   U7862 : BUF_X1 port map( A => n10305, Z => n10298);
   U7863 : BUF_X1 port map( A => n10305, Z => n10299);
   U7864 : BUF_X1 port map( A => n10305, Z => n10300);
   U7865 : BUF_X1 port map( A => n10305, Z => n10301);
   U7866 : BUF_X1 port map( A => n10305, Z => n10302);
   U7867 : BUF_X1 port map( A => n10314, Z => n10307);
   U7868 : BUF_X1 port map( A => n10314, Z => n10308);
   U7869 : BUF_X1 port map( A => n10314, Z => n10309);
   U7870 : BUF_X1 port map( A => n10314, Z => n10310);
   U7871 : BUF_X1 port map( A => n10314, Z => n10311);
   U7872 : BUF_X1 port map( A => n10323, Z => n10316);
   U7873 : BUF_X1 port map( A => n10323, Z => n10317);
   U7874 : BUF_X1 port map( A => n10323, Z => n10318);
   U7875 : BUF_X1 port map( A => n10323, Z => n10319);
   U7876 : BUF_X1 port map( A => n10323, Z => n10320);
   U7877 : BUF_X1 port map( A => n10332, Z => n10325);
   U7878 : BUF_X1 port map( A => n10332, Z => n10326);
   U7879 : BUF_X1 port map( A => n10332, Z => n10327);
   U7880 : BUF_X1 port map( A => n10332, Z => n10328);
   U7881 : BUF_X1 port map( A => n10332, Z => n10329);
   U7882 : BUF_X1 port map( A => n10332, Z => n10330);
   U7883 : BUF_X1 port map( A => n10341, Z => n10334);
   U7884 : BUF_X1 port map( A => n10341, Z => n10335);
   U7885 : BUF_X1 port map( A => n10341, Z => n10336);
   U7886 : BUF_X1 port map( A => n10341, Z => n10337);
   U7887 : BUF_X1 port map( A => n10341, Z => n10338);
   U7888 : BUF_X1 port map( A => n10341, Z => n10339);
   U7889 : BUF_X1 port map( A => n10350, Z => n10343);
   U7890 : BUF_X1 port map( A => n10350, Z => n10344);
   U7891 : BUF_X1 port map( A => n10350, Z => n10345);
   U7892 : BUF_X1 port map( A => n10350, Z => n10346);
   U7893 : BUF_X1 port map( A => n10350, Z => n10347);
   U7894 : BUF_X1 port map( A => n10350, Z => n10348);
   U7895 : BUF_X1 port map( A => n10359, Z => n10352);
   U7896 : BUF_X1 port map( A => n10359, Z => n10353);
   U7897 : BUF_X1 port map( A => n10359, Z => n10354);
   U7898 : BUF_X1 port map( A => n10359, Z => n10355);
   U7899 : BUF_X1 port map( A => n10359, Z => n10356);
   U7900 : BUF_X1 port map( A => n10359, Z => n10357);
   U7901 : BUF_X1 port map( A => n10368, Z => n10361);
   U7902 : BUF_X1 port map( A => n10368, Z => n10362);
   U7903 : BUF_X1 port map( A => n10368, Z => n10363);
   U7904 : BUF_X1 port map( A => n10368, Z => n10364);
   U7905 : BUF_X1 port map( A => n10368, Z => n10365);
   U7906 : BUF_X1 port map( A => n10368, Z => n10366);
   U7907 : BUF_X1 port map( A => n10377, Z => n10370);
   U7908 : BUF_X1 port map( A => n10377, Z => n10371);
   U7909 : BUF_X1 port map( A => n10377, Z => n10372);
   U7910 : BUF_X1 port map( A => n10377, Z => n10373);
   U7911 : BUF_X1 port map( A => n10377, Z => n10374);
   U7912 : BUF_X1 port map( A => n10377, Z => n10375);
   U7913 : BUF_X1 port map( A => n10386, Z => n10379);
   U7914 : BUF_X1 port map( A => n10386, Z => n10380);
   U7915 : BUF_X1 port map( A => n10386, Z => n10381);
   U7916 : BUF_X1 port map( A => n10386, Z => n10382);
   U7917 : BUF_X1 port map( A => n10386, Z => n10383);
   U7918 : BUF_X1 port map( A => n10386, Z => n10384);
   U7919 : BUF_X1 port map( A => n10395, Z => n10388);
   U7920 : BUF_X1 port map( A => n10395, Z => n10389);
   U7921 : BUF_X1 port map( A => n10395, Z => n10390);
   U7922 : BUF_X1 port map( A => n10395, Z => n10391);
   U7923 : BUF_X1 port map( A => n10395, Z => n10392);
   U7924 : BUF_X1 port map( A => n10395, Z => n10393);
   U7925 : BUF_X1 port map( A => n10404, Z => n10397);
   U7926 : BUF_X1 port map( A => n10404, Z => n10398);
   U7927 : BUF_X1 port map( A => n10404, Z => n10399);
   U7928 : BUF_X1 port map( A => n10404, Z => n10400);
   U7929 : BUF_X1 port map( A => n10404, Z => n10401);
   U7930 : BUF_X1 port map( A => n10404, Z => n10402);
   U7931 : BUF_X1 port map( A => n10413, Z => n10406);
   U7932 : BUF_X1 port map( A => n10413, Z => n10407);
   U7933 : BUF_X1 port map( A => n10413, Z => n10408);
   U7934 : BUF_X1 port map( A => n10413, Z => n10409);
   U7935 : BUF_X1 port map( A => n10413, Z => n10410);
   U7936 : BUF_X1 port map( A => n10413, Z => n10411);
   U7937 : BUF_X1 port map( A => n10422, Z => n10415);
   U7938 : BUF_X1 port map( A => n10422, Z => n10416);
   U7939 : BUF_X1 port map( A => n10422, Z => n10417);
   U7940 : BUF_X1 port map( A => n10422, Z => n10418);
   U7941 : BUF_X1 port map( A => n10422, Z => n10419);
   U7942 : BUF_X1 port map( A => n10422, Z => n10420);
   U7943 : BUF_X1 port map( A => n10161, Z => n10160);
   U7944 : BUF_X1 port map( A => n10170, Z => n10169);
   U7945 : BUF_X1 port map( A => n10179, Z => n10178);
   U7946 : BUF_X1 port map( A => n10188, Z => n10187);
   U7947 : BUF_X1 port map( A => n10197, Z => n10196);
   U7948 : BUF_X1 port map( A => n10206, Z => n10205);
   U7949 : BUF_X1 port map( A => n10215, Z => n10214);
   U7950 : BUF_X1 port map( A => n10224, Z => n10223);
   U7951 : BUF_X1 port map( A => n10233, Z => n10232);
   U7952 : BUF_X1 port map( A => n10242, Z => n10241);
   U7953 : BUF_X1 port map( A => n10251, Z => n10250);
   U7954 : BUF_X1 port map( A => n10260, Z => n10259);
   U7955 : BUF_X1 port map( A => n10269, Z => n10268);
   U7956 : BUF_X1 port map( A => n10278, Z => n10277);
   U7957 : BUF_X1 port map( A => n10296, Z => n10295);
   U7958 : BUF_X1 port map( A => n10305, Z => n10304);
   U7959 : BUF_X1 port map( A => n10314, Z => n10313);
   U7960 : BUF_X1 port map( A => n10323, Z => n10322);
   U7961 : BUF_X1 port map( A => n10332, Z => n10331);
   U7962 : BUF_X1 port map( A => n10341, Z => n10340);
   U7963 : BUF_X1 port map( A => n10350, Z => n10349);
   U7964 : BUF_X1 port map( A => n10359, Z => n10358);
   U7965 : BUF_X1 port map( A => n10368, Z => n10367);
   U7966 : BUF_X1 port map( A => n10377, Z => n10376);
   U7967 : BUF_X1 port map( A => n10386, Z => n10385);
   U7968 : BUF_X1 port map( A => n10395, Z => n10394);
   U7969 : BUF_X1 port map( A => n10404, Z => n10403);
   U7970 : BUF_X1 port map( A => n10413, Z => n10412);
   U7971 : BUF_X1 port map( A => n10422, Z => n10421);
   U7972 : INV_X1 port map( A => n8745, ZN => n10524);
   U7973 : OAI21_X1 port map( B1 => n8777, B2 => n8778, A => n10533, ZN => 
                           n8745);
   U7974 : INV_X1 port map( A => n8801, ZN => n10287);
   U7975 : OAI21_X1 port map( B1 => n8778, B2 => n8802, A => n10531, ZN => 
                           n8801);
   U7976 : INV_X1 port map( A => n10142, ZN => n10152);
   U7977 : OAI22_X1 port map( A1 => n10158, A2 => n10497, B1 => n8820, B2 => 
                           n8684, ZN => n1236);
   U7978 : OAI22_X1 port map( A1 => n10159, A2 => n10500, B1 => n8820, B2 => 
                           n8683, ZN => n1237);
   U7979 : OAI22_X1 port map( A1 => n10159, A2 => n10503, B1 => n8820, B2 => 
                           n8682, ZN => n1238);
   U7980 : OAI22_X1 port map( A1 => n10159, A2 => n10506, B1 => n8820, B2 => 
                           n8681, ZN => n1239);
   U7981 : OAI22_X1 port map( A1 => n10159, A2 => n10509, B1 => n8820, B2 => 
                           n8680, ZN => n1240);
   U7982 : OAI22_X1 port map( A1 => n10159, A2 => n10512, B1 => n8820, B2 => 
                           n8679, ZN => n1241);
   U7983 : OAI22_X1 port map( A1 => n10160, A2 => n10515, B1 => n8820, B2 => 
                           n8678, ZN => n1242);
   U7984 : OAI22_X1 port map( A1 => n10160, A2 => n10527, B1 => n8820, B2 => 
                           n8677, ZN => n1243);
   U7985 : OAI22_X1 port map( A1 => n10167, A2 => n10497, B1 => n8819, B2 => 
                           n8652, ZN => n1268);
   U7986 : OAI22_X1 port map( A1 => n10168, A2 => n10500, B1 => n8819, B2 => 
                           n8651, ZN => n1269);
   U7987 : OAI22_X1 port map( A1 => n10168, A2 => n10503, B1 => n8819, B2 => 
                           n8650, ZN => n1270);
   U7988 : OAI22_X1 port map( A1 => n10168, A2 => n10506, B1 => n8819, B2 => 
                           n8649, ZN => n1271);
   U7989 : OAI22_X1 port map( A1 => n10168, A2 => n10509, B1 => n8819, B2 => 
                           n8648, ZN => n1272);
   U7990 : OAI22_X1 port map( A1 => n10168, A2 => n10512, B1 => n8819, B2 => 
                           n8647, ZN => n1273);
   U7991 : OAI22_X1 port map( A1 => n10169, A2 => n10515, B1 => n8819, B2 => 
                           n8646, ZN => n1274);
   U7992 : OAI22_X1 port map( A1 => n10169, A2 => n10527, B1 => n8819, B2 => 
                           n8645, ZN => n1275);
   U7993 : OAI22_X1 port map( A1 => n10176, A2 => n10497, B1 => n8817, B2 => 
                           n8620, ZN => n1300);
   U7994 : OAI22_X1 port map( A1 => n10177, A2 => n10500, B1 => n8817, B2 => 
                           n8619, ZN => n1301);
   U7995 : OAI22_X1 port map( A1 => n10177, A2 => n10503, B1 => n8817, B2 => 
                           n8618, ZN => n1302);
   U7996 : OAI22_X1 port map( A1 => n10177, A2 => n10506, B1 => n8817, B2 => 
                           n8617, ZN => n1303);
   U7997 : OAI22_X1 port map( A1 => n10177, A2 => n10509, B1 => n8817, B2 => 
                           n8616, ZN => n1304);
   U7998 : OAI22_X1 port map( A1 => n10177, A2 => n10512, B1 => n8817, B2 => 
                           n8615, ZN => n1305);
   U7999 : OAI22_X1 port map( A1 => n10178, A2 => n10515, B1 => n8817, B2 => 
                           n8614, ZN => n1306);
   U8000 : OAI22_X1 port map( A1 => n10178, A2 => n10527, B1 => n8817, B2 => 
                           n8613, ZN => n1307);
   U8001 : OAI22_X1 port map( A1 => n10185, A2 => n10497, B1 => n8816, B2 => 
                           n8588, ZN => n1332);
   U8002 : OAI22_X1 port map( A1 => n10186, A2 => n10500, B1 => n8816, B2 => 
                           n8587, ZN => n1333);
   U8003 : OAI22_X1 port map( A1 => n10186, A2 => n10503, B1 => n8816, B2 => 
                           n8586, ZN => n1334);
   U8004 : OAI22_X1 port map( A1 => n10186, A2 => n10506, B1 => n8816, B2 => 
                           n8585, ZN => n1335);
   U8005 : OAI22_X1 port map( A1 => n10186, A2 => n10509, B1 => n8816, B2 => 
                           n8584, ZN => n1336);
   U8006 : OAI22_X1 port map( A1 => n10186, A2 => n10512, B1 => n8816, B2 => 
                           n8583, ZN => n1337);
   U8007 : OAI22_X1 port map( A1 => n10187, A2 => n10515, B1 => n8816, B2 => 
                           n8582, ZN => n1338);
   U8008 : OAI22_X1 port map( A1 => n10187, A2 => n10527, B1 => n8816, B2 => 
                           n8581, ZN => n1339);
   U8009 : OAI22_X1 port map( A1 => n10194, A2 => n10497, B1 => n8815, B2 => 
                           n8556, ZN => n1364);
   U8010 : OAI22_X1 port map( A1 => n10195, A2 => n10500, B1 => n8815, B2 => 
                           n8555, ZN => n1365);
   U8011 : OAI22_X1 port map( A1 => n10195, A2 => n10503, B1 => n8815, B2 => 
                           n8554, ZN => n1366);
   U8012 : OAI22_X1 port map( A1 => n10195, A2 => n10506, B1 => n8815, B2 => 
                           n8553, ZN => n1367);
   U8013 : OAI22_X1 port map( A1 => n10195, A2 => n10509, B1 => n8815, B2 => 
                           n8552, ZN => n1368);
   U8014 : OAI22_X1 port map( A1 => n10195, A2 => n10512, B1 => n8815, B2 => 
                           n8551, ZN => n1369);
   U8015 : OAI22_X1 port map( A1 => n10196, A2 => n10515, B1 => n8815, B2 => 
                           n8550, ZN => n1370);
   U8016 : OAI22_X1 port map( A1 => n10196, A2 => n10527, B1 => n8815, B2 => 
                           n8549, ZN => n1371);
   U8017 : OAI22_X1 port map( A1 => n10203, A2 => n10497, B1 => n8814, B2 => 
                           n8524, ZN => n1396);
   U8018 : OAI22_X1 port map( A1 => n10204, A2 => n10500, B1 => n8814, B2 => 
                           n8523, ZN => n1397);
   U8019 : OAI22_X1 port map( A1 => n10204, A2 => n10503, B1 => n8814, B2 => 
                           n8522, ZN => n1398);
   U8020 : OAI22_X1 port map( A1 => n10204, A2 => n10506, B1 => n8814, B2 => 
                           n8521, ZN => n1399);
   U8021 : OAI22_X1 port map( A1 => n10204, A2 => n10509, B1 => n8814, B2 => 
                           n8520, ZN => n1400);
   U8022 : OAI22_X1 port map( A1 => n10204, A2 => n10512, B1 => n8814, B2 => 
                           n8519, ZN => n1401);
   U8023 : OAI22_X1 port map( A1 => n10205, A2 => n10515, B1 => n8814, B2 => 
                           n8518, ZN => n1402);
   U8024 : OAI22_X1 port map( A1 => n10205, A2 => n10527, B1 => n8814, B2 => 
                           n8517, ZN => n1403);
   U8025 : OAI22_X1 port map( A1 => n10212, A2 => n10497, B1 => n8812, B2 => 
                           n8492, ZN => n1428);
   U8026 : OAI22_X1 port map( A1 => n10213, A2 => n10500, B1 => n8812, B2 => 
                           n8491, ZN => n1429);
   U8027 : OAI22_X1 port map( A1 => n10213, A2 => n10503, B1 => n8812, B2 => 
                           n8490, ZN => n1430);
   U8028 : OAI22_X1 port map( A1 => n10213, A2 => n10506, B1 => n8812, B2 => 
                           n8489, ZN => n1431);
   U8029 : OAI22_X1 port map( A1 => n10213, A2 => n10509, B1 => n8812, B2 => 
                           n8488, ZN => n1432);
   U8030 : OAI22_X1 port map( A1 => n10213, A2 => n10512, B1 => n8812, B2 => 
                           n8487, ZN => n1433);
   U8031 : OAI22_X1 port map( A1 => n10214, A2 => n10515, B1 => n8812, B2 => 
                           n8486, ZN => n1434);
   U8032 : OAI22_X1 port map( A1 => n10214, A2 => n10527, B1 => n8812, B2 => 
                           n8485, ZN => n1435);
   U8033 : OAI22_X1 port map( A1 => n10221, A2 => n10496, B1 => n8811, B2 => 
                           n8460, ZN => n1460);
   U8034 : OAI22_X1 port map( A1 => n10222, A2 => n10499, B1 => n8811, B2 => 
                           n8459, ZN => n1461);
   U8035 : OAI22_X1 port map( A1 => n10222, A2 => n10502, B1 => n8811, B2 => 
                           n8458, ZN => n1462);
   U8036 : OAI22_X1 port map( A1 => n10222, A2 => n10505, B1 => n8811, B2 => 
                           n8457, ZN => n1463);
   U8037 : OAI22_X1 port map( A1 => n10222, A2 => n10508, B1 => n8811, B2 => 
                           n8456, ZN => n1464);
   U8038 : OAI22_X1 port map( A1 => n10222, A2 => n10511, B1 => n8811, B2 => 
                           n8455, ZN => n1465);
   U8039 : OAI22_X1 port map( A1 => n10223, A2 => n10514, B1 => n8811, B2 => 
                           n8454, ZN => n1466);
   U8040 : OAI22_X1 port map( A1 => n10223, A2 => n10526, B1 => n8811, B2 => 
                           n8453, ZN => n1467);
   U8041 : OAI22_X1 port map( A1 => n10230, A2 => n10496, B1 => n8810, B2 => 
                           n8428, ZN => n1492);
   U8042 : OAI22_X1 port map( A1 => n10231, A2 => n10499, B1 => n8810, B2 => 
                           n8427, ZN => n1493);
   U8043 : OAI22_X1 port map( A1 => n10231, A2 => n10502, B1 => n8810, B2 => 
                           n8426, ZN => n1494);
   U8044 : OAI22_X1 port map( A1 => n10231, A2 => n10505, B1 => n8810, B2 => 
                           n8425, ZN => n1495);
   U8045 : OAI22_X1 port map( A1 => n10231, A2 => n10508, B1 => n8810, B2 => 
                           n8424, ZN => n1496);
   U8046 : OAI22_X1 port map( A1 => n10231, A2 => n10511, B1 => n8810, B2 => 
                           n8423, ZN => n1497);
   U8047 : OAI22_X1 port map( A1 => n10232, A2 => n10514, B1 => n8810, B2 => 
                           n8422, ZN => n1498);
   U8048 : OAI22_X1 port map( A1 => n10232, A2 => n10526, B1 => n8810, B2 => 
                           n8421, ZN => n1499);
   U8049 : OAI22_X1 port map( A1 => n10239, A2 => n10496, B1 => n8809, B2 => 
                           n8396, ZN => n1524);
   U8050 : OAI22_X1 port map( A1 => n10240, A2 => n10499, B1 => n8809, B2 => 
                           n8395, ZN => n1525);
   U8051 : OAI22_X1 port map( A1 => n10240, A2 => n10502, B1 => n8809, B2 => 
                           n8394, ZN => n1526);
   U8052 : OAI22_X1 port map( A1 => n10240, A2 => n10505, B1 => n8809, B2 => 
                           n8393, ZN => n1527);
   U8053 : OAI22_X1 port map( A1 => n10240, A2 => n10508, B1 => n8809, B2 => 
                           n8392, ZN => n1528);
   U8054 : OAI22_X1 port map( A1 => n10240, A2 => n10511, B1 => n8809, B2 => 
                           n8391, ZN => n1529);
   U8055 : OAI22_X1 port map( A1 => n10241, A2 => n10514, B1 => n8809, B2 => 
                           n8390, ZN => n1530);
   U8056 : OAI22_X1 port map( A1 => n10241, A2 => n10526, B1 => n8809, B2 => 
                           n8389, ZN => n1531);
   U8057 : OAI22_X1 port map( A1 => n10248, A2 => n10496, B1 => n8807, B2 => 
                           n8364, ZN => n1556);
   U8058 : OAI22_X1 port map( A1 => n10249, A2 => n10499, B1 => n8807, B2 => 
                           n8363, ZN => n1557);
   U8059 : OAI22_X1 port map( A1 => n10249, A2 => n10502, B1 => n8807, B2 => 
                           n8362, ZN => n1558);
   U8060 : OAI22_X1 port map( A1 => n10249, A2 => n10505, B1 => n8807, B2 => 
                           n8361, ZN => n1559);
   U8061 : OAI22_X1 port map( A1 => n10249, A2 => n10508, B1 => n8807, B2 => 
                           n8360, ZN => n1560);
   U8062 : OAI22_X1 port map( A1 => n10249, A2 => n10511, B1 => n8807, B2 => 
                           n8359, ZN => n1561);
   U8063 : OAI22_X1 port map( A1 => n10250, A2 => n10514, B1 => n8807, B2 => 
                           n8358, ZN => n1562);
   U8064 : OAI22_X1 port map( A1 => n10250, A2 => n10526, B1 => n8807, B2 => 
                           n8357, ZN => n1563);
   U8065 : OAI22_X1 port map( A1 => n10257, A2 => n10496, B1 => n8805, B2 => 
                           n8332, ZN => n1588);
   U8066 : OAI22_X1 port map( A1 => n10258, A2 => n10499, B1 => n8805, B2 => 
                           n8331, ZN => n1589);
   U8067 : OAI22_X1 port map( A1 => n10258, A2 => n10502, B1 => n8805, B2 => 
                           n8330, ZN => n1590);
   U8068 : OAI22_X1 port map( A1 => n10258, A2 => n10505, B1 => n8805, B2 => 
                           n8329, ZN => n1591);
   U8069 : OAI22_X1 port map( A1 => n10258, A2 => n10508, B1 => n8805, B2 => 
                           n8328, ZN => n1592);
   U8070 : OAI22_X1 port map( A1 => n10258, A2 => n10511, B1 => n8805, B2 => 
                           n8327, ZN => n1593);
   U8071 : OAI22_X1 port map( A1 => n10259, A2 => n10514, B1 => n8805, B2 => 
                           n8326, ZN => n1594);
   U8072 : OAI22_X1 port map( A1 => n10259, A2 => n10526, B1 => n8805, B2 => 
                           n8325, ZN => n1595);
   U8073 : OAI22_X1 port map( A1 => n10266, A2 => n10496, B1 => n8804, B2 => 
                           n8300, ZN => n1620);
   U8074 : OAI22_X1 port map( A1 => n10267, A2 => n10499, B1 => n8804, B2 => 
                           n8299, ZN => n1621);
   U8075 : OAI22_X1 port map( A1 => n10267, A2 => n10502, B1 => n8804, B2 => 
                           n8298, ZN => n1622);
   U8076 : OAI22_X1 port map( A1 => n10267, A2 => n10505, B1 => n8804, B2 => 
                           n8297, ZN => n1623);
   U8077 : OAI22_X1 port map( A1 => n10267, A2 => n10508, B1 => n8804, B2 => 
                           n8296, ZN => n1624);
   U8078 : OAI22_X1 port map( A1 => n10267, A2 => n10511, B1 => n8804, B2 => 
                           n8295, ZN => n1625);
   U8079 : OAI22_X1 port map( A1 => n10268, A2 => n10514, B1 => n8804, B2 => 
                           n8294, ZN => n1626);
   U8080 : OAI22_X1 port map( A1 => n10268, A2 => n10526, B1 => n8804, B2 => 
                           n8293, ZN => n1627);
   U8081 : OAI22_X1 port map( A1 => n10275, A2 => n10496, B1 => n8803, B2 => 
                           n8268, ZN => n1652);
   U8082 : OAI22_X1 port map( A1 => n10276, A2 => n10499, B1 => n8803, B2 => 
                           n8267, ZN => n1653);
   U8083 : OAI22_X1 port map( A1 => n10276, A2 => n10502, B1 => n8803, B2 => 
                           n8266, ZN => n1654);
   U8084 : OAI22_X1 port map( A1 => n10276, A2 => n10505, B1 => n8803, B2 => 
                           n8265, ZN => n1655);
   U8085 : OAI22_X1 port map( A1 => n10276, A2 => n10508, B1 => n8803, B2 => 
                           n8264, ZN => n1656);
   U8086 : OAI22_X1 port map( A1 => n10276, A2 => n10511, B1 => n8803, B2 => 
                           n8263, ZN => n1657);
   U8087 : OAI22_X1 port map( A1 => n10277, A2 => n10514, B1 => n8803, B2 => 
                           n8262, ZN => n1658);
   U8088 : OAI22_X1 port map( A1 => n10277, A2 => n10526, B1 => n8803, B2 => 
                           n8261, ZN => n1659);
   U8089 : OAI22_X1 port map( A1 => n10284, A2 => n10496, B1 => n8801, B2 => 
                           n8236, ZN => n1684);
   U8090 : OAI22_X1 port map( A1 => n10285, A2 => n10499, B1 => n8801, B2 => 
                           n8235, ZN => n1685);
   U8091 : OAI22_X1 port map( A1 => n10285, A2 => n10502, B1 => n8801, B2 => 
                           n8234, ZN => n1686);
   U8092 : OAI22_X1 port map( A1 => n10285, A2 => n10505, B1 => n8801, B2 => 
                           n8233, ZN => n1687);
   U8093 : OAI22_X1 port map( A1 => n10285, A2 => n10508, B1 => n8801, B2 => 
                           n8232, ZN => n1688);
   U8094 : OAI22_X1 port map( A1 => n10285, A2 => n10511, B1 => n8801, B2 => 
                           n8231, ZN => n1689);
   U8095 : OAI22_X1 port map( A1 => n10286, A2 => n10514, B1 => n8801, B2 => 
                           n8230, ZN => n1690);
   U8096 : OAI22_X1 port map( A1 => n10286, A2 => n10526, B1 => n8801, B2 => 
                           n8229, ZN => n1691);
   U8097 : OAI22_X1 port map( A1 => n10154, A2 => n10425, B1 => n10153, B2 => 
                           n8708, ZN => n1212);
   U8098 : OAI22_X1 port map( A1 => n10154, A2 => n10428, B1 => n10153, B2 => 
                           n8707, ZN => n1213);
   U8099 : OAI22_X1 port map( A1 => n10154, A2 => n10431, B1 => n10153, B2 => 
                           n8706, ZN => n1214);
   U8100 : OAI22_X1 port map( A1 => n10154, A2 => n10434, B1 => n10153, B2 => 
                           n8705, ZN => n1215);
   U8101 : OAI22_X1 port map( A1 => n10154, A2 => n10437, B1 => n10153, B2 => 
                           n8704, ZN => n1216);
   U8102 : OAI22_X1 port map( A1 => n10155, A2 => n10440, B1 => n10153, B2 => 
                           n8703, ZN => n1217);
   U8103 : OAI22_X1 port map( A1 => n10155, A2 => n10443, B1 => n10153, B2 => 
                           n8702, ZN => n1218);
   U8104 : OAI22_X1 port map( A1 => n10155, A2 => n10446, B1 => n10153, B2 => 
                           n8701, ZN => n1219);
   U8105 : OAI22_X1 port map( A1 => n10155, A2 => n10449, B1 => n10153, B2 => 
                           n8700, ZN => n1220);
   U8106 : OAI22_X1 port map( A1 => n10155, A2 => n10452, B1 => n10153, B2 => 
                           n8699, ZN => n1221);
   U8107 : OAI22_X1 port map( A1 => n10156, A2 => n10455, B1 => n10153, B2 => 
                           n8698, ZN => n1222);
   U8108 : OAI22_X1 port map( A1 => n10156, A2 => n10458, B1 => n10153, B2 => 
                           n8697, ZN => n1223);
   U8109 : OAI22_X1 port map( A1 => n10156, A2 => n10461, B1 => n8820, B2 => 
                           n8696, ZN => n1224);
   U8110 : OAI22_X1 port map( A1 => n10156, A2 => n10464, B1 => n8820, B2 => 
                           n8695, ZN => n1225);
   U8111 : OAI22_X1 port map( A1 => n10156, A2 => n10467, B1 => n8820, B2 => 
                           n8694, ZN => n1226);
   U8112 : OAI22_X1 port map( A1 => n10157, A2 => n10470, B1 => n10153, B2 => 
                           n8693, ZN => n1227);
   U8113 : OAI22_X1 port map( A1 => n10157, A2 => n10473, B1 => n10153, B2 => 
                           n8692, ZN => n1228);
   U8114 : OAI22_X1 port map( A1 => n10157, A2 => n10476, B1 => n10153, B2 => 
                           n8691, ZN => n1229);
   U8115 : OAI22_X1 port map( A1 => n10157, A2 => n10479, B1 => n10153, B2 => 
                           n8690, ZN => n1230);
   U8116 : OAI22_X1 port map( A1 => n10157, A2 => n10482, B1 => n10153, B2 => 
                           n8689, ZN => n1231);
   U8117 : OAI22_X1 port map( A1 => n10158, A2 => n10485, B1 => n10153, B2 => 
                           n8688, ZN => n1232);
   U8118 : OAI22_X1 port map( A1 => n10158, A2 => n10488, B1 => n10153, B2 => 
                           n8687, ZN => n1233);
   U8119 : OAI22_X1 port map( A1 => n10158, A2 => n10491, B1 => n10153, B2 => 
                           n8686, ZN => n1234);
   U8120 : OAI22_X1 port map( A1 => n10158, A2 => n10494, B1 => n10153, B2 => 
                           n8685, ZN => n1235);
   U8121 : OAI22_X1 port map( A1 => n10163, A2 => n10425, B1 => n10162, B2 => 
                           n8676, ZN => n1244);
   U8122 : OAI22_X1 port map( A1 => n10163, A2 => n10428, B1 => n10162, B2 => 
                           n8675, ZN => n1245);
   U8123 : OAI22_X1 port map( A1 => n10163, A2 => n10431, B1 => n10162, B2 => 
                           n8674, ZN => n1246);
   U8124 : OAI22_X1 port map( A1 => n10163, A2 => n10434, B1 => n10162, B2 => 
                           n8673, ZN => n1247);
   U8125 : OAI22_X1 port map( A1 => n10163, A2 => n10437, B1 => n10162, B2 => 
                           n8672, ZN => n1248);
   U8126 : OAI22_X1 port map( A1 => n10164, A2 => n10440, B1 => n10162, B2 => 
                           n8671, ZN => n1249);
   U8127 : OAI22_X1 port map( A1 => n10164, A2 => n10443, B1 => n10162, B2 => 
                           n8670, ZN => n1250);
   U8128 : OAI22_X1 port map( A1 => n10164, A2 => n10446, B1 => n10162, B2 => 
                           n8669, ZN => n1251);
   U8129 : OAI22_X1 port map( A1 => n10164, A2 => n10449, B1 => n10162, B2 => 
                           n8668, ZN => n1252);
   U8130 : OAI22_X1 port map( A1 => n10164, A2 => n10452, B1 => n10162, B2 => 
                           n8667, ZN => n1253);
   U8131 : OAI22_X1 port map( A1 => n10165, A2 => n10455, B1 => n10162, B2 => 
                           n8666, ZN => n1254);
   U8132 : OAI22_X1 port map( A1 => n10165, A2 => n10458, B1 => n10162, B2 => 
                           n8665, ZN => n1255);
   U8133 : OAI22_X1 port map( A1 => n10165, A2 => n10461, B1 => n8819, B2 => 
                           n8664, ZN => n1256);
   U8134 : OAI22_X1 port map( A1 => n10165, A2 => n10464, B1 => n8819, B2 => 
                           n8663, ZN => n1257);
   U8135 : OAI22_X1 port map( A1 => n10165, A2 => n10467, B1 => n8819, B2 => 
                           n8662, ZN => n1258);
   U8136 : OAI22_X1 port map( A1 => n10166, A2 => n10470, B1 => n10162, B2 => 
                           n8661, ZN => n1259);
   U8137 : OAI22_X1 port map( A1 => n10166, A2 => n10473, B1 => n10162, B2 => 
                           n8660, ZN => n1260);
   U8138 : OAI22_X1 port map( A1 => n10166, A2 => n10476, B1 => n10162, B2 => 
                           n8659, ZN => n1261);
   U8139 : OAI22_X1 port map( A1 => n10166, A2 => n10479, B1 => n10162, B2 => 
                           n8658, ZN => n1262);
   U8140 : OAI22_X1 port map( A1 => n10166, A2 => n10482, B1 => n10162, B2 => 
                           n8657, ZN => n1263);
   U8141 : OAI22_X1 port map( A1 => n10167, A2 => n10485, B1 => n10162, B2 => 
                           n8656, ZN => n1264);
   U8142 : OAI22_X1 port map( A1 => n10167, A2 => n10488, B1 => n10162, B2 => 
                           n8655, ZN => n1265);
   U8143 : OAI22_X1 port map( A1 => n10167, A2 => n10491, B1 => n10162, B2 => 
                           n8654, ZN => n1266);
   U8144 : OAI22_X1 port map( A1 => n10167, A2 => n10494, B1 => n10162, B2 => 
                           n8653, ZN => n1267);
   U8145 : OAI22_X1 port map( A1 => n10172, A2 => n10425, B1 => n10171, B2 => 
                           n8644, ZN => n1276);
   U8146 : OAI22_X1 port map( A1 => n10172, A2 => n10428, B1 => n10171, B2 => 
                           n8643, ZN => n1277);
   U8147 : OAI22_X1 port map( A1 => n10172, A2 => n10431, B1 => n10171, B2 => 
                           n8642, ZN => n1278);
   U8148 : OAI22_X1 port map( A1 => n10172, A2 => n10434, B1 => n10171, B2 => 
                           n8641, ZN => n1279);
   U8149 : OAI22_X1 port map( A1 => n10172, A2 => n10437, B1 => n10171, B2 => 
                           n8640, ZN => n1280);
   U8150 : OAI22_X1 port map( A1 => n10173, A2 => n10440, B1 => n10171, B2 => 
                           n8639, ZN => n1281);
   U8151 : OAI22_X1 port map( A1 => n10173, A2 => n10443, B1 => n10171, B2 => 
                           n8638, ZN => n1282);
   U8152 : OAI22_X1 port map( A1 => n10173, A2 => n10446, B1 => n10171, B2 => 
                           n8637, ZN => n1283);
   U8153 : OAI22_X1 port map( A1 => n10173, A2 => n10449, B1 => n10171, B2 => 
                           n8636, ZN => n1284);
   U8154 : OAI22_X1 port map( A1 => n10173, A2 => n10452, B1 => n10171, B2 => 
                           n8635, ZN => n1285);
   U8155 : OAI22_X1 port map( A1 => n10174, A2 => n10455, B1 => n10171, B2 => 
                           n8634, ZN => n1286);
   U8156 : OAI22_X1 port map( A1 => n10174, A2 => n10458, B1 => n10171, B2 => 
                           n8633, ZN => n1287);
   U8157 : OAI22_X1 port map( A1 => n10174, A2 => n10461, B1 => n8817, B2 => 
                           n8632, ZN => n1288);
   U8158 : OAI22_X1 port map( A1 => n10174, A2 => n10464, B1 => n8817, B2 => 
                           n8631, ZN => n1289);
   U8159 : OAI22_X1 port map( A1 => n10174, A2 => n10467, B1 => n8817, B2 => 
                           n8630, ZN => n1290);
   U8160 : OAI22_X1 port map( A1 => n10175, A2 => n10470, B1 => n10171, B2 => 
                           n8629, ZN => n1291);
   U8161 : OAI22_X1 port map( A1 => n10175, A2 => n10473, B1 => n10171, B2 => 
                           n8628, ZN => n1292);
   U8162 : OAI22_X1 port map( A1 => n10175, A2 => n10476, B1 => n10171, B2 => 
                           n8627, ZN => n1293);
   U8163 : OAI22_X1 port map( A1 => n10175, A2 => n10479, B1 => n10171, B2 => 
                           n8626, ZN => n1294);
   U8164 : OAI22_X1 port map( A1 => n10175, A2 => n10482, B1 => n10171, B2 => 
                           n8625, ZN => n1295);
   U8165 : OAI22_X1 port map( A1 => n10176, A2 => n10485, B1 => n10171, B2 => 
                           n8624, ZN => n1296);
   U8166 : OAI22_X1 port map( A1 => n10176, A2 => n10488, B1 => n10171, B2 => 
                           n8623, ZN => n1297);
   U8167 : OAI22_X1 port map( A1 => n10176, A2 => n10491, B1 => n10171, B2 => 
                           n8622, ZN => n1298);
   U8168 : OAI22_X1 port map( A1 => n10176, A2 => n10494, B1 => n10171, B2 => 
                           n8621, ZN => n1299);
   U8169 : OAI22_X1 port map( A1 => n10181, A2 => n10425, B1 => n10180, B2 => 
                           n8612, ZN => n1308);
   U8170 : OAI22_X1 port map( A1 => n10181, A2 => n10428, B1 => n10180, B2 => 
                           n8611, ZN => n1309);
   U8171 : OAI22_X1 port map( A1 => n10181, A2 => n10431, B1 => n10180, B2 => 
                           n8610, ZN => n1310);
   U8172 : OAI22_X1 port map( A1 => n10181, A2 => n10434, B1 => n10180, B2 => 
                           n8609, ZN => n1311);
   U8173 : OAI22_X1 port map( A1 => n10181, A2 => n10437, B1 => n10180, B2 => 
                           n8608, ZN => n1312);
   U8174 : OAI22_X1 port map( A1 => n10182, A2 => n10440, B1 => n10180, B2 => 
                           n8607, ZN => n1313);
   U8175 : OAI22_X1 port map( A1 => n10182, A2 => n10443, B1 => n10180, B2 => 
                           n8606, ZN => n1314);
   U8176 : OAI22_X1 port map( A1 => n10182, A2 => n10446, B1 => n10180, B2 => 
                           n8605, ZN => n1315);
   U8177 : OAI22_X1 port map( A1 => n10182, A2 => n10449, B1 => n10180, B2 => 
                           n8604, ZN => n1316);
   U8178 : OAI22_X1 port map( A1 => n10182, A2 => n10452, B1 => n10180, B2 => 
                           n8603, ZN => n1317);
   U8179 : OAI22_X1 port map( A1 => n10183, A2 => n10455, B1 => n10180, B2 => 
                           n8602, ZN => n1318);
   U8180 : OAI22_X1 port map( A1 => n10183, A2 => n10458, B1 => n10180, B2 => 
                           n8601, ZN => n1319);
   U8181 : OAI22_X1 port map( A1 => n10183, A2 => n10461, B1 => n8816, B2 => 
                           n8600, ZN => n1320);
   U8182 : OAI22_X1 port map( A1 => n10183, A2 => n10464, B1 => n8816, B2 => 
                           n8599, ZN => n1321);
   U8183 : OAI22_X1 port map( A1 => n10183, A2 => n10467, B1 => n8816, B2 => 
                           n8598, ZN => n1322);
   U8184 : OAI22_X1 port map( A1 => n10184, A2 => n10470, B1 => n10180, B2 => 
                           n8597, ZN => n1323);
   U8185 : OAI22_X1 port map( A1 => n10184, A2 => n10473, B1 => n10180, B2 => 
                           n8596, ZN => n1324);
   U8186 : OAI22_X1 port map( A1 => n10184, A2 => n10476, B1 => n10180, B2 => 
                           n8595, ZN => n1325);
   U8187 : OAI22_X1 port map( A1 => n10184, A2 => n10479, B1 => n10180, B2 => 
                           n8594, ZN => n1326);
   U8188 : OAI22_X1 port map( A1 => n10184, A2 => n10482, B1 => n10180, B2 => 
                           n8593, ZN => n1327);
   U8189 : OAI22_X1 port map( A1 => n10185, A2 => n10485, B1 => n10180, B2 => 
                           n8592, ZN => n1328);
   U8190 : OAI22_X1 port map( A1 => n10185, A2 => n10488, B1 => n10180, B2 => 
                           n8591, ZN => n1329);
   U8191 : OAI22_X1 port map( A1 => n10185, A2 => n10491, B1 => n10180, B2 => 
                           n8590, ZN => n1330);
   U8192 : OAI22_X1 port map( A1 => n10185, A2 => n10494, B1 => n10180, B2 => 
                           n8589, ZN => n1331);
   U8193 : OAI22_X1 port map( A1 => n10190, A2 => n10425, B1 => n10189, B2 => 
                           n8580, ZN => n1340);
   U8194 : OAI22_X1 port map( A1 => n10190, A2 => n10428, B1 => n10189, B2 => 
                           n8579, ZN => n1341);
   U8195 : OAI22_X1 port map( A1 => n10190, A2 => n10431, B1 => n10189, B2 => 
                           n8578, ZN => n1342);
   U8196 : OAI22_X1 port map( A1 => n10190, A2 => n10434, B1 => n10189, B2 => 
                           n8577, ZN => n1343);
   U8197 : OAI22_X1 port map( A1 => n10190, A2 => n10437, B1 => n10189, B2 => 
                           n8576, ZN => n1344);
   U8198 : OAI22_X1 port map( A1 => n10191, A2 => n10440, B1 => n10189, B2 => 
                           n8575, ZN => n1345);
   U8199 : OAI22_X1 port map( A1 => n10191, A2 => n10443, B1 => n10189, B2 => 
                           n8574, ZN => n1346);
   U8200 : OAI22_X1 port map( A1 => n10191, A2 => n10446, B1 => n10189, B2 => 
                           n8573, ZN => n1347);
   U8201 : OAI22_X1 port map( A1 => n10191, A2 => n10449, B1 => n10189, B2 => 
                           n8572, ZN => n1348);
   U8202 : OAI22_X1 port map( A1 => n10191, A2 => n10452, B1 => n10189, B2 => 
                           n8571, ZN => n1349);
   U8203 : OAI22_X1 port map( A1 => n10192, A2 => n10455, B1 => n10189, B2 => 
                           n8570, ZN => n1350);
   U8204 : OAI22_X1 port map( A1 => n10192, A2 => n10458, B1 => n10189, B2 => 
                           n8569, ZN => n1351);
   U8205 : OAI22_X1 port map( A1 => n10192, A2 => n10461, B1 => n8815, B2 => 
                           n8568, ZN => n1352);
   U8206 : OAI22_X1 port map( A1 => n10192, A2 => n10464, B1 => n8815, B2 => 
                           n8567, ZN => n1353);
   U8207 : OAI22_X1 port map( A1 => n10192, A2 => n10467, B1 => n8815, B2 => 
                           n8566, ZN => n1354);
   U8208 : OAI22_X1 port map( A1 => n10193, A2 => n10470, B1 => n10189, B2 => 
                           n8565, ZN => n1355);
   U8209 : OAI22_X1 port map( A1 => n10193, A2 => n10473, B1 => n10189, B2 => 
                           n8564, ZN => n1356);
   U8210 : OAI22_X1 port map( A1 => n10193, A2 => n10476, B1 => n10189, B2 => 
                           n8563, ZN => n1357);
   U8211 : OAI22_X1 port map( A1 => n10193, A2 => n10479, B1 => n10189, B2 => 
                           n8562, ZN => n1358);
   U8212 : OAI22_X1 port map( A1 => n10193, A2 => n10482, B1 => n10189, B2 => 
                           n8561, ZN => n1359);
   U8213 : OAI22_X1 port map( A1 => n10194, A2 => n10485, B1 => n10189, B2 => 
                           n8560, ZN => n1360);
   U8214 : OAI22_X1 port map( A1 => n10194, A2 => n10488, B1 => n10189, B2 => 
                           n8559, ZN => n1361);
   U8215 : OAI22_X1 port map( A1 => n10194, A2 => n10491, B1 => n10189, B2 => 
                           n8558, ZN => n1362);
   U8216 : OAI22_X1 port map( A1 => n10194, A2 => n10494, B1 => n10189, B2 => 
                           n8557, ZN => n1363);
   U8217 : OAI22_X1 port map( A1 => n10199, A2 => n10425, B1 => n10198, B2 => 
                           n8548, ZN => n1372);
   U8218 : OAI22_X1 port map( A1 => n10199, A2 => n10428, B1 => n10198, B2 => 
                           n8547, ZN => n1373);
   U8219 : OAI22_X1 port map( A1 => n10199, A2 => n10431, B1 => n10198, B2 => 
                           n8546, ZN => n1374);
   U8220 : OAI22_X1 port map( A1 => n10199, A2 => n10434, B1 => n10198, B2 => 
                           n8545, ZN => n1375);
   U8221 : OAI22_X1 port map( A1 => n10199, A2 => n10437, B1 => n10198, B2 => 
                           n8544, ZN => n1376);
   U8222 : OAI22_X1 port map( A1 => n10200, A2 => n10440, B1 => n10198, B2 => 
                           n8543, ZN => n1377);
   U8223 : OAI22_X1 port map( A1 => n10200, A2 => n10443, B1 => n10198, B2 => 
                           n8542, ZN => n1378);
   U8224 : OAI22_X1 port map( A1 => n10200, A2 => n10446, B1 => n10198, B2 => 
                           n8541, ZN => n1379);
   U8225 : OAI22_X1 port map( A1 => n10200, A2 => n10449, B1 => n10198, B2 => 
                           n8540, ZN => n1380);
   U8226 : OAI22_X1 port map( A1 => n10200, A2 => n10452, B1 => n10198, B2 => 
                           n8539, ZN => n1381);
   U8227 : OAI22_X1 port map( A1 => n10201, A2 => n10455, B1 => n10198, B2 => 
                           n8538, ZN => n1382);
   U8228 : OAI22_X1 port map( A1 => n10201, A2 => n10458, B1 => n10198, B2 => 
                           n8537, ZN => n1383);
   U8229 : OAI22_X1 port map( A1 => n10201, A2 => n10461, B1 => n8814, B2 => 
                           n8536, ZN => n1384);
   U8230 : OAI22_X1 port map( A1 => n10201, A2 => n10464, B1 => n8814, B2 => 
                           n8535, ZN => n1385);
   U8231 : OAI22_X1 port map( A1 => n10201, A2 => n10467, B1 => n8814, B2 => 
                           n8534, ZN => n1386);
   U8232 : OAI22_X1 port map( A1 => n10202, A2 => n10470, B1 => n10198, B2 => 
                           n8533, ZN => n1387);
   U8233 : OAI22_X1 port map( A1 => n10202, A2 => n10473, B1 => n10198, B2 => 
                           n8532, ZN => n1388);
   U8234 : OAI22_X1 port map( A1 => n10202, A2 => n10476, B1 => n10198, B2 => 
                           n8531, ZN => n1389);
   U8235 : OAI22_X1 port map( A1 => n10202, A2 => n10479, B1 => n10198, B2 => 
                           n8530, ZN => n1390);
   U8236 : OAI22_X1 port map( A1 => n10202, A2 => n10482, B1 => n10198, B2 => 
                           n8529, ZN => n1391);
   U8237 : OAI22_X1 port map( A1 => n10203, A2 => n10485, B1 => n10198, B2 => 
                           n8528, ZN => n1392);
   U8238 : OAI22_X1 port map( A1 => n10203, A2 => n10488, B1 => n10198, B2 => 
                           n8527, ZN => n1393);
   U8239 : OAI22_X1 port map( A1 => n10203, A2 => n10491, B1 => n10198, B2 => 
                           n8526, ZN => n1394);
   U8240 : OAI22_X1 port map( A1 => n10203, A2 => n10494, B1 => n10198, B2 => 
                           n8525, ZN => n1395);
   U8241 : OAI22_X1 port map( A1 => n10208, A2 => n10425, B1 => n10207, B2 => 
                           n8516, ZN => n1404);
   U8242 : OAI22_X1 port map( A1 => n10208, A2 => n10428, B1 => n10207, B2 => 
                           n8515, ZN => n1405);
   U8243 : OAI22_X1 port map( A1 => n10208, A2 => n10431, B1 => n10207, B2 => 
                           n8514, ZN => n1406);
   U8244 : OAI22_X1 port map( A1 => n10208, A2 => n10434, B1 => n10207, B2 => 
                           n8513, ZN => n1407);
   U8245 : OAI22_X1 port map( A1 => n10208, A2 => n10437, B1 => n10207, B2 => 
                           n8512, ZN => n1408);
   U8246 : OAI22_X1 port map( A1 => n10209, A2 => n10440, B1 => n10207, B2 => 
                           n8511, ZN => n1409);
   U8247 : OAI22_X1 port map( A1 => n10209, A2 => n10443, B1 => n10207, B2 => 
                           n8510, ZN => n1410);
   U8248 : OAI22_X1 port map( A1 => n10209, A2 => n10446, B1 => n10207, B2 => 
                           n8509, ZN => n1411);
   U8249 : OAI22_X1 port map( A1 => n10209, A2 => n10449, B1 => n10207, B2 => 
                           n8508, ZN => n1412);
   U8250 : OAI22_X1 port map( A1 => n10209, A2 => n10452, B1 => n10207, B2 => 
                           n8507, ZN => n1413);
   U8251 : OAI22_X1 port map( A1 => n10210, A2 => n10455, B1 => n10207, B2 => 
                           n8506, ZN => n1414);
   U8252 : OAI22_X1 port map( A1 => n10210, A2 => n10458, B1 => n10207, B2 => 
                           n8505, ZN => n1415);
   U8253 : OAI22_X1 port map( A1 => n10210, A2 => n10461, B1 => n8812, B2 => 
                           n8504, ZN => n1416);
   U8254 : OAI22_X1 port map( A1 => n10210, A2 => n10464, B1 => n8812, B2 => 
                           n8503, ZN => n1417);
   U8255 : OAI22_X1 port map( A1 => n10210, A2 => n10467, B1 => n8812, B2 => 
                           n8502, ZN => n1418);
   U8256 : OAI22_X1 port map( A1 => n10211, A2 => n10470, B1 => n10207, B2 => 
                           n8501, ZN => n1419);
   U8257 : OAI22_X1 port map( A1 => n10211, A2 => n10473, B1 => n10207, B2 => 
                           n8500, ZN => n1420);
   U8258 : OAI22_X1 port map( A1 => n10211, A2 => n10476, B1 => n10207, B2 => 
                           n8499, ZN => n1421);
   U8259 : OAI22_X1 port map( A1 => n10211, A2 => n10479, B1 => n10207, B2 => 
                           n8498, ZN => n1422);
   U8260 : OAI22_X1 port map( A1 => n10211, A2 => n10482, B1 => n10207, B2 => 
                           n8497, ZN => n1423);
   U8261 : OAI22_X1 port map( A1 => n10212, A2 => n10485, B1 => n10207, B2 => 
                           n8496, ZN => n1424);
   U8262 : OAI22_X1 port map( A1 => n10212, A2 => n10488, B1 => n10207, B2 => 
                           n8495, ZN => n1425);
   U8263 : OAI22_X1 port map( A1 => n10212, A2 => n10491, B1 => n10207, B2 => 
                           n8494, ZN => n1426);
   U8264 : OAI22_X1 port map( A1 => n10212, A2 => n10494, B1 => n10207, B2 => 
                           n8493, ZN => n1427);
   U8265 : OAI22_X1 port map( A1 => n10217, A2 => n10424, B1 => n10216, B2 => 
                           n8484, ZN => n1436);
   U8266 : OAI22_X1 port map( A1 => n10217, A2 => n10427, B1 => n10216, B2 => 
                           n8483, ZN => n1437);
   U8267 : OAI22_X1 port map( A1 => n10217, A2 => n10430, B1 => n10216, B2 => 
                           n8482, ZN => n1438);
   U8268 : OAI22_X1 port map( A1 => n10217, A2 => n10433, B1 => n10216, B2 => 
                           n8481, ZN => n1439);
   U8269 : OAI22_X1 port map( A1 => n10217, A2 => n10436, B1 => n10216, B2 => 
                           n8480, ZN => n1440);
   U8270 : OAI22_X1 port map( A1 => n10218, A2 => n10439, B1 => n10216, B2 => 
                           n8479, ZN => n1441);
   U8271 : OAI22_X1 port map( A1 => n10218, A2 => n10442, B1 => n10216, B2 => 
                           n8478, ZN => n1442);
   U8272 : OAI22_X1 port map( A1 => n10218, A2 => n10445, B1 => n10216, B2 => 
                           n8477, ZN => n1443);
   U8273 : OAI22_X1 port map( A1 => n10218, A2 => n10448, B1 => n10216, B2 => 
                           n8476, ZN => n1444);
   U8274 : OAI22_X1 port map( A1 => n10218, A2 => n10451, B1 => n10216, B2 => 
                           n8475, ZN => n1445);
   U8275 : OAI22_X1 port map( A1 => n10219, A2 => n10454, B1 => n10216, B2 => 
                           n8474, ZN => n1446);
   U8276 : OAI22_X1 port map( A1 => n10219, A2 => n10457, B1 => n10216, B2 => 
                           n8473, ZN => n1447);
   U8277 : OAI22_X1 port map( A1 => n10219, A2 => n10460, B1 => n8811, B2 => 
                           n8472, ZN => n1448);
   U8278 : OAI22_X1 port map( A1 => n10219, A2 => n10463, B1 => n8811, B2 => 
                           n8471, ZN => n1449);
   U8279 : OAI22_X1 port map( A1 => n10219, A2 => n10466, B1 => n8811, B2 => 
                           n8470, ZN => n1450);
   U8280 : OAI22_X1 port map( A1 => n10220, A2 => n10469, B1 => n10216, B2 => 
                           n8469, ZN => n1451);
   U8281 : OAI22_X1 port map( A1 => n10220, A2 => n10472, B1 => n10216, B2 => 
                           n8468, ZN => n1452);
   U8282 : OAI22_X1 port map( A1 => n10220, A2 => n10475, B1 => n10216, B2 => 
                           n8467, ZN => n1453);
   U8283 : OAI22_X1 port map( A1 => n10220, A2 => n10478, B1 => n10216, B2 => 
                           n8466, ZN => n1454);
   U8284 : OAI22_X1 port map( A1 => n10220, A2 => n10481, B1 => n10216, B2 => 
                           n8465, ZN => n1455);
   U8285 : OAI22_X1 port map( A1 => n10221, A2 => n10484, B1 => n10216, B2 => 
                           n8464, ZN => n1456);
   U8286 : OAI22_X1 port map( A1 => n10221, A2 => n10487, B1 => n10216, B2 => 
                           n8463, ZN => n1457);
   U8287 : OAI22_X1 port map( A1 => n10221, A2 => n10490, B1 => n10216, B2 => 
                           n8462, ZN => n1458);
   U8288 : OAI22_X1 port map( A1 => n10221, A2 => n10493, B1 => n10216, B2 => 
                           n8461, ZN => n1459);
   U8289 : OAI22_X1 port map( A1 => n10226, A2 => n10424, B1 => n10225, B2 => 
                           n8452, ZN => n1468);
   U8290 : OAI22_X1 port map( A1 => n10226, A2 => n10427, B1 => n10225, B2 => 
                           n8451, ZN => n1469);
   U8291 : OAI22_X1 port map( A1 => n10226, A2 => n10430, B1 => n10225, B2 => 
                           n8450, ZN => n1470);
   U8292 : OAI22_X1 port map( A1 => n10226, A2 => n10433, B1 => n10225, B2 => 
                           n8449, ZN => n1471);
   U8293 : OAI22_X1 port map( A1 => n10226, A2 => n10436, B1 => n10225, B2 => 
                           n8448, ZN => n1472);
   U8294 : OAI22_X1 port map( A1 => n10227, A2 => n10439, B1 => n10225, B2 => 
                           n8447, ZN => n1473);
   U8295 : OAI22_X1 port map( A1 => n10227, A2 => n10442, B1 => n10225, B2 => 
                           n8446, ZN => n1474);
   U8296 : OAI22_X1 port map( A1 => n10227, A2 => n10445, B1 => n10225, B2 => 
                           n8445, ZN => n1475);
   U8297 : OAI22_X1 port map( A1 => n10227, A2 => n10448, B1 => n10225, B2 => 
                           n8444, ZN => n1476);
   U8298 : OAI22_X1 port map( A1 => n10227, A2 => n10451, B1 => n10225, B2 => 
                           n8443, ZN => n1477);
   U8299 : OAI22_X1 port map( A1 => n10228, A2 => n10454, B1 => n10225, B2 => 
                           n8442, ZN => n1478);
   U8300 : OAI22_X1 port map( A1 => n10228, A2 => n10457, B1 => n10225, B2 => 
                           n8441, ZN => n1479);
   U8301 : OAI22_X1 port map( A1 => n10228, A2 => n10460, B1 => n8810, B2 => 
                           n8440, ZN => n1480);
   U8302 : OAI22_X1 port map( A1 => n10228, A2 => n10463, B1 => n8810, B2 => 
                           n8439, ZN => n1481);
   U8303 : OAI22_X1 port map( A1 => n10228, A2 => n10466, B1 => n8810, B2 => 
                           n8438, ZN => n1482);
   U8304 : OAI22_X1 port map( A1 => n10229, A2 => n10469, B1 => n10225, B2 => 
                           n8437, ZN => n1483);
   U8305 : OAI22_X1 port map( A1 => n10229, A2 => n10472, B1 => n10225, B2 => 
                           n8436, ZN => n1484);
   U8306 : OAI22_X1 port map( A1 => n10229, A2 => n10475, B1 => n10225, B2 => 
                           n8435, ZN => n1485);
   U8307 : OAI22_X1 port map( A1 => n10229, A2 => n10478, B1 => n10225, B2 => 
                           n8434, ZN => n1486);
   U8308 : OAI22_X1 port map( A1 => n10229, A2 => n10481, B1 => n10225, B2 => 
                           n8433, ZN => n1487);
   U8309 : OAI22_X1 port map( A1 => n10230, A2 => n10484, B1 => n10225, B2 => 
                           n8432, ZN => n1488);
   U8310 : OAI22_X1 port map( A1 => n10230, A2 => n10487, B1 => n10225, B2 => 
                           n8431, ZN => n1489);
   U8311 : OAI22_X1 port map( A1 => n10230, A2 => n10490, B1 => n10225, B2 => 
                           n8430, ZN => n1490);
   U8312 : OAI22_X1 port map( A1 => n10230, A2 => n10493, B1 => n10225, B2 => 
                           n8429, ZN => n1491);
   U8313 : OAI22_X1 port map( A1 => n10235, A2 => n10424, B1 => n10234, B2 => 
                           n8420, ZN => n1500);
   U8314 : OAI22_X1 port map( A1 => n10235, A2 => n10427, B1 => n10234, B2 => 
                           n8419, ZN => n1501);
   U8315 : OAI22_X1 port map( A1 => n10235, A2 => n10430, B1 => n10234, B2 => 
                           n8418, ZN => n1502);
   U8316 : OAI22_X1 port map( A1 => n10235, A2 => n10433, B1 => n10234, B2 => 
                           n8417, ZN => n1503);
   U8317 : OAI22_X1 port map( A1 => n10235, A2 => n10436, B1 => n10234, B2 => 
                           n8416, ZN => n1504);
   U8318 : OAI22_X1 port map( A1 => n10236, A2 => n10439, B1 => n10234, B2 => 
                           n8415, ZN => n1505);
   U8319 : OAI22_X1 port map( A1 => n10236, A2 => n10442, B1 => n10234, B2 => 
                           n8414, ZN => n1506);
   U8320 : OAI22_X1 port map( A1 => n10236, A2 => n10445, B1 => n10234, B2 => 
                           n8413, ZN => n1507);
   U8321 : OAI22_X1 port map( A1 => n10236, A2 => n10448, B1 => n10234, B2 => 
                           n8412, ZN => n1508);
   U8322 : OAI22_X1 port map( A1 => n10236, A2 => n10451, B1 => n10234, B2 => 
                           n8411, ZN => n1509);
   U8323 : OAI22_X1 port map( A1 => n10237, A2 => n10454, B1 => n10234, B2 => 
                           n8410, ZN => n1510);
   U8324 : OAI22_X1 port map( A1 => n10237, A2 => n10457, B1 => n10234, B2 => 
                           n8409, ZN => n1511);
   U8325 : OAI22_X1 port map( A1 => n10237, A2 => n10460, B1 => n8809, B2 => 
                           n8408, ZN => n1512);
   U8326 : OAI22_X1 port map( A1 => n10237, A2 => n10463, B1 => n8809, B2 => 
                           n8407, ZN => n1513);
   U8327 : OAI22_X1 port map( A1 => n10237, A2 => n10466, B1 => n8809, B2 => 
                           n8406, ZN => n1514);
   U8328 : OAI22_X1 port map( A1 => n10238, A2 => n10469, B1 => n10234, B2 => 
                           n8405, ZN => n1515);
   U8329 : OAI22_X1 port map( A1 => n10238, A2 => n10472, B1 => n10234, B2 => 
                           n8404, ZN => n1516);
   U8330 : OAI22_X1 port map( A1 => n10238, A2 => n10475, B1 => n10234, B2 => 
                           n8403, ZN => n1517);
   U8331 : OAI22_X1 port map( A1 => n10238, A2 => n10478, B1 => n10234, B2 => 
                           n8402, ZN => n1518);
   U8332 : OAI22_X1 port map( A1 => n10238, A2 => n10481, B1 => n10234, B2 => 
                           n8401, ZN => n1519);
   U8333 : OAI22_X1 port map( A1 => n10239, A2 => n10484, B1 => n10234, B2 => 
                           n8400, ZN => n1520);
   U8334 : OAI22_X1 port map( A1 => n10239, A2 => n10487, B1 => n10234, B2 => 
                           n8399, ZN => n1521);
   U8335 : OAI22_X1 port map( A1 => n10239, A2 => n10490, B1 => n10234, B2 => 
                           n8398, ZN => n1522);
   U8336 : OAI22_X1 port map( A1 => n10239, A2 => n10493, B1 => n10234, B2 => 
                           n8397, ZN => n1523);
   U8337 : OAI22_X1 port map( A1 => n10244, A2 => n10424, B1 => n10243, B2 => 
                           n8388, ZN => n1532);
   U8338 : OAI22_X1 port map( A1 => n10244, A2 => n10427, B1 => n10243, B2 => 
                           n8387, ZN => n1533);
   U8339 : OAI22_X1 port map( A1 => n10244, A2 => n10430, B1 => n10243, B2 => 
                           n8386, ZN => n1534);
   U8340 : OAI22_X1 port map( A1 => n10244, A2 => n10433, B1 => n10243, B2 => 
                           n8385, ZN => n1535);
   U8341 : OAI22_X1 port map( A1 => n10244, A2 => n10436, B1 => n10243, B2 => 
                           n8384, ZN => n1536);
   U8342 : OAI22_X1 port map( A1 => n10245, A2 => n10439, B1 => n10243, B2 => 
                           n8383, ZN => n1537);
   U8343 : OAI22_X1 port map( A1 => n10245, A2 => n10442, B1 => n10243, B2 => 
                           n8382, ZN => n1538);
   U8344 : OAI22_X1 port map( A1 => n10245, A2 => n10445, B1 => n10243, B2 => 
                           n8381, ZN => n1539);
   U8345 : OAI22_X1 port map( A1 => n10245, A2 => n10448, B1 => n10243, B2 => 
                           n8380, ZN => n1540);
   U8346 : OAI22_X1 port map( A1 => n10245, A2 => n10451, B1 => n10243, B2 => 
                           n8379, ZN => n1541);
   U8347 : OAI22_X1 port map( A1 => n10246, A2 => n10454, B1 => n10243, B2 => 
                           n8378, ZN => n1542);
   U8348 : OAI22_X1 port map( A1 => n10246, A2 => n10457, B1 => n10243, B2 => 
                           n8377, ZN => n1543);
   U8349 : OAI22_X1 port map( A1 => n10246, A2 => n10460, B1 => n8807, B2 => 
                           n8376, ZN => n1544);
   U8350 : OAI22_X1 port map( A1 => n10246, A2 => n10463, B1 => n8807, B2 => 
                           n8375, ZN => n1545);
   U8351 : OAI22_X1 port map( A1 => n10246, A2 => n10466, B1 => n8807, B2 => 
                           n8374, ZN => n1546);
   U8352 : OAI22_X1 port map( A1 => n10247, A2 => n10469, B1 => n10243, B2 => 
                           n8373, ZN => n1547);
   U8353 : OAI22_X1 port map( A1 => n10247, A2 => n10472, B1 => n10243, B2 => 
                           n8372, ZN => n1548);
   U8354 : OAI22_X1 port map( A1 => n10247, A2 => n10475, B1 => n10243, B2 => 
                           n8371, ZN => n1549);
   U8355 : OAI22_X1 port map( A1 => n10247, A2 => n10478, B1 => n10243, B2 => 
                           n8370, ZN => n1550);
   U8356 : OAI22_X1 port map( A1 => n10247, A2 => n10481, B1 => n10243, B2 => 
                           n8369, ZN => n1551);
   U8357 : OAI22_X1 port map( A1 => n10248, A2 => n10484, B1 => n10243, B2 => 
                           n8368, ZN => n1552);
   U8358 : OAI22_X1 port map( A1 => n10248, A2 => n10487, B1 => n10243, B2 => 
                           n8367, ZN => n1553);
   U8359 : OAI22_X1 port map( A1 => n10248, A2 => n10490, B1 => n10243, B2 => 
                           n8366, ZN => n1554);
   U8360 : OAI22_X1 port map( A1 => n10248, A2 => n10493, B1 => n10243, B2 => 
                           n8365, ZN => n1555);
   U8361 : OAI22_X1 port map( A1 => n10253, A2 => n10424, B1 => n10252, B2 => 
                           n8356, ZN => n1564);
   U8362 : OAI22_X1 port map( A1 => n10253, A2 => n10427, B1 => n10252, B2 => 
                           n8355, ZN => n1565);
   U8363 : OAI22_X1 port map( A1 => n10253, A2 => n10430, B1 => n10252, B2 => 
                           n8354, ZN => n1566);
   U8364 : OAI22_X1 port map( A1 => n10253, A2 => n10433, B1 => n10252, B2 => 
                           n8353, ZN => n1567);
   U8365 : OAI22_X1 port map( A1 => n10253, A2 => n10436, B1 => n10252, B2 => 
                           n8352, ZN => n1568);
   U8366 : OAI22_X1 port map( A1 => n10254, A2 => n10439, B1 => n10252, B2 => 
                           n8351, ZN => n1569);
   U8367 : OAI22_X1 port map( A1 => n10254, A2 => n10442, B1 => n10252, B2 => 
                           n8350, ZN => n1570);
   U8368 : OAI22_X1 port map( A1 => n10254, A2 => n10445, B1 => n10252, B2 => 
                           n8349, ZN => n1571);
   U8369 : OAI22_X1 port map( A1 => n10254, A2 => n10448, B1 => n10252, B2 => 
                           n8348, ZN => n1572);
   U8370 : OAI22_X1 port map( A1 => n10254, A2 => n10451, B1 => n10252, B2 => 
                           n8347, ZN => n1573);
   U8371 : OAI22_X1 port map( A1 => n10255, A2 => n10454, B1 => n10252, B2 => 
                           n8346, ZN => n1574);
   U8372 : OAI22_X1 port map( A1 => n10255, A2 => n10457, B1 => n10252, B2 => 
                           n8345, ZN => n1575);
   U8373 : OAI22_X1 port map( A1 => n10255, A2 => n10460, B1 => n8805, B2 => 
                           n8344, ZN => n1576);
   U8374 : OAI22_X1 port map( A1 => n10255, A2 => n10463, B1 => n8805, B2 => 
                           n8343, ZN => n1577);
   U8375 : OAI22_X1 port map( A1 => n10255, A2 => n10466, B1 => n8805, B2 => 
                           n8342, ZN => n1578);
   U8376 : OAI22_X1 port map( A1 => n10256, A2 => n10469, B1 => n10252, B2 => 
                           n8341, ZN => n1579);
   U8377 : OAI22_X1 port map( A1 => n10256, A2 => n10472, B1 => n10252, B2 => 
                           n8340, ZN => n1580);
   U8378 : OAI22_X1 port map( A1 => n10256, A2 => n10475, B1 => n10252, B2 => 
                           n8339, ZN => n1581);
   U8379 : OAI22_X1 port map( A1 => n10256, A2 => n10478, B1 => n10252, B2 => 
                           n8338, ZN => n1582);
   U8380 : OAI22_X1 port map( A1 => n10256, A2 => n10481, B1 => n10252, B2 => 
                           n8337, ZN => n1583);
   U8381 : OAI22_X1 port map( A1 => n10257, A2 => n10484, B1 => n10252, B2 => 
                           n8336, ZN => n1584);
   U8382 : OAI22_X1 port map( A1 => n10257, A2 => n10487, B1 => n10252, B2 => 
                           n8335, ZN => n1585);
   U8383 : OAI22_X1 port map( A1 => n10257, A2 => n10490, B1 => n10252, B2 => 
                           n8334, ZN => n1586);
   U8384 : OAI22_X1 port map( A1 => n10257, A2 => n10493, B1 => n10252, B2 => 
                           n8333, ZN => n1587);
   U8385 : OAI22_X1 port map( A1 => n10262, A2 => n10424, B1 => n10261, B2 => 
                           n8324, ZN => n1596);
   U8386 : OAI22_X1 port map( A1 => n10262, A2 => n10427, B1 => n10261, B2 => 
                           n8323, ZN => n1597);
   U8387 : OAI22_X1 port map( A1 => n10262, A2 => n10430, B1 => n10261, B2 => 
                           n8322, ZN => n1598);
   U8388 : OAI22_X1 port map( A1 => n10262, A2 => n10433, B1 => n10261, B2 => 
                           n8321, ZN => n1599);
   U8389 : OAI22_X1 port map( A1 => n10262, A2 => n10436, B1 => n10261, B2 => 
                           n8320, ZN => n1600);
   U8390 : OAI22_X1 port map( A1 => n10263, A2 => n10439, B1 => n10261, B2 => 
                           n8319, ZN => n1601);
   U8391 : OAI22_X1 port map( A1 => n10263, A2 => n10442, B1 => n10261, B2 => 
                           n8318, ZN => n1602);
   U8392 : OAI22_X1 port map( A1 => n10263, A2 => n10445, B1 => n10261, B2 => 
                           n8317, ZN => n1603);
   U8393 : OAI22_X1 port map( A1 => n10263, A2 => n10448, B1 => n10261, B2 => 
                           n8316, ZN => n1604);
   U8394 : OAI22_X1 port map( A1 => n10263, A2 => n10451, B1 => n10261, B2 => 
                           n8315, ZN => n1605);
   U8395 : OAI22_X1 port map( A1 => n10264, A2 => n10454, B1 => n10261, B2 => 
                           n8314, ZN => n1606);
   U8396 : OAI22_X1 port map( A1 => n10264, A2 => n10457, B1 => n10261, B2 => 
                           n8313, ZN => n1607);
   U8397 : OAI22_X1 port map( A1 => n10264, A2 => n10460, B1 => n8804, B2 => 
                           n8312, ZN => n1608);
   U8398 : OAI22_X1 port map( A1 => n10264, A2 => n10463, B1 => n8804, B2 => 
                           n8311, ZN => n1609);
   U8399 : OAI22_X1 port map( A1 => n10264, A2 => n10466, B1 => n8804, B2 => 
                           n8310, ZN => n1610);
   U8400 : OAI22_X1 port map( A1 => n10265, A2 => n10469, B1 => n10261, B2 => 
                           n8309, ZN => n1611);
   U8401 : OAI22_X1 port map( A1 => n10265, A2 => n10472, B1 => n10261, B2 => 
                           n8308, ZN => n1612);
   U8402 : OAI22_X1 port map( A1 => n10265, A2 => n10475, B1 => n10261, B2 => 
                           n8307, ZN => n1613);
   U8403 : OAI22_X1 port map( A1 => n10265, A2 => n10478, B1 => n10261, B2 => 
                           n8306, ZN => n1614);
   U8404 : OAI22_X1 port map( A1 => n10265, A2 => n10481, B1 => n10261, B2 => 
                           n8305, ZN => n1615);
   U8405 : OAI22_X1 port map( A1 => n10266, A2 => n10484, B1 => n10261, B2 => 
                           n8304, ZN => n1616);
   U8406 : OAI22_X1 port map( A1 => n10266, A2 => n10487, B1 => n10261, B2 => 
                           n8303, ZN => n1617);
   U8407 : OAI22_X1 port map( A1 => n10266, A2 => n10490, B1 => n10261, B2 => 
                           n8302, ZN => n1618);
   U8408 : OAI22_X1 port map( A1 => n10266, A2 => n10493, B1 => n10261, B2 => 
                           n8301, ZN => n1619);
   U8409 : OAI22_X1 port map( A1 => n10271, A2 => n10424, B1 => n10270, B2 => 
                           n8292, ZN => n1628);
   U8410 : OAI22_X1 port map( A1 => n10271, A2 => n10427, B1 => n10270, B2 => 
                           n8291, ZN => n1629);
   U8411 : OAI22_X1 port map( A1 => n10271, A2 => n10430, B1 => n10270, B2 => 
                           n8290, ZN => n1630);
   U8412 : OAI22_X1 port map( A1 => n10271, A2 => n10433, B1 => n10270, B2 => 
                           n8289, ZN => n1631);
   U8413 : OAI22_X1 port map( A1 => n10271, A2 => n10436, B1 => n10270, B2 => 
                           n8288, ZN => n1632);
   U8414 : OAI22_X1 port map( A1 => n10272, A2 => n10439, B1 => n10270, B2 => 
                           n8287, ZN => n1633);
   U8415 : OAI22_X1 port map( A1 => n10272, A2 => n10442, B1 => n10270, B2 => 
                           n8286, ZN => n1634);
   U8416 : OAI22_X1 port map( A1 => n10272, A2 => n10445, B1 => n10270, B2 => 
                           n8285, ZN => n1635);
   U8417 : OAI22_X1 port map( A1 => n10272, A2 => n10448, B1 => n10270, B2 => 
                           n8284, ZN => n1636);
   U8418 : OAI22_X1 port map( A1 => n10272, A2 => n10451, B1 => n10270, B2 => 
                           n8283, ZN => n1637);
   U8419 : OAI22_X1 port map( A1 => n10273, A2 => n10454, B1 => n10270, B2 => 
                           n8282, ZN => n1638);
   U8420 : OAI22_X1 port map( A1 => n10273, A2 => n10457, B1 => n10270, B2 => 
                           n8281, ZN => n1639);
   U8421 : OAI22_X1 port map( A1 => n10273, A2 => n10460, B1 => n8803, B2 => 
                           n8280, ZN => n1640);
   U8422 : OAI22_X1 port map( A1 => n10273, A2 => n10463, B1 => n8803, B2 => 
                           n8279, ZN => n1641);
   U8423 : OAI22_X1 port map( A1 => n10273, A2 => n10466, B1 => n8803, B2 => 
                           n8278, ZN => n1642);
   U8424 : OAI22_X1 port map( A1 => n10274, A2 => n10469, B1 => n10270, B2 => 
                           n8277, ZN => n1643);
   U8425 : OAI22_X1 port map( A1 => n10274, A2 => n10472, B1 => n10270, B2 => 
                           n8276, ZN => n1644);
   U8426 : OAI22_X1 port map( A1 => n10274, A2 => n10475, B1 => n10270, B2 => 
                           n8275, ZN => n1645);
   U8427 : OAI22_X1 port map( A1 => n10274, A2 => n10478, B1 => n10270, B2 => 
                           n8274, ZN => n1646);
   U8428 : OAI22_X1 port map( A1 => n10274, A2 => n10481, B1 => n10270, B2 => 
                           n8273, ZN => n1647);
   U8429 : OAI22_X1 port map( A1 => n10275, A2 => n10484, B1 => n10270, B2 => 
                           n8272, ZN => n1648);
   U8430 : OAI22_X1 port map( A1 => n10275, A2 => n10487, B1 => n10270, B2 => 
                           n8271, ZN => n1649);
   U8431 : OAI22_X1 port map( A1 => n10275, A2 => n10490, B1 => n10270, B2 => 
                           n8270, ZN => n1650);
   U8432 : OAI22_X1 port map( A1 => n10275, A2 => n10493, B1 => n10270, B2 => 
                           n8269, ZN => n1651);
   U8433 : OAI22_X1 port map( A1 => n10280, A2 => n10424, B1 => n10279, B2 => 
                           n8260, ZN => n1660);
   U8434 : OAI22_X1 port map( A1 => n10280, A2 => n10427, B1 => n10279, B2 => 
                           n8259, ZN => n1661);
   U8435 : OAI22_X1 port map( A1 => n10280, A2 => n10430, B1 => n10279, B2 => 
                           n8258, ZN => n1662);
   U8436 : OAI22_X1 port map( A1 => n10280, A2 => n10433, B1 => n10279, B2 => 
                           n8257, ZN => n1663);
   U8437 : OAI22_X1 port map( A1 => n10280, A2 => n10436, B1 => n10279, B2 => 
                           n8256, ZN => n1664);
   U8438 : OAI22_X1 port map( A1 => n10281, A2 => n10439, B1 => n10279, B2 => 
                           n8255, ZN => n1665);
   U8439 : OAI22_X1 port map( A1 => n10281, A2 => n10442, B1 => n10279, B2 => 
                           n8254, ZN => n1666);
   U8440 : OAI22_X1 port map( A1 => n10281, A2 => n10445, B1 => n10279, B2 => 
                           n8253, ZN => n1667);
   U8441 : OAI22_X1 port map( A1 => n10281, A2 => n10448, B1 => n10279, B2 => 
                           n8252, ZN => n1668);
   U8442 : OAI22_X1 port map( A1 => n10281, A2 => n10451, B1 => n10279, B2 => 
                           n8251, ZN => n1669);
   U8443 : OAI22_X1 port map( A1 => n10282, A2 => n10454, B1 => n10279, B2 => 
                           n8250, ZN => n1670);
   U8444 : OAI22_X1 port map( A1 => n10282, A2 => n10457, B1 => n10279, B2 => 
                           n8249, ZN => n1671);
   U8445 : OAI22_X1 port map( A1 => n10282, A2 => n10460, B1 => n8801, B2 => 
                           n8248, ZN => n1672);
   U8446 : OAI22_X1 port map( A1 => n10282, A2 => n10463, B1 => n8801, B2 => 
                           n8247, ZN => n1673);
   U8447 : OAI22_X1 port map( A1 => n10282, A2 => n10466, B1 => n8801, B2 => 
                           n8246, ZN => n1674);
   U8448 : OAI22_X1 port map( A1 => n10283, A2 => n10469, B1 => n10279, B2 => 
                           n8245, ZN => n1675);
   U8449 : OAI22_X1 port map( A1 => n10283, A2 => n10472, B1 => n10279, B2 => 
                           n8244, ZN => n1676);
   U8450 : OAI22_X1 port map( A1 => n10283, A2 => n10475, B1 => n10279, B2 => 
                           n8243, ZN => n1677);
   U8451 : OAI22_X1 port map( A1 => n10283, A2 => n10478, B1 => n10279, B2 => 
                           n8242, ZN => n1678);
   U8452 : OAI22_X1 port map( A1 => n10283, A2 => n10481, B1 => n10279, B2 => 
                           n8241, ZN => n1679);
   U8453 : OAI22_X1 port map( A1 => n10284, A2 => n10484, B1 => n10279, B2 => 
                           n8240, ZN => n1680);
   U8454 : OAI22_X1 port map( A1 => n10284, A2 => n10487, B1 => n10279, B2 => 
                           n8239, ZN => n1681);
   U8455 : OAI22_X1 port map( A1 => n10284, A2 => n10490, B1 => n10279, B2 => 
                           n8238, ZN => n1682);
   U8456 : OAI22_X1 port map( A1 => n10284, A2 => n10493, B1 => n10279, B2 => 
                           n8237, ZN => n1683);
   U8457 : OAI22_X1 port map( A1 => n8821, A2 => n8709, B1 => n10143, B2 => 
                           n10425, ZN => n1180);
   U8458 : AND4_X1 port map( A1 => n8888, A2 => n8889, A3 => n8890, A4 => n8891
                           , ZN => n8824);
   U8459 : OAI21_X1 port map( B1 => n8904, B2 => n8905, A => n10022, ZN => 
                           n8888);
   U8460 : OAI21_X1 port map( B1 => n8900, B2 => n8901, A => n10025, ZN => 
                           n8889);
   U8461 : OAI21_X1 port map( B1 => n8896, B2 => n8897, A => n10028, ZN => 
                           n8890);
   U8462 : AND4_X1 port map( A1 => n8856, A2 => n8857, A3 => n8858, A4 => n8859
                           , ZN => n8822);
   U8463 : OAI21_X1 port map( B1 => n8883, B2 => n8884, A => n10022, ZN => 
                           n8856);
   U8464 : OAI21_X1 port map( B1 => n8878, B2 => n8879, A => n10025, ZN => 
                           n8857);
   U8465 : OAI21_X1 port map( B1 => n8873, B2 => n8874, A => n10028, ZN => 
                           n8858);
   U8466 : AND4_X1 port map( A1 => n9488, A2 => n9489, A3 => n9490, A4 => n9491
                           , ZN => n8854);
   U8467 : OAI21_X1 port map( B1 => n9504, B2 => n9505, A => n10020, ZN => 
                           n9488);
   U8468 : OAI21_X1 port map( B1 => n9500, B2 => n9501, A => n10023, ZN => 
                           n9489);
   U8469 : OAI21_X1 port map( B1 => n9496, B2 => n9497, A => n10026, ZN => 
                           n9490);
   U8470 : AND4_X1 port map( A1 => n9468, A2 => n9469, A3 => n9470, A4 => n9471
                           , ZN => n8853);
   U8471 : OAI21_X1 port map( B1 => n9484, B2 => n9485, A => n10020, ZN => 
                           n9468);
   U8472 : OAI21_X1 port map( B1 => n9480, B2 => n9481, A => n10023, ZN => 
                           n9469);
   U8473 : OAI21_X1 port map( B1 => n9476, B2 => n9477, A => n10026, ZN => 
                           n9470);
   U8474 : AND4_X1 port map( A1 => n9448, A2 => n9449, A3 => n9450, A4 => n9451
                           , ZN => n8852);
   U8475 : OAI21_X1 port map( B1 => n9464, B2 => n9465, A => n10020, ZN => 
                           n9448);
   U8476 : OAI21_X1 port map( B1 => n9460, B2 => n9461, A => n10023, ZN => 
                           n9449);
   U8477 : OAI21_X1 port map( B1 => n9456, B2 => n9457, A => n10026, ZN => 
                           n9450);
   U8478 : AND4_X1 port map( A1 => n9428, A2 => n9429, A3 => n9430, A4 => n9431
                           , ZN => n8851);
   U8479 : OAI21_X1 port map( B1 => n9444, B2 => n9445, A => n10020, ZN => 
                           n9428);
   U8480 : OAI21_X1 port map( B1 => n9440, B2 => n9441, A => n10023, ZN => 
                           n9429);
   U8481 : OAI21_X1 port map( B1 => n9436, B2 => n9437, A => n10026, ZN => 
                           n9430);
   U8482 : AND4_X1 port map( A1 => n9408, A2 => n9409, A3 => n9410, A4 => n9411
                           , ZN => n8850);
   U8483 : OAI21_X1 port map( B1 => n9424, B2 => n9425, A => n10020, ZN => 
                           n9408);
   U8484 : OAI21_X1 port map( B1 => n9420, B2 => n9421, A => n10023, ZN => 
                           n9409);
   U8485 : OAI21_X1 port map( B1 => n9416, B2 => n9417, A => n10026, ZN => 
                           n9410);
   U8486 : AND4_X1 port map( A1 => n9388, A2 => n9389, A3 => n9390, A4 => n9391
                           , ZN => n8849);
   U8487 : OAI21_X1 port map( B1 => n9404, B2 => n9405, A => n10020, ZN => 
                           n9388);
   U8488 : OAI21_X1 port map( B1 => n9400, B2 => n9401, A => n10023, ZN => 
                           n9389);
   U8489 : OAI21_X1 port map( B1 => n9396, B2 => n9397, A => n10026, ZN => 
                           n9390);
   U8490 : AND4_X1 port map( A1 => n9368, A2 => n9369, A3 => n9370, A4 => n9371
                           , ZN => n8848);
   U8491 : OAI21_X1 port map( B1 => n9384, B2 => n9385, A => n10020, ZN => 
                           n9368);
   U8492 : OAI21_X1 port map( B1 => n9380, B2 => n9381, A => n10023, ZN => 
                           n9369);
   U8493 : OAI21_X1 port map( B1 => n9376, B2 => n9377, A => n10026, ZN => 
                           n9370);
   U8494 : AND4_X1 port map( A1 => n9348, A2 => n9349, A3 => n9350, A4 => n9351
                           , ZN => n8847);
   U8495 : OAI21_X1 port map( B1 => n9364, B2 => n9365, A => n10020, ZN => 
                           n9348);
   U8496 : OAI21_X1 port map( B1 => n9360, B2 => n9361, A => n10023, ZN => 
                           n9349);
   U8497 : OAI21_X1 port map( B1 => n9356, B2 => n9357, A => n10026, ZN => 
                           n9350);
   U8498 : AND4_X1 port map( A1 => n9328, A2 => n9329, A3 => n9330, A4 => n9331
                           , ZN => n8846);
   U8499 : OAI21_X1 port map( B1 => n9344, B2 => n9345, A => n10020, ZN => 
                           n9328);
   U8500 : OAI21_X1 port map( B1 => n9340, B2 => n9341, A => n10023, ZN => 
                           n9329);
   U8501 : OAI21_X1 port map( B1 => n9336, B2 => n9337, A => n10026, ZN => 
                           n9330);
   U8502 : AND4_X1 port map( A1 => n9308, A2 => n9309, A3 => n9310, A4 => n9311
                           , ZN => n8845);
   U8503 : OAI21_X1 port map( B1 => n9324, B2 => n9325, A => n10020, ZN => 
                           n9308);
   U8504 : OAI21_X1 port map( B1 => n9320, B2 => n9321, A => n10023, ZN => 
                           n9309);
   U8505 : OAI21_X1 port map( B1 => n9316, B2 => n9317, A => n10026, ZN => 
                           n9310);
   U8506 : AND4_X1 port map( A1 => n9288, A2 => n9289, A3 => n9290, A4 => n9291
                           , ZN => n8844);
   U8507 : OAI21_X1 port map( B1 => n9304, B2 => n9305, A => n10020, ZN => 
                           n9288);
   U8508 : OAI21_X1 port map( B1 => n9300, B2 => n9301, A => n10023, ZN => 
                           n9289);
   U8509 : OAI21_X1 port map( B1 => n9296, B2 => n9297, A => n10026, ZN => 
                           n9290);
   U8510 : AND4_X1 port map( A1 => n9268, A2 => n9269, A3 => n9270, A4 => n9271
                           , ZN => n8843);
   U8511 : OAI21_X1 port map( B1 => n9284, B2 => n9285, A => n10020, ZN => 
                           n9268);
   U8512 : OAI21_X1 port map( B1 => n9280, B2 => n9281, A => n10023, ZN => 
                           n9269);
   U8513 : OAI21_X1 port map( B1 => n9276, B2 => n9277, A => n10026, ZN => 
                           n9270);
   U8514 : AND4_X1 port map( A1 => n9248, A2 => n9249, A3 => n9250, A4 => n9251
                           , ZN => n8842);
   U8515 : OAI21_X1 port map( B1 => n9264, B2 => n9265, A => n10021, ZN => 
                           n9248);
   U8516 : OAI21_X1 port map( B1 => n9260, B2 => n9261, A => n10024, ZN => 
                           n9249);
   U8517 : OAI21_X1 port map( B1 => n9256, B2 => n9257, A => n10027, ZN => 
                           n9250);
   U8518 : AND4_X1 port map( A1 => n9228, A2 => n9229, A3 => n9230, A4 => n9231
                           , ZN => n8841);
   U8519 : OAI21_X1 port map( B1 => n9244, B2 => n9245, A => n10021, ZN => 
                           n9228);
   U8520 : OAI21_X1 port map( B1 => n9240, B2 => n9241, A => n10024, ZN => 
                           n9229);
   U8521 : OAI21_X1 port map( B1 => n9236, B2 => n9237, A => n10027, ZN => 
                           n9230);
   U8522 : AND4_X1 port map( A1 => n9208, A2 => n9209, A3 => n9210, A4 => n9211
                           , ZN => n8840);
   U8523 : OAI21_X1 port map( B1 => n9224, B2 => n9225, A => n10021, ZN => 
                           n9208);
   U8524 : OAI21_X1 port map( B1 => n9220, B2 => n9221, A => n10024, ZN => 
                           n9209);
   U8525 : OAI21_X1 port map( B1 => n9216, B2 => n9217, A => n10027, ZN => 
                           n9210);
   U8526 : AND4_X1 port map( A1 => n9188, A2 => n9189, A3 => n9190, A4 => n9191
                           , ZN => n8839);
   U8527 : OAI21_X1 port map( B1 => n9204, B2 => n9205, A => n10021, ZN => 
                           n9188);
   U8528 : OAI21_X1 port map( B1 => n9200, B2 => n9201, A => n10024, ZN => 
                           n9189);
   U8529 : OAI21_X1 port map( B1 => n9196, B2 => n9197, A => n10027, ZN => 
                           n9190);
   U8530 : AND4_X1 port map( A1 => n9168, A2 => n9169, A3 => n9170, A4 => n9171
                           , ZN => n8838);
   U8531 : OAI21_X1 port map( B1 => n9184, B2 => n9185, A => n10021, ZN => 
                           n9168);
   U8532 : OAI21_X1 port map( B1 => n9180, B2 => n9181, A => n10024, ZN => 
                           n9169);
   U8533 : OAI21_X1 port map( B1 => n9176, B2 => n9177, A => n10027, ZN => 
                           n9170);
   U8534 : AND4_X1 port map( A1 => n9148, A2 => n9149, A3 => n9150, A4 => n9151
                           , ZN => n8837);
   U8535 : OAI21_X1 port map( B1 => n9164, B2 => n9165, A => n10021, ZN => 
                           n9148);
   U8536 : OAI21_X1 port map( B1 => n9160, B2 => n9161, A => n10024, ZN => 
                           n9149);
   U8537 : OAI21_X1 port map( B1 => n9156, B2 => n9157, A => n10027, ZN => 
                           n9150);
   U8538 : AND4_X1 port map( A1 => n9128, A2 => n9129, A3 => n9130, A4 => n9131
                           , ZN => n8836);
   U8539 : OAI21_X1 port map( B1 => n9144, B2 => n9145, A => n10021, ZN => 
                           n9128);
   U8540 : OAI21_X1 port map( B1 => n9140, B2 => n9141, A => n10024, ZN => 
                           n9129);
   U8541 : OAI21_X1 port map( B1 => n9136, B2 => n9137, A => n10027, ZN => 
                           n9130);
   U8542 : AND4_X1 port map( A1 => n9108, A2 => n9109, A3 => n9110, A4 => n9111
                           , ZN => n8835);
   U8543 : OAI21_X1 port map( B1 => n9124, B2 => n9125, A => n10021, ZN => 
                           n9108);
   U8544 : OAI21_X1 port map( B1 => n9120, B2 => n9121, A => n10024, ZN => 
                           n9109);
   U8545 : OAI21_X1 port map( B1 => n9116, B2 => n9117, A => n10027, ZN => 
                           n9110);
   U8546 : AND4_X1 port map( A1 => n9088, A2 => n9089, A3 => n9090, A4 => n9091
                           , ZN => n8834);
   U8547 : OAI21_X1 port map( B1 => n9104, B2 => n9105, A => n10021, ZN => 
                           n9088);
   U8548 : OAI21_X1 port map( B1 => n9100, B2 => n9101, A => n10024, ZN => 
                           n9089);
   U8549 : OAI21_X1 port map( B1 => n9096, B2 => n9097, A => n10027, ZN => 
                           n9090);
   U8550 : AND4_X1 port map( A1 => n9068, A2 => n9069, A3 => n9070, A4 => n9071
                           , ZN => n8833);
   U8551 : OAI21_X1 port map( B1 => n9084, B2 => n9085, A => n10021, ZN => 
                           n9068);
   U8552 : OAI21_X1 port map( B1 => n9080, B2 => n9081, A => n10024, ZN => 
                           n9069);
   U8553 : OAI21_X1 port map( B1 => n9076, B2 => n9077, A => n10027, ZN => 
                           n9070);
   U8554 : AND4_X1 port map( A1 => n9048, A2 => n9049, A3 => n9050, A4 => n9051
                           , ZN => n8832);
   U8555 : OAI21_X1 port map( B1 => n9064, B2 => n9065, A => n10021, ZN => 
                           n9048);
   U8556 : OAI21_X1 port map( B1 => n9060, B2 => n9061, A => n10024, ZN => 
                           n9049);
   U8557 : OAI21_X1 port map( B1 => n9056, B2 => n9057, A => n10027, ZN => 
                           n9050);
   U8558 : AND4_X1 port map( A1 => n9028, A2 => n9029, A3 => n9030, A4 => n9031
                           , ZN => n8831);
   U8559 : OAI21_X1 port map( B1 => n9044, B2 => n9045, A => n10021, ZN => 
                           n9028);
   U8560 : OAI21_X1 port map( B1 => n9040, B2 => n9041, A => n10024, ZN => 
                           n9029);
   U8561 : OAI21_X1 port map( B1 => n9036, B2 => n9037, A => n10027, ZN => 
                           n9030);
   U8562 : AND4_X1 port map( A1 => n9008, A2 => n9009, A3 => n9010, A4 => n9011
                           , ZN => n8830);
   U8563 : OAI21_X1 port map( B1 => n9024, B2 => n9025, A => n10022, ZN => 
                           n9008);
   U8564 : OAI21_X1 port map( B1 => n9020, B2 => n9021, A => n10025, ZN => 
                           n9009);
   U8565 : OAI21_X1 port map( B1 => n9016, B2 => n9017, A => n10028, ZN => 
                           n9010);
   U8566 : AND4_X1 port map( A1 => n8988, A2 => n8989, A3 => n8990, A4 => n8991
                           , ZN => n8829);
   U8567 : OAI21_X1 port map( B1 => n9004, B2 => n9005, A => n10022, ZN => 
                           n8988);
   U8568 : OAI21_X1 port map( B1 => n9000, B2 => n9001, A => n10025, ZN => 
                           n8989);
   U8569 : OAI21_X1 port map( B1 => n8996, B2 => n8997, A => n10028, ZN => 
                           n8990);
   U8570 : AND4_X1 port map( A1 => n8968, A2 => n8969, A3 => n8970, A4 => n8971
                           , ZN => n8828);
   U8571 : OAI21_X1 port map( B1 => n8984, B2 => n8985, A => n10022, ZN => 
                           n8968);
   U8572 : OAI21_X1 port map( B1 => n8980, B2 => n8981, A => n10025, ZN => 
                           n8969);
   U8573 : OAI21_X1 port map( B1 => n8976, B2 => n8977, A => n10028, ZN => 
                           n8970);
   U8574 : AND4_X1 port map( A1 => n8948, A2 => n8949, A3 => n8950, A4 => n8951
                           , ZN => n8827);
   U8575 : OAI21_X1 port map( B1 => n8964, B2 => n8965, A => n10022, ZN => 
                           n8948);
   U8576 : OAI21_X1 port map( B1 => n8960, B2 => n8961, A => n10025, ZN => 
                           n8949);
   U8577 : OAI21_X1 port map( B1 => n8956, B2 => n8957, A => n10028, ZN => 
                           n8950);
   U8578 : AND4_X1 port map( A1 => n8928, A2 => n8929, A3 => n8930, A4 => n8931
                           , ZN => n8826);
   U8579 : OAI21_X1 port map( B1 => n8944, B2 => n8945, A => n10022, ZN => 
                           n8928);
   U8580 : OAI21_X1 port map( B1 => n8940, B2 => n8941, A => n10025, ZN => 
                           n8929);
   U8581 : OAI21_X1 port map( B1 => n8936, B2 => n8937, A => n10028, ZN => 
                           n8930);
   U8582 : AND4_X1 port map( A1 => n8908, A2 => n8909, A3 => n8910, A4 => n8911
                           , ZN => n8825);
   U8583 : OAI21_X1 port map( B1 => n8924, B2 => n8925, A => n10022, ZN => 
                           n8908);
   U8584 : OAI21_X1 port map( B1 => n8920, B2 => n8921, A => n10025, ZN => 
                           n8909);
   U8585 : OAI21_X1 port map( B1 => n8916, B2 => n8917, A => n10028, ZN => 
                           n8910);
   U8586 : NAND2_X1 port map( A1 => n7745, A2 => n7746, ZN => n8778);
   U8587 : BUF_X1 port map( A => n8862, Z => n10133);
   U8588 : BUF_X1 port map( A => n8875, Z => n10026);
   U8589 : BUF_X1 port map( A => n8880, Z => n10023);
   U8590 : BUF_X1 port map( A => n8862, Z => n10134);
   U8591 : BUF_X1 port map( A => n8875, Z => n10027);
   U8592 : BUF_X1 port map( A => n8880, Z => n10024);
   U8593 : BUF_X1 port map( A => n7741, Z => n10532);
   U8594 : BUF_X1 port map( A => n7741, Z => n10531);
   U8595 : BUF_X1 port map( A => n7741, Z => n10529);
   U8596 : BUF_X1 port map( A => n7741, Z => n10528);
   U8597 : BUF_X1 port map( A => n8752, Z => n10496);
   U8598 : BUF_X1 port map( A => n8751, Z => n10499);
   U8599 : BUF_X1 port map( A => n8750, Z => n10502);
   U8600 : BUF_X1 port map( A => n8749, Z => n10505);
   U8601 : BUF_X1 port map( A => n8748, Z => n10508);
   U8602 : BUF_X1 port map( A => n8747, Z => n10511);
   U8603 : BUF_X1 port map( A => n8746, Z => n10514);
   U8604 : BUF_X1 port map( A => n8744, Z => n10526);
   U8605 : BUF_X1 port map( A => n8776, Z => n10424);
   U8606 : BUF_X1 port map( A => n8775, Z => n10427);
   U8607 : BUF_X1 port map( A => n8774, Z => n10430);
   U8608 : BUF_X1 port map( A => n8773, Z => n10433);
   U8609 : BUF_X1 port map( A => n8772, Z => n10436);
   U8610 : BUF_X1 port map( A => n8771, Z => n10439);
   U8611 : BUF_X1 port map( A => n8770, Z => n10442);
   U8612 : BUF_X1 port map( A => n8769, Z => n10445);
   U8613 : BUF_X1 port map( A => n8768, Z => n10448);
   U8614 : BUF_X1 port map( A => n8767, Z => n10451);
   U8615 : BUF_X1 port map( A => n8766, Z => n10454);
   U8616 : BUF_X1 port map( A => n8765, Z => n10457);
   U8617 : BUF_X1 port map( A => n8764, Z => n10460);
   U8618 : BUF_X1 port map( A => n8763, Z => n10463);
   U8619 : BUF_X1 port map( A => n8762, Z => n10466);
   U8620 : BUF_X1 port map( A => n8761, Z => n10469);
   U8621 : BUF_X1 port map( A => n8760, Z => n10472);
   U8622 : BUF_X1 port map( A => n8759, Z => n10475);
   U8623 : BUF_X1 port map( A => n8758, Z => n10478);
   U8624 : BUF_X1 port map( A => n8757, Z => n10481);
   U8625 : BUF_X1 port map( A => n8756, Z => n10484);
   U8626 : BUF_X1 port map( A => n8755, Z => n10487);
   U8627 : BUF_X1 port map( A => n8754, Z => n10490);
   U8628 : BUF_X1 port map( A => n8753, Z => n10493);
   U8629 : BUF_X1 port map( A => n8776, Z => n10423);
   U8630 : BUF_X1 port map( A => n8775, Z => n10426);
   U8631 : BUF_X1 port map( A => n8774, Z => n10429);
   U8632 : BUF_X1 port map( A => n8773, Z => n10432);
   U8633 : BUF_X1 port map( A => n8772, Z => n10435);
   U8634 : BUF_X1 port map( A => n8771, Z => n10438);
   U8635 : BUF_X1 port map( A => n8770, Z => n10441);
   U8636 : BUF_X1 port map( A => n8769, Z => n10444);
   U8637 : BUF_X1 port map( A => n8768, Z => n10447);
   U8638 : BUF_X1 port map( A => n8767, Z => n10450);
   U8639 : BUF_X1 port map( A => n8766, Z => n10453);
   U8640 : BUF_X1 port map( A => n8765, Z => n10456);
   U8641 : BUF_X1 port map( A => n8764, Z => n10459);
   U8642 : BUF_X1 port map( A => n8763, Z => n10462);
   U8643 : BUF_X1 port map( A => n8762, Z => n10465);
   U8644 : BUF_X1 port map( A => n8761, Z => n10468);
   U8645 : BUF_X1 port map( A => n8760, Z => n10471);
   U8646 : BUF_X1 port map( A => n8759, Z => n10474);
   U8647 : BUF_X1 port map( A => n8758, Z => n10477);
   U8648 : BUF_X1 port map( A => n8757, Z => n10480);
   U8649 : BUF_X1 port map( A => n8756, Z => n10483);
   U8650 : BUF_X1 port map( A => n8755, Z => n10486);
   U8651 : BUF_X1 port map( A => n8754, Z => n10489);
   U8652 : BUF_X1 port map( A => n8753, Z => n10492);
   U8653 : BUF_X1 port map( A => n8752, Z => n10495);
   U8654 : BUF_X1 port map( A => n8751, Z => n10498);
   U8655 : BUF_X1 port map( A => n8750, Z => n10501);
   U8656 : BUF_X1 port map( A => n8749, Z => n10504);
   U8657 : BUF_X1 port map( A => n8748, Z => n10507);
   U8658 : BUF_X1 port map( A => n8747, Z => n10510);
   U8659 : BUF_X1 port map( A => n8746, Z => n10513);
   U8660 : BUF_X1 port map( A => n8744, Z => n10525);
   U8661 : BUF_X1 port map( A => n7741, Z => n10530);
   U8662 : BUF_X1 port map( A => n8855, Z => n10136);
   U8663 : BUF_X1 port map( A => n8855, Z => n10137);
   U8664 : BUF_X1 port map( A => n8823, Z => n10139);
   U8665 : BUF_X1 port map( A => n8823, Z => n10140);
   U8666 : BUF_X1 port map( A => n8776, Z => n10425);
   U8667 : BUF_X1 port map( A => n8775, Z => n10428);
   U8668 : BUF_X1 port map( A => n8774, Z => n10431);
   U8669 : BUF_X1 port map( A => n8773, Z => n10434);
   U8670 : BUF_X1 port map( A => n8772, Z => n10437);
   U8671 : BUF_X1 port map( A => n8771, Z => n10440);
   U8672 : BUF_X1 port map( A => n8770, Z => n10443);
   U8673 : BUF_X1 port map( A => n8769, Z => n10446);
   U8674 : BUF_X1 port map( A => n8768, Z => n10449);
   U8675 : BUF_X1 port map( A => n8767, Z => n10452);
   U8676 : BUF_X1 port map( A => n8766, Z => n10455);
   U8677 : BUF_X1 port map( A => n8765, Z => n10458);
   U8678 : BUF_X1 port map( A => n8764, Z => n10461);
   U8679 : BUF_X1 port map( A => n8763, Z => n10464);
   U8680 : BUF_X1 port map( A => n8762, Z => n10467);
   U8681 : BUF_X1 port map( A => n8761, Z => n10470);
   U8682 : BUF_X1 port map( A => n8760, Z => n10473);
   U8683 : BUF_X1 port map( A => n8759, Z => n10476);
   U8684 : BUF_X1 port map( A => n8758, Z => n10479);
   U8685 : BUF_X1 port map( A => n8757, Z => n10482);
   U8686 : BUF_X1 port map( A => n8756, Z => n10485);
   U8687 : BUF_X1 port map( A => n8755, Z => n10488);
   U8688 : BUF_X1 port map( A => n8754, Z => n10491);
   U8689 : BUF_X1 port map( A => n8753, Z => n10494);
   U8690 : BUF_X1 port map( A => n8752, Z => n10497);
   U8691 : BUF_X1 port map( A => n8751, Z => n10500);
   U8692 : BUF_X1 port map( A => n8750, Z => n10503);
   U8693 : BUF_X1 port map( A => n8749, Z => n10506);
   U8694 : BUF_X1 port map( A => n8748, Z => n10509);
   U8695 : BUF_X1 port map( A => n8747, Z => n10512);
   U8696 : BUF_X1 port map( A => n8746, Z => n10515);
   U8697 : BUF_X1 port map( A => n8744, Z => n10527);
   U8698 : BUF_X1 port map( A => n8855, Z => n10138);
   U8699 : BUF_X1 port map( A => n8823, Z => n10141);
   U8700 : BUF_X1 port map( A => n8862, Z => n10135);
   U8701 : BUF_X1 port map( A => n8875, Z => n10028);
   U8702 : BUF_X1 port map( A => n8880, Z => n10025);
   U8703 : BUF_X1 port map( A => n8866, Z => n10094);
   U8704 : BUF_X1 port map( A => n8867, Z => n10081);
   U8705 : BUF_X1 port map( A => n8871, Z => n10042);
   U8706 : BUF_X1 port map( A => n8872, Z => n10029);
   U8707 : BUF_X1 port map( A => n8864, Z => n10107);
   U8708 : BUF_X1 port map( A => n8863, Z => n10120);
   U8709 : BUF_X1 port map( A => n8869, Z => n10055);
   U8710 : BUF_X1 port map( A => n8868, Z => n10068);
   U8711 : NOR2_X1 port map( A1 => n7750, A2 => n7749, ZN => n8885);
   U8712 : BUF_X1 port map( A => n8866, Z => n10095);
   U8713 : BUF_X1 port map( A => n8867, Z => n10082);
   U8714 : BUF_X1 port map( A => n8871, Z => n10043);
   U8715 : BUF_X1 port map( A => n8872, Z => n10030);
   U8716 : BUF_X1 port map( A => n8864, Z => n10108);
   U8717 : BUF_X1 port map( A => n8863, Z => n10121);
   U8718 : BUF_X1 port map( A => n8869, Z => n10056);
   U8719 : BUF_X1 port map( A => n8868, Z => n10069);
   U8720 : BUF_X1 port map( A => n8821, Z => n10142);
   U8721 : OAI21_X1 port map( B1 => n8784, B2 => n8818, A => n10532, ZN => 
                           n8821);
   U8722 : INV_X1 port map( A => n8783, ZN => n10404);
   U8723 : OAI21_X1 port map( B1 => n8777, B2 => n8784, A => n10532, ZN => 
                           n8783);
   U8724 : INV_X1 port map( A => n8781, ZN => n10413);
   U8725 : OAI21_X1 port map( B1 => n8777, B2 => n8782, A => n10532, ZN => 
                           n8781);
   U8726 : INV_X1 port map( A => n8779, ZN => n10422);
   U8727 : OAI21_X1 port map( B1 => n8777, B2 => n8780, A => n10533, ZN => 
                           n8779);
   U8728 : INV_X1 port map( A => n8820, ZN => n10161);
   U8729 : OAI21_X1 port map( B1 => n8782, B2 => n8818, A => n10530, ZN => 
                           n8820);
   U8730 : INV_X1 port map( A => n8819, ZN => n10170);
   U8731 : OAI21_X1 port map( B1 => n8780, B2 => n8818, A => n10530, ZN => 
                           n8819);
   U8732 : INV_X1 port map( A => n8817, ZN => n10179);
   U8733 : OAI21_X1 port map( B1 => n8778, B2 => n8818, A => n10530, ZN => 
                           n8817);
   U8734 : INV_X1 port map( A => n8816, ZN => n10188);
   U8735 : OAI21_X1 port map( B1 => n8784, B2 => n8813, A => n10531, ZN => 
                           n8816);
   U8736 : INV_X1 port map( A => n8815, ZN => n10197);
   U8737 : OAI21_X1 port map( B1 => n8782, B2 => n8813, A => n10530, ZN => 
                           n8815);
   U8738 : INV_X1 port map( A => n8814, ZN => n10206);
   U8739 : OAI21_X1 port map( B1 => n8780, B2 => n8813, A => n10531, ZN => 
                           n8814);
   U8740 : INV_X1 port map( A => n8812, ZN => n10215);
   U8741 : OAI21_X1 port map( B1 => n8778, B2 => n8813, A => n10531, ZN => 
                           n8812);
   U8742 : INV_X1 port map( A => n8811, ZN => n10224);
   U8743 : OAI21_X1 port map( B1 => n8784, B2 => n8808, A => n10531, ZN => 
                           n8811);
   U8744 : INV_X1 port map( A => n8810, ZN => n10233);
   U8745 : OAI21_X1 port map( B1 => n8782, B2 => n8808, A => n10531, ZN => 
                           n8810);
   U8746 : INV_X1 port map( A => n8809, ZN => n10242);
   U8747 : OAI21_X1 port map( B1 => n8780, B2 => n8808, A => n10531, ZN => 
                           n8809);
   U8748 : INV_X1 port map( A => n8807, ZN => n10251);
   U8749 : OAI21_X1 port map( B1 => n8778, B2 => n8808, A => n10531, ZN => 
                           n8807);
   U8750 : INV_X1 port map( A => n8805, ZN => n10260);
   U8751 : OAI21_X1 port map( B1 => n8784, B2 => n8802, A => n10531, ZN => 
                           n8805);
   U8752 : INV_X1 port map( A => n8804, ZN => n10269);
   U8753 : OAI21_X1 port map( B1 => n8782, B2 => n8802, A => n10531, ZN => 
                           n8804);
   U8754 : INV_X1 port map( A => n8803, ZN => n10278);
   U8755 : OAI21_X1 port map( B1 => n8780, B2 => n8802, A => n10531, ZN => 
                           n8803);
   U8756 : INV_X1 port map( A => n8800, ZN => n10296);
   U8757 : OAI21_X1 port map( B1 => n8784, B2 => n8797, A => n10531, ZN => 
                           n8800);
   U8758 : INV_X1 port map( A => n8799, ZN => n10305);
   U8759 : OAI21_X1 port map( B1 => n8782, B2 => n8797, A => n10531, ZN => 
                           n8799);
   U8760 : INV_X1 port map( A => n8798, ZN => n10314);
   U8761 : OAI21_X1 port map( B1 => n8780, B2 => n8797, A => n10532, ZN => 
                           n8798);
   U8762 : INV_X1 port map( A => n8796, ZN => n10323);
   U8763 : OAI21_X1 port map( B1 => n8778, B2 => n8797, A => n10532, ZN => 
                           n8796);
   U8764 : INV_X1 port map( A => n8795, ZN => n10332);
   U8765 : OAI21_X1 port map( B1 => n8784, B2 => n8792, A => n10532, ZN => 
                           n8795);
   U8766 : INV_X1 port map( A => n8794, ZN => n10341);
   U8767 : OAI21_X1 port map( B1 => n8782, B2 => n8792, A => n10532, ZN => 
                           n8794);
   U8768 : INV_X1 port map( A => n8793, ZN => n10350);
   U8769 : OAI21_X1 port map( B1 => n8780, B2 => n8792, A => n10532, ZN => 
                           n8793);
   U8770 : INV_X1 port map( A => n8791, ZN => n10359);
   U8771 : OAI21_X1 port map( B1 => n8778, B2 => n8792, A => n10532, ZN => 
                           n8791);
   U8772 : INV_X1 port map( A => n8790, ZN => n10368);
   U8773 : OAI21_X1 port map( B1 => n8784, B2 => n8787, A => n10532, ZN => 
                           n8790);
   U8774 : INV_X1 port map( A => n8789, ZN => n10377);
   U8775 : OAI21_X1 port map( B1 => n8782, B2 => n8787, A => n10532, ZN => 
                           n8789);
   U8776 : INV_X1 port map( A => n8788, ZN => n10386);
   U8777 : OAI21_X1 port map( B1 => n8780, B2 => n8787, A => n10532, ZN => 
                           n8788);
   U8778 : INV_X1 port map( A => n8786, ZN => n10395);
   U8779 : OAI21_X1 port map( B1 => n8778, B2 => n8787, A => n10532, ZN => 
                           n8786);
   U8780 : OAI21_X1 port map( B1 => n8892, B2 => n8893, A => n10135, ZN => 
                           n8891);
   U8781 : OAI221_X1 port map( B1 => n8550, B2 => n10080, C1 => n8294, C2 => 
                           n10067, A => n8895, ZN => n8892);
   U8782 : OAI221_X1 port map( B1 => n8678, B2 => n10132, C1 => n8422, C2 => 
                           n10119, A => n8894, ZN => n8893);
   U8783 : AOI22_X1 port map( A1 => n10054, A2 => n9548, B1 => n10041, B2 => 
                           n9600, ZN => n8895);
   U8784 : OAI21_X1 port map( B1 => n8860, B2 => n8861, A => n10135, ZN => 
                           n8859);
   U8785 : OAI221_X1 port map( B1 => n8549, B2 => n10080, C1 => n8293, C2 => 
                           n10067, A => n8870, ZN => n8860);
   U8786 : OAI221_X1 port map( B1 => n8677, B2 => n10132, C1 => n8421, C2 => 
                           n10119, A => n8865, ZN => n8861);
   U8787 : AOI22_X1 port map( A1 => n10054, A2 => n9549, B1 => n10041, B2 => 
                           n9601, ZN => n8870);
   U8788 : OAI221_X1 port map( B1 => n6712, B2 => n10122, C1 => n8483, C2 => 
                           n10109, A => n9486, ZN => n9485);
   U8789 : AOI22_X1 port map( A1 => n10096, A2 => n9613, B1 => n10083, B2 => 
                           n9757, ZN => n9486);
   U8790 : OAI221_X1 port map( B1 => n6711, B2 => n10122, C1 => n8482, C2 => 
                           n10109, A => n9466, ZN => n9465);
   U8791 : AOI22_X1 port map( A1 => n10096, A2 => n9614, B1 => n10083, B2 => 
                           n9758, ZN => n9466);
   U8792 : OAI221_X1 port map( B1 => n6710, B2 => n10123, C1 => n8481, C2 => 
                           n10110, A => n9446, ZN => n9445);
   U8793 : AOI22_X1 port map( A1 => n10097, A2 => n9615, B1 => n10084, B2 => 
                           n9759, ZN => n9446);
   U8794 : OAI221_X1 port map( B1 => n6709, B2 => n10123, C1 => n8480, C2 => 
                           n10110, A => n9426, ZN => n9425);
   U8795 : AOI22_X1 port map( A1 => n10097, A2 => n9616, B1 => n10084, B2 => 
                           n9760, ZN => n9426);
   U8796 : OAI221_X1 port map( B1 => n6708, B2 => n10123, C1 => n8479, C2 => 
                           n10110, A => n9406, ZN => n9405);
   U8797 : AOI22_X1 port map( A1 => n10097, A2 => n9617, B1 => n10084, B2 => 
                           n9761, ZN => n9406);
   U8798 : OAI221_X1 port map( B1 => n6707, B2 => n10124, C1 => n8478, C2 => 
                           n10111, A => n9386, ZN => n9385);
   U8799 : AOI22_X1 port map( A1 => n10098, A2 => n9618, B1 => n10085, B2 => 
                           n9762, ZN => n9386);
   U8800 : OAI221_X1 port map( B1 => n6706, B2 => n10124, C1 => n8477, C2 => 
                           n10111, A => n9366, ZN => n9365);
   U8801 : AOI22_X1 port map( A1 => n10098, A2 => n9619, B1 => n10085, B2 => 
                           n9763, ZN => n9366);
   U8802 : OAI221_X1 port map( B1 => n6705, B2 => n10124, C1 => n8476, C2 => 
                           n10111, A => n9346, ZN => n9345);
   U8803 : AOI22_X1 port map( A1 => n10098, A2 => n9620, B1 => n10085, B2 => 
                           n9764, ZN => n9346);
   U8804 : OAI221_X1 port map( B1 => n6704, B2 => n10125, C1 => n8475, C2 => 
                           n10112, A => n9326, ZN => n9325);
   U8805 : AOI22_X1 port map( A1 => n10099, A2 => n9621, B1 => n10086, B2 => 
                           n9765, ZN => n9326);
   U8806 : OAI221_X1 port map( B1 => n6703, B2 => n10125, C1 => n8474, C2 => 
                           n10112, A => n9306, ZN => n9305);
   U8807 : AOI22_X1 port map( A1 => n10099, A2 => n9622, B1 => n10086, B2 => 
                           n9766, ZN => n9306);
   U8808 : OAI221_X1 port map( B1 => n6702, B2 => n10125, C1 => n8473, C2 => 
                           n10112, A => n9286, ZN => n9285);
   U8809 : AOI22_X1 port map( A1 => n10099, A2 => n9623, B1 => n10086, B2 => 
                           n9767, ZN => n9286);
   U8810 : OAI221_X1 port map( B1 => n6701, B2 => n10126, C1 => n8472, C2 => 
                           n10113, A => n9266, ZN => n9265);
   U8811 : AOI22_X1 port map( A1 => n10100, A2 => n9624, B1 => n10087, B2 => 
                           n9768, ZN => n9266);
   U8812 : OAI221_X1 port map( B1 => n6700, B2 => n10126, C1 => n8471, C2 => 
                           n10113, A => n9246, ZN => n9245);
   U8813 : AOI22_X1 port map( A1 => n10100, A2 => n9625, B1 => n10087, B2 => 
                           n9769, ZN => n9246);
   U8814 : OAI221_X1 port map( B1 => n6699, B2 => n10126, C1 => n8470, C2 => 
                           n10113, A => n9226, ZN => n9225);
   U8815 : AOI22_X1 port map( A1 => n10100, A2 => n9626, B1 => n10087, B2 => 
                           n9770, ZN => n9226);
   U8816 : OAI221_X1 port map( B1 => n6698, B2 => n10127, C1 => n8469, C2 => 
                           n10114, A => n9206, ZN => n9205);
   U8817 : AOI22_X1 port map( A1 => n10101, A2 => n9627, B1 => n10088, B2 => 
                           n9771, ZN => n9206);
   U8818 : OAI221_X1 port map( B1 => n6697, B2 => n10127, C1 => n8468, C2 => 
                           n10114, A => n9186, ZN => n9185);
   U8819 : AOI22_X1 port map( A1 => n10101, A2 => n9628, B1 => n10088, B2 => 
                           n9772, ZN => n9186);
   U8820 : OAI221_X1 port map( B1 => n6696, B2 => n10127, C1 => n8467, C2 => 
                           n10114, A => n9166, ZN => n9165);
   U8821 : AOI22_X1 port map( A1 => n10101, A2 => n9629, B1 => n10088, B2 => 
                           n9773, ZN => n9166);
   U8822 : OAI221_X1 port map( B1 => n6695, B2 => n10128, C1 => n8466, C2 => 
                           n10115, A => n9146, ZN => n9145);
   U8823 : AOI22_X1 port map( A1 => n10102, A2 => n9630, B1 => n10089, B2 => 
                           n9774, ZN => n9146);
   U8824 : OAI221_X1 port map( B1 => n6694, B2 => n10128, C1 => n8465, C2 => 
                           n10115, A => n9126, ZN => n9125);
   U8825 : AOI22_X1 port map( A1 => n10102, A2 => n9631, B1 => n10089, B2 => 
                           n9775, ZN => n9126);
   U8826 : OAI221_X1 port map( B1 => n6693, B2 => n10128, C1 => n8464, C2 => 
                           n10115, A => n9106, ZN => n9105);
   U8827 : AOI22_X1 port map( A1 => n10102, A2 => n9632, B1 => n10089, B2 => 
                           n9776, ZN => n9106);
   U8828 : OAI221_X1 port map( B1 => n6692, B2 => n10129, C1 => n8463, C2 => 
                           n10116, A => n9086, ZN => n9085);
   U8829 : AOI22_X1 port map( A1 => n10103, A2 => n9633, B1 => n10090, B2 => 
                           n9777, ZN => n9086);
   U8830 : OAI221_X1 port map( B1 => n6691, B2 => n10129, C1 => n8462, C2 => 
                           n10116, A => n9066, ZN => n9065);
   U8831 : AOI22_X1 port map( A1 => n10103, A2 => n9634, B1 => n10090, B2 => 
                           n9778, ZN => n9066);
   U8832 : OAI221_X1 port map( B1 => n6690, B2 => n10129, C1 => n8461, C2 => 
                           n10116, A => n9046, ZN => n9045);
   U8833 : AOI22_X1 port map( A1 => n10103, A2 => n9635, B1 => n10090, B2 => 
                           n9779, ZN => n9046);
   U8834 : OAI221_X1 port map( B1 => n6689, B2 => n10130, C1 => n8460, C2 => 
                           n10117, A => n9026, ZN => n9025);
   U8835 : AOI22_X1 port map( A1 => n10104, A2 => n9508, B1 => n10091, B2 => 
                           n9560, ZN => n9026);
   U8836 : OAI221_X1 port map( B1 => n6688, B2 => n10130, C1 => n8459, C2 => 
                           n10117, A => n9006, ZN => n9005);
   U8837 : AOI22_X1 port map( A1 => n10104, A2 => n9509, B1 => n10091, B2 => 
                           n9561, ZN => n9006);
   U8838 : OAI221_X1 port map( B1 => n6687, B2 => n10130, C1 => n8458, C2 => 
                           n10117, A => n8986, ZN => n8985);
   U8839 : AOI22_X1 port map( A1 => n10104, A2 => n9510, B1 => n10091, B2 => 
                           n9562, ZN => n8986);
   U8840 : OAI221_X1 port map( B1 => n6686, B2 => n10131, C1 => n8457, C2 => 
                           n10118, A => n8966, ZN => n8965);
   U8841 : AOI22_X1 port map( A1 => n10105, A2 => n9511, B1 => n10092, B2 => 
                           n9563, ZN => n8966);
   U8842 : OAI221_X1 port map( B1 => n6685, B2 => n10131, C1 => n8456, C2 => 
                           n10118, A => n8946, ZN => n8945);
   U8843 : AOI22_X1 port map( A1 => n10105, A2 => n9512, B1 => n10092, B2 => 
                           n9564, ZN => n8946);
   U8844 : OAI221_X1 port map( B1 => n6684, B2 => n10131, C1 => n8455, C2 => 
                           n10118, A => n8926, ZN => n8925);
   U8845 : AOI22_X1 port map( A1 => n10105, A2 => n9513, B1 => n10092, B2 => 
                           n9565, ZN => n8926);
   U8846 : OAI221_X1 port map( B1 => n8676, B2 => n10122, C1 => n8420, C2 => 
                           n10109, A => n9498, ZN => n9497);
   U8847 : AOI22_X1 port map( A1 => n10096, A2 => n9660, B1 => n10083, B2 => 
                           n9804, ZN => n9498);
   U8848 : OAI221_X1 port map( B1 => n8644, B2 => n10122, C1 => n8388, C2 => 
                           n10109, A => n9502, ZN => n9501);
   U8849 : AOI22_X1 port map( A1 => n10096, A2 => n9902, B1 => n10083, B2 => 
                           n9903, ZN => n9502);
   U8850 : OAI221_X1 port map( B1 => n8709, B2 => n10122, C1 => n8484, C2 => 
                           n10109, A => n9506, ZN => n9505);
   U8851 : AOI22_X1 port map( A1 => n10096, A2 => n9612, B1 => n10083, B2 => 
                           n9756, ZN => n9506);
   U8852 : OAI221_X1 port map( B1 => n8675, B2 => n10122, C1 => n8419, C2 => 
                           n10109, A => n9478, ZN => n9477);
   U8853 : AOI22_X1 port map( A1 => n10096, A2 => n9661, B1 => n10083, B2 => 
                           n9805, ZN => n9478);
   U8854 : OAI221_X1 port map( B1 => n8643, B2 => n10122, C1 => n8387, C2 => 
                           n10109, A => n9482, ZN => n9481);
   U8855 : AOI22_X1 port map( A1 => n10096, A2 => n9906, B1 => n10083, B2 => 
                           n9907, ZN => n9482);
   U8856 : OAI221_X1 port map( B1 => n8674, B2 => n10122, C1 => n8418, C2 => 
                           n10109, A => n9458, ZN => n9457);
   U8857 : AOI22_X1 port map( A1 => n10096, A2 => n9662, B1 => n10083, B2 => 
                           n9806, ZN => n9458);
   U8858 : OAI221_X1 port map( B1 => n8642, B2 => n10122, C1 => n8386, C2 => 
                           n10109, A => n9462, ZN => n9461);
   U8859 : AOI22_X1 port map( A1 => n10096, A2 => n9910, B1 => n10083, B2 => 
                           n9911, ZN => n9462);
   U8860 : OAI221_X1 port map( B1 => n8673, B2 => n10123, C1 => n8417, C2 => 
                           n10110, A => n9438, ZN => n9437);
   U8861 : AOI22_X1 port map( A1 => n10097, A2 => n9663, B1 => n10084, B2 => 
                           n9807, ZN => n9438);
   U8862 : OAI221_X1 port map( B1 => n8641, B2 => n10123, C1 => n8385, C2 => 
                           n10110, A => n9442, ZN => n9441);
   U8863 : AOI22_X1 port map( A1 => n10097, A2 => n9914, B1 => n10084, B2 => 
                           n9915, ZN => n9442);
   U8864 : OAI221_X1 port map( B1 => n8672, B2 => n10123, C1 => n8416, C2 => 
                           n10110, A => n9418, ZN => n9417);
   U8865 : AOI22_X1 port map( A1 => n10097, A2 => n9664, B1 => n10084, B2 => 
                           n9808, ZN => n9418);
   U8866 : OAI221_X1 port map( B1 => n8640, B2 => n10123, C1 => n8384, C2 => 
                           n10110, A => n9422, ZN => n9421);
   U8867 : AOI22_X1 port map( A1 => n10097, A2 => n9918, B1 => n10084, B2 => 
                           n9919, ZN => n9422);
   U8868 : OAI221_X1 port map( B1 => n8671, B2 => n10123, C1 => n8415, C2 => 
                           n10110, A => n9398, ZN => n9397);
   U8869 : AOI22_X1 port map( A1 => n10097, A2 => n9665, B1 => n10084, B2 => 
                           n9809, ZN => n9398);
   U8870 : OAI221_X1 port map( B1 => n8639, B2 => n10123, C1 => n8383, C2 => 
                           n10110, A => n9402, ZN => n9401);
   U8871 : AOI22_X1 port map( A1 => n10097, A2 => n9922, B1 => n10084, B2 => 
                           n9923, ZN => n9402);
   U8872 : OAI221_X1 port map( B1 => n8670, B2 => n10124, C1 => n8414, C2 => 
                           n10111, A => n9378, ZN => n9377);
   U8873 : AOI22_X1 port map( A1 => n10098, A2 => n9666, B1 => n10085, B2 => 
                           n9810, ZN => n9378);
   U8874 : OAI221_X1 port map( B1 => n8638, B2 => n10124, C1 => n8382, C2 => 
                           n10111, A => n9382, ZN => n9381);
   U8875 : AOI22_X1 port map( A1 => n10098, A2 => n9926, B1 => n10085, B2 => 
                           n9927, ZN => n9382);
   U8876 : OAI221_X1 port map( B1 => n8669, B2 => n10124, C1 => n8413, C2 => 
                           n10111, A => n9358, ZN => n9357);
   U8877 : AOI22_X1 port map( A1 => n10098, A2 => n9667, B1 => n10085, B2 => 
                           n9811, ZN => n9358);
   U8878 : OAI221_X1 port map( B1 => n8637, B2 => n10124, C1 => n8381, C2 => 
                           n10111, A => n9362, ZN => n9361);
   U8879 : AOI22_X1 port map( A1 => n10098, A2 => n9930, B1 => n10085, B2 => 
                           n9931, ZN => n9362);
   U8880 : OAI221_X1 port map( B1 => n8668, B2 => n10124, C1 => n8412, C2 => 
                           n10111, A => n9338, ZN => n9337);
   U8881 : AOI22_X1 port map( A1 => n10098, A2 => n9668, B1 => n10085, B2 => 
                           n9812, ZN => n9338);
   U8882 : OAI221_X1 port map( B1 => n8636, B2 => n10124, C1 => n8380, C2 => 
                           n10111, A => n9342, ZN => n9341);
   U8883 : AOI22_X1 port map( A1 => n10098, A2 => n9934, B1 => n10085, B2 => 
                           n9935, ZN => n9342);
   U8884 : OAI221_X1 port map( B1 => n8667, B2 => n10125, C1 => n8411, C2 => 
                           n10112, A => n9318, ZN => n9317);
   U8885 : AOI22_X1 port map( A1 => n10099, A2 => n9669, B1 => n10086, B2 => 
                           n9813, ZN => n9318);
   U8886 : OAI221_X1 port map( B1 => n8635, B2 => n10125, C1 => n8379, C2 => 
                           n10112, A => n9322, ZN => n9321);
   U8887 : AOI22_X1 port map( A1 => n10099, A2 => n9938, B1 => n10086, B2 => 
                           n9939, ZN => n9322);
   U8888 : OAI221_X1 port map( B1 => n8666, B2 => n10125, C1 => n8410, C2 => 
                           n10112, A => n9298, ZN => n9297);
   U8889 : AOI22_X1 port map( A1 => n10099, A2 => n9670, B1 => n10086, B2 => 
                           n9814, ZN => n9298);
   U8890 : OAI221_X1 port map( B1 => n8634, B2 => n10125, C1 => n8378, C2 => 
                           n10112, A => n9302, ZN => n9301);
   U8891 : AOI22_X1 port map( A1 => n10099, A2 => n9942, B1 => n10086, B2 => 
                           n9943, ZN => n9302);
   U8892 : OAI221_X1 port map( B1 => n8665, B2 => n10125, C1 => n8409, C2 => 
                           n10112, A => n9278, ZN => n9277);
   U8893 : AOI22_X1 port map( A1 => n10099, A2 => n9671, B1 => n10086, B2 => 
                           n9815, ZN => n9278);
   U8894 : OAI221_X1 port map( B1 => n8633, B2 => n10125, C1 => n8377, C2 => 
                           n10112, A => n9282, ZN => n9281);
   U8895 : AOI22_X1 port map( A1 => n10099, A2 => n9946, B1 => n10086, B2 => 
                           n9947, ZN => n9282);
   U8896 : OAI221_X1 port map( B1 => n8664, B2 => n10126, C1 => n8408, C2 => 
                           n10113, A => n9258, ZN => n9257);
   U8897 : AOI22_X1 port map( A1 => n10100, A2 => n9672, B1 => n10087, B2 => 
                           n9816, ZN => n9258);
   U8898 : OAI221_X1 port map( B1 => n8632, B2 => n10126, C1 => n8376, C2 => 
                           n10113, A => n9262, ZN => n9261);
   U8899 : AOI22_X1 port map( A1 => n10100, A2 => n9950, B1 => n10087, B2 => 
                           n9951, ZN => n9262);
   U8900 : OAI221_X1 port map( B1 => n8663, B2 => n10126, C1 => n8407, C2 => 
                           n10113, A => n9238, ZN => n9237);
   U8901 : AOI22_X1 port map( A1 => n10100, A2 => n9673, B1 => n10087, B2 => 
                           n9817, ZN => n9238);
   U8902 : OAI221_X1 port map( B1 => n8631, B2 => n10126, C1 => n8375, C2 => 
                           n10113, A => n9242, ZN => n9241);
   U8903 : AOI22_X1 port map( A1 => n10100, A2 => n9954, B1 => n10087, B2 => 
                           n9955, ZN => n9242);
   U8904 : OAI221_X1 port map( B1 => n8662, B2 => n10126, C1 => n8406, C2 => 
                           n10113, A => n9218, ZN => n9217);
   U8905 : AOI22_X1 port map( A1 => n10100, A2 => n9674, B1 => n10087, B2 => 
                           n9818, ZN => n9218);
   U8906 : OAI221_X1 port map( B1 => n8630, B2 => n10126, C1 => n8374, C2 => 
                           n10113, A => n9222, ZN => n9221);
   U8907 : AOI22_X1 port map( A1 => n10100, A2 => n9958, B1 => n10087, B2 => 
                           n9959, ZN => n9222);
   U8908 : OAI221_X1 port map( B1 => n8661, B2 => n10127, C1 => n8405, C2 => 
                           n10114, A => n9198, ZN => n9197);
   U8909 : AOI22_X1 port map( A1 => n10101, A2 => n9675, B1 => n10088, B2 => 
                           n9819, ZN => n9198);
   U8910 : OAI221_X1 port map( B1 => n8629, B2 => n10127, C1 => n8373, C2 => 
                           n10114, A => n9202, ZN => n9201);
   U8911 : AOI22_X1 port map( A1 => n10101, A2 => n9962, B1 => n10088, B2 => 
                           n9963, ZN => n9202);
   U8912 : OAI221_X1 port map( B1 => n8660, B2 => n10127, C1 => n8404, C2 => 
                           n10114, A => n9178, ZN => n9177);
   U8913 : AOI22_X1 port map( A1 => n10101, A2 => n9676, B1 => n10088, B2 => 
                           n9820, ZN => n9178);
   U8914 : OAI221_X1 port map( B1 => n8628, B2 => n10127, C1 => n8372, C2 => 
                           n10114, A => n9182, ZN => n9181);
   U8915 : AOI22_X1 port map( A1 => n10101, A2 => n9966, B1 => n10088, B2 => 
                           n9967, ZN => n9182);
   U8916 : OAI221_X1 port map( B1 => n8659, B2 => n10127, C1 => n8403, C2 => 
                           n10114, A => n9158, ZN => n9157);
   U8917 : AOI22_X1 port map( A1 => n10101, A2 => n9677, B1 => n10088, B2 => 
                           n9821, ZN => n9158);
   U8918 : OAI221_X1 port map( B1 => n8627, B2 => n10127, C1 => n8371, C2 => 
                           n10114, A => n9162, ZN => n9161);
   U8919 : AOI22_X1 port map( A1 => n10101, A2 => n9970, B1 => n10088, B2 => 
                           n9971, ZN => n9162);
   U8920 : OAI221_X1 port map( B1 => n8658, B2 => n10128, C1 => n8402, C2 => 
                           n10115, A => n9138, ZN => n9137);
   U8921 : AOI22_X1 port map( A1 => n10102, A2 => n9678, B1 => n10089, B2 => 
                           n9822, ZN => n9138);
   U8922 : OAI221_X1 port map( B1 => n8626, B2 => n10128, C1 => n8370, C2 => 
                           n10115, A => n9142, ZN => n9141);
   U8923 : AOI22_X1 port map( A1 => n10102, A2 => n9974, B1 => n10089, B2 => 
                           n9975, ZN => n9142);
   U8924 : OAI221_X1 port map( B1 => n8657, B2 => n10128, C1 => n8401, C2 => 
                           n10115, A => n9118, ZN => n9117);
   U8925 : AOI22_X1 port map( A1 => n10102, A2 => n9679, B1 => n10089, B2 => 
                           n9823, ZN => n9118);
   U8926 : OAI221_X1 port map( B1 => n8625, B2 => n10128, C1 => n8369, C2 => 
                           n10115, A => n9122, ZN => n9121);
   U8927 : AOI22_X1 port map( A1 => n10102, A2 => n9978, B1 => n10089, B2 => 
                           n9979, ZN => n9122);
   U8928 : OAI221_X1 port map( B1 => n8656, B2 => n10128, C1 => n8400, C2 => 
                           n10115, A => n9098, ZN => n9097);
   U8929 : AOI22_X1 port map( A1 => n10102, A2 => n9680, B1 => n10089, B2 => 
                           n9824, ZN => n9098);
   U8930 : OAI221_X1 port map( B1 => n8624, B2 => n10128, C1 => n8368, C2 => 
                           n10115, A => n9102, ZN => n9101);
   U8931 : AOI22_X1 port map( A1 => n10102, A2 => n9982, B1 => n10089, B2 => 
                           n9983, ZN => n9102);
   U8932 : OAI221_X1 port map( B1 => n8655, B2 => n10129, C1 => n8399, C2 => 
                           n10116, A => n9078, ZN => n9077);
   U8933 : AOI22_X1 port map( A1 => n10103, A2 => n9681, B1 => n10090, B2 => 
                           n9825, ZN => n9078);
   U8934 : OAI221_X1 port map( B1 => n8623, B2 => n10129, C1 => n8367, C2 => 
                           n10116, A => n9082, ZN => n9081);
   U8935 : AOI22_X1 port map( A1 => n10103, A2 => n9986, B1 => n10090, B2 => 
                           n9987, ZN => n9082);
   U8936 : OAI221_X1 port map( B1 => n8654, B2 => n10129, C1 => n8398, C2 => 
                           n10116, A => n9058, ZN => n9057);
   U8937 : AOI22_X1 port map( A1 => n10103, A2 => n9682, B1 => n10090, B2 => 
                           n9826, ZN => n9058);
   U8938 : OAI221_X1 port map( B1 => n8622, B2 => n10129, C1 => n8366, C2 => 
                           n10116, A => n9062, ZN => n9061);
   U8939 : AOI22_X1 port map( A1 => n10103, A2 => n9990, B1 => n10090, B2 => 
                           n9991, ZN => n9062);
   U8940 : OAI221_X1 port map( B1 => n8653, B2 => n10129, C1 => n8397, C2 => 
                           n10116, A => n9038, ZN => n9037);
   U8941 : AOI22_X1 port map( A1 => n10103, A2 => n9683, B1 => n10090, B2 => 
                           n9827, ZN => n9038);
   U8942 : OAI221_X1 port map( B1 => n8621, B2 => n10129, C1 => n8365, C2 => 
                           n10116, A => n9042, ZN => n9041);
   U8943 : AOI22_X1 port map( A1 => n10103, A2 => n9994, B1 => n10090, B2 => 
                           n9995, ZN => n9042);
   U8944 : OAI221_X1 port map( B1 => n8652, B2 => n10130, C1 => n8396, C2 => 
                           n10117, A => n9018, ZN => n9017);
   U8945 : AOI22_X1 port map( A1 => n10104, A2 => n9524, B1 => n10091, B2 => 
                           n9576, ZN => n9018);
   U8946 : OAI221_X1 port map( B1 => n8620, B2 => n10130, C1 => n8364, C2 => 
                           n10117, A => n9022, ZN => n9021);
   U8947 : AOI22_X1 port map( A1 => n10104, A2 => n9998, B1 => n10091, B2 => 
                           n9999, ZN => n9022);
   U8948 : OAI221_X1 port map( B1 => n8651, B2 => n10130, C1 => n8395, C2 => 
                           n10117, A => n8998, ZN => n8997);
   U8949 : AOI22_X1 port map( A1 => n10104, A2 => n9525, B1 => n10091, B2 => 
                           n9577, ZN => n8998);
   U8950 : OAI221_X1 port map( B1 => n8619, B2 => n10130, C1 => n8363, C2 => 
                           n10117, A => n9002, ZN => n9001);
   U8951 : AOI22_X1 port map( A1 => n10104, A2 => n10002, B1 => n10091, B2 => 
                           n10003, ZN => n9002);
   U8952 : OAI221_X1 port map( B1 => n8650, B2 => n10130, C1 => n8394, C2 => 
                           n10117, A => n8978, ZN => n8977);
   U8953 : AOI22_X1 port map( A1 => n10104, A2 => n9526, B1 => n10091, B2 => 
                           n9578, ZN => n8978);
   U8954 : OAI221_X1 port map( B1 => n8618, B2 => n10130, C1 => n8362, C2 => 
                           n10117, A => n8982, ZN => n8981);
   U8955 : AOI22_X1 port map( A1 => n10104, A2 => n10006, B1 => n10091, B2 => 
                           n10007, ZN => n8982);
   U8956 : OAI221_X1 port map( B1 => n8649, B2 => n10131, C1 => n8393, C2 => 
                           n10118, A => n8958, ZN => n8957);
   U8957 : AOI22_X1 port map( A1 => n10105, A2 => n9527, B1 => n10092, B2 => 
                           n9579, ZN => n8958);
   U8958 : OAI221_X1 port map( B1 => n8617, B2 => n10131, C1 => n8361, C2 => 
                           n10118, A => n8962, ZN => n8961);
   U8959 : AOI22_X1 port map( A1 => n10105, A2 => n10010, B1 => n10092, B2 => 
                           n10011, ZN => n8962);
   U8960 : OAI221_X1 port map( B1 => n8648, B2 => n10131, C1 => n8392, C2 => 
                           n10118, A => n8938, ZN => n8937);
   U8961 : AOI22_X1 port map( A1 => n10105, A2 => n9528, B1 => n10092, B2 => 
                           n9580, ZN => n8938);
   U8962 : OAI221_X1 port map( B1 => n8616, B2 => n10131, C1 => n8360, C2 => 
                           n10118, A => n8942, ZN => n8941);
   U8963 : AOI22_X1 port map( A1 => n10105, A2 => n10014, B1 => n10092, B2 => 
                           n10015, ZN => n8942);
   U8964 : OAI221_X1 port map( B1 => n8647, B2 => n10131, C1 => n8391, C2 => 
                           n10118, A => n8918, ZN => n8917);
   U8965 : AOI22_X1 port map( A1 => n10105, A2 => n9529, B1 => n10092, B2 => 
                           n9581, ZN => n8918);
   U8966 : OAI221_X1 port map( B1 => n8615, B2 => n10131, C1 => n8359, C2 => 
                           n10118, A => n8922, ZN => n8921);
   U8967 : AOI22_X1 port map( A1 => n10105, A2 => n10018, B1 => n10092, B2 => 
                           n10019, ZN => n8922);
   U8968 : OAI21_X1 port map( B1 => n9492, B2 => n9493, A => n10133, ZN => 
                           n9491);
   U8969 : OAI221_X1 port map( B1 => n8580, B2 => n10070, C1 => n8324, C2 => 
                           n10057, A => n9495, ZN => n9492);
   U8970 : OAI221_X1 port map( B1 => n8708, B2 => n10122, C1 => n8452, C2 => 
                           n10109, A => n9494, ZN => n9493);
   U8971 : AOI22_X1 port map( A1 => n10044, A2 => n9708, B1 => n10031, B2 => 
                           n9852, ZN => n9495);
   U8972 : OAI21_X1 port map( B1 => n9472, B2 => n9473, A => n10133, ZN => 
                           n9471);
   U8973 : OAI221_X1 port map( B1 => n8579, B2 => n10070, C1 => n8323, C2 => 
                           n10057, A => n9475, ZN => n9472);
   U8974 : OAI221_X1 port map( B1 => n8707, B2 => n10122, C1 => n8451, C2 => 
                           n10109, A => n9474, ZN => n9473);
   U8975 : AOI22_X1 port map( A1 => n10044, A2 => n9709, B1 => n10031, B2 => 
                           n9853, ZN => n9475);
   U8976 : OAI21_X1 port map( B1 => n9452, B2 => n9453, A => n10133, ZN => 
                           n9451);
   U8977 : OAI221_X1 port map( B1 => n8578, B2 => n10070, C1 => n8322, C2 => 
                           n10057, A => n9455, ZN => n9452);
   U8978 : OAI221_X1 port map( B1 => n8706, B2 => n10122, C1 => n8450, C2 => 
                           n10109, A => n9454, ZN => n9453);
   U8979 : AOI22_X1 port map( A1 => n10044, A2 => n9710, B1 => n10031, B2 => 
                           n9854, ZN => n9455);
   U8980 : OAI21_X1 port map( B1 => n9432, B2 => n9433, A => n10133, ZN => 
                           n9431);
   U8981 : OAI221_X1 port map( B1 => n8577, B2 => n10071, C1 => n8321, C2 => 
                           n10058, A => n9435, ZN => n9432);
   U8982 : OAI221_X1 port map( B1 => n8705, B2 => n10123, C1 => n8449, C2 => 
                           n10110, A => n9434, ZN => n9433);
   U8983 : AOI22_X1 port map( A1 => n10045, A2 => n9711, B1 => n10032, B2 => 
                           n9855, ZN => n9435);
   U8984 : OAI21_X1 port map( B1 => n9412, B2 => n9413, A => n10133, ZN => 
                           n9411);
   U8985 : OAI221_X1 port map( B1 => n8576, B2 => n10071, C1 => n8320, C2 => 
                           n10058, A => n9415, ZN => n9412);
   U8986 : OAI221_X1 port map( B1 => n8704, B2 => n10123, C1 => n8448, C2 => 
                           n10110, A => n9414, ZN => n9413);
   U8987 : AOI22_X1 port map( A1 => n10045, A2 => n9712, B1 => n10032, B2 => 
                           n9856, ZN => n9415);
   U8988 : OAI21_X1 port map( B1 => n9392, B2 => n9393, A => n10133, ZN => 
                           n9391);
   U8989 : OAI221_X1 port map( B1 => n8575, B2 => n10071, C1 => n8319, C2 => 
                           n10058, A => n9395, ZN => n9392);
   U8990 : OAI221_X1 port map( B1 => n8703, B2 => n10123, C1 => n8447, C2 => 
                           n10110, A => n9394, ZN => n9393);
   U8991 : AOI22_X1 port map( A1 => n10045, A2 => n9713, B1 => n10032, B2 => 
                           n9857, ZN => n9395);
   U8992 : OAI21_X1 port map( B1 => n9372, B2 => n9373, A => n10133, ZN => 
                           n9371);
   U8993 : OAI221_X1 port map( B1 => n8574, B2 => n10072, C1 => n8318, C2 => 
                           n10059, A => n9375, ZN => n9372);
   U8994 : OAI221_X1 port map( B1 => n8702, B2 => n10124, C1 => n8446, C2 => 
                           n10111, A => n9374, ZN => n9373);
   U8995 : AOI22_X1 port map( A1 => n10046, A2 => n9714, B1 => n10033, B2 => 
                           n9858, ZN => n9375);
   U8996 : OAI21_X1 port map( B1 => n9352, B2 => n9353, A => n10133, ZN => 
                           n9351);
   U8997 : OAI221_X1 port map( B1 => n8573, B2 => n10072, C1 => n8317, C2 => 
                           n10059, A => n9355, ZN => n9352);
   U8998 : OAI221_X1 port map( B1 => n8701, B2 => n10124, C1 => n8445, C2 => 
                           n10111, A => n9354, ZN => n9353);
   U8999 : AOI22_X1 port map( A1 => n10046, A2 => n9715, B1 => n10033, B2 => 
                           n9859, ZN => n9355);
   U9000 : OAI21_X1 port map( B1 => n9332, B2 => n9333, A => n10133, ZN => 
                           n9331);
   U9001 : OAI221_X1 port map( B1 => n8572, B2 => n10072, C1 => n8316, C2 => 
                           n10059, A => n9335, ZN => n9332);
   U9002 : OAI221_X1 port map( B1 => n8700, B2 => n10124, C1 => n8444, C2 => 
                           n10111, A => n9334, ZN => n9333);
   U9003 : AOI22_X1 port map( A1 => n10046, A2 => n9716, B1 => n10033, B2 => 
                           n9860, ZN => n9335);
   U9004 : OAI21_X1 port map( B1 => n9312, B2 => n9313, A => n10133, ZN => 
                           n9311);
   U9005 : OAI221_X1 port map( B1 => n8571, B2 => n10073, C1 => n8315, C2 => 
                           n10060, A => n9315, ZN => n9312);
   U9006 : OAI221_X1 port map( B1 => n8699, B2 => n10125, C1 => n8443, C2 => 
                           n10112, A => n9314, ZN => n9313);
   U9007 : AOI22_X1 port map( A1 => n10047, A2 => n9717, B1 => n10034, B2 => 
                           n9861, ZN => n9315);
   U9008 : OAI21_X1 port map( B1 => n9292, B2 => n9293, A => n10133, ZN => 
                           n9291);
   U9009 : OAI221_X1 port map( B1 => n8570, B2 => n10073, C1 => n8314, C2 => 
                           n10060, A => n9295, ZN => n9292);
   U9010 : OAI221_X1 port map( B1 => n8698, B2 => n10125, C1 => n8442, C2 => 
                           n10112, A => n9294, ZN => n9293);
   U9011 : AOI22_X1 port map( A1 => n10047, A2 => n9718, B1 => n10034, B2 => 
                           n9862, ZN => n9295);
   U9012 : OAI21_X1 port map( B1 => n9272, B2 => n9273, A => n10133, ZN => 
                           n9271);
   U9013 : OAI221_X1 port map( B1 => n8569, B2 => n10073, C1 => n8313, C2 => 
                           n10060, A => n9275, ZN => n9272);
   U9014 : OAI221_X1 port map( B1 => n8697, B2 => n10125, C1 => n8441, C2 => 
                           n10112, A => n9274, ZN => n9273);
   U9015 : AOI22_X1 port map( A1 => n10047, A2 => n9719, B1 => n10034, B2 => 
                           n9863, ZN => n9275);
   U9016 : OAI21_X1 port map( B1 => n9252, B2 => n9253, A => n10134, ZN => 
                           n9251);
   U9017 : OAI221_X1 port map( B1 => n8568, B2 => n10074, C1 => n8312, C2 => 
                           n10061, A => n9255, ZN => n9252);
   U9018 : OAI221_X1 port map( B1 => n8696, B2 => n10126, C1 => n8440, C2 => 
                           n10113, A => n9254, ZN => n9253);
   U9019 : AOI22_X1 port map( A1 => n10048, A2 => n9720, B1 => n10035, B2 => 
                           n9864, ZN => n9255);
   U9020 : OAI21_X1 port map( B1 => n9232, B2 => n9233, A => n10134, ZN => 
                           n9231);
   U9021 : OAI221_X1 port map( B1 => n8567, B2 => n10074, C1 => n8311, C2 => 
                           n10061, A => n9235, ZN => n9232);
   U9022 : OAI221_X1 port map( B1 => n8695, B2 => n10126, C1 => n8439, C2 => 
                           n10113, A => n9234, ZN => n9233);
   U9023 : AOI22_X1 port map( A1 => n10048, A2 => n9721, B1 => n10035, B2 => 
                           n9865, ZN => n9235);
   U9024 : OAI21_X1 port map( B1 => n9212, B2 => n9213, A => n10134, ZN => 
                           n9211);
   U9025 : OAI221_X1 port map( B1 => n8566, B2 => n10074, C1 => n8310, C2 => 
                           n10061, A => n9215, ZN => n9212);
   U9026 : OAI221_X1 port map( B1 => n8694, B2 => n10126, C1 => n8438, C2 => 
                           n10113, A => n9214, ZN => n9213);
   U9027 : AOI22_X1 port map( A1 => n10048, A2 => n9722, B1 => n10035, B2 => 
                           n9866, ZN => n9215);
   U9028 : OAI21_X1 port map( B1 => n9192, B2 => n9193, A => n10134, ZN => 
                           n9191);
   U9029 : OAI221_X1 port map( B1 => n8565, B2 => n10075, C1 => n8309, C2 => 
                           n10062, A => n9195, ZN => n9192);
   U9030 : OAI221_X1 port map( B1 => n8693, B2 => n10127, C1 => n8437, C2 => 
                           n10114, A => n9194, ZN => n9193);
   U9031 : AOI22_X1 port map( A1 => n10049, A2 => n9723, B1 => n10036, B2 => 
                           n9867, ZN => n9195);
   U9032 : OAI21_X1 port map( B1 => n9172, B2 => n9173, A => n10134, ZN => 
                           n9171);
   U9033 : OAI221_X1 port map( B1 => n8564, B2 => n10075, C1 => n8308, C2 => 
                           n10062, A => n9175, ZN => n9172);
   U9034 : OAI221_X1 port map( B1 => n8692, B2 => n10127, C1 => n8436, C2 => 
                           n10114, A => n9174, ZN => n9173);
   U9035 : AOI22_X1 port map( A1 => n10049, A2 => n9724, B1 => n10036, B2 => 
                           n9868, ZN => n9175);
   U9036 : OAI21_X1 port map( B1 => n9152, B2 => n9153, A => n10134, ZN => 
                           n9151);
   U9037 : OAI221_X1 port map( B1 => n8563, B2 => n10075, C1 => n8307, C2 => 
                           n10062, A => n9155, ZN => n9152);
   U9038 : OAI221_X1 port map( B1 => n8691, B2 => n10127, C1 => n8435, C2 => 
                           n10114, A => n9154, ZN => n9153);
   U9039 : AOI22_X1 port map( A1 => n10049, A2 => n9725, B1 => n10036, B2 => 
                           n9869, ZN => n9155);
   U9040 : OAI21_X1 port map( B1 => n9012, B2 => n9013, A => n10135, ZN => 
                           n9011);
   U9041 : OAI221_X1 port map( B1 => n8556, B2 => n10078, C1 => n8300, C2 => 
                           n10065, A => n9015, ZN => n9012);
   U9042 : OAI221_X1 port map( B1 => n8684, B2 => n10130, C1 => n8428, C2 => 
                           n10117, A => n9014, ZN => n9013);
   U9043 : AOI22_X1 port map( A1 => n10052, A2 => n9542, B1 => n10039, B2 => 
                           n9594, ZN => n9015);
   U9044 : OAI21_X1 port map( B1 => n8992, B2 => n8993, A => n10135, ZN => 
                           n8991);
   U9045 : OAI221_X1 port map( B1 => n8555, B2 => n10078, C1 => n8299, C2 => 
                           n10065, A => n8995, ZN => n8992);
   U9046 : OAI221_X1 port map( B1 => n8683, B2 => n10130, C1 => n8427, C2 => 
                           n10117, A => n8994, ZN => n8993);
   U9047 : AOI22_X1 port map( A1 => n10052, A2 => n9543, B1 => n10039, B2 => 
                           n9595, ZN => n8995);
   U9048 : OAI21_X1 port map( B1 => n8972, B2 => n8973, A => n10135, ZN => 
                           n8971);
   U9049 : OAI221_X1 port map( B1 => n8554, B2 => n10078, C1 => n8298, C2 => 
                           n10065, A => n8975, ZN => n8972);
   U9050 : OAI221_X1 port map( B1 => n8682, B2 => n10130, C1 => n8426, C2 => 
                           n10117, A => n8974, ZN => n8973);
   U9051 : AOI22_X1 port map( A1 => n10052, A2 => n9544, B1 => n10039, B2 => 
                           n9596, ZN => n8975);
   U9052 : OAI21_X1 port map( B1 => n8952, B2 => n8953, A => n10135, ZN => 
                           n8951);
   U9053 : OAI221_X1 port map( B1 => n8553, B2 => n10079, C1 => n8297, C2 => 
                           n10066, A => n8955, ZN => n8952);
   U9054 : OAI221_X1 port map( B1 => n8681, B2 => n10131, C1 => n8425, C2 => 
                           n10118, A => n8954, ZN => n8953);
   U9055 : AOI22_X1 port map( A1 => n10053, A2 => n9545, B1 => n10040, B2 => 
                           n9597, ZN => n8955);
   U9056 : OAI21_X1 port map( B1 => n8932, B2 => n8933, A => n10135, ZN => 
                           n8931);
   U9057 : OAI221_X1 port map( B1 => n8552, B2 => n10079, C1 => n8296, C2 => 
                           n10066, A => n8935, ZN => n8932);
   U9058 : OAI221_X1 port map( B1 => n8680, B2 => n10131, C1 => n8424, C2 => 
                           n10118, A => n8934, ZN => n8933);
   U9059 : AOI22_X1 port map( A1 => n10053, A2 => n9546, B1 => n10040, B2 => 
                           n9598, ZN => n8935);
   U9060 : OAI21_X1 port map( B1 => n8912, B2 => n8913, A => n10135, ZN => 
                           n8911);
   U9061 : OAI221_X1 port map( B1 => n8551, B2 => n10079, C1 => n8295, C2 => 
                           n10066, A => n8915, ZN => n8912);
   U9062 : OAI221_X1 port map( B1 => n8679, B2 => n10131, C1 => n8423, C2 => 
                           n10118, A => n8914, ZN => n8913);
   U9063 : AOI22_X1 port map( A1 => n10053, A2 => n9547, B1 => n10040, B2 => 
                           n9599, ZN => n8915);
   U9064 : AOI22_X1 port map( A1 => n10106, A2 => n9522, B1 => n10093, B2 => 
                           n9574, ZN => n8894);
   U9065 : AOI22_X1 port map( A1 => n10106, A2 => n9523, B1 => n10093, B2 => 
                           n9575, ZN => n8865);
   U9066 : OAI221_X1 port map( B1 => n8646, B2 => n10132, C1 => n8390, C2 => 
                           n10119, A => n8898, ZN => n8897);
   U9067 : AOI22_X1 port map( A1 => n10106, A2 => n9530, B1 => n10093, B2 => 
                           n9582, ZN => n8898);
   U9068 : OAI221_X1 port map( B1 => n8518, B2 => n10080, C1 => n8262, C2 => 
                           n10067, A => n8899, ZN => n8896);
   U9069 : AOI22_X1 port map( A1 => n10054, A2 => n9556, B1 => n10041, B2 => 
                           n9608, ZN => n8899);
   U9070 : OAI221_X1 port map( B1 => n8614, B2 => n10132, C1 => n8358, C2 => 
                           n10119, A => n8902, ZN => n8901);
   U9071 : AOI22_X1 port map( A1 => n10106, A2 => n9532, B1 => n10093, B2 => 
                           n9584, ZN => n8902);
   U9072 : OAI221_X1 port map( B1 => n8486, B2 => n10080, C1 => n8230, C2 => 
                           n10067, A => n8903, ZN => n8900);
   U9073 : AOI22_X1 port map( A1 => n10054, A2 => n9558, B1 => n10041, B2 => 
                           n9610, ZN => n8903);
   U9074 : OAI221_X1 port map( B1 => n6683, B2 => n10132, C1 => n8454, C2 => 
                           n10119, A => n8906, ZN => n8905);
   U9075 : AOI22_X1 port map( A1 => n10106, A2 => n9514, B1 => n10093, B2 => 
                           n9566, ZN => n8906);
   U9076 : OAI221_X1 port map( B1 => n8582, B2 => n10080, C1 => n8326, C2 => 
                           n10067, A => n8907, ZN => n8904);
   U9077 : AOI22_X1 port map( A1 => n10054, A2 => n9540, B1 => n10041, B2 => 
                           n9592, ZN => n8907);
   U9078 : OAI221_X1 port map( B1 => n8645, B2 => n10132, C1 => n8389, C2 => 
                           n10119, A => n8876, ZN => n8874);
   U9079 : AOI22_X1 port map( A1 => n10106, A2 => n9531, B1 => n10093, B2 => 
                           n9583, ZN => n8876);
   U9080 : OAI221_X1 port map( B1 => n8517, B2 => n10080, C1 => n8261, C2 => 
                           n10067, A => n8877, ZN => n8873);
   U9081 : AOI22_X1 port map( A1 => n10054, A2 => n9557, B1 => n10041, B2 => 
                           n9609, ZN => n8877);
   U9082 : OAI221_X1 port map( B1 => n8613, B2 => n10132, C1 => n8357, C2 => 
                           n10119, A => n8881, ZN => n8879);
   U9083 : AOI22_X1 port map( A1 => n10106, A2 => n9533, B1 => n10093, B2 => 
                           n9585, ZN => n8881);
   U9084 : OAI221_X1 port map( B1 => n8485, B2 => n10080, C1 => n8229, C2 => 
                           n10067, A => n8882, ZN => n8878);
   U9085 : AOI22_X1 port map( A1 => n10054, A2 => n9559, B1 => n10041, B2 => 
                           n9611, ZN => n8882);
   U9086 : OAI221_X1 port map( B1 => n6682, B2 => n10132, C1 => n8453, C2 => 
                           n10119, A => n8886, ZN => n8884);
   U9087 : AOI22_X1 port map( A1 => n10106, A2 => n9515, B1 => n10093, B2 => 
                           n9567, ZN => n8886);
   U9088 : OAI221_X1 port map( B1 => n8581, B2 => n10080, C1 => n8325, C2 => 
                           n10067, A => n8887, ZN => n8883);
   U9089 : AOI22_X1 port map( A1 => n10054, A2 => n9541, B1 => n10041, B2 => 
                           n9593, ZN => n8887);
   U9090 : OAI22_X1 port map( A1 => n10331, A2 => n10513, B1 => n8795, B2 => 
                           n8743, ZN => n1850);
   U9091 : OAI22_X1 port map( A1 => n10331, A2 => n10525, B1 => n8795, B2 => 
                           n8742, ZN => n1851);
   U9092 : OAI22_X1 port map( A1 => n10320, A2 => n10496, B1 => n8796, B2 => 
                           n8741, ZN => n1812);
   U9093 : OAI22_X1 port map( A1 => n10321, A2 => n10499, B1 => n8796, B2 => 
                           n8740, ZN => n1813);
   U9094 : OAI22_X1 port map( A1 => n10321, A2 => n10502, B1 => n8796, B2 => 
                           n8739, ZN => n1814);
   U9095 : OAI22_X1 port map( A1 => n10321, A2 => n10505, B1 => n8796, B2 => 
                           n8738, ZN => n1815);
   U9096 : OAI22_X1 port map( A1 => n10321, A2 => n10508, B1 => n8796, B2 => 
                           n8737, ZN => n1816);
   U9097 : OAI22_X1 port map( A1 => n10321, A2 => n10511, B1 => n8796, B2 => 
                           n8736, ZN => n1817);
   U9098 : OAI22_X1 port map( A1 => n10322, A2 => n10514, B1 => n8796, B2 => 
                           n8735, ZN => n1818);
   U9099 : OAI22_X1 port map( A1 => n10322, A2 => n10526, B1 => n8796, B2 => 
                           n8734, ZN => n1819);
   U9100 : OAI22_X1 port map( A1 => n10311, A2 => n10496, B1 => n8798, B2 => 
                           n8733, ZN => n1780);
   U9101 : OAI22_X1 port map( A1 => n10312, A2 => n10499, B1 => n8798, B2 => 
                           n8732, ZN => n1781);
   U9102 : OAI22_X1 port map( A1 => n10312, A2 => n10502, B1 => n8798, B2 => 
                           n8731, ZN => n1782);
   U9103 : OAI22_X1 port map( A1 => n10312, A2 => n10505, B1 => n8798, B2 => 
                           n8730, ZN => n1783);
   U9104 : OAI22_X1 port map( A1 => n10312, A2 => n10508, B1 => n8798, B2 => 
                           n8729, ZN => n1784);
   U9105 : OAI22_X1 port map( A1 => n10312, A2 => n10511, B1 => n8798, B2 => 
                           n8728, ZN => n1785);
   U9106 : OAI22_X1 port map( A1 => n10313, A2 => n10514, B1 => n8798, B2 => 
                           n8727, ZN => n1786);
   U9107 : OAI22_X1 port map( A1 => n10313, A2 => n10526, B1 => n8798, B2 => 
                           n8726, ZN => n1787);
   U9108 : OAI22_X1 port map( A1 => n10302, A2 => n10496, B1 => n8799, B2 => 
                           n8725, ZN => n1748);
   U9109 : OAI22_X1 port map( A1 => n10303, A2 => n10499, B1 => n8799, B2 => 
                           n8724, ZN => n1749);
   U9110 : OAI22_X1 port map( A1 => n10303, A2 => n10502, B1 => n8799, B2 => 
                           n8723, ZN => n1750);
   U9111 : OAI22_X1 port map( A1 => n10303, A2 => n10505, B1 => n8799, B2 => 
                           n8722, ZN => n1751);
   U9112 : OAI22_X1 port map( A1 => n10303, A2 => n10508, B1 => n8799, B2 => 
                           n8721, ZN => n1752);
   U9113 : OAI22_X1 port map( A1 => n10303, A2 => n10511, B1 => n8799, B2 => 
                           n8720, ZN => n1753);
   U9114 : OAI22_X1 port map( A1 => n10304, A2 => n10514, B1 => n8799, B2 => 
                           n8719, ZN => n1754);
   U9115 : OAI22_X1 port map( A1 => n10304, A2 => n10526, B1 => n8799, B2 => 
                           n8718, ZN => n1755);
   U9116 : OAI22_X1 port map( A1 => n10293, A2 => n10496, B1 => n8800, B2 => 
                           n8717, ZN => n1716);
   U9117 : OAI22_X1 port map( A1 => n10294, A2 => n10499, B1 => n8800, B2 => 
                           n8716, ZN => n1717);
   U9118 : OAI22_X1 port map( A1 => n10294, A2 => n10502, B1 => n8800, B2 => 
                           n8715, ZN => n1718);
   U9119 : OAI22_X1 port map( A1 => n10294, A2 => n10505, B1 => n8800, B2 => 
                           n8714, ZN => n1719);
   U9120 : OAI22_X1 port map( A1 => n10294, A2 => n10508, B1 => n8800, B2 => 
                           n8713, ZN => n1720);
   U9121 : OAI22_X1 port map( A1 => n10294, A2 => n10511, B1 => n8800, B2 => 
                           n8712, ZN => n1721);
   U9122 : OAI22_X1 port map( A1 => n10295, A2 => n10514, B1 => n8800, B2 => 
                           n8711, ZN => n1722);
   U9123 : OAI22_X1 port map( A1 => n10295, A2 => n10526, B1 => n8800, B2 => 
                           n8710, ZN => n1723);
   U9124 : OAI22_X1 port map( A1 => n10329, A2 => n10495, B1 => n8795, B2 => 
                           n8108, ZN => n1844);
   U9125 : OAI22_X1 port map( A1 => n10330, A2 => n10498, B1 => n8795, B2 => 
                           n8107, ZN => n1845);
   U9126 : OAI22_X1 port map( A1 => n10330, A2 => n10501, B1 => n8795, B2 => 
                           n8106, ZN => n1846);
   U9127 : OAI22_X1 port map( A1 => n10330, A2 => n10504, B1 => n8795, B2 => 
                           n8105, ZN => n1847);
   U9128 : OAI22_X1 port map( A1 => n10330, A2 => n10507, B1 => n8795, B2 => 
                           n8104, ZN => n1848);
   U9129 : OAI22_X1 port map( A1 => n10330, A2 => n10510, B1 => n8795, B2 => 
                           n8103, ZN => n1849);
   U9130 : OAI22_X1 port map( A1 => n10338, A2 => n10495, B1 => n8794, B2 => 
                           n8078, ZN => n1876);
   U9131 : OAI22_X1 port map( A1 => n10339, A2 => n10498, B1 => n8794, B2 => 
                           n8077, ZN => n1877);
   U9132 : OAI22_X1 port map( A1 => n10339, A2 => n10501, B1 => n8794, B2 => 
                           n8076, ZN => n1878);
   U9133 : OAI22_X1 port map( A1 => n10339, A2 => n10504, B1 => n8794, B2 => 
                           n8075, ZN => n1879);
   U9134 : OAI22_X1 port map( A1 => n10339, A2 => n10507, B1 => n8794, B2 => 
                           n8074, ZN => n1880);
   U9135 : OAI22_X1 port map( A1 => n10339, A2 => n10510, B1 => n8794, B2 => 
                           n8073, ZN => n1881);
   U9136 : OAI22_X1 port map( A1 => n10340, A2 => n10513, B1 => n8794, B2 => 
                           n8072, ZN => n1882);
   U9137 : OAI22_X1 port map( A1 => n10340, A2 => n10525, B1 => n8794, B2 => 
                           n8071, ZN => n1883);
   U9138 : OAI22_X1 port map( A1 => n10347, A2 => n10495, B1 => n8793, B2 => 
                           n8046, ZN => n1908);
   U9139 : OAI22_X1 port map( A1 => n10348, A2 => n10498, B1 => n8793, B2 => 
                           n8045, ZN => n1909);
   U9140 : OAI22_X1 port map( A1 => n10348, A2 => n10501, B1 => n8793, B2 => 
                           n8044, ZN => n1910);
   U9141 : OAI22_X1 port map( A1 => n10348, A2 => n10504, B1 => n8793, B2 => 
                           n8043, ZN => n1911);
   U9142 : OAI22_X1 port map( A1 => n10348, A2 => n10507, B1 => n8793, B2 => 
                           n8042, ZN => n1912);
   U9143 : OAI22_X1 port map( A1 => n10348, A2 => n10510, B1 => n8793, B2 => 
                           n8041, ZN => n1913);
   U9144 : OAI22_X1 port map( A1 => n10349, A2 => n10513, B1 => n8793, B2 => 
                           n8040, ZN => n1914);
   U9145 : OAI22_X1 port map( A1 => n10349, A2 => n10525, B1 => n8793, B2 => 
                           n8039, ZN => n1915);
   U9146 : OAI22_X1 port map( A1 => n10356, A2 => n10495, B1 => n8791, B2 => 
                           n8014, ZN => n1940);
   U9147 : OAI22_X1 port map( A1 => n10357, A2 => n10498, B1 => n8791, B2 => 
                           n8013, ZN => n1941);
   U9148 : OAI22_X1 port map( A1 => n10357, A2 => n10501, B1 => n8791, B2 => 
                           n8012, ZN => n1942);
   U9149 : OAI22_X1 port map( A1 => n10357, A2 => n10504, B1 => n8791, B2 => 
                           n8011, ZN => n1943);
   U9150 : OAI22_X1 port map( A1 => n10357, A2 => n10507, B1 => n8791, B2 => 
                           n8010, ZN => n1944);
   U9151 : OAI22_X1 port map( A1 => n10357, A2 => n10510, B1 => n8791, B2 => 
                           n8009, ZN => n1945);
   U9152 : OAI22_X1 port map( A1 => n10358, A2 => n10513, B1 => n8791, B2 => 
                           n8008, ZN => n1946);
   U9153 : OAI22_X1 port map( A1 => n10358, A2 => n10525, B1 => n8791, B2 => 
                           n8007, ZN => n1947);
   U9154 : OAI22_X1 port map( A1 => n10365, A2 => n10495, B1 => n8790, B2 => 
                           n7982, ZN => n1972);
   U9155 : OAI22_X1 port map( A1 => n10366, A2 => n10498, B1 => n8790, B2 => 
                           n7981, ZN => n1973);
   U9156 : OAI22_X1 port map( A1 => n10366, A2 => n10501, B1 => n8790, B2 => 
                           n7980, ZN => n1974);
   U9157 : OAI22_X1 port map( A1 => n10366, A2 => n10504, B1 => n8790, B2 => 
                           n7979, ZN => n1975);
   U9158 : OAI22_X1 port map( A1 => n10366, A2 => n10507, B1 => n8790, B2 => 
                           n7978, ZN => n1976);
   U9159 : OAI22_X1 port map( A1 => n10366, A2 => n10510, B1 => n8790, B2 => 
                           n7977, ZN => n1977);
   U9160 : OAI22_X1 port map( A1 => n10367, A2 => n10513, B1 => n8790, B2 => 
                           n7976, ZN => n1978);
   U9161 : OAI22_X1 port map( A1 => n10367, A2 => n10525, B1 => n8790, B2 => 
                           n7975, ZN => n1979);
   U9162 : OAI22_X1 port map( A1 => n10374, A2 => n10495, B1 => n8789, B2 => 
                           n7950, ZN => n2004);
   U9163 : OAI22_X1 port map( A1 => n10375, A2 => n10498, B1 => n8789, B2 => 
                           n7949, ZN => n2005);
   U9164 : OAI22_X1 port map( A1 => n10375, A2 => n10501, B1 => n8789, B2 => 
                           n7948, ZN => n2006);
   U9165 : OAI22_X1 port map( A1 => n10375, A2 => n10504, B1 => n8789, B2 => 
                           n7947, ZN => n2007);
   U9166 : OAI22_X1 port map( A1 => n10375, A2 => n10507, B1 => n8789, B2 => 
                           n7946, ZN => n2008);
   U9167 : OAI22_X1 port map( A1 => n10375, A2 => n10510, B1 => n8789, B2 => 
                           n7945, ZN => n2009);
   U9168 : OAI22_X1 port map( A1 => n10376, A2 => n10513, B1 => n8789, B2 => 
                           n7944, ZN => n2010);
   U9169 : OAI22_X1 port map( A1 => n10376, A2 => n10525, B1 => n8789, B2 => 
                           n7943, ZN => n2011);
   U9170 : OAI22_X1 port map( A1 => n10383, A2 => n10495, B1 => n8788, B2 => 
                           n7918, ZN => n2036);
   U9171 : OAI22_X1 port map( A1 => n10384, A2 => n10498, B1 => n8788, B2 => 
                           n7917, ZN => n2037);
   U9172 : OAI22_X1 port map( A1 => n10384, A2 => n10501, B1 => n8788, B2 => 
                           n7916, ZN => n2038);
   U9173 : OAI22_X1 port map( A1 => n10384, A2 => n10504, B1 => n8788, B2 => 
                           n7915, ZN => n2039);
   U9174 : OAI22_X1 port map( A1 => n10384, A2 => n10507, B1 => n8788, B2 => 
                           n7914, ZN => n2040);
   U9175 : OAI22_X1 port map( A1 => n10384, A2 => n10510, B1 => n8788, B2 => 
                           n7913, ZN => n2041);
   U9176 : OAI22_X1 port map( A1 => n10385, A2 => n10513, B1 => n8788, B2 => 
                           n7912, ZN => n2042);
   U9177 : OAI22_X1 port map( A1 => n10385, A2 => n10525, B1 => n8788, B2 => 
                           n7911, ZN => n2043);
   U9178 : OAI22_X1 port map( A1 => n10392, A2 => n10495, B1 => n8786, B2 => 
                           n7886, ZN => n2068);
   U9179 : OAI22_X1 port map( A1 => n10393, A2 => n10498, B1 => n8786, B2 => 
                           n7885, ZN => n2069);
   U9180 : OAI22_X1 port map( A1 => n10393, A2 => n10501, B1 => n8786, B2 => 
                           n7884, ZN => n2070);
   U9181 : OAI22_X1 port map( A1 => n10393, A2 => n10504, B1 => n8786, B2 => 
                           n7883, ZN => n2071);
   U9182 : OAI22_X1 port map( A1 => n10393, A2 => n10507, B1 => n8786, B2 => 
                           n7882, ZN => n2072);
   U9183 : OAI22_X1 port map( A1 => n10393, A2 => n10510, B1 => n8786, B2 => 
                           n7881, ZN => n2073);
   U9184 : OAI22_X1 port map( A1 => n10394, A2 => n10513, B1 => n8786, B2 => 
                           n7880, ZN => n2074);
   U9185 : OAI22_X1 port map( A1 => n10394, A2 => n10525, B1 => n8786, B2 => 
                           n7879, ZN => n2075);
   U9186 : OAI22_X1 port map( A1 => n10401, A2 => n10495, B1 => n8783, B2 => 
                           n7854, ZN => n2100);
   U9187 : OAI22_X1 port map( A1 => n10402, A2 => n10498, B1 => n8783, B2 => 
                           n7853, ZN => n2101);
   U9188 : OAI22_X1 port map( A1 => n10402, A2 => n10501, B1 => n8783, B2 => 
                           n7852, ZN => n2102);
   U9189 : OAI22_X1 port map( A1 => n10402, A2 => n10504, B1 => n8783, B2 => 
                           n7851, ZN => n2103);
   U9190 : OAI22_X1 port map( A1 => n10402, A2 => n10507, B1 => n8783, B2 => 
                           n7850, ZN => n2104);
   U9191 : OAI22_X1 port map( A1 => n10402, A2 => n10510, B1 => n8783, B2 => 
                           n7849, ZN => n2105);
   U9192 : OAI22_X1 port map( A1 => n10403, A2 => n10513, B1 => n8783, B2 => 
                           n7848, ZN => n2106);
   U9193 : OAI22_X1 port map( A1 => n10403, A2 => n10525, B1 => n8783, B2 => 
                           n7847, ZN => n2107);
   U9194 : OAI22_X1 port map( A1 => n10410, A2 => n10495, B1 => n8781, B2 => 
                           n7822, ZN => n2132);
   U9195 : OAI22_X1 port map( A1 => n10411, A2 => n10498, B1 => n8781, B2 => 
                           n7821, ZN => n2133);
   U9196 : OAI22_X1 port map( A1 => n10411, A2 => n10501, B1 => n8781, B2 => 
                           n7820, ZN => n2134);
   U9197 : OAI22_X1 port map( A1 => n10411, A2 => n10504, B1 => n8781, B2 => 
                           n7819, ZN => n2135);
   U9198 : OAI22_X1 port map( A1 => n10411, A2 => n10507, B1 => n8781, B2 => 
                           n7818, ZN => n2136);
   U9199 : OAI22_X1 port map( A1 => n10411, A2 => n10510, B1 => n8781, B2 => 
                           n7817, ZN => n2137);
   U9200 : OAI22_X1 port map( A1 => n10412, A2 => n10513, B1 => n8781, B2 => 
                           n7816, ZN => n2138);
   U9201 : OAI22_X1 port map( A1 => n10412, A2 => n10525, B1 => n8781, B2 => 
                           n7815, ZN => n2139);
   U9202 : OAI22_X1 port map( A1 => n10419, A2 => n10495, B1 => n8779, B2 => 
                           n7790, ZN => n2164);
   U9203 : OAI22_X1 port map( A1 => n10420, A2 => n10498, B1 => n8779, B2 => 
                           n7789, ZN => n2165);
   U9204 : OAI22_X1 port map( A1 => n10420, A2 => n10501, B1 => n8779, B2 => 
                           n7788, ZN => n2166);
   U9205 : OAI22_X1 port map( A1 => n10420, A2 => n10504, B1 => n8779, B2 => 
                           n7787, ZN => n2167);
   U9206 : OAI22_X1 port map( A1 => n10420, A2 => n10507, B1 => n8779, B2 => 
                           n7786, ZN => n2168);
   U9207 : OAI22_X1 port map( A1 => n10420, A2 => n10510, B1 => n8779, B2 => 
                           n7785, ZN => n2169);
   U9208 : OAI22_X1 port map( A1 => n10421, A2 => n10513, B1 => n8779, B2 => 
                           n7784, ZN => n2170);
   U9209 : OAI22_X1 port map( A1 => n10421, A2 => n10525, B1 => n8779, B2 => 
                           n7783, ZN => n2171);
   U9210 : OAI22_X1 port map( A1 => n10521, A2 => n10495, B1 => n8745, B2 => 
                           n7758, ZN => n2196);
   U9211 : OAI22_X1 port map( A1 => n10522, A2 => n10498, B1 => n8745, B2 => 
                           n7757, ZN => n2197);
   U9212 : OAI22_X1 port map( A1 => n10522, A2 => n10501, B1 => n8745, B2 => 
                           n7756, ZN => n2198);
   U9213 : OAI22_X1 port map( A1 => n10522, A2 => n10504, B1 => n8745, B2 => 
                           n7755, ZN => n2199);
   U9214 : OAI22_X1 port map( A1 => n10522, A2 => n10507, B1 => n8745, B2 => 
                           n7754, ZN => n2200);
   U9215 : OAI22_X1 port map( A1 => n10522, A2 => n10510, B1 => n8745, B2 => 
                           n7753, ZN => n2201);
   U9216 : OAI22_X1 port map( A1 => n10523, A2 => n10513, B1 => n8745, B2 => 
                           n7752, ZN => n2202);
   U9217 : OAI22_X1 port map( A1 => n10523, A2 => n10525, B1 => n8745, B2 => 
                           n7751, ZN => n2203);
   U9218 : AOI22_X1 port map( A1 => n10096, A2 => n9636, B1 => n10083, B2 => 
                           n9780, ZN => n9494);
   U9219 : AOI22_X1 port map( A1 => n10096, A2 => n9637, B1 => n10083, B2 => 
                           n9781, ZN => n9474);
   U9220 : AOI22_X1 port map( A1 => n10096, A2 => n9638, B1 => n10083, B2 => 
                           n9782, ZN => n9454);
   U9221 : AOI22_X1 port map( A1 => n10097, A2 => n9639, B1 => n10084, B2 => 
                           n9783, ZN => n9434);
   U9222 : AOI22_X1 port map( A1 => n10097, A2 => n9640, B1 => n10084, B2 => 
                           n9784, ZN => n9414);
   U9223 : AOI22_X1 port map( A1 => n10097, A2 => n9641, B1 => n10084, B2 => 
                           n9785, ZN => n9394);
   U9224 : AOI22_X1 port map( A1 => n10098, A2 => n9642, B1 => n10085, B2 => 
                           n9786, ZN => n9374);
   U9225 : AOI22_X1 port map( A1 => n10098, A2 => n9643, B1 => n10085, B2 => 
                           n9787, ZN => n9354);
   U9226 : AOI22_X1 port map( A1 => n10098, A2 => n9644, B1 => n10085, B2 => 
                           n9788, ZN => n9334);
   U9227 : AOI22_X1 port map( A1 => n10099, A2 => n9645, B1 => n10086, B2 => 
                           n9789, ZN => n9314);
   U9228 : AOI22_X1 port map( A1 => n10099, A2 => n9646, B1 => n10086, B2 => 
                           n9790, ZN => n9294);
   U9229 : AOI22_X1 port map( A1 => n10099, A2 => n9647, B1 => n10086, B2 => 
                           n9791, ZN => n9274);
   U9230 : AOI22_X1 port map( A1 => n10100, A2 => n9648, B1 => n10087, B2 => 
                           n9792, ZN => n9254);
   U9231 : AOI22_X1 port map( A1 => n10100, A2 => n9649, B1 => n10087, B2 => 
                           n9793, ZN => n9234);
   U9232 : AOI22_X1 port map( A1 => n10100, A2 => n9650, B1 => n10087, B2 => 
                           n9794, ZN => n9214);
   U9233 : AOI22_X1 port map( A1 => n10101, A2 => n9651, B1 => n10088, B2 => 
                           n9795, ZN => n9194);
   U9234 : AOI22_X1 port map( A1 => n10101, A2 => n9652, B1 => n10088, B2 => 
                           n9796, ZN => n9174);
   U9235 : AOI22_X1 port map( A1 => n10101, A2 => n9653, B1 => n10088, B2 => 
                           n9797, ZN => n9154);
   U9236 : AOI22_X1 port map( A1 => n10102, A2 => n9654, B1 => n10089, B2 => 
                           n9798, ZN => n9134);
   U9237 : AOI22_X1 port map( A1 => n10102, A2 => n9655, B1 => n10089, B2 => 
                           n9799, ZN => n9114);
   U9238 : AOI22_X1 port map( A1 => n10102, A2 => n9656, B1 => n10089, B2 => 
                           n9800, ZN => n9094);
   U9239 : AOI22_X1 port map( A1 => n10103, A2 => n9657, B1 => n10090, B2 => 
                           n9801, ZN => n9074);
   U9240 : AOI22_X1 port map( A1 => n10103, A2 => n9658, B1 => n10090, B2 => 
                           n9802, ZN => n9054);
   U9241 : AOI22_X1 port map( A1 => n10103, A2 => n9659, B1 => n10090, B2 => 
                           n9803, ZN => n9034);
   U9242 : AOI22_X1 port map( A1 => n10104, A2 => n9516, B1 => n10091, B2 => 
                           n9568, ZN => n9014);
   U9243 : AOI22_X1 port map( A1 => n10104, A2 => n9517, B1 => n10091, B2 => 
                           n9569, ZN => n8994);
   U9244 : AOI22_X1 port map( A1 => n10104, A2 => n9518, B1 => n10091, B2 => 
                           n9570, ZN => n8974);
   U9245 : AOI22_X1 port map( A1 => n10105, A2 => n9519, B1 => n10092, B2 => 
                           n9571, ZN => n8954);
   U9246 : AOI22_X1 port map( A1 => n10105, A2 => n9520, B1 => n10092, B2 => 
                           n9572, ZN => n8934);
   U9247 : AOI22_X1 port map( A1 => n10105, A2 => n9521, B1 => n10092, B2 => 
                           n9573, ZN => n8914);
   U9248 : OAI221_X1 port map( B1 => n8548, B2 => n10070, C1 => n8292, C2 => 
                           n10057, A => n9499, ZN => n9496);
   U9249 : AOI22_X1 port map( A1 => n10044, A2 => n9732, B1 => n10031, B2 => 
                           n9876, ZN => n9499);
   U9250 : OAI221_X1 port map( B1 => n8516, B2 => n10070, C1 => n8260, C2 => 
                           n10057, A => n9503, ZN => n9500);
   U9251 : AOI22_X1 port map( A1 => n10044, A2 => n9900, B1 => n10031, B2 => 
                           n9901, ZN => n9503);
   U9252 : OAI221_X1 port map( B1 => n8612, B2 => n10070, C1 => n8356, C2 => 
                           n10057, A => n9507, ZN => n9504);
   U9253 : AOI22_X1 port map( A1 => n10044, A2 => n9684, B1 => n10031, B2 => 
                           n9828, ZN => n9507);
   U9254 : OAI221_X1 port map( B1 => n8547, B2 => n10070, C1 => n8291, C2 => 
                           n10057, A => n9479, ZN => n9476);
   U9255 : AOI22_X1 port map( A1 => n10044, A2 => n9733, B1 => n10031, B2 => 
                           n9877, ZN => n9479);
   U9256 : OAI221_X1 port map( B1 => n8515, B2 => n10070, C1 => n8259, C2 => 
                           n10057, A => n9483, ZN => n9480);
   U9257 : AOI22_X1 port map( A1 => n10044, A2 => n9904, B1 => n10031, B2 => 
                           n9905, ZN => n9483);
   U9258 : OAI221_X1 port map( B1 => n8611, B2 => n10070, C1 => n8355, C2 => 
                           n10057, A => n9487, ZN => n9484);
   U9259 : AOI22_X1 port map( A1 => n10044, A2 => n9685, B1 => n10031, B2 => 
                           n9829, ZN => n9487);
   U9260 : OAI221_X1 port map( B1 => n8546, B2 => n10070, C1 => n8290, C2 => 
                           n10057, A => n9459, ZN => n9456);
   U9261 : AOI22_X1 port map( A1 => n10044, A2 => n9734, B1 => n10031, B2 => 
                           n9878, ZN => n9459);
   U9262 : OAI221_X1 port map( B1 => n8514, B2 => n10070, C1 => n8258, C2 => 
                           n10057, A => n9463, ZN => n9460);
   U9263 : AOI22_X1 port map( A1 => n10044, A2 => n9908, B1 => n10031, B2 => 
                           n9909, ZN => n9463);
   U9264 : OAI221_X1 port map( B1 => n8610, B2 => n10070, C1 => n8354, C2 => 
                           n10057, A => n9467, ZN => n9464);
   U9265 : AOI22_X1 port map( A1 => n10044, A2 => n9686, B1 => n10031, B2 => 
                           n9830, ZN => n9467);
   U9266 : OAI221_X1 port map( B1 => n8545, B2 => n10071, C1 => n8289, C2 => 
                           n10058, A => n9439, ZN => n9436);
   U9267 : AOI22_X1 port map( A1 => n10045, A2 => n9735, B1 => n10032, B2 => 
                           n9879, ZN => n9439);
   U9268 : OAI221_X1 port map( B1 => n8513, B2 => n10071, C1 => n8257, C2 => 
                           n10058, A => n9443, ZN => n9440);
   U9269 : AOI22_X1 port map( A1 => n10045, A2 => n9912, B1 => n10032, B2 => 
                           n9913, ZN => n9443);
   U9270 : OAI221_X1 port map( B1 => n8609, B2 => n10071, C1 => n8353, C2 => 
                           n10058, A => n9447, ZN => n9444);
   U9271 : AOI22_X1 port map( A1 => n10045, A2 => n9687, B1 => n10032, B2 => 
                           n9831, ZN => n9447);
   U9272 : OAI221_X1 port map( B1 => n8544, B2 => n10071, C1 => n8288, C2 => 
                           n10058, A => n9419, ZN => n9416);
   U9273 : AOI22_X1 port map( A1 => n10045, A2 => n9736, B1 => n10032, B2 => 
                           n9880, ZN => n9419);
   U9274 : OAI221_X1 port map( B1 => n8512, B2 => n10071, C1 => n8256, C2 => 
                           n10058, A => n9423, ZN => n9420);
   U9275 : AOI22_X1 port map( A1 => n10045, A2 => n9916, B1 => n10032, B2 => 
                           n9917, ZN => n9423);
   U9276 : OAI221_X1 port map( B1 => n8608, B2 => n10071, C1 => n8352, C2 => 
                           n10058, A => n9427, ZN => n9424);
   U9277 : AOI22_X1 port map( A1 => n10045, A2 => n9688, B1 => n10032, B2 => 
                           n9832, ZN => n9427);
   U9278 : OAI221_X1 port map( B1 => n8543, B2 => n10071, C1 => n8287, C2 => 
                           n10058, A => n9399, ZN => n9396);
   U9279 : AOI22_X1 port map( A1 => n10045, A2 => n9737, B1 => n10032, B2 => 
                           n9881, ZN => n9399);
   U9280 : OAI221_X1 port map( B1 => n8511, B2 => n10071, C1 => n8255, C2 => 
                           n10058, A => n9403, ZN => n9400);
   U9281 : AOI22_X1 port map( A1 => n10045, A2 => n9920, B1 => n10032, B2 => 
                           n9921, ZN => n9403);
   U9282 : OAI221_X1 port map( B1 => n8607, B2 => n10071, C1 => n8351, C2 => 
                           n10058, A => n9407, ZN => n9404);
   U9283 : AOI22_X1 port map( A1 => n10045, A2 => n9689, B1 => n10032, B2 => 
                           n9833, ZN => n9407);
   U9284 : OAI221_X1 port map( B1 => n8542, B2 => n10072, C1 => n8286, C2 => 
                           n10059, A => n9379, ZN => n9376);
   U9285 : AOI22_X1 port map( A1 => n10046, A2 => n9738, B1 => n10033, B2 => 
                           n9882, ZN => n9379);
   U9286 : OAI221_X1 port map( B1 => n8510, B2 => n10072, C1 => n8254, C2 => 
                           n10059, A => n9383, ZN => n9380);
   U9287 : AOI22_X1 port map( A1 => n10046, A2 => n9924, B1 => n10033, B2 => 
                           n9925, ZN => n9383);
   U9288 : OAI221_X1 port map( B1 => n8606, B2 => n10072, C1 => n8350, C2 => 
                           n10059, A => n9387, ZN => n9384);
   U9289 : AOI22_X1 port map( A1 => n10046, A2 => n9690, B1 => n10033, B2 => 
                           n9834, ZN => n9387);
   U9290 : OAI221_X1 port map( B1 => n8541, B2 => n10072, C1 => n8285, C2 => 
                           n10059, A => n9359, ZN => n9356);
   U9291 : AOI22_X1 port map( A1 => n10046, A2 => n9739, B1 => n10033, B2 => 
                           n9883, ZN => n9359);
   U9292 : OAI221_X1 port map( B1 => n8509, B2 => n10072, C1 => n8253, C2 => 
                           n10059, A => n9363, ZN => n9360);
   U9293 : AOI22_X1 port map( A1 => n10046, A2 => n9928, B1 => n10033, B2 => 
                           n9929, ZN => n9363);
   U9294 : OAI221_X1 port map( B1 => n8605, B2 => n10072, C1 => n8349, C2 => 
                           n10059, A => n9367, ZN => n9364);
   U9295 : AOI22_X1 port map( A1 => n10046, A2 => n9691, B1 => n10033, B2 => 
                           n9835, ZN => n9367);
   U9296 : OAI221_X1 port map( B1 => n8540, B2 => n10072, C1 => n8284, C2 => 
                           n10059, A => n9339, ZN => n9336);
   U9297 : AOI22_X1 port map( A1 => n10046, A2 => n9740, B1 => n10033, B2 => 
                           n9884, ZN => n9339);
   U9298 : OAI221_X1 port map( B1 => n8508, B2 => n10072, C1 => n8252, C2 => 
                           n10059, A => n9343, ZN => n9340);
   U9299 : AOI22_X1 port map( A1 => n10046, A2 => n9932, B1 => n10033, B2 => 
                           n9933, ZN => n9343);
   U9300 : OAI221_X1 port map( B1 => n8604, B2 => n10072, C1 => n8348, C2 => 
                           n10059, A => n9347, ZN => n9344);
   U9301 : AOI22_X1 port map( A1 => n10046, A2 => n9692, B1 => n10033, B2 => 
                           n9836, ZN => n9347);
   U9302 : OAI221_X1 port map( B1 => n8539, B2 => n10073, C1 => n8283, C2 => 
                           n10060, A => n9319, ZN => n9316);
   U9303 : AOI22_X1 port map( A1 => n10047, A2 => n9741, B1 => n10034, B2 => 
                           n9885, ZN => n9319);
   U9304 : OAI221_X1 port map( B1 => n8507, B2 => n10073, C1 => n8251, C2 => 
                           n10060, A => n9323, ZN => n9320);
   U9305 : AOI22_X1 port map( A1 => n10047, A2 => n9936, B1 => n10034, B2 => 
                           n9937, ZN => n9323);
   U9306 : OAI221_X1 port map( B1 => n8603, B2 => n10073, C1 => n8347, C2 => 
                           n10060, A => n9327, ZN => n9324);
   U9307 : AOI22_X1 port map( A1 => n10047, A2 => n9693, B1 => n10034, B2 => 
                           n9837, ZN => n9327);
   U9308 : OAI221_X1 port map( B1 => n8538, B2 => n10073, C1 => n8282, C2 => 
                           n10060, A => n9299, ZN => n9296);
   U9309 : AOI22_X1 port map( A1 => n10047, A2 => n9742, B1 => n10034, B2 => 
                           n9886, ZN => n9299);
   U9310 : OAI221_X1 port map( B1 => n8506, B2 => n10073, C1 => n8250, C2 => 
                           n10060, A => n9303, ZN => n9300);
   U9311 : AOI22_X1 port map( A1 => n10047, A2 => n9940, B1 => n10034, B2 => 
                           n9941, ZN => n9303);
   U9312 : OAI221_X1 port map( B1 => n8602, B2 => n10073, C1 => n8346, C2 => 
                           n10060, A => n9307, ZN => n9304);
   U9313 : AOI22_X1 port map( A1 => n10047, A2 => n9694, B1 => n10034, B2 => 
                           n9838, ZN => n9307);
   U9314 : OAI221_X1 port map( B1 => n8537, B2 => n10073, C1 => n8281, C2 => 
                           n10060, A => n9279, ZN => n9276);
   U9315 : AOI22_X1 port map( A1 => n10047, A2 => n9743, B1 => n10034, B2 => 
                           n9887, ZN => n9279);
   U9316 : OAI221_X1 port map( B1 => n8505, B2 => n10073, C1 => n8249, C2 => 
                           n10060, A => n9283, ZN => n9280);
   U9317 : AOI22_X1 port map( A1 => n10047, A2 => n9944, B1 => n10034, B2 => 
                           n9945, ZN => n9283);
   U9318 : OAI221_X1 port map( B1 => n8601, B2 => n10073, C1 => n8345, C2 => 
                           n10060, A => n9287, ZN => n9284);
   U9319 : AOI22_X1 port map( A1 => n10047, A2 => n9695, B1 => n10034, B2 => 
                           n9839, ZN => n9287);
   U9320 : OAI221_X1 port map( B1 => n8536, B2 => n10074, C1 => n8280, C2 => 
                           n10061, A => n9259, ZN => n9256);
   U9321 : AOI22_X1 port map( A1 => n10048, A2 => n9744, B1 => n10035, B2 => 
                           n9888, ZN => n9259);
   U9322 : OAI221_X1 port map( B1 => n8504, B2 => n10074, C1 => n8248, C2 => 
                           n10061, A => n9263, ZN => n9260);
   U9323 : AOI22_X1 port map( A1 => n10048, A2 => n9948, B1 => n10035, B2 => 
                           n9949, ZN => n9263);
   U9324 : OAI221_X1 port map( B1 => n8600, B2 => n10074, C1 => n8344, C2 => 
                           n10061, A => n9267, ZN => n9264);
   U9325 : AOI22_X1 port map( A1 => n10048, A2 => n9696, B1 => n10035, B2 => 
                           n9840, ZN => n9267);
   U9326 : OAI221_X1 port map( B1 => n8535, B2 => n10074, C1 => n8279, C2 => 
                           n10061, A => n9239, ZN => n9236);
   U9327 : AOI22_X1 port map( A1 => n10048, A2 => n9745, B1 => n10035, B2 => 
                           n9889, ZN => n9239);
   U9328 : OAI221_X1 port map( B1 => n8503, B2 => n10074, C1 => n8247, C2 => 
                           n10061, A => n9243, ZN => n9240);
   U9329 : AOI22_X1 port map( A1 => n10048, A2 => n9952, B1 => n10035, B2 => 
                           n9953, ZN => n9243);
   U9330 : OAI221_X1 port map( B1 => n8599, B2 => n10074, C1 => n8343, C2 => 
                           n10061, A => n9247, ZN => n9244);
   U9331 : AOI22_X1 port map( A1 => n10048, A2 => n9697, B1 => n10035, B2 => 
                           n9841, ZN => n9247);
   U9332 : OAI221_X1 port map( B1 => n8534, B2 => n10074, C1 => n8278, C2 => 
                           n10061, A => n9219, ZN => n9216);
   U9333 : AOI22_X1 port map( A1 => n10048, A2 => n9746, B1 => n10035, B2 => 
                           n9890, ZN => n9219);
   U9334 : OAI221_X1 port map( B1 => n8502, B2 => n10074, C1 => n8246, C2 => 
                           n10061, A => n9223, ZN => n9220);
   U9335 : AOI22_X1 port map( A1 => n10048, A2 => n9956, B1 => n10035, B2 => 
                           n9957, ZN => n9223);
   U9336 : OAI221_X1 port map( B1 => n8598, B2 => n10074, C1 => n8342, C2 => 
                           n10061, A => n9227, ZN => n9224);
   U9337 : AOI22_X1 port map( A1 => n10048, A2 => n9698, B1 => n10035, B2 => 
                           n9842, ZN => n9227);
   U9338 : OAI221_X1 port map( B1 => n8533, B2 => n10075, C1 => n8277, C2 => 
                           n10062, A => n9199, ZN => n9196);
   U9339 : AOI22_X1 port map( A1 => n10049, A2 => n9747, B1 => n10036, B2 => 
                           n9891, ZN => n9199);
   U9340 : OAI221_X1 port map( B1 => n8501, B2 => n10075, C1 => n8245, C2 => 
                           n10062, A => n9203, ZN => n9200);
   U9341 : AOI22_X1 port map( A1 => n10049, A2 => n9960, B1 => n10036, B2 => 
                           n9961, ZN => n9203);
   U9342 : OAI221_X1 port map( B1 => n8597, B2 => n10075, C1 => n8341, C2 => 
                           n10062, A => n9207, ZN => n9204);
   U9343 : AOI22_X1 port map( A1 => n10049, A2 => n9699, B1 => n10036, B2 => 
                           n9843, ZN => n9207);
   U9344 : OAI221_X1 port map( B1 => n8532, B2 => n10075, C1 => n8276, C2 => 
                           n10062, A => n9179, ZN => n9176);
   U9345 : AOI22_X1 port map( A1 => n10049, A2 => n9748, B1 => n10036, B2 => 
                           n9892, ZN => n9179);
   U9346 : OAI221_X1 port map( B1 => n8500, B2 => n10075, C1 => n8244, C2 => 
                           n10062, A => n9183, ZN => n9180);
   U9347 : AOI22_X1 port map( A1 => n10049, A2 => n9964, B1 => n10036, B2 => 
                           n9965, ZN => n9183);
   U9348 : OAI221_X1 port map( B1 => n8596, B2 => n10075, C1 => n8340, C2 => 
                           n10062, A => n9187, ZN => n9184);
   U9349 : AOI22_X1 port map( A1 => n10049, A2 => n9700, B1 => n10036, B2 => 
                           n9844, ZN => n9187);
   U9350 : OAI221_X1 port map( B1 => n8531, B2 => n10075, C1 => n8275, C2 => 
                           n10062, A => n9159, ZN => n9156);
   U9351 : AOI22_X1 port map( A1 => n10049, A2 => n9749, B1 => n10036, B2 => 
                           n9893, ZN => n9159);
   U9352 : OAI221_X1 port map( B1 => n8499, B2 => n10075, C1 => n8243, C2 => 
                           n10062, A => n9163, ZN => n9160);
   U9353 : AOI22_X1 port map( A1 => n10049, A2 => n9968, B1 => n10036, B2 => 
                           n9969, ZN => n9163);
   U9354 : OAI221_X1 port map( B1 => n8595, B2 => n10075, C1 => n8339, C2 => 
                           n10062, A => n9167, ZN => n9164);
   U9355 : AOI22_X1 port map( A1 => n10049, A2 => n9701, B1 => n10036, B2 => 
                           n9845, ZN => n9167);
   U9356 : OAI221_X1 port map( B1 => n8530, B2 => n10076, C1 => n8274, C2 => 
                           n10063, A => n9139, ZN => n9136);
   U9357 : AOI22_X1 port map( A1 => n10050, A2 => n9750, B1 => n10037, B2 => 
                           n9894, ZN => n9139);
   U9358 : OAI221_X1 port map( B1 => n8498, B2 => n10076, C1 => n8242, C2 => 
                           n10063, A => n9143, ZN => n9140);
   U9359 : AOI22_X1 port map( A1 => n10050, A2 => n9972, B1 => n10037, B2 => 
                           n9973, ZN => n9143);
   U9360 : OAI221_X1 port map( B1 => n8594, B2 => n10076, C1 => n8338, C2 => 
                           n10063, A => n9147, ZN => n9144);
   U9361 : AOI22_X1 port map( A1 => n10050, A2 => n9702, B1 => n10037, B2 => 
                           n9846, ZN => n9147);
   U9362 : OAI221_X1 port map( B1 => n8529, B2 => n10076, C1 => n8273, C2 => 
                           n10063, A => n9119, ZN => n9116);
   U9363 : AOI22_X1 port map( A1 => n10050, A2 => n9751, B1 => n10037, B2 => 
                           n9895, ZN => n9119);
   U9364 : OAI221_X1 port map( B1 => n8497, B2 => n10076, C1 => n8241, C2 => 
                           n10063, A => n9123, ZN => n9120);
   U9365 : AOI22_X1 port map( A1 => n10050, A2 => n9976, B1 => n10037, B2 => 
                           n9977, ZN => n9123);
   U9366 : OAI221_X1 port map( B1 => n8593, B2 => n10076, C1 => n8337, C2 => 
                           n10063, A => n9127, ZN => n9124);
   U9367 : AOI22_X1 port map( A1 => n10050, A2 => n9703, B1 => n10037, B2 => 
                           n9847, ZN => n9127);
   U9368 : OAI221_X1 port map( B1 => n8528, B2 => n10076, C1 => n8272, C2 => 
                           n10063, A => n9099, ZN => n9096);
   U9369 : AOI22_X1 port map( A1 => n10050, A2 => n9752, B1 => n10037, B2 => 
                           n9896, ZN => n9099);
   U9370 : OAI221_X1 port map( B1 => n8496, B2 => n10076, C1 => n8240, C2 => 
                           n10063, A => n9103, ZN => n9100);
   U9371 : AOI22_X1 port map( A1 => n10050, A2 => n9980, B1 => n10037, B2 => 
                           n9981, ZN => n9103);
   U9372 : OAI221_X1 port map( B1 => n8592, B2 => n10076, C1 => n8336, C2 => 
                           n10063, A => n9107, ZN => n9104);
   U9373 : AOI22_X1 port map( A1 => n10050, A2 => n9704, B1 => n10037, B2 => 
                           n9848, ZN => n9107);
   U9374 : OAI221_X1 port map( B1 => n8527, B2 => n10077, C1 => n8271, C2 => 
                           n10064, A => n9079, ZN => n9076);
   U9375 : AOI22_X1 port map( A1 => n10051, A2 => n9753, B1 => n10038, B2 => 
                           n9897, ZN => n9079);
   U9376 : OAI221_X1 port map( B1 => n8495, B2 => n10077, C1 => n8239, C2 => 
                           n10064, A => n9083, ZN => n9080);
   U9377 : AOI22_X1 port map( A1 => n10051, A2 => n9984, B1 => n10038, B2 => 
                           n9985, ZN => n9083);
   U9378 : OAI221_X1 port map( B1 => n8591, B2 => n10077, C1 => n8335, C2 => 
                           n10064, A => n9087, ZN => n9084);
   U9379 : AOI22_X1 port map( A1 => n10051, A2 => n9705, B1 => n10038, B2 => 
                           n9849, ZN => n9087);
   U9380 : OAI221_X1 port map( B1 => n8526, B2 => n10077, C1 => n8270, C2 => 
                           n10064, A => n9059, ZN => n9056);
   U9381 : AOI22_X1 port map( A1 => n10051, A2 => n9754, B1 => n10038, B2 => 
                           n9898, ZN => n9059);
   U9382 : OAI221_X1 port map( B1 => n8494, B2 => n10077, C1 => n8238, C2 => 
                           n10064, A => n9063, ZN => n9060);
   U9383 : AOI22_X1 port map( A1 => n10051, A2 => n9988, B1 => n10038, B2 => 
                           n9989, ZN => n9063);
   U9384 : OAI221_X1 port map( B1 => n8590, B2 => n10077, C1 => n8334, C2 => 
                           n10064, A => n9067, ZN => n9064);
   U9385 : AOI22_X1 port map( A1 => n10051, A2 => n9706, B1 => n10038, B2 => 
                           n9850, ZN => n9067);
   U9386 : OAI221_X1 port map( B1 => n8525, B2 => n10077, C1 => n8269, C2 => 
                           n10064, A => n9039, ZN => n9036);
   U9387 : AOI22_X1 port map( A1 => n10051, A2 => n9755, B1 => n10038, B2 => 
                           n9899, ZN => n9039);
   U9388 : OAI221_X1 port map( B1 => n8493, B2 => n10077, C1 => n8237, C2 => 
                           n10064, A => n9043, ZN => n9040);
   U9389 : AOI22_X1 port map( A1 => n10051, A2 => n9992, B1 => n10038, B2 => 
                           n9993, ZN => n9043);
   U9390 : OAI221_X1 port map( B1 => n8589, B2 => n10077, C1 => n8333, C2 => 
                           n10064, A => n9047, ZN => n9044);
   U9391 : AOI22_X1 port map( A1 => n10051, A2 => n9707, B1 => n10038, B2 => 
                           n9851, ZN => n9047);
   U9392 : OAI221_X1 port map( B1 => n8524, B2 => n10078, C1 => n8268, C2 => 
                           n10065, A => n9019, ZN => n9016);
   U9393 : AOI22_X1 port map( A1 => n10052, A2 => n9550, B1 => n10039, B2 => 
                           n9602, ZN => n9019);
   U9394 : OAI221_X1 port map( B1 => n8492, B2 => n10078, C1 => n8236, C2 => 
                           n10065, A => n9023, ZN => n9020);
   U9395 : AOI22_X1 port map( A1 => n10052, A2 => n9996, B1 => n10039, B2 => 
                           n9997, ZN => n9023);
   U9396 : OAI221_X1 port map( B1 => n8588, B2 => n10078, C1 => n8332, C2 => 
                           n10065, A => n9027, ZN => n9024);
   U9397 : AOI22_X1 port map( A1 => n10052, A2 => n9534, B1 => n10039, B2 => 
                           n9586, ZN => n9027);
   U9398 : OAI221_X1 port map( B1 => n8523, B2 => n10078, C1 => n8267, C2 => 
                           n10065, A => n8999, ZN => n8996);
   U9399 : AOI22_X1 port map( A1 => n10052, A2 => n9551, B1 => n10039, B2 => 
                           n9603, ZN => n8999);
   U9400 : OAI221_X1 port map( B1 => n8491, B2 => n10078, C1 => n8235, C2 => 
                           n10065, A => n9003, ZN => n9000);
   U9401 : AOI22_X1 port map( A1 => n10052, A2 => n10000, B1 => n10039, B2 => 
                           n10001, ZN => n9003);
   U9402 : OAI221_X1 port map( B1 => n8587, B2 => n10078, C1 => n8331, C2 => 
                           n10065, A => n9007, ZN => n9004);
   U9403 : AOI22_X1 port map( A1 => n10052, A2 => n9535, B1 => n10039, B2 => 
                           n9587, ZN => n9007);
   U9404 : OAI221_X1 port map( B1 => n8522, B2 => n10078, C1 => n8266, C2 => 
                           n10065, A => n8979, ZN => n8976);
   U9405 : AOI22_X1 port map( A1 => n10052, A2 => n9552, B1 => n10039, B2 => 
                           n9604, ZN => n8979);
   U9406 : OAI221_X1 port map( B1 => n8490, B2 => n10078, C1 => n8234, C2 => 
                           n10065, A => n8983, ZN => n8980);
   U9407 : AOI22_X1 port map( A1 => n10052, A2 => n10004, B1 => n10039, B2 => 
                           n10005, ZN => n8983);
   U9408 : OAI221_X1 port map( B1 => n8586, B2 => n10078, C1 => n8330, C2 => 
                           n10065, A => n8987, ZN => n8984);
   U9409 : AOI22_X1 port map( A1 => n10052, A2 => n9536, B1 => n10039, B2 => 
                           n9588, ZN => n8987);
   U9410 : OAI221_X1 port map( B1 => n8521, B2 => n10079, C1 => n8265, C2 => 
                           n10066, A => n8959, ZN => n8956);
   U9411 : AOI22_X1 port map( A1 => n10053, A2 => n9553, B1 => n10040, B2 => 
                           n9605, ZN => n8959);
   U9412 : OAI221_X1 port map( B1 => n8489, B2 => n10079, C1 => n8233, C2 => 
                           n10066, A => n8963, ZN => n8960);
   U9413 : AOI22_X1 port map( A1 => n10053, A2 => n10008, B1 => n10040, B2 => 
                           n10009, ZN => n8963);
   U9414 : OAI221_X1 port map( B1 => n8585, B2 => n10079, C1 => n8329, C2 => 
                           n10066, A => n8967, ZN => n8964);
   U9415 : AOI22_X1 port map( A1 => n10053, A2 => n9537, B1 => n10040, B2 => 
                           n9589, ZN => n8967);
   U9416 : OAI221_X1 port map( B1 => n8520, B2 => n10079, C1 => n8264, C2 => 
                           n10066, A => n8939, ZN => n8936);
   U9417 : AOI22_X1 port map( A1 => n10053, A2 => n9554, B1 => n10040, B2 => 
                           n9606, ZN => n8939);
   U9418 : OAI221_X1 port map( B1 => n8488, B2 => n10079, C1 => n8232, C2 => 
                           n10066, A => n8943, ZN => n8940);
   U9419 : AOI22_X1 port map( A1 => n10053, A2 => n10012, B1 => n10040, B2 => 
                           n10013, ZN => n8943);
   U9420 : OAI221_X1 port map( B1 => n8584, B2 => n10079, C1 => n8328, C2 => 
                           n10066, A => n8947, ZN => n8944);
   U9421 : AOI22_X1 port map( A1 => n10053, A2 => n9538, B1 => n10040, B2 => 
                           n9590, ZN => n8947);
   U9422 : OAI221_X1 port map( B1 => n8519, B2 => n10079, C1 => n8263, C2 => 
                           n10066, A => n8919, ZN => n8916);
   U9423 : AOI22_X1 port map( A1 => n10053, A2 => n9555, B1 => n10040, B2 => 
                           n9607, ZN => n8919);
   U9424 : OAI221_X1 port map( B1 => n8487, B2 => n10079, C1 => n8231, C2 => 
                           n10066, A => n8923, ZN => n8920);
   U9425 : AOI22_X1 port map( A1 => n10053, A2 => n10016, B1 => n10040, B2 => 
                           n10017, ZN => n8923);
   U9426 : OAI221_X1 port map( B1 => n8583, B2 => n10079, C1 => n8327, C2 => 
                           n10066, A => n8927, ZN => n8924);
   U9427 : AOI22_X1 port map( A1 => n10053, A2 => n9539, B1 => n10040, B2 => 
                           n9591, ZN => n8927);
   U9428 : OAI22_X1 port map( A1 => n10361, A2 => n10423, B1 => n10360, B2 => 
                           n8006, ZN => n1948);
   U9429 : OAI22_X1 port map( A1 => n10361, A2 => n10426, B1 => n10360, B2 => 
                           n8005, ZN => n1949);
   U9430 : OAI22_X1 port map( A1 => n10361, A2 => n10429, B1 => n10360, B2 => 
                           n8004, ZN => n1950);
   U9431 : OAI22_X1 port map( A1 => n10361, A2 => n10432, B1 => n10360, B2 => 
                           n8003, ZN => n1951);
   U9432 : OAI22_X1 port map( A1 => n10361, A2 => n10435, B1 => n10360, B2 => 
                           n8002, ZN => n1952);
   U9433 : OAI22_X1 port map( A1 => n10362, A2 => n10438, B1 => n10360, B2 => 
                           n8001, ZN => n1953);
   U9434 : OAI22_X1 port map( A1 => n10362, A2 => n10441, B1 => n10360, B2 => 
                           n8000, ZN => n1954);
   U9435 : OAI22_X1 port map( A1 => n10362, A2 => n10444, B1 => n10360, B2 => 
                           n7999, ZN => n1955);
   U9436 : OAI22_X1 port map( A1 => n10362, A2 => n10447, B1 => n10360, B2 => 
                           n7998, ZN => n1956);
   U9437 : OAI22_X1 port map( A1 => n10362, A2 => n10450, B1 => n10360, B2 => 
                           n7997, ZN => n1957);
   U9438 : OAI22_X1 port map( A1 => n10363, A2 => n10453, B1 => n10360, B2 => 
                           n7996, ZN => n1958);
   U9439 : OAI22_X1 port map( A1 => n10363, A2 => n10456, B1 => n10360, B2 => 
                           n7995, ZN => n1959);
   U9440 : OAI22_X1 port map( A1 => n10363, A2 => n10459, B1 => n8790, B2 => 
                           n7994, ZN => n1960);
   U9441 : OAI22_X1 port map( A1 => n10363, A2 => n10462, B1 => n8790, B2 => 
                           n7993, ZN => n1961);
   U9442 : OAI22_X1 port map( A1 => n10363, A2 => n10465, B1 => n8790, B2 => 
                           n7992, ZN => n1962);
   U9443 : OAI22_X1 port map( A1 => n10364, A2 => n10468, B1 => n10360, B2 => 
                           n7991, ZN => n1963);
   U9444 : OAI22_X1 port map( A1 => n10364, A2 => n10471, B1 => n10360, B2 => 
                           n7990, ZN => n1964);
   U9445 : OAI22_X1 port map( A1 => n10364, A2 => n10474, B1 => n10360, B2 => 
                           n7989, ZN => n1965);
   U9446 : OAI22_X1 port map( A1 => n10364, A2 => n10477, B1 => n10360, B2 => 
                           n7988, ZN => n1966);
   U9447 : OAI22_X1 port map( A1 => n10364, A2 => n10480, B1 => n10360, B2 => 
                           n7987, ZN => n1967);
   U9448 : OAI22_X1 port map( A1 => n10365, A2 => n10483, B1 => n10360, B2 => 
                           n7986, ZN => n1968);
   U9449 : OAI22_X1 port map( A1 => n10365, A2 => n10486, B1 => n10360, B2 => 
                           n7985, ZN => n1969);
   U9450 : OAI22_X1 port map( A1 => n10365, A2 => n10489, B1 => n10360, B2 => 
                           n7984, ZN => n1970);
   U9451 : OAI22_X1 port map( A1 => n10365, A2 => n10492, B1 => n10360, B2 => 
                           n7983, ZN => n1971);
   U9452 : OAI22_X1 port map( A1 => n10370, A2 => n10423, B1 => n10369, B2 => 
                           n7974, ZN => n1980);
   U9453 : OAI22_X1 port map( A1 => n10370, A2 => n10426, B1 => n10369, B2 => 
                           n7973, ZN => n1981);
   U9454 : OAI22_X1 port map( A1 => n10370, A2 => n10429, B1 => n10369, B2 => 
                           n7972, ZN => n1982);
   U9455 : OAI22_X1 port map( A1 => n10370, A2 => n10432, B1 => n10369, B2 => 
                           n7971, ZN => n1983);
   U9456 : OAI22_X1 port map( A1 => n10370, A2 => n10435, B1 => n10369, B2 => 
                           n7970, ZN => n1984);
   U9457 : OAI22_X1 port map( A1 => n10371, A2 => n10438, B1 => n10369, B2 => 
                           n7969, ZN => n1985);
   U9458 : OAI22_X1 port map( A1 => n10371, A2 => n10441, B1 => n10369, B2 => 
                           n7968, ZN => n1986);
   U9459 : OAI22_X1 port map( A1 => n10371, A2 => n10444, B1 => n10369, B2 => 
                           n7967, ZN => n1987);
   U9460 : OAI22_X1 port map( A1 => n10371, A2 => n10447, B1 => n10369, B2 => 
                           n7966, ZN => n1988);
   U9461 : OAI22_X1 port map( A1 => n10371, A2 => n10450, B1 => n10369, B2 => 
                           n7965, ZN => n1989);
   U9462 : OAI22_X1 port map( A1 => n10372, A2 => n10453, B1 => n10369, B2 => 
                           n7964, ZN => n1990);
   U9463 : OAI22_X1 port map( A1 => n10372, A2 => n10456, B1 => n10369, B2 => 
                           n7963, ZN => n1991);
   U9464 : OAI22_X1 port map( A1 => n10372, A2 => n10459, B1 => n8789, B2 => 
                           n7962, ZN => n1992);
   U9465 : OAI22_X1 port map( A1 => n10372, A2 => n10462, B1 => n8789, B2 => 
                           n7961, ZN => n1993);
   U9466 : OAI22_X1 port map( A1 => n10372, A2 => n10465, B1 => n8789, B2 => 
                           n7960, ZN => n1994);
   U9467 : OAI22_X1 port map( A1 => n10373, A2 => n10468, B1 => n10369, B2 => 
                           n7959, ZN => n1995);
   U9468 : OAI22_X1 port map( A1 => n10373, A2 => n10471, B1 => n10369, B2 => 
                           n7958, ZN => n1996);
   U9469 : OAI22_X1 port map( A1 => n10373, A2 => n10474, B1 => n10369, B2 => 
                           n7957, ZN => n1997);
   U9470 : OAI22_X1 port map( A1 => n10373, A2 => n10477, B1 => n10369, B2 => 
                           n7956, ZN => n1998);
   U9471 : OAI22_X1 port map( A1 => n10373, A2 => n10480, B1 => n10369, B2 => 
                           n7955, ZN => n1999);
   U9472 : OAI22_X1 port map( A1 => n10374, A2 => n10483, B1 => n10369, B2 => 
                           n7954, ZN => n2000);
   U9473 : OAI22_X1 port map( A1 => n10374, A2 => n10486, B1 => n10369, B2 => 
                           n7953, ZN => n2001);
   U9474 : OAI22_X1 port map( A1 => n10374, A2 => n10489, B1 => n10369, B2 => 
                           n7952, ZN => n2002);
   U9475 : OAI22_X1 port map( A1 => n10374, A2 => n10492, B1 => n10369, B2 => 
                           n7951, ZN => n2003);
   U9476 : OAI22_X1 port map( A1 => n10379, A2 => n10423, B1 => n10378, B2 => 
                           n7942, ZN => n2012);
   U9477 : OAI22_X1 port map( A1 => n10379, A2 => n10426, B1 => n10378, B2 => 
                           n7941, ZN => n2013);
   U9478 : OAI22_X1 port map( A1 => n10379, A2 => n10429, B1 => n10378, B2 => 
                           n7940, ZN => n2014);
   U9479 : OAI22_X1 port map( A1 => n10379, A2 => n10432, B1 => n10378, B2 => 
                           n7939, ZN => n2015);
   U9480 : OAI22_X1 port map( A1 => n10379, A2 => n10435, B1 => n10378, B2 => 
                           n7938, ZN => n2016);
   U9481 : OAI22_X1 port map( A1 => n10380, A2 => n10438, B1 => n10378, B2 => 
                           n7937, ZN => n2017);
   U9482 : OAI22_X1 port map( A1 => n10380, A2 => n10441, B1 => n10378, B2 => 
                           n7936, ZN => n2018);
   U9483 : OAI22_X1 port map( A1 => n10380, A2 => n10444, B1 => n10378, B2 => 
                           n7935, ZN => n2019);
   U9484 : OAI22_X1 port map( A1 => n10380, A2 => n10447, B1 => n10378, B2 => 
                           n7934, ZN => n2020);
   U9485 : OAI22_X1 port map( A1 => n10380, A2 => n10450, B1 => n10378, B2 => 
                           n7933, ZN => n2021);
   U9486 : OAI22_X1 port map( A1 => n10381, A2 => n10453, B1 => n10378, B2 => 
                           n7932, ZN => n2022);
   U9487 : OAI22_X1 port map( A1 => n10381, A2 => n10456, B1 => n10378, B2 => 
                           n7931, ZN => n2023);
   U9488 : OAI22_X1 port map( A1 => n10381, A2 => n10459, B1 => n8788, B2 => 
                           n7930, ZN => n2024);
   U9489 : OAI22_X1 port map( A1 => n10381, A2 => n10462, B1 => n8788, B2 => 
                           n7929, ZN => n2025);
   U9490 : OAI22_X1 port map( A1 => n10381, A2 => n10465, B1 => n8788, B2 => 
                           n7928, ZN => n2026);
   U9491 : OAI22_X1 port map( A1 => n10382, A2 => n10468, B1 => n10378, B2 => 
                           n7927, ZN => n2027);
   U9492 : OAI22_X1 port map( A1 => n10382, A2 => n10471, B1 => n10378, B2 => 
                           n7926, ZN => n2028);
   U9493 : OAI22_X1 port map( A1 => n10382, A2 => n10474, B1 => n10378, B2 => 
                           n7925, ZN => n2029);
   U9494 : OAI22_X1 port map( A1 => n10382, A2 => n10477, B1 => n10378, B2 => 
                           n7924, ZN => n2030);
   U9495 : OAI22_X1 port map( A1 => n10382, A2 => n10480, B1 => n10378, B2 => 
                           n7923, ZN => n2031);
   U9496 : OAI22_X1 port map( A1 => n10383, A2 => n10483, B1 => n10378, B2 => 
                           n7922, ZN => n2032);
   U9497 : OAI22_X1 port map( A1 => n10383, A2 => n10486, B1 => n10378, B2 => 
                           n7921, ZN => n2033);
   U9498 : OAI22_X1 port map( A1 => n10383, A2 => n10489, B1 => n10378, B2 => 
                           n7920, ZN => n2034);
   U9499 : OAI22_X1 port map( A1 => n10383, A2 => n10492, B1 => n10378, B2 => 
                           n7919, ZN => n2035);
   U9500 : OAI22_X1 port map( A1 => n10388, A2 => n10423, B1 => n10387, B2 => 
                           n7910, ZN => n2044);
   U9501 : OAI22_X1 port map( A1 => n10388, A2 => n10426, B1 => n10387, B2 => 
                           n7909, ZN => n2045);
   U9502 : OAI22_X1 port map( A1 => n10388, A2 => n10429, B1 => n10387, B2 => 
                           n7908, ZN => n2046);
   U9503 : OAI22_X1 port map( A1 => n10388, A2 => n10432, B1 => n10387, B2 => 
                           n7907, ZN => n2047);
   U9504 : OAI22_X1 port map( A1 => n10388, A2 => n10435, B1 => n10387, B2 => 
                           n7906, ZN => n2048);
   U9505 : OAI22_X1 port map( A1 => n10389, A2 => n10438, B1 => n10387, B2 => 
                           n7905, ZN => n2049);
   U9506 : OAI22_X1 port map( A1 => n10389, A2 => n10441, B1 => n10387, B2 => 
                           n7904, ZN => n2050);
   U9507 : OAI22_X1 port map( A1 => n10389, A2 => n10444, B1 => n10387, B2 => 
                           n7903, ZN => n2051);
   U9508 : OAI22_X1 port map( A1 => n10389, A2 => n10447, B1 => n10387, B2 => 
                           n7902, ZN => n2052);
   U9509 : OAI22_X1 port map( A1 => n10389, A2 => n10450, B1 => n10387, B2 => 
                           n7901, ZN => n2053);
   U9510 : OAI22_X1 port map( A1 => n10390, A2 => n10453, B1 => n10387, B2 => 
                           n7900, ZN => n2054);
   U9511 : OAI22_X1 port map( A1 => n10390, A2 => n10456, B1 => n10387, B2 => 
                           n7899, ZN => n2055);
   U9512 : OAI22_X1 port map( A1 => n10390, A2 => n10459, B1 => n8786, B2 => 
                           n7898, ZN => n2056);
   U9513 : OAI22_X1 port map( A1 => n10390, A2 => n10462, B1 => n8786, B2 => 
                           n7897, ZN => n2057);
   U9514 : OAI22_X1 port map( A1 => n10390, A2 => n10465, B1 => n8786, B2 => 
                           n7896, ZN => n2058);
   U9515 : OAI22_X1 port map( A1 => n10391, A2 => n10468, B1 => n10387, B2 => 
                           n7895, ZN => n2059);
   U9516 : OAI22_X1 port map( A1 => n10391, A2 => n10471, B1 => n10387, B2 => 
                           n7894, ZN => n2060);
   U9517 : OAI22_X1 port map( A1 => n10391, A2 => n10474, B1 => n10387, B2 => 
                           n7893, ZN => n2061);
   U9518 : OAI22_X1 port map( A1 => n10391, A2 => n10477, B1 => n10387, B2 => 
                           n7892, ZN => n2062);
   U9519 : OAI22_X1 port map( A1 => n10391, A2 => n10480, B1 => n10387, B2 => 
                           n7891, ZN => n2063);
   U9520 : OAI22_X1 port map( A1 => n10392, A2 => n10483, B1 => n10387, B2 => 
                           n7890, ZN => n2064);
   U9521 : OAI22_X1 port map( A1 => n10392, A2 => n10486, B1 => n10387, B2 => 
                           n7889, ZN => n2065);
   U9522 : OAI22_X1 port map( A1 => n10392, A2 => n10489, B1 => n10387, B2 => 
                           n7888, ZN => n2066);
   U9523 : OAI22_X1 port map( A1 => n10392, A2 => n10492, B1 => n10387, B2 => 
                           n7887, ZN => n2067);
   U9524 : OAI22_X1 port map( A1 => n10397, A2 => n10423, B1 => n10396, B2 => 
                           n7878, ZN => n2076);
   U9525 : OAI22_X1 port map( A1 => n10397, A2 => n10426, B1 => n10396, B2 => 
                           n7877, ZN => n2077);
   U9526 : OAI22_X1 port map( A1 => n10397, A2 => n10429, B1 => n10396, B2 => 
                           n7876, ZN => n2078);
   U9527 : OAI22_X1 port map( A1 => n10397, A2 => n10432, B1 => n10396, B2 => 
                           n7875, ZN => n2079);
   U9528 : OAI22_X1 port map( A1 => n10397, A2 => n10435, B1 => n10396, B2 => 
                           n7874, ZN => n2080);
   U9529 : OAI22_X1 port map( A1 => n10398, A2 => n10438, B1 => n10396, B2 => 
                           n7873, ZN => n2081);
   U9530 : OAI22_X1 port map( A1 => n10398, A2 => n10441, B1 => n10396, B2 => 
                           n7872, ZN => n2082);
   U9531 : OAI22_X1 port map( A1 => n10398, A2 => n10444, B1 => n10396, B2 => 
                           n7871, ZN => n2083);
   U9532 : OAI22_X1 port map( A1 => n10398, A2 => n10447, B1 => n10396, B2 => 
                           n7870, ZN => n2084);
   U9533 : OAI22_X1 port map( A1 => n10398, A2 => n10450, B1 => n10396, B2 => 
                           n7869, ZN => n2085);
   U9534 : OAI22_X1 port map( A1 => n10399, A2 => n10453, B1 => n10396, B2 => 
                           n7868, ZN => n2086);
   U9535 : OAI22_X1 port map( A1 => n10399, A2 => n10456, B1 => n10396, B2 => 
                           n7867, ZN => n2087);
   U9536 : OAI22_X1 port map( A1 => n10399, A2 => n10459, B1 => n8783, B2 => 
                           n7866, ZN => n2088);
   U9537 : OAI22_X1 port map( A1 => n10399, A2 => n10462, B1 => n8783, B2 => 
                           n7865, ZN => n2089);
   U9538 : OAI22_X1 port map( A1 => n10399, A2 => n10465, B1 => n8783, B2 => 
                           n7864, ZN => n2090);
   U9539 : OAI22_X1 port map( A1 => n10400, A2 => n10468, B1 => n10396, B2 => 
                           n7863, ZN => n2091);
   U9540 : OAI22_X1 port map( A1 => n10400, A2 => n10471, B1 => n10396, B2 => 
                           n7862, ZN => n2092);
   U9541 : OAI22_X1 port map( A1 => n10400, A2 => n10474, B1 => n10396, B2 => 
                           n7861, ZN => n2093);
   U9542 : OAI22_X1 port map( A1 => n10400, A2 => n10477, B1 => n10396, B2 => 
                           n7860, ZN => n2094);
   U9543 : OAI22_X1 port map( A1 => n10400, A2 => n10480, B1 => n10396, B2 => 
                           n7859, ZN => n2095);
   U9544 : OAI22_X1 port map( A1 => n10401, A2 => n10483, B1 => n10396, B2 => 
                           n7858, ZN => n2096);
   U9545 : OAI22_X1 port map( A1 => n10401, A2 => n10486, B1 => n10396, B2 => 
                           n7857, ZN => n2097);
   U9546 : OAI22_X1 port map( A1 => n10401, A2 => n10489, B1 => n10396, B2 => 
                           n7856, ZN => n2098);
   U9547 : OAI22_X1 port map( A1 => n10401, A2 => n10492, B1 => n10396, B2 => 
                           n7855, ZN => n2099);
   U9548 : OAI22_X1 port map( A1 => n10406, A2 => n10423, B1 => n10405, B2 => 
                           n7846, ZN => n2108);
   U9549 : OAI22_X1 port map( A1 => n10406, A2 => n10426, B1 => n10405, B2 => 
                           n7845, ZN => n2109);
   U9550 : OAI22_X1 port map( A1 => n10406, A2 => n10429, B1 => n10405, B2 => 
                           n7844, ZN => n2110);
   U9551 : OAI22_X1 port map( A1 => n10406, A2 => n10432, B1 => n10405, B2 => 
                           n7843, ZN => n2111);
   U9552 : OAI22_X1 port map( A1 => n10406, A2 => n10435, B1 => n10405, B2 => 
                           n7842, ZN => n2112);
   U9553 : OAI22_X1 port map( A1 => n10407, A2 => n10438, B1 => n10405, B2 => 
                           n7841, ZN => n2113);
   U9554 : OAI22_X1 port map( A1 => n10407, A2 => n10441, B1 => n10405, B2 => 
                           n7840, ZN => n2114);
   U9555 : OAI22_X1 port map( A1 => n10407, A2 => n10444, B1 => n10405, B2 => 
                           n7839, ZN => n2115);
   U9556 : OAI22_X1 port map( A1 => n10407, A2 => n10447, B1 => n10405, B2 => 
                           n7838, ZN => n2116);
   U9557 : OAI22_X1 port map( A1 => n10407, A2 => n10450, B1 => n10405, B2 => 
                           n7837, ZN => n2117);
   U9558 : OAI22_X1 port map( A1 => n10408, A2 => n10453, B1 => n10405, B2 => 
                           n7836, ZN => n2118);
   U9559 : OAI22_X1 port map( A1 => n10408, A2 => n10456, B1 => n10405, B2 => 
                           n7835, ZN => n2119);
   U9560 : OAI22_X1 port map( A1 => n10408, A2 => n10459, B1 => n8781, B2 => 
                           n7834, ZN => n2120);
   U9561 : OAI22_X1 port map( A1 => n10408, A2 => n10462, B1 => n8781, B2 => 
                           n7833, ZN => n2121);
   U9562 : OAI22_X1 port map( A1 => n10408, A2 => n10465, B1 => n8781, B2 => 
                           n7832, ZN => n2122);
   U9563 : OAI22_X1 port map( A1 => n10409, A2 => n10468, B1 => n10405, B2 => 
                           n7831, ZN => n2123);
   U9564 : OAI22_X1 port map( A1 => n10409, A2 => n10471, B1 => n10405, B2 => 
                           n7830, ZN => n2124);
   U9565 : OAI22_X1 port map( A1 => n10409, A2 => n10474, B1 => n10405, B2 => 
                           n7829, ZN => n2125);
   U9566 : OAI22_X1 port map( A1 => n10409, A2 => n10477, B1 => n10405, B2 => 
                           n7828, ZN => n2126);
   U9567 : OAI22_X1 port map( A1 => n10409, A2 => n10480, B1 => n10405, B2 => 
                           n7827, ZN => n2127);
   U9568 : OAI22_X1 port map( A1 => n10410, A2 => n10483, B1 => n10405, B2 => 
                           n7826, ZN => n2128);
   U9569 : OAI22_X1 port map( A1 => n10410, A2 => n10486, B1 => n10405, B2 => 
                           n7825, ZN => n2129);
   U9570 : OAI22_X1 port map( A1 => n10410, A2 => n10489, B1 => n10405, B2 => 
                           n7824, ZN => n2130);
   U9571 : OAI22_X1 port map( A1 => n10410, A2 => n10492, B1 => n10405, B2 => 
                           n7823, ZN => n2131);
   U9572 : OAI22_X1 port map( A1 => n10415, A2 => n10423, B1 => n10414, B2 => 
                           n7814, ZN => n2140);
   U9573 : OAI22_X1 port map( A1 => n10415, A2 => n10426, B1 => n10414, B2 => 
                           n7813, ZN => n2141);
   U9574 : OAI22_X1 port map( A1 => n10415, A2 => n10429, B1 => n10414, B2 => 
                           n7812, ZN => n2142);
   U9575 : OAI22_X1 port map( A1 => n10415, A2 => n10432, B1 => n10414, B2 => 
                           n7811, ZN => n2143);
   U9576 : OAI22_X1 port map( A1 => n10415, A2 => n10435, B1 => n10414, B2 => 
                           n7810, ZN => n2144);
   U9577 : OAI22_X1 port map( A1 => n10416, A2 => n10438, B1 => n10414, B2 => 
                           n7809, ZN => n2145);
   U9578 : OAI22_X1 port map( A1 => n10416, A2 => n10441, B1 => n10414, B2 => 
                           n7808, ZN => n2146);
   U9579 : OAI22_X1 port map( A1 => n10416, A2 => n10444, B1 => n10414, B2 => 
                           n7807, ZN => n2147);
   U9580 : OAI22_X1 port map( A1 => n10416, A2 => n10447, B1 => n10414, B2 => 
                           n7806, ZN => n2148);
   U9581 : OAI22_X1 port map( A1 => n10416, A2 => n10450, B1 => n10414, B2 => 
                           n7805, ZN => n2149);
   U9582 : OAI22_X1 port map( A1 => n10417, A2 => n10453, B1 => n10414, B2 => 
                           n7804, ZN => n2150);
   U9583 : OAI22_X1 port map( A1 => n10417, A2 => n10456, B1 => n10414, B2 => 
                           n7803, ZN => n2151);
   U9584 : OAI22_X1 port map( A1 => n10417, A2 => n10459, B1 => n8779, B2 => 
                           n7802, ZN => n2152);
   U9585 : OAI22_X1 port map( A1 => n10417, A2 => n10462, B1 => n8779, B2 => 
                           n7801, ZN => n2153);
   U9586 : OAI22_X1 port map( A1 => n10417, A2 => n10465, B1 => n8779, B2 => 
                           n7800, ZN => n2154);
   U9587 : OAI22_X1 port map( A1 => n10418, A2 => n10468, B1 => n10414, B2 => 
                           n7799, ZN => n2155);
   U9588 : OAI22_X1 port map( A1 => n10418, A2 => n10471, B1 => n10414, B2 => 
                           n7798, ZN => n2156);
   U9589 : OAI22_X1 port map( A1 => n10418, A2 => n10474, B1 => n10414, B2 => 
                           n7797, ZN => n2157);
   U9590 : OAI22_X1 port map( A1 => n10418, A2 => n10477, B1 => n10414, B2 => 
                           n7796, ZN => n2158);
   U9591 : OAI22_X1 port map( A1 => n10418, A2 => n10480, B1 => n10414, B2 => 
                           n7795, ZN => n2159);
   U9592 : OAI22_X1 port map( A1 => n10419, A2 => n10483, B1 => n10414, B2 => 
                           n7794, ZN => n2160);
   U9593 : OAI22_X1 port map( A1 => n10419, A2 => n10486, B1 => n10414, B2 => 
                           n7793, ZN => n2161);
   U9594 : OAI22_X1 port map( A1 => n10419, A2 => n10489, B1 => n10414, B2 => 
                           n7792, ZN => n2162);
   U9595 : OAI22_X1 port map( A1 => n10419, A2 => n10492, B1 => n10414, B2 => 
                           n7791, ZN => n2163);
   U9596 : OAI22_X1 port map( A1 => n10517, A2 => n10423, B1 => n10516, B2 => 
                           n7782, ZN => n2172);
   U9597 : OAI22_X1 port map( A1 => n10517, A2 => n10426, B1 => n10516, B2 => 
                           n7781, ZN => n2173);
   U9598 : OAI22_X1 port map( A1 => n10517, A2 => n10429, B1 => n10516, B2 => 
                           n7780, ZN => n2174);
   U9599 : OAI22_X1 port map( A1 => n10517, A2 => n10432, B1 => n10516, B2 => 
                           n7779, ZN => n2175);
   U9600 : OAI22_X1 port map( A1 => n10517, A2 => n10435, B1 => n10516, B2 => 
                           n7778, ZN => n2176);
   U9601 : OAI22_X1 port map( A1 => n10518, A2 => n10438, B1 => n10516, B2 => 
                           n7777, ZN => n2177);
   U9602 : OAI22_X1 port map( A1 => n10518, A2 => n10441, B1 => n10516, B2 => 
                           n7776, ZN => n2178);
   U9603 : OAI22_X1 port map( A1 => n10518, A2 => n10444, B1 => n10516, B2 => 
                           n7775, ZN => n2179);
   U9604 : OAI22_X1 port map( A1 => n10518, A2 => n10447, B1 => n10516, B2 => 
                           n7774, ZN => n2180);
   U9605 : OAI22_X1 port map( A1 => n10518, A2 => n10450, B1 => n10516, B2 => 
                           n7773, ZN => n2181);
   U9606 : OAI22_X1 port map( A1 => n10519, A2 => n10453, B1 => n10516, B2 => 
                           n7772, ZN => n2182);
   U9607 : OAI22_X1 port map( A1 => n10519, A2 => n10456, B1 => n10516, B2 => 
                           n7771, ZN => n2183);
   U9608 : OAI22_X1 port map( A1 => n10519, A2 => n10459, B1 => n8745, B2 => 
                           n7770, ZN => n2184);
   U9609 : OAI22_X1 port map( A1 => n10519, A2 => n10462, B1 => n8745, B2 => 
                           n7769, ZN => n2185);
   U9610 : OAI22_X1 port map( A1 => n10519, A2 => n10465, B1 => n8745, B2 => 
                           n7768, ZN => n2186);
   U9611 : OAI22_X1 port map( A1 => n10520, A2 => n10468, B1 => n10516, B2 => 
                           n7767, ZN => n2187);
   U9612 : OAI22_X1 port map( A1 => n10520, A2 => n10471, B1 => n10516, B2 => 
                           n7766, ZN => n2188);
   U9613 : OAI22_X1 port map( A1 => n10520, A2 => n10474, B1 => n10516, B2 => 
                           n7765, ZN => n2189);
   U9614 : OAI22_X1 port map( A1 => n10520, A2 => n10477, B1 => n10516, B2 => 
                           n7764, ZN => n2190);
   U9615 : OAI22_X1 port map( A1 => n10520, A2 => n10480, B1 => n10516, B2 => 
                           n7763, ZN => n2191);
   U9616 : OAI22_X1 port map( A1 => n10521, A2 => n10483, B1 => n10516, B2 => 
                           n7762, ZN => n2192);
   U9617 : OAI22_X1 port map( A1 => n10521, A2 => n10486, B1 => n10516, B2 => 
                           n7761, ZN => n2193);
   U9618 : OAI22_X1 port map( A1 => n10521, A2 => n10489, B1 => n10516, B2 => 
                           n7760, ZN => n2194);
   U9619 : OAI22_X1 port map( A1 => n10521, A2 => n10492, B1 => n10516, B2 => 
                           n7759, ZN => n2195);
   U9620 : OAI22_X1 port map( A1 => n6712, A2 => n10142, B1 => n10143, B2 => 
                           n10428, ZN => n1181);
   U9621 : OAI22_X1 port map( A1 => n6711, A2 => n8821, B1 => n10143, B2 => 
                           n10431, ZN => n1182);
   U9622 : OAI22_X1 port map( A1 => n6710, A2 => n10142, B1 => n10143, B2 => 
                           n10434, ZN => n1183);
   U9623 : OAI22_X1 port map( A1 => n6709, A2 => n8821, B1 => n10144, B2 => 
                           n10437, ZN => n1184);
   U9624 : OAI22_X1 port map( A1 => n6708, A2 => n10142, B1 => n10144, B2 => 
                           n10440, ZN => n1185);
   U9625 : OAI22_X1 port map( A1 => n6707, A2 => n8821, B1 => n10144, B2 => 
                           n10443, ZN => n1186);
   U9626 : OAI22_X1 port map( A1 => n6706, A2 => n10142, B1 => n10144, B2 => 
                           n10446, ZN => n1187);
   U9627 : OAI22_X1 port map( A1 => n6705, A2 => n8821, B1 => n10145, B2 => 
                           n10449, ZN => n1188);
   U9628 : OAI22_X1 port map( A1 => n6704, A2 => n10142, B1 => n10145, B2 => 
                           n10452, ZN => n1189);
   U9629 : OAI22_X1 port map( A1 => n6703, A2 => n10142, B1 => n10145, B2 => 
                           n10455, ZN => n1190);
   U9630 : OAI22_X1 port map( A1 => n6702, A2 => n10142, B1 => n10145, B2 => 
                           n10458, ZN => n1191);
   U9631 : OAI22_X1 port map( A1 => n6701, A2 => n10142, B1 => n10146, B2 => 
                           n10461, ZN => n1192);
   U9632 : OAI22_X1 port map( A1 => n6700, A2 => n10142, B1 => n10146, B2 => 
                           n10464, ZN => n1193);
   U9633 : OAI22_X1 port map( A1 => n6699, A2 => n10142, B1 => n10146, B2 => 
                           n10467, ZN => n1194);
   U9634 : OAI22_X1 port map( A1 => n6698, A2 => n10142, B1 => n10146, B2 => 
                           n10470, ZN => n1195);
   U9635 : OAI22_X1 port map( A1 => n6697, A2 => n10142, B1 => n10147, B2 => 
                           n10473, ZN => n1196);
   U9636 : OAI22_X1 port map( A1 => n6696, A2 => n10142, B1 => n10147, B2 => 
                           n10476, ZN => n1197);
   U9637 : OAI22_X1 port map( A1 => n6695, A2 => n10142, B1 => n10147, B2 => 
                           n10479, ZN => n1198);
   U9638 : OAI22_X1 port map( A1 => n6694, A2 => n10142, B1 => n10147, B2 => 
                           n10482, ZN => n1199);
   U9639 : OAI22_X1 port map( A1 => n6693, A2 => n8821, B1 => n10148, B2 => 
                           n10485, ZN => n1200);
   U9640 : OAI22_X1 port map( A1 => n6692, A2 => n10142, B1 => n10148, B2 => 
                           n10488, ZN => n1201);
   U9641 : OAI22_X1 port map( A1 => n6691, A2 => n8821, B1 => n10148, B2 => 
                           n10491, ZN => n1202);
   U9642 : OAI22_X1 port map( A1 => n6690, A2 => n10142, B1 => n10148, B2 => 
                           n10494, ZN => n1203);
   U9643 : OAI22_X1 port map( A1 => n6689, A2 => n8821, B1 => n10149, B2 => 
                           n10497, ZN => n1204);
   U9644 : OAI22_X1 port map( A1 => n6688, A2 => n10142, B1 => n10149, B2 => 
                           n10500, ZN => n1205);
   U9645 : OAI22_X1 port map( A1 => n6687, A2 => n8821, B1 => n10149, B2 => 
                           n10503, ZN => n1206);
   U9646 : OAI22_X1 port map( A1 => n6686, A2 => n10142, B1 => n10149, B2 => 
                           n10506, ZN => n1207);
   U9647 : OAI22_X1 port map( A1 => n6685, A2 => n8821, B1 => n10150, B2 => 
                           n10509, ZN => n1208);
   U9648 : OAI22_X1 port map( A1 => n6684, A2 => n10142, B1 => n10150, B2 => 
                           n10512, ZN => n1209);
   U9649 : OAI22_X1 port map( A1 => n6683, A2 => n8821, B1 => n10150, B2 => 
                           n10515, ZN => n1210);
   U9650 : OAI22_X1 port map( A1 => n6682, A2 => n10142, B1 => n10150, B2 => 
                           n10527, ZN => n1211);
   U9651 : OAI21_X1 port map( B1 => n9132, B2 => n9133, A => n10134, ZN => 
                           n9131);
   U9652 : OAI221_X1 port map( B1 => n8562, B2 => n10076, C1 => n8306, C2 => 
                           n10063, A => n9135, ZN => n9132);
   U9653 : OAI221_X1 port map( B1 => n8690, B2 => n10128, C1 => n8434, C2 => 
                           n10115, A => n9134, ZN => n9133);
   U9654 : AOI22_X1 port map( A1 => n10050, A2 => n9726, B1 => n10037, B2 => 
                           n9870, ZN => n9135);
   U9655 : OAI21_X1 port map( B1 => n9112, B2 => n9113, A => n10134, ZN => 
                           n9111);
   U9656 : OAI221_X1 port map( B1 => n8561, B2 => n10076, C1 => n8305, C2 => 
                           n10063, A => n9115, ZN => n9112);
   U9657 : OAI221_X1 port map( B1 => n8689, B2 => n10128, C1 => n8433, C2 => 
                           n10115, A => n9114, ZN => n9113);
   U9658 : AOI22_X1 port map( A1 => n10050, A2 => n9727, B1 => n10037, B2 => 
                           n9871, ZN => n9115);
   U9659 : OAI21_X1 port map( B1 => n9092, B2 => n9093, A => n10134, ZN => 
                           n9091);
   U9660 : OAI221_X1 port map( B1 => n8560, B2 => n10076, C1 => n8304, C2 => 
                           n10063, A => n9095, ZN => n9092);
   U9661 : OAI221_X1 port map( B1 => n8688, B2 => n10128, C1 => n8432, C2 => 
                           n10115, A => n9094, ZN => n9093);
   U9662 : AOI22_X1 port map( A1 => n10050, A2 => n9728, B1 => n10037, B2 => 
                           n9872, ZN => n9095);
   U9663 : OAI21_X1 port map( B1 => n9072, B2 => n9073, A => n10134, ZN => 
                           n9071);
   U9664 : OAI221_X1 port map( B1 => n8559, B2 => n10077, C1 => n8303, C2 => 
                           n10064, A => n9075, ZN => n9072);
   U9665 : OAI221_X1 port map( B1 => n8687, B2 => n10129, C1 => n8431, C2 => 
                           n10116, A => n9074, ZN => n9073);
   U9666 : AOI22_X1 port map( A1 => n10051, A2 => n9729, B1 => n10038, B2 => 
                           n9873, ZN => n9075);
   U9667 : OAI21_X1 port map( B1 => n9052, B2 => n9053, A => n10134, ZN => 
                           n9051);
   U9668 : OAI221_X1 port map( B1 => n8558, B2 => n10077, C1 => n8302, C2 => 
                           n10064, A => n9055, ZN => n9052);
   U9669 : OAI221_X1 port map( B1 => n8686, B2 => n10129, C1 => n8430, C2 => 
                           n10116, A => n9054, ZN => n9053);
   U9670 : AOI22_X1 port map( A1 => n10051, A2 => n9730, B1 => n10038, B2 => 
                           n9874, ZN => n9055);
   U9671 : OAI21_X1 port map( B1 => n9032, B2 => n9033, A => n10134, ZN => 
                           n9031);
   U9672 : OAI221_X1 port map( B1 => n8557, B2 => n10077, C1 => n8301, C2 => 
                           n10064, A => n9035, ZN => n9032);
   U9673 : OAI221_X1 port map( B1 => n8685, B2 => n10129, C1 => n8429, C2 => 
                           n10116, A => n9034, ZN => n9033);
   U9674 : AOI22_X1 port map( A1 => n10051, A2 => n9731, B1 => n10038, B2 => 
                           n9875, ZN => n9035);
   U9675 : OAI22_X1 port map( A1 => n10289, A2 => n10424, B1 => n10288, B2 => 
                           n8228, ZN => n1692);
   U9676 : OAI22_X1 port map( A1 => n10289, A2 => n10427, B1 => n10288, B2 => 
                           n8227, ZN => n1693);
   U9677 : OAI22_X1 port map( A1 => n10289, A2 => n10430, B1 => n10288, B2 => 
                           n8226, ZN => n1694);
   U9678 : OAI22_X1 port map( A1 => n10289, A2 => n10433, B1 => n10288, B2 => 
                           n8225, ZN => n1695);
   U9679 : OAI22_X1 port map( A1 => n10289, A2 => n10436, B1 => n10288, B2 => 
                           n8224, ZN => n1696);
   U9680 : OAI22_X1 port map( A1 => n10290, A2 => n10439, B1 => n10288, B2 => 
                           n8223, ZN => n1697);
   U9681 : OAI22_X1 port map( A1 => n10290, A2 => n10442, B1 => n10288, B2 => 
                           n8222, ZN => n1698);
   U9682 : OAI22_X1 port map( A1 => n10290, A2 => n10445, B1 => n10288, B2 => 
                           n8221, ZN => n1699);
   U9683 : OAI22_X1 port map( A1 => n10290, A2 => n10448, B1 => n10288, B2 => 
                           n8220, ZN => n1700);
   U9684 : OAI22_X1 port map( A1 => n10290, A2 => n10451, B1 => n10288, B2 => 
                           n8219, ZN => n1701);
   U9685 : OAI22_X1 port map( A1 => n10291, A2 => n10454, B1 => n10288, B2 => 
                           n8218, ZN => n1702);
   U9686 : OAI22_X1 port map( A1 => n10291, A2 => n10457, B1 => n10288, B2 => 
                           n8217, ZN => n1703);
   U9687 : OAI22_X1 port map( A1 => n10291, A2 => n10460, B1 => n8800, B2 => 
                           n8216, ZN => n1704);
   U9688 : OAI22_X1 port map( A1 => n10291, A2 => n10463, B1 => n8800, B2 => 
                           n8215, ZN => n1705);
   U9689 : OAI22_X1 port map( A1 => n10291, A2 => n10466, B1 => n8800, B2 => 
                           n8214, ZN => n1706);
   U9690 : OAI22_X1 port map( A1 => n10292, A2 => n10469, B1 => n10288, B2 => 
                           n8213, ZN => n1707);
   U9691 : OAI22_X1 port map( A1 => n10292, A2 => n10472, B1 => n10288, B2 => 
                           n8212, ZN => n1708);
   U9692 : OAI22_X1 port map( A1 => n10292, A2 => n10475, B1 => n10288, B2 => 
                           n8211, ZN => n1709);
   U9693 : OAI22_X1 port map( A1 => n10292, A2 => n10478, B1 => n10288, B2 => 
                           n8210, ZN => n1710);
   U9694 : OAI22_X1 port map( A1 => n10292, A2 => n10481, B1 => n10288, B2 => 
                           n8209, ZN => n1711);
   U9695 : OAI22_X1 port map( A1 => n10293, A2 => n10484, B1 => n10288, B2 => 
                           n8208, ZN => n1712);
   U9696 : OAI22_X1 port map( A1 => n10293, A2 => n10487, B1 => n10288, B2 => 
                           n8207, ZN => n1713);
   U9697 : OAI22_X1 port map( A1 => n10293, A2 => n10490, B1 => n10288, B2 => 
                           n8206, ZN => n1714);
   U9698 : OAI22_X1 port map( A1 => n10293, A2 => n10493, B1 => n10288, B2 => 
                           n8205, ZN => n1715);
   U9699 : OAI22_X1 port map( A1 => n10298, A2 => n10424, B1 => n10297, B2 => 
                           n8204, ZN => n1724);
   U9700 : OAI22_X1 port map( A1 => n10298, A2 => n10427, B1 => n10297, B2 => 
                           n8203, ZN => n1725);
   U9701 : OAI22_X1 port map( A1 => n10298, A2 => n10430, B1 => n10297, B2 => 
                           n8202, ZN => n1726);
   U9702 : OAI22_X1 port map( A1 => n10298, A2 => n10433, B1 => n10297, B2 => 
                           n8201, ZN => n1727);
   U9703 : OAI22_X1 port map( A1 => n10298, A2 => n10436, B1 => n10297, B2 => 
                           n8200, ZN => n1728);
   U9704 : OAI22_X1 port map( A1 => n10299, A2 => n10439, B1 => n10297, B2 => 
                           n8199, ZN => n1729);
   U9705 : OAI22_X1 port map( A1 => n10299, A2 => n10442, B1 => n10297, B2 => 
                           n8198, ZN => n1730);
   U9706 : OAI22_X1 port map( A1 => n10299, A2 => n10445, B1 => n10297, B2 => 
                           n8197, ZN => n1731);
   U9707 : OAI22_X1 port map( A1 => n10299, A2 => n10448, B1 => n10297, B2 => 
                           n8196, ZN => n1732);
   U9708 : OAI22_X1 port map( A1 => n10299, A2 => n10451, B1 => n10297, B2 => 
                           n8195, ZN => n1733);
   U9709 : OAI22_X1 port map( A1 => n10300, A2 => n10454, B1 => n10297, B2 => 
                           n8194, ZN => n1734);
   U9710 : OAI22_X1 port map( A1 => n10300, A2 => n10457, B1 => n10297, B2 => 
                           n8193, ZN => n1735);
   U9711 : OAI22_X1 port map( A1 => n10300, A2 => n10460, B1 => n8799, B2 => 
                           n8192, ZN => n1736);
   U9712 : OAI22_X1 port map( A1 => n10300, A2 => n10463, B1 => n8799, B2 => 
                           n8191, ZN => n1737);
   U9713 : OAI22_X1 port map( A1 => n10300, A2 => n10466, B1 => n8799, B2 => 
                           n8190, ZN => n1738);
   U9714 : OAI22_X1 port map( A1 => n10301, A2 => n10469, B1 => n10297, B2 => 
                           n8189, ZN => n1739);
   U9715 : OAI22_X1 port map( A1 => n10301, A2 => n10472, B1 => n10297, B2 => 
                           n8188, ZN => n1740);
   U9716 : OAI22_X1 port map( A1 => n10301, A2 => n10475, B1 => n10297, B2 => 
                           n8187, ZN => n1741);
   U9717 : OAI22_X1 port map( A1 => n10301, A2 => n10478, B1 => n10297, B2 => 
                           n8186, ZN => n1742);
   U9718 : OAI22_X1 port map( A1 => n10301, A2 => n10481, B1 => n10297, B2 => 
                           n8185, ZN => n1743);
   U9719 : OAI22_X1 port map( A1 => n10302, A2 => n10484, B1 => n10297, B2 => 
                           n8184, ZN => n1744);
   U9720 : OAI22_X1 port map( A1 => n10302, A2 => n10487, B1 => n10297, B2 => 
                           n8183, ZN => n1745);
   U9721 : OAI22_X1 port map( A1 => n10302, A2 => n10490, B1 => n10297, B2 => 
                           n8182, ZN => n1746);
   U9722 : OAI22_X1 port map( A1 => n10302, A2 => n10493, B1 => n10297, B2 => 
                           n8181, ZN => n1747);
   U9723 : OAI22_X1 port map( A1 => n10307, A2 => n10424, B1 => n10306, B2 => 
                           n8180, ZN => n1756);
   U9724 : OAI22_X1 port map( A1 => n10307, A2 => n10427, B1 => n10306, B2 => 
                           n8179, ZN => n1757);
   U9725 : OAI22_X1 port map( A1 => n10307, A2 => n10430, B1 => n10306, B2 => 
                           n8178, ZN => n1758);
   U9726 : OAI22_X1 port map( A1 => n10307, A2 => n10433, B1 => n10306, B2 => 
                           n8177, ZN => n1759);
   U9727 : OAI22_X1 port map( A1 => n10307, A2 => n10436, B1 => n10306, B2 => 
                           n8176, ZN => n1760);
   U9728 : OAI22_X1 port map( A1 => n10308, A2 => n10439, B1 => n10306, B2 => 
                           n8175, ZN => n1761);
   U9729 : OAI22_X1 port map( A1 => n10308, A2 => n10442, B1 => n10306, B2 => 
                           n8174, ZN => n1762);
   U9730 : OAI22_X1 port map( A1 => n10308, A2 => n10445, B1 => n10306, B2 => 
                           n8173, ZN => n1763);
   U9731 : OAI22_X1 port map( A1 => n10308, A2 => n10448, B1 => n10306, B2 => 
                           n8172, ZN => n1764);
   U9732 : OAI22_X1 port map( A1 => n10308, A2 => n10451, B1 => n10306, B2 => 
                           n8171, ZN => n1765);
   U9733 : OAI22_X1 port map( A1 => n10309, A2 => n10454, B1 => n10306, B2 => 
                           n8170, ZN => n1766);
   U9734 : OAI22_X1 port map( A1 => n10309, A2 => n10457, B1 => n10306, B2 => 
                           n8169, ZN => n1767);
   U9735 : OAI22_X1 port map( A1 => n10309, A2 => n10460, B1 => n8798, B2 => 
                           n8168, ZN => n1768);
   U9736 : OAI22_X1 port map( A1 => n10309, A2 => n10463, B1 => n8798, B2 => 
                           n8167, ZN => n1769);
   U9737 : OAI22_X1 port map( A1 => n10309, A2 => n10466, B1 => n8798, B2 => 
                           n8166, ZN => n1770);
   U9738 : OAI22_X1 port map( A1 => n10310, A2 => n10469, B1 => n10306, B2 => 
                           n8165, ZN => n1771);
   U9739 : OAI22_X1 port map( A1 => n10310, A2 => n10472, B1 => n10306, B2 => 
                           n8164, ZN => n1772);
   U9740 : OAI22_X1 port map( A1 => n10310, A2 => n10475, B1 => n10306, B2 => 
                           n8163, ZN => n1773);
   U9741 : OAI22_X1 port map( A1 => n10310, A2 => n10478, B1 => n10306, B2 => 
                           n8162, ZN => n1774);
   U9742 : OAI22_X1 port map( A1 => n10310, A2 => n10481, B1 => n10306, B2 => 
                           n8161, ZN => n1775);
   U9743 : OAI22_X1 port map( A1 => n10311, A2 => n10484, B1 => n10306, B2 => 
                           n8160, ZN => n1776);
   U9744 : OAI22_X1 port map( A1 => n10311, A2 => n10487, B1 => n10306, B2 => 
                           n8159, ZN => n1777);
   U9745 : OAI22_X1 port map( A1 => n10311, A2 => n10490, B1 => n10306, B2 => 
                           n8158, ZN => n1778);
   U9746 : OAI22_X1 port map( A1 => n10311, A2 => n10493, B1 => n10306, B2 => 
                           n8157, ZN => n1779);
   U9747 : OAI22_X1 port map( A1 => n10316, A2 => n10424, B1 => n10315, B2 => 
                           n8156, ZN => n1788);
   U9748 : OAI22_X1 port map( A1 => n10316, A2 => n10427, B1 => n10315, B2 => 
                           n8155, ZN => n1789);
   U9749 : OAI22_X1 port map( A1 => n10316, A2 => n10430, B1 => n10315, B2 => 
                           n8154, ZN => n1790);
   U9750 : OAI22_X1 port map( A1 => n10316, A2 => n10433, B1 => n10315, B2 => 
                           n8153, ZN => n1791);
   U9751 : OAI22_X1 port map( A1 => n10316, A2 => n10436, B1 => n10315, B2 => 
                           n8152, ZN => n1792);
   U9752 : OAI22_X1 port map( A1 => n10317, A2 => n10439, B1 => n10315, B2 => 
                           n8151, ZN => n1793);
   U9753 : OAI22_X1 port map( A1 => n10317, A2 => n10442, B1 => n10315, B2 => 
                           n8150, ZN => n1794);
   U9754 : OAI22_X1 port map( A1 => n10317, A2 => n10445, B1 => n10315, B2 => 
                           n8149, ZN => n1795);
   U9755 : OAI22_X1 port map( A1 => n10317, A2 => n10448, B1 => n10315, B2 => 
                           n8148, ZN => n1796);
   U9756 : OAI22_X1 port map( A1 => n10317, A2 => n10451, B1 => n10315, B2 => 
                           n8147, ZN => n1797);
   U9757 : OAI22_X1 port map( A1 => n10318, A2 => n10454, B1 => n10315, B2 => 
                           n8146, ZN => n1798);
   U9758 : OAI22_X1 port map( A1 => n10318, A2 => n10457, B1 => n10315, B2 => 
                           n8145, ZN => n1799);
   U9759 : OAI22_X1 port map( A1 => n10318, A2 => n10460, B1 => n8796, B2 => 
                           n8144, ZN => n1800);
   U9760 : OAI22_X1 port map( A1 => n10318, A2 => n10463, B1 => n8796, B2 => 
                           n8143, ZN => n1801);
   U9761 : OAI22_X1 port map( A1 => n10318, A2 => n10466, B1 => n8796, B2 => 
                           n8142, ZN => n1802);
   U9762 : OAI22_X1 port map( A1 => n10319, A2 => n10469, B1 => n10315, B2 => 
                           n8141, ZN => n1803);
   U9763 : OAI22_X1 port map( A1 => n10319, A2 => n10472, B1 => n10315, B2 => 
                           n8140, ZN => n1804);
   U9764 : OAI22_X1 port map( A1 => n10319, A2 => n10475, B1 => n10315, B2 => 
                           n8139, ZN => n1805);
   U9765 : OAI22_X1 port map( A1 => n10319, A2 => n10478, B1 => n10315, B2 => 
                           n8138, ZN => n1806);
   U9766 : OAI22_X1 port map( A1 => n10319, A2 => n10481, B1 => n10315, B2 => 
                           n8137, ZN => n1807);
   U9767 : OAI22_X1 port map( A1 => n10320, A2 => n10484, B1 => n10315, B2 => 
                           n8136, ZN => n1808);
   U9768 : OAI22_X1 port map( A1 => n10320, A2 => n10487, B1 => n10315, B2 => 
                           n8135, ZN => n1809);
   U9769 : OAI22_X1 port map( A1 => n10320, A2 => n10490, B1 => n10315, B2 => 
                           n8134, ZN => n1810);
   U9770 : OAI22_X1 port map( A1 => n10320, A2 => n10493, B1 => n10315, B2 => 
                           n8133, ZN => n1811);
   U9771 : OAI22_X1 port map( A1 => n10325, A2 => n10423, B1 => n10324, B2 => 
                           n8132, ZN => n1820);
   U9772 : OAI22_X1 port map( A1 => n10325, A2 => n10426, B1 => n10324, B2 => 
                           n8131, ZN => n1821);
   U9773 : OAI22_X1 port map( A1 => n10325, A2 => n10429, B1 => n10324, B2 => 
                           n8130, ZN => n1822);
   U9774 : OAI22_X1 port map( A1 => n10325, A2 => n10432, B1 => n10324, B2 => 
                           n8129, ZN => n1823);
   U9775 : OAI22_X1 port map( A1 => n10325, A2 => n10435, B1 => n10324, B2 => 
                           n8128, ZN => n1824);
   U9776 : OAI22_X1 port map( A1 => n10326, A2 => n10438, B1 => n10324, B2 => 
                           n8127, ZN => n1825);
   U9777 : OAI22_X1 port map( A1 => n10326, A2 => n10441, B1 => n10324, B2 => 
                           n8126, ZN => n1826);
   U9778 : OAI22_X1 port map( A1 => n10326, A2 => n10444, B1 => n10324, B2 => 
                           n8125, ZN => n1827);
   U9779 : OAI22_X1 port map( A1 => n10326, A2 => n10447, B1 => n10324, B2 => 
                           n8124, ZN => n1828);
   U9780 : OAI22_X1 port map( A1 => n10326, A2 => n10450, B1 => n10324, B2 => 
                           n8123, ZN => n1829);
   U9781 : OAI22_X1 port map( A1 => n10327, A2 => n10453, B1 => n10324, B2 => 
                           n8122, ZN => n1830);
   U9782 : OAI22_X1 port map( A1 => n10327, A2 => n10456, B1 => n10324, B2 => 
                           n8121, ZN => n1831);
   U9783 : OAI22_X1 port map( A1 => n10327, A2 => n10459, B1 => n8795, B2 => 
                           n8120, ZN => n1832);
   U9784 : OAI22_X1 port map( A1 => n10327, A2 => n10462, B1 => n8795, B2 => 
                           n8119, ZN => n1833);
   U9785 : OAI22_X1 port map( A1 => n10327, A2 => n10465, B1 => n8795, B2 => 
                           n8118, ZN => n1834);
   U9786 : OAI22_X1 port map( A1 => n10328, A2 => n10468, B1 => n10324, B2 => 
                           n8117, ZN => n1835);
   U9787 : OAI22_X1 port map( A1 => n10328, A2 => n10471, B1 => n10324, B2 => 
                           n8116, ZN => n1836);
   U9788 : OAI22_X1 port map( A1 => n10328, A2 => n10474, B1 => n10324, B2 => 
                           n8115, ZN => n1837);
   U9789 : OAI22_X1 port map( A1 => n10328, A2 => n10477, B1 => n10324, B2 => 
                           n8114, ZN => n1838);
   U9790 : OAI22_X1 port map( A1 => n10328, A2 => n10480, B1 => n10324, B2 => 
                           n8113, ZN => n1839);
   U9791 : OAI22_X1 port map( A1 => n10329, A2 => n10483, B1 => n10324, B2 => 
                           n8112, ZN => n1840);
   U9792 : OAI22_X1 port map( A1 => n10329, A2 => n10486, B1 => n10324, B2 => 
                           n8111, ZN => n1841);
   U9793 : OAI22_X1 port map( A1 => n10329, A2 => n10489, B1 => n10324, B2 => 
                           n8110, ZN => n1842);
   U9794 : OAI22_X1 port map( A1 => n10329, A2 => n10492, B1 => n10324, B2 => 
                           n8109, ZN => n1843);
   U9795 : OAI22_X1 port map( A1 => n10334, A2 => n10423, B1 => n10333, B2 => 
                           n8102, ZN => n1852);
   U9796 : OAI22_X1 port map( A1 => n10334, A2 => n10426, B1 => n10333, B2 => 
                           n8101, ZN => n1853);
   U9797 : OAI22_X1 port map( A1 => n10334, A2 => n10429, B1 => n10333, B2 => 
                           n8100, ZN => n1854);
   U9798 : OAI22_X1 port map( A1 => n10334, A2 => n10432, B1 => n10333, B2 => 
                           n8099, ZN => n1855);
   U9799 : OAI22_X1 port map( A1 => n10334, A2 => n10435, B1 => n10333, B2 => 
                           n8098, ZN => n1856);
   U9800 : OAI22_X1 port map( A1 => n10335, A2 => n10438, B1 => n10333, B2 => 
                           n8097, ZN => n1857);
   U9801 : OAI22_X1 port map( A1 => n10335, A2 => n10441, B1 => n10333, B2 => 
                           n8096, ZN => n1858);
   U9802 : OAI22_X1 port map( A1 => n10335, A2 => n10444, B1 => n10333, B2 => 
                           n8095, ZN => n1859);
   U9803 : OAI22_X1 port map( A1 => n10335, A2 => n10447, B1 => n10333, B2 => 
                           n8094, ZN => n1860);
   U9804 : OAI22_X1 port map( A1 => n10335, A2 => n10450, B1 => n10333, B2 => 
                           n8093, ZN => n1861);
   U9805 : OAI22_X1 port map( A1 => n10336, A2 => n10453, B1 => n10333, B2 => 
                           n8092, ZN => n1862);
   U9806 : OAI22_X1 port map( A1 => n10336, A2 => n10456, B1 => n10333, B2 => 
                           n8091, ZN => n1863);
   U9807 : OAI22_X1 port map( A1 => n10336, A2 => n10459, B1 => n8794, B2 => 
                           n8090, ZN => n1864);
   U9808 : OAI22_X1 port map( A1 => n10336, A2 => n10462, B1 => n8794, B2 => 
                           n8089, ZN => n1865);
   U9809 : OAI22_X1 port map( A1 => n10336, A2 => n10465, B1 => n8794, B2 => 
                           n8088, ZN => n1866);
   U9810 : OAI22_X1 port map( A1 => n10337, A2 => n10468, B1 => n10333, B2 => 
                           n8087, ZN => n1867);
   U9811 : OAI22_X1 port map( A1 => n10337, A2 => n10471, B1 => n10333, B2 => 
                           n8086, ZN => n1868);
   U9812 : OAI22_X1 port map( A1 => n10337, A2 => n10474, B1 => n10333, B2 => 
                           n8085, ZN => n1869);
   U9813 : OAI22_X1 port map( A1 => n10337, A2 => n10477, B1 => n10333, B2 => 
                           n8084, ZN => n1870);
   U9814 : OAI22_X1 port map( A1 => n10337, A2 => n10480, B1 => n10333, B2 => 
                           n8083, ZN => n1871);
   U9815 : OAI22_X1 port map( A1 => n10338, A2 => n10483, B1 => n10333, B2 => 
                           n8082, ZN => n1872);
   U9816 : OAI22_X1 port map( A1 => n10338, A2 => n10486, B1 => n10333, B2 => 
                           n8081, ZN => n1873);
   U9817 : OAI22_X1 port map( A1 => n10338, A2 => n10489, B1 => n10333, B2 => 
                           n8080, ZN => n1874);
   U9818 : OAI22_X1 port map( A1 => n10338, A2 => n10492, B1 => n10333, B2 => 
                           n8079, ZN => n1875);
   U9819 : OAI22_X1 port map( A1 => n10343, A2 => n10423, B1 => n10342, B2 => 
                           n8070, ZN => n1884);
   U9820 : OAI22_X1 port map( A1 => n10343, A2 => n10426, B1 => n10342, B2 => 
                           n8069, ZN => n1885);
   U9821 : OAI22_X1 port map( A1 => n10343, A2 => n10429, B1 => n10342, B2 => 
                           n8068, ZN => n1886);
   U9822 : OAI22_X1 port map( A1 => n10343, A2 => n10432, B1 => n10342, B2 => 
                           n8067, ZN => n1887);
   U9823 : OAI22_X1 port map( A1 => n10343, A2 => n10435, B1 => n10342, B2 => 
                           n8066, ZN => n1888);
   U9824 : OAI22_X1 port map( A1 => n10344, A2 => n10438, B1 => n10342, B2 => 
                           n8065, ZN => n1889);
   U9825 : OAI22_X1 port map( A1 => n10344, A2 => n10441, B1 => n10342, B2 => 
                           n8064, ZN => n1890);
   U9826 : OAI22_X1 port map( A1 => n10344, A2 => n10444, B1 => n10342, B2 => 
                           n8063, ZN => n1891);
   U9827 : OAI22_X1 port map( A1 => n10344, A2 => n10447, B1 => n10342, B2 => 
                           n8062, ZN => n1892);
   U9828 : OAI22_X1 port map( A1 => n10344, A2 => n10450, B1 => n10342, B2 => 
                           n8061, ZN => n1893);
   U9829 : OAI22_X1 port map( A1 => n10345, A2 => n10453, B1 => n10342, B2 => 
                           n8060, ZN => n1894);
   U9830 : OAI22_X1 port map( A1 => n10345, A2 => n10456, B1 => n10342, B2 => 
                           n8059, ZN => n1895);
   U9831 : OAI22_X1 port map( A1 => n10345, A2 => n10459, B1 => n8793, B2 => 
                           n8058, ZN => n1896);
   U9832 : OAI22_X1 port map( A1 => n10345, A2 => n10462, B1 => n8793, B2 => 
                           n8057, ZN => n1897);
   U9833 : OAI22_X1 port map( A1 => n10345, A2 => n10465, B1 => n8793, B2 => 
                           n8056, ZN => n1898);
   U9834 : OAI22_X1 port map( A1 => n10346, A2 => n10468, B1 => n10342, B2 => 
                           n8055, ZN => n1899);
   U9835 : OAI22_X1 port map( A1 => n10346, A2 => n10471, B1 => n10342, B2 => 
                           n8054, ZN => n1900);
   U9836 : OAI22_X1 port map( A1 => n10346, A2 => n10474, B1 => n10342, B2 => 
                           n8053, ZN => n1901);
   U9837 : OAI22_X1 port map( A1 => n10346, A2 => n10477, B1 => n10342, B2 => 
                           n8052, ZN => n1902);
   U9838 : OAI22_X1 port map( A1 => n10346, A2 => n10480, B1 => n10342, B2 => 
                           n8051, ZN => n1903);
   U9839 : OAI22_X1 port map( A1 => n10347, A2 => n10483, B1 => n10342, B2 => 
                           n8050, ZN => n1904);
   U9840 : OAI22_X1 port map( A1 => n10347, A2 => n10486, B1 => n10342, B2 => 
                           n8049, ZN => n1905);
   U9841 : OAI22_X1 port map( A1 => n10347, A2 => n10489, B1 => n10342, B2 => 
                           n8048, ZN => n1906);
   U9842 : OAI22_X1 port map( A1 => n10347, A2 => n10492, B1 => n10342, B2 => 
                           n8047, ZN => n1907);
   U9843 : OAI22_X1 port map( A1 => n10352, A2 => n10423, B1 => n10351, B2 => 
                           n8038, ZN => n1916);
   U9844 : OAI22_X1 port map( A1 => n10352, A2 => n10426, B1 => n10351, B2 => 
                           n8037, ZN => n1917);
   U9845 : OAI22_X1 port map( A1 => n10352, A2 => n10429, B1 => n10351, B2 => 
                           n8036, ZN => n1918);
   U9846 : OAI22_X1 port map( A1 => n10352, A2 => n10432, B1 => n10351, B2 => 
                           n8035, ZN => n1919);
   U9847 : OAI22_X1 port map( A1 => n10352, A2 => n10435, B1 => n10351, B2 => 
                           n8034, ZN => n1920);
   U9848 : OAI22_X1 port map( A1 => n10353, A2 => n10438, B1 => n10351, B2 => 
                           n8033, ZN => n1921);
   U9849 : OAI22_X1 port map( A1 => n10353, A2 => n10441, B1 => n10351, B2 => 
                           n8032, ZN => n1922);
   U9850 : OAI22_X1 port map( A1 => n10353, A2 => n10444, B1 => n10351, B2 => 
                           n8031, ZN => n1923);
   U9851 : OAI22_X1 port map( A1 => n10353, A2 => n10447, B1 => n10351, B2 => 
                           n8030, ZN => n1924);
   U9852 : OAI22_X1 port map( A1 => n10353, A2 => n10450, B1 => n10351, B2 => 
                           n8029, ZN => n1925);
   U9853 : OAI22_X1 port map( A1 => n10354, A2 => n10453, B1 => n10351, B2 => 
                           n8028, ZN => n1926);
   U9854 : OAI22_X1 port map( A1 => n10354, A2 => n10456, B1 => n10351, B2 => 
                           n8027, ZN => n1927);
   U9855 : OAI22_X1 port map( A1 => n10354, A2 => n10459, B1 => n8791, B2 => 
                           n8026, ZN => n1928);
   U9856 : OAI22_X1 port map( A1 => n10354, A2 => n10462, B1 => n8791, B2 => 
                           n8025, ZN => n1929);
   U9857 : OAI22_X1 port map( A1 => n10354, A2 => n10465, B1 => n8791, B2 => 
                           n8024, ZN => n1930);
   U9858 : OAI22_X1 port map( A1 => n10355, A2 => n10468, B1 => n10351, B2 => 
                           n8023, ZN => n1931);
   U9859 : OAI22_X1 port map( A1 => n10355, A2 => n10471, B1 => n10351, B2 => 
                           n8022, ZN => n1932);
   U9860 : OAI22_X1 port map( A1 => n10355, A2 => n10474, B1 => n10351, B2 => 
                           n8021, ZN => n1933);
   U9861 : OAI22_X1 port map( A1 => n10355, A2 => n10477, B1 => n10351, B2 => 
                           n8020, ZN => n1934);
   U9862 : OAI22_X1 port map( A1 => n10355, A2 => n10480, B1 => n10351, B2 => 
                           n8019, ZN => n1935);
   U9863 : OAI22_X1 port map( A1 => n10356, A2 => n10483, B1 => n10351, B2 => 
                           n8018, ZN => n1936);
   U9864 : OAI22_X1 port map( A1 => n10356, A2 => n10486, B1 => n10351, B2 => 
                           n8017, ZN => n1937);
   U9865 : OAI22_X1 port map( A1 => n10356, A2 => n10489, B1 => n10351, B2 => 
                           n8016, ZN => n1938);
   U9866 : OAI22_X1 port map( A1 => n10356, A2 => n10492, B1 => n10351, B2 => 
                           n8015, ZN => n1939);
   U9867 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n8784);
   U9868 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n7746, ZN => n8782);
   U9869 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n7745, ZN => n8780);
   U9870 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(2), ZN => n8872);
   U9871 : NOR3_X1 port map( A1 => n7747, A2 => ADD_RD1(4), A3 => n7748, ZN => 
                           n8866);
   U9872 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n7748, 
                           ZN => n8867);
   U9873 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => ADD_RD1(4), A3 => n7747, 
                           ZN => n8871);
   U9874 : INV_X1 port map( A => RESET, ZN => n7741);
   U9875 : NOR2_X1 port map( A1 => n7749, A2 => ADD_RD1(0), ZN => n8862);
   U9876 : NOR2_X1 port map( A1 => n7750, A2 => ADD_RD1(1), ZN => n8875);
   U9877 : NOR2_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(1), ZN => n8880);
   U9878 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n10529, ZN => n8769);
   U9879 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n10529, ZN => n8767);
   U9880 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n10529, ZN => n8766);
   U9881 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n10529, ZN => n8765);
   U9882 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n10529, ZN => n8764);
   U9883 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n10529, ZN => n8763);
   U9884 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n10529, ZN => n8762);
   U9885 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n10529, ZN => n8761);
   U9886 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n10529, ZN => n8760);
   U9887 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n10529, ZN => n8759);
   U9888 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n10529, ZN => n8758);
   U9889 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n10529, ZN => n8757);
   U9890 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n10528, ZN => n8756);
   U9891 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n10528, ZN => n8755);
   U9892 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n10528, ZN => n8754);
   U9893 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n10528, ZN => n8753);
   U9894 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n10528, ZN => n8752);
   U9895 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n10528, ZN => n8751);
   U9896 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n10528, ZN => n8750);
   U9897 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n10528, ZN => n8749);
   U9898 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n10528, ZN => n8748);
   U9899 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n10528, ZN => n8747);
   U9900 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n10528, ZN => n8746);
   U9901 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n10528, ZN => n8744);
   U9902 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n10530, ZN => n8776);
   U9903 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n10530, ZN => n8775);
   U9904 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n10530, ZN => n8774);
   U9905 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n10530, ZN => n8773);
   U9906 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n10530, ZN => n8772);
   U9907 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n10530, ZN => n8771);
   U9908 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n10530, ZN => n8770);
   U9909 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n10530, ZN => n8768);
   U9910 : INV_X1 port map( A => ADD_RD1(2), ZN => n7748);
   U9911 : INV_X1 port map( A => ADD_RD1(3), ZN => n7747);
   U9912 : AND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => ADD_WR(4), ZN => 
                           n8806);
   U9913 : AND3_X1 port map( A1 => ENABLE, A2 => n7742, A3 => WR, ZN => n8785);
   U9914 : INV_X1 port map( A => ADD_WR(4), ZN => n7742);
   U9915 : INV_X1 port map( A => ADD_WR(3), ZN => n7743);
   U9916 : INV_X1 port map( A => ADD_WR(2), ZN => n7744);
   U9917 : INV_X1 port map( A => ADD_WR(0), ZN => n7746);
   U9918 : INV_X1 port map( A => ADD_RD1(1), ZN => n7749);
   U9919 : INV_X1 port map( A => ADD_RD1(0), ZN => n7750);
   U9920 : INV_X1 port map( A => ADD_WR(1), ZN => n7745);
   U9921 : CLKBUF_X1 port map( A => n10030, Z => n10041);
   U9922 : CLKBUF_X1 port map( A => n10043, Z => n10054);
   U9923 : CLKBUF_X1 port map( A => n10056, Z => n10067);
   U9924 : CLKBUF_X1 port map( A => n10069, Z => n10080);
   U9925 : CLKBUF_X1 port map( A => n10082, Z => n10093);
   U9926 : CLKBUF_X1 port map( A => n10095, Z => n10106);
   U9927 : CLKBUF_X1 port map( A => n10108, Z => n10119);
   U9928 : CLKBUF_X1 port map( A => n10121, Z => n10132);
   U9929 : CLKBUF_X1 port map( A => n7741, Z => n10533);

end SYN_behavioural;
