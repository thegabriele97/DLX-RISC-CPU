
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_mux21_generic_NBIT16 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_mux21_generic_NBIT16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_47 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_47;

architecture SYN_arch1 of nd2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_46 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_46;

architecture SYN_arch1 of nd2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_45 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_45;

architecture SYN_arch1 of nd2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_44 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_44;

architecture SYN_arch1 of nd2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_43 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_43;

architecture SYN_arch1 of nd2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_42 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_42;

architecture SYN_arch1 of nd2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_41 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_41;

architecture SYN_arch1 of nd2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_40 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_40;

architecture SYN_arch1 of nd2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_39 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_39;

architecture SYN_arch1 of nd2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_38 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_38;

architecture SYN_arch1 of nd2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_37 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_37;

architecture SYN_arch1 of nd2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_36 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_36;

architecture SYN_arch1 of nd2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_35 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_35;

architecture SYN_arch1 of nd2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_34 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_34;

architecture SYN_arch1 of nd2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_33 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_33;

architecture SYN_arch1 of nd2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_32 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_32;

architecture SYN_arch1 of nd2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_31 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_31;

architecture SYN_arch1 of nd2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_30 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_30;

architecture SYN_arch1 of nd2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_29 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_29;

architecture SYN_arch1 of nd2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_28 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_28;

architecture SYN_arch1 of nd2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_27 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_27;

architecture SYN_arch1 of nd2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_26 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_26;

architecture SYN_arch1 of nd2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_25 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_25;

architecture SYN_arch1 of nd2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_24 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_24;

architecture SYN_arch1 of nd2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_23 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_23;

architecture SYN_arch1 of nd2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_22 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_22;

architecture SYN_arch1 of nd2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_21 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_21;

architecture SYN_arch1 of nd2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_20 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_20;

architecture SYN_arch1 of nd2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_19 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_19;

architecture SYN_arch1 of nd2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_18 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_18;

architecture SYN_arch1 of nd2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_17 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_17;

architecture SYN_arch1 of nd2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_16 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_16;

architecture SYN_arch1 of nd2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_15 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_15;

architecture SYN_arch1 of nd2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_14 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_14;

architecture SYN_arch1 of nd2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_13 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_13;

architecture SYN_arch1 of nd2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_12 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_12;

architecture SYN_arch1 of nd2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_11 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_11;

architecture SYN_arch1 of nd2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_10 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_10;

architecture SYN_arch1 of nd2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_9 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_9;

architecture SYN_arch1 of nd2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_8 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_8;

architecture SYN_arch1 of nd2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_7 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_7;

architecture SYN_arch1 of nd2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_6 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_6;

architecture SYN_arch1 of nd2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_5 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_5;

architecture SYN_arch1 of nd2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_4 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_4;

architecture SYN_arch1 of nd2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_3 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_3;

architecture SYN_arch1 of nd2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_2 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_2;

architecture SYN_arch1 of nd2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_1 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_1;

architecture SYN_arch1 of nd2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_15 is

   port( a : in std_logic;  y : out std_logic);

end iv_15;

architecture SYN_behavioural of iv_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_14 is

   port( a : in std_logic;  y : out std_logic);

end iv_14;

architecture SYN_behavioural of iv_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_13 is

   port( a : in std_logic;  y : out std_logic);

end iv_13;

architecture SYN_behavioural of iv_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_12 is

   port( a : in std_logic;  y : out std_logic);

end iv_12;

architecture SYN_behavioural of iv_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_11 is

   port( a : in std_logic;  y : out std_logic);

end iv_11;

architecture SYN_behavioural of iv_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_10 is

   port( a : in std_logic;  y : out std_logic);

end iv_10;

architecture SYN_behavioural of iv_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_9 is

   port( a : in std_logic;  y : out std_logic);

end iv_9;

architecture SYN_behavioural of iv_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_8 is

   port( a : in std_logic;  y : out std_logic);

end iv_8;

architecture SYN_behavioural of iv_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_7 is

   port( a : in std_logic;  y : out std_logic);

end iv_7;

architecture SYN_behavioural of iv_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_6 is

   port( a : in std_logic;  y : out std_logic);

end iv_6;

architecture SYN_behavioural of iv_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_5 is

   port( a : in std_logic;  y : out std_logic);

end iv_5;

architecture SYN_behavioural of iv_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_4 is

   port( a : in std_logic;  y : out std_logic);

end iv_4;

architecture SYN_behavioural of iv_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_3 is

   port( a : in std_logic;  y : out std_logic);

end iv_3;

architecture SYN_behavioural of iv_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_2 is

   port( a : in std_logic;  y : out std_logic);

end iv_2;

architecture SYN_behavioural of iv_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_1 is

   port( a : in std_logic;  y : out std_logic);

end iv_1;

architecture SYN_behavioural of iv_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_generic_NBIT16_2 is

   port( a, b : in std_logic_vector (15 downto 0);  y : out std_logic_vector 
         (15 downto 0));

end nd2_generic_NBIT16_2;

architecture SYN_structural of nd2_generic_NBIT16_2 is

   component nd2_17
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_18
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_19
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_20
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_21
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_22
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_23
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_24
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_25
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_26
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_27
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_28
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_29
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_30
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_31
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_32
      port( a, b : in std_logic;  y : out std_logic);
   end component;

begin
   
   ndi_0 : nd2_32 port map( a => a(0), b => b(0), y => y(0));
   ndi_1 : nd2_31 port map( a => a(1), b => b(1), y => y(1));
   ndi_2 : nd2_30 port map( a => a(2), b => b(2), y => y(2));
   ndi_3 : nd2_29 port map( a => a(3), b => b(3), y => y(3));
   ndi_4 : nd2_28 port map( a => a(4), b => b(4), y => y(4));
   ndi_5 : nd2_27 port map( a => a(5), b => b(5), y => y(5));
   ndi_6 : nd2_26 port map( a => a(6), b => b(6), y => y(6));
   ndi_7 : nd2_25 port map( a => a(7), b => b(7), y => y(7));
   ndi_8 : nd2_24 port map( a => a(8), b => b(8), y => y(8));
   ndi_9 : nd2_23 port map( a => a(9), b => b(9), y => y(9));
   ndi_10 : nd2_22 port map( a => a(10), b => b(10), y => y(10));
   ndi_11 : nd2_21 port map( a => a(11), b => b(11), y => y(11));
   ndi_12 : nd2_20 port map( a => a(12), b => b(12), y => y(12));
   ndi_13 : nd2_19 port map( a => a(13), b => b(13), y => y(13));
   ndi_14 : nd2_18 port map( a => a(14), b => b(14), y => y(14));
   ndi_15 : nd2_17 port map( a => a(15), b => b(15), y => y(15));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_generic_NBIT16_1 is

   port( a, b : in std_logic_vector (15 downto 0);  y : out std_logic_vector 
         (15 downto 0));

end nd2_generic_NBIT16_1;

architecture SYN_structural of nd2_generic_NBIT16_1 is

   component nd2_1
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_2
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_3
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_4
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_5
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_6
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_7
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_8
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_9
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_10
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_11
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_12
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_13
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_14
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_15
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_16
      port( a, b : in std_logic;  y : out std_logic);
   end component;

begin
   
   ndi_0 : nd2_16 port map( a => a(0), b => b(0), y => y(0));
   ndi_1 : nd2_15 port map( a => a(1), b => b(1), y => y(1));
   ndi_2 : nd2_14 port map( a => a(2), b => b(2), y => y(2));
   ndi_3 : nd2_13 port map( a => a(3), b => b(3), y => y(3));
   ndi_4 : nd2_12 port map( a => a(4), b => b(4), y => y(4));
   ndi_5 : nd2_11 port map( a => a(5), b => b(5), y => y(5));
   ndi_6 : nd2_10 port map( a => a(6), b => b(6), y => y(6));
   ndi_7 : nd2_9 port map( a => a(7), b => b(7), y => y(7));
   ndi_8 : nd2_8 port map( a => a(8), b => b(8), y => y(8));
   ndi_9 : nd2_7 port map( a => a(9), b => b(9), y => y(9));
   ndi_10 : nd2_6 port map( a => a(10), b => b(10), y => y(10));
   ndi_11 : nd2_5 port map( a => a(11), b => b(11), y => y(11));
   ndi_12 : nd2_4 port map( a => a(12), b => b(12), y => y(12));
   ndi_13 : nd2_3 port map( a => a(13), b => b(13), y => y(13));
   ndi_14 : nd2_2 port map( a => a(14), b => b(14), y => y(14));
   ndi_15 : nd2_1 port map( a => a(15), b => b(15), y => y(15));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_0 is

   port( a, b : in std_logic;  y : out std_logic);

end nd2_0;

architecture SYN_arch1 of nd2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => y);

end SYN_arch1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_0 is

   port( a : in std_logic;  y : out std_logic);

end iv_0;

architecture SYN_behavioural of iv_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => y);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity nd2_generic_NBIT16_0 is

   port( a, b : in std_logic_vector (15 downto 0);  y : out std_logic_vector 
         (15 downto 0));

end nd2_generic_NBIT16_0;

architecture SYN_structural of nd2_generic_NBIT16_0 is

   component nd2_33
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_34
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_35
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_36
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_37
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_38
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_39
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_40
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_41
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_42
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_43
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_44
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_45
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_46
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_47
      port( a, b : in std_logic;  y : out std_logic);
   end component;
   
   component nd2_0
      port( a, b : in std_logic;  y : out std_logic);
   end component;

begin
   
   ndi_0 : nd2_0 port map( a => a(0), b => b(0), y => y(0));
   ndi_1 : nd2_47 port map( a => a(1), b => b(1), y => y(1));
   ndi_2 : nd2_46 port map( a => a(2), b => b(2), y => y(2));
   ndi_3 : nd2_45 port map( a => a(3), b => b(3), y => y(3));
   ndi_4 : nd2_44 port map( a => a(4), b => b(4), y => y(4));
   ndi_5 : nd2_43 port map( a => a(5), b => b(5), y => y(5));
   ndi_6 : nd2_42 port map( a => a(6), b => b(6), y => y(6));
   ndi_7 : nd2_41 port map( a => a(7), b => b(7), y => y(7));
   ndi_8 : nd2_40 port map( a => a(8), b => b(8), y => y(8));
   ndi_9 : nd2_39 port map( a => a(9), b => b(9), y => y(9));
   ndi_10 : nd2_38 port map( a => a(10), b => b(10), y => y(10));
   ndi_11 : nd2_37 port map( a => a(11), b => b(11), y => y(11));
   ndi_12 : nd2_36 port map( a => a(12), b => b(12), y => y(12));
   ndi_13 : nd2_35 port map( a => a(13), b => b(13), y => y(13));
   ndi_14 : nd2_34 port map( a => a(14), b => b(14), y => y(14));
   ndi_15 : nd2_33 port map( a => a(15), b => b(15), y => y(15));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity iv_generic_NBIT16 is

   port( a : in std_logic_vector (15 downto 0);  y : out std_logic_vector (15 
         downto 0));

end iv_generic_NBIT16;

architecture SYN_structural of iv_generic_NBIT16 is

   component iv_1
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_2
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_3
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_4
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_5
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_6
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_7
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_8
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_9
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_10
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_11
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_12
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_13
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_14
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_15
      port( a : in std_logic;  y : out std_logic);
   end component;
   
   component iv_0
      port( a : in std_logic;  y : out std_logic);
   end component;

begin
   
   ivi_0 : iv_0 port map( a => a(0), y => y(0));
   ivi_1 : iv_15 port map( a => a(1), y => y(1));
   ivi_2 : iv_14 port map( a => a(2), y => y(2));
   ivi_3 : iv_13 port map( a => a(3), y => y(3));
   ivi_4 : iv_12 port map( a => a(4), y => y(4));
   ivi_5 : iv_11 port map( a => a(5), y => y(5));
   ivi_6 : iv_10 port map( a => a(6), y => y(6));
   ivi_7 : iv_9 port map( a => a(7), y => y(7));
   ivi_8 : iv_8 port map( a => a(8), y => y(8));
   ivi_9 : iv_7 port map( a => a(9), y => y(9));
   ivi_10 : iv_6 port map( a => a(10), y => y(10));
   ivi_11 : iv_5 port map( a => a(11), y => y(11));
   ivi_12 : iv_4 port map( a => a(12), y => y(12));
   ivi_13 : iv_3 port map( a => a(13), y => y(13));
   ivi_14 : iv_2 port map( a => a(14), y => y(14));
   ivi_15 : iv_1 port map( a => a(15), y => y(15));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_mux21_generic_NBIT16.all;

entity mux21_generic_NBIT16 is

   port( a, b : in std_logic_vector (15 downto 0);  s : in std_logic;  y : out 
         std_logic_vector (15 downto 0));

end mux21_generic_NBIT16;

architecture SYN_structural of mux21_generic_NBIT16 is

   component nd2_generic_NBIT16_1
      port( a, b : in std_logic_vector (15 downto 0);  y : out std_logic_vector
            (15 downto 0));
   end component;
   
   component nd2_generic_NBIT16_2
      port( a, b : in std_logic_vector (15 downto 0);  y : out std_logic_vector
            (15 downto 0));
   end component;
   
   component nd2_generic_NBIT16_0
      port( a, b : in std_logic_vector (15 downto 0);  y : out std_logic_vector
            (15 downto 0));
   end component;
   
   component iv_generic_NBIT16
      port( a : in std_logic_vector (15 downto 0);  y : out std_logic_vector 
            (15 downto 0));
   end component;
   
   signal sb_15_port, sb_14_port, sb_13_port, sb_12_port, sb_11_port, 
      sb_10_port, sb_9_port, sb_8_port, sb_7_port, sb_6_port, sb_5_port, 
      sb_4_port, sb_3_port, sb_2_port, sb_1_port, sb_0_port, y1_15_port, 
      y1_14_port, y1_13_port, y1_12_port, y1_11_port, y1_10_port, y1_9_port, 
      y1_8_port, y1_7_port, y1_6_port, y1_5_port, y1_4_port, y1_3_port, 
      y1_2_port, y1_1_port, y1_0_port, y2_15_port, y2_14_port, y2_13_port, 
      y2_12_port, y2_11_port, y2_10_port, y2_9_port, y2_8_port, y2_7_port, 
      y2_6_port, y2_5_port, y2_4_port, y2_3_port, y2_2_port, y2_1_port, 
      y2_0_port : std_logic;

begin
   
   UIV : iv_generic_NBIT16 port map( a(15) => s, a(14) => s, a(13) => s, a(12) 
                           => s, a(11) => s, a(10) => s, a(9) => s, a(8) => s, 
                           a(7) => s, a(6) => s, a(5) => s, a(4) => s, a(3) => 
                           s, a(2) => s, a(1) => s, a(0) => s, y(15) => 
                           sb_15_port, y(14) => sb_14_port, y(13) => sb_13_port
                           , y(12) => sb_12_port, y(11) => sb_11_port, y(10) =>
                           sb_10_port, y(9) => sb_9_port, y(8) => sb_8_port, 
                           y(7) => sb_7_port, y(6) => sb_6_port, y(5) => 
                           sb_5_port, y(4) => sb_4_port, y(3) => sb_3_port, 
                           y(2) => sb_2_port, y(1) => sb_1_port, y(0) => 
                           sb_0_port);
   UND1 : nd2_generic_NBIT16_0 port map( a(15) => a(15), a(14) => a(14), a(13) 
                           => a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(15) => s, b(14) => s, b(13) => s, b(12) => s, 
                           b(11) => s, b(10) => s, b(9) => s, b(8) => s, b(7) 
                           => s, b(6) => s, b(5) => s, b(4) => s, b(3) => s, 
                           b(2) => s, b(1) => s, b(0) => s, y(15) => y1_15_port
                           , y(14) => y1_14_port, y(13) => y1_13_port, y(12) =>
                           y1_12_port, y(11) => y1_11_port, y(10) => y1_10_port
                           , y(9) => y1_9_port, y(8) => y1_8_port, y(7) => 
                           y1_7_port, y(6) => y1_6_port, y(5) => y1_5_port, 
                           y(4) => y1_4_port, y(3) => y1_3_port, y(2) => 
                           y1_2_port, y(1) => y1_1_port, y(0) => y1_0_port);
   UND2 : nd2_generic_NBIT16_2 port map( a(15) => b(15), a(14) => b(14), a(13) 
                           => b(13), a(12) => b(12), a(11) => b(11), a(10) => 
                           b(10), a(9) => b(9), a(8) => b(8), a(7) => b(7), 
                           a(6) => b(6), a(5) => b(5), a(4) => b(4), a(3) => 
                           b(3), a(2) => b(2), a(1) => b(1), a(0) => b(0), 
                           b(15) => sb_15_port, b(14) => sb_14_port, b(13) => 
                           sb_13_port, b(12) => sb_12_port, b(11) => sb_11_port
                           , b(10) => sb_10_port, b(9) => sb_9_port, b(8) => 
                           sb_8_port, b(7) => sb_7_port, b(6) => sb_6_port, 
                           b(5) => sb_5_port, b(4) => sb_4_port, b(3) => 
                           sb_3_port, b(2) => sb_2_port, b(1) => sb_1_port, 
                           b(0) => sb_0_port, y(15) => y2_15_port, y(14) => 
                           y2_14_port, y(13) => y2_13_port, y(12) => y2_12_port
                           , y(11) => y2_11_port, y(10) => y2_10_port, y(9) => 
                           y2_9_port, y(8) => y2_8_port, y(7) => y2_7_port, 
                           y(6) => y2_6_port, y(5) => y2_5_port, y(4) => 
                           y2_4_port, y(3) => y2_3_port, y(2) => y2_2_port, 
                           y(1) => y2_1_port, y(0) => y2_0_port);
   UND3 : nd2_generic_NBIT16_1 port map( a(15) => y1_15_port, a(14) => 
                           y1_14_port, a(13) => y1_13_port, a(12) => y1_12_port
                           , a(11) => y1_11_port, a(10) => y1_10_port, a(9) => 
                           y1_9_port, a(8) => y1_8_port, a(7) => y1_7_port, 
                           a(6) => y1_6_port, a(5) => y1_5_port, a(4) => 
                           y1_4_port, a(3) => y1_3_port, a(2) => y1_2_port, 
                           a(1) => y1_1_port, a(0) => y1_0_port, b(15) => 
                           y2_15_port, b(14) => y2_14_port, b(13) => y2_13_port
                           , b(12) => y2_12_port, b(11) => y2_11_port, b(10) =>
                           y2_10_port, b(9) => y2_9_port, b(8) => y2_8_port, 
                           b(7) => y2_7_port, b(6) => y2_6_port, b(5) => 
                           y2_5_port, b(4) => y2_4_port, b(3) => y2_3_port, 
                           b(2) => y2_2_port, b(1) => y2_1_port, b(0) => 
                           y2_0_port, y(15) => y(15), y(14) => y(14), y(13) => 
                           y(13), y(12) => y(12), y(11) => y(11), y(10) => 
                           y(10), y(9) => y(9), y(8) => y(8), y(7) => y(7), 
                           y(6) => y(6), y(5) => y(5), y(4) => y(4), y(3) => 
                           y(3), y(2) => y(2), y(1) => y(1), y(0) => y(0));

end SYN_structural;
