library ieee;

package constants is

    constant numBit         : integer := 4;
    constant numBitXBlock   : integer := 1;

end package;