.subckt ND2HS A B Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:38:12 2001
*** spice backannotate
XMN0 net15 A gnd gnd ENHSGP_BS3JU W=0.640U L=0.130U 
+  AD=0.061P AS=0.305P PD=0.190U PS=2.870U 
XMN1 Z B net15 gnd ENHSGP_BS3JU W=0.640U L=0.130U 
+  AD=0.218P AS=0.061P PD=1.320U PS=0.190U 
XMP0 Z A vdd vdd EPHSGP_BS3JU W=0.770U L=0.130U 
+  AD=0.192P AS=0.471P PD=1.130U PS=4.130U 
XMP1 Z B vdd vdd EPHSGP_BS3JU W=0.770U L=0.130U 
+  AS=0.471P AD=0.192P PS=4.130U PD=1.130U 
C1 vdd gnd 0.142ff
C2 gnd gnd 0.897ff
C4 Z gnd 0.108ff
C5 A gnd 0.129ff
C6 B gnd 0.132ff
C1-2 vdd gnd 0.132ff
C1-4 vdd Z 0.018ff
C1-5 vdd A 0.002ff
C1-6 vdd B 0.002ff
C2-4 gnd Z 0.178ff
C2-5 gnd A 0.067ff
C2-6 gnd B 0.063ff
C4-5 Z A 0.099ff
C4-6 Z B 0.132ff
C5-6 A B 0.131ff
*
*
*
.ends ND2HS

.subckt ND2HSX8 A B Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:39:37 2001
*** spice backannotate
XMN7 net132 A gnd gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AD=0.160P AS=0.531P PD=0.250U PS=2.110U 
XMN6 Z B net132 gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AD=0.243P AS=0.160P PD=0.380U PS=0.250U 
XMN4 Z B net140 gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AS=0.150P AD=0.243P PS=0.235U PD=0.380U 
XMN5 net140 A gnd gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AS=0.243P AD=0.150P PS=0.380U PD=0.235U 
XMN2 net148 A gnd gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AD=0.150P AS=0.243P PD=0.235U PS=0.380U 
XMN3 Z B net148 gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AD=0.243P AS=0.150P PD=0.380U PS=0.235U 
XMN1 Z B net156 gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AS=0.150P AD=0.243P PS=0.235U PD=0.380U 
XMN0 net156 A gnd gnd ENHSGP_BS3JU W=1.280U L=0.130U 
+  AS=0.435P AD=0.150P PS=1.960U PD=0.235U 
XMP7 Z A vdd vdd EPHSGP_BS3JU W=2.050U L=0.130U 
+  AD=0.482P AS=0.674P PD=0.470U PS=2.810U 
XMP6 Z B vdd vdd EPHSGP_BS3JU W=2.050U L=0.130U 
+  AS=0.482P AD=0.482P PS=0.470U PD=0.470U 
XMP6_2 Z B vdd vdd EPHSGP_BS3JU W=2.050U L=0.130U 
+  AD=0.482P AS=0.482P PD=0.470U PS=0.470U 
XMP7_2 Z A vdd vdd EPHSGP_BS3JU W=2.050U L=0.130U 
+  AS=0.482P AD=0.482P PS=0.470U PD=0.470U 
XMP6_3 Z B vdd vdd EPHSGP_BS3JU W=2.050U L=0.130U 
+  AD=0.482P AS=0.482P PD=0.470U PS=0.470U 
XMP7_3 Z A vdd vdd EPHSGP_BS3JU W=2.050U L=0.130U 
+  AS=0.674P AD=0.482P PS=2.810U PD=0.470U 
C1 vdd gnd 0.341ff
C2 gnd gnd 1.486ff
C4 Z gnd 0.213ff
C8 A gnd 0.398ff
C9 B gnd 0.300ff
C1-2 vdd gnd 0.409ff
C1-8 vdd A 0.112ff
C1-9 vdd B 0.102ff
C2-4 gnd Z 0.602ff
C2-8 gnd A 0.475ff
C2-9 gnd B 0.341ff
C4-8 Z A 0.414ff
C4-9 Z B 0.243ff
C8-9 A B 0.825ff
*
*
*
.ends ND2HSX8

.subckt ND2LL A B Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:38:12 2001
*** spice backannotate
XMN0 net15 A gnd gnd ENLLGP_BS3JU W=0.640U L=0.130U 
+  AD=0.061P AS=0.305P PD=0.190U PS=2.870U 
XMN1 Z B net15 gnd ENLLGP_BS3JU W=0.640U L=0.130U 
+  AD=0.218P AS=0.061P PD=1.320U PS=0.190U 
XMP0 Z A vdd vdd EPLLGP_BS3JU W=0.770U L=0.130U 
+  AD=0.192P AS=0.471P PD=1.130U PS=4.130U 
XMP1 Z B vdd vdd EPLLGP_BS3JU W=0.770U L=0.130U 
+  AS=0.471P AD=0.192P PS=4.130U PD=1.130U 
C1 vdd gnd 0.142ff
C2 gnd gnd 0.897ff
C4 Z gnd 0.108ff
C5 A gnd 0.129ff
C6 B gnd 0.132ff
C1-2 vdd gnd 0.132ff
C1-4 vdd Z 0.018ff
C1-5 vdd A 0.002ff
C1-6 vdd B 0.002ff
C2-4 gnd Z 0.178ff
C2-5 gnd A 0.067ff
C2-6 gnd B 0.063ff
C4-5 Z A 0.099ff
C4-6 Z B 0.132ff
C5-6 A B 0.131ff
*
*
*
.ends ND2LL

.subckt ND2LLX8 A B Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:39:37 2001
*** spice backannotate
XMN7 net132 A gnd gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AD=0.160P AS=0.531P PD=0.250U PS=2.110U 
XMN6 Z B net132 gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AD=0.243P AS=0.160P PD=0.380U PS=0.250U 
XMN4 Z B net140 gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AS=0.150P AD=0.243P PS=0.235U PD=0.380U 
XMN5 net140 A gnd gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AS=0.243P AD=0.150P PS=0.380U PD=0.235U 
XMN2 net148 A gnd gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AD=0.150P AS=0.243P PD=0.235U PS=0.380U 
XMN3 Z B net148 gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AD=0.243P AS=0.150P PD=0.380U PS=0.235U 
XMN1 Z B net156 gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AS=0.150P AD=0.243P PS=0.235U PD=0.380U 
XMN0 net156 A gnd gnd ENLLGP_BS3JU W=1.280U L=0.130U 
+  AS=0.435P AD=0.150P PS=1.960U PD=0.235U 
XMP7 Z A vdd vdd EPLLGP_BS3JU W=2.050U L=0.130U 
+  AD=0.482P AS=0.674P PD=0.470U PS=2.810U 
XMP6 Z B vdd vdd EPLLGP_BS3JU W=2.050U L=0.130U 
+  AS=0.482P AD=0.482P PS=0.470U PD=0.470U 
XMP6_2 Z B vdd vdd EPLLGP_BS3JU W=2.050U L=0.130U 
+  AD=0.482P AS=0.482P PD=0.470U PS=0.470U 
XMP7_2 Z A vdd vdd EPLLGP_BS3JU W=2.050U L=0.130U 
+  AS=0.482P AD=0.482P PS=0.470U PD=0.470U 
XMP6_3 Z B vdd vdd EPLLGP_BS3JU W=2.050U L=0.130U 
+  AD=0.482P AS=0.482P PD=0.470U PS=0.470U 
XMP7_3 Z A vdd vdd EPLLGP_BS3JU W=2.050U L=0.130U 
+  AS=0.674P AD=0.482P PS=2.810U PD=0.470U 
C1 vdd gnd 0.341ff
C2 gnd gnd 1.486ff
C4 Z gnd 0.213ff
C8 A gnd 0.398ff
C9 B gnd 0.300ff
C1-2 vdd gnd 0.409ff
C1-8 vdd A 0.112ff
C1-9 vdd B 0.102ff
C2-4 gnd Z 0.602ff
C2-8 gnd A 0.475ff
C2-9 gnd B 0.341ff
C4-8 Z A 0.414ff
C4-9 Z B 0.243ff
C8-9 A B 0.825ff
*
*
*
.ends ND2LLX8


.subckt IVHS A Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:05:54 2001
*** spice backannotate
XMN0 Z A gnd gnd ENHSGP_BS3JU W=0.585U L=0.130U 
+  AD=0.216P AS=0.426P PD=1.325U PS=2.725U 
XMP0 Z A vdd vdd EPHSGP_BS3JU W=1.050U L=0.130U 
+  AD=0.389P AS=0.734P PD=1.790U PS=4.090U 
C1 vdd gnd 0.147ff
C2 gnd gnd 0.929ff
C3 Z gnd 0.072ff
C4 A gnd 0.167ff
C1-2 vdd gnd 0.136ff
C1-4 vdd A 0.002ff
C2-3 gnd Z 0.110ff
C2-4 gnd A 0.098ff
C3-4 Z A 0.061ff
*
*
*
.ends IVHS

.subckt IVHSX8 A Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:08:32 2001
*** spice backannotate
XMN3 Z A gnd gnd ENHSGP_BS3JU W=1.170U L=0.130U 
+  AD=0.257P AS=0.433P PD=0.440U PS=1.910U 
XMN3_2 Z A gnd gnd ENHSGP_BS3JU W=1.170U L=0.130U 
+  AS=0.257P AD=0.257P PS=0.440U PD=0.440U 
XMN3_3 Z A gnd gnd ENHSGP_BS3JU W=1.170U L=0.130U 
+  AD=0.257P AS=0.257P PD=0.440U PS=0.440U 
XMN3_4 Z A gnd gnd ENHSGP_BS3JU W=1.170U L=0.130U 
+  AS=0.433P AD=0.257P PS=1.910U PD=0.440U 
XMP3 Z A vdd vdd EPHSGP_BS3JU W=2.100U L=0.130U 
+  AD=0.462P AS=0.777P PD=0.440U PS=2.840U 
XMP3_2 Z A vdd vdd EPHSGP_BS3JU W=2.100U L=0.130U 
+  AS=0.462P AD=0.462P PS=0.440U PD=0.440U 
XMP3_3 Z A vdd vdd EPHSGP_BS3JU W=2.100U L=0.130U 
+  AD=0.462P AS=0.462P PD=0.440U PS=0.440U 
XMP3_4 Z A vdd vdd EPHSGP_BS3JU W=2.100U L=0.130U 
+  AS=0.777P AD=0.462P PS=2.840U PD=0.440U 
C1 vdd gnd 0.263ff
C2 gnd gnd 1.247ff
C3 Z gnd 0.160ff
C4 A gnd 0.414ff
C1-2 vdd gnd 0.309ff
C1-3 vdd Z 0.007ff
C1-4 vdd A 0.168ff
C2-3 gnd Z 0.523ff
C2-4 gnd A 0.315ff
C3-4 Z A 0.473ff
*
*
*
.ends IVHSX8

.subckt IVHSA A Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:05:54 2001
*** spice backannotate
XMN0 Z A gnd gnd ENHSGP_BS3JU W=2.585U L=0.130U 
+  AD=0.916P AS=1.56P PD=1.825U PS=2.725U 
XMP0 Z A vdd vdd EPHSGP_BS3JU W=4.050U L=0.130U 
+  AD=1.4P AS=2.634P PD=2.790U PS=4.090U 
C1 vdd gnd 0.147ff
C2 vdd gnd 0.929ff
C3 Z gnd 0.072ff
C4 A gnd 0.167ff
C1-2 vdd gnd 0.136ff
C1-4 vdd A 0.002ff
C2-3 gnd Z 0.110ff
C2-4 gnd A 0.098ff
C3-4 Z A 0.061ff
*
*
*
.ends IVHSA


.subckt IVLL A Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:05:54 2001
*** spice backannotate
XMN0 Z A gnd gnd ENLLGP_BS3JU W=0.585U L=0.130U 
+  AD=0.216P AS=0.426P PD=1.325U PS=2.725U 
XMP0 Z A vdd vdd EPLLGP_BS3JU W=1.050U L=0.130U 
+  AD=0.389P AS=0.734P PD=1.790U PS=4.090U 
C1 vdd gnd 0.147ff
C2 gnd gnd 0.929ff
C3 Z gnd 0.072ff
C4 A gnd 0.167ff
C1-2 vdd gnd 0.136ff
C1-4 vdd A 0.002ff
C2-3 gnd Z 0.110ff
C2-4 gnd A 0.098ff
C3-4 Z A 0.061ff
*
*
*
.ends IVLL



.subckt NR2HS A B Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:54:55 2001
*** spice backannotate
XMN0 Z A gnd gnd ENHSGP_BS3JU W=0.340U L=0.130U 
+  AD=0.116P AS=0.323P PD=0.995U PS=3.445U 
XMN1 Z B gnd gnd ENHSGP_BS3JU W=0.340U L=0.130U 
+  AS=0.323P AD=0.116P PS=3.445U PD=0.995U 
XMP0 net028 A vdd vdd EPHSGP_BS3JU W=1.050U L=0.130U 
+  AD=0.131P AS=0.689P PD=0.250U PS=4.990U 
XMP1 Z B net028 vdd EPHSGP_BS3JU W=1.050U L=0.130U 
+  AD=0.423P AS=0.131P PD=3.180U PS=0.250U 
C1 vdd gnd 0.135ff
C2 gnd gnd 0.899ff
C3 Z gnd 0.135ff
C5 A gnd 0.117ff
C6 B gnd 0.117ff
C1-2 vdd gnd 0.125ff
C1-3 vdd Z 0.048ff
C1-5 vdd A 0.002ff
C2-3 gnd Z 0.211ff
C2-5 gnd A 0.059ff
C2-6 gnd B 0.058ff
C3-5 Z A 0.105ff
C3-6 Z B 0.109ff
C5-6 A B 0.104ff
*
*
*
.ends NR2HS

.subckt NR2LL A B Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 23:54:55 2001
*** spice backannotate
XMN0 Z A gnd gnd ENLLGP_BS3JU W=0.340U L=0.130U 
+  AD=0.116P AS=0.323P PD=0.995U PS=3.445U 
XMN1 Z B gnd gnd ENLLGP_BS3JU W=0.340U L=0.130U 
+  AS=0.323P AD=0.116P PS=3.445U PD=0.995U 
XMP0 net028 A vdd vdd EPLLGP_BS3JU W=1.050U L=0.130U 
+  AD=0.131P AS=0.689P PD=0.250U PS=4.990U 
XMP1 Z B net028 vdd EPLLGP_BS3JU W=1.050U L=0.130U 
+  AD=0.423P AS=0.131P PD=3.180U PS=0.250U 
C1 vdd gnd 0.135ff
C2 gnd gnd 0.899ff
C3 Z gnd 0.135ff
C5 A gnd 0.117ff
C6 B gnd 0.117ff
C1-2 vdd gnd 0.125ff
C1-3 vdd Z 0.048ff
C1-5 vdd A 0.002ff
C2-3 gnd Z 0.211ff
C2-5 gnd A 0.059ff
C2-6 gnd B 0.058ff
C3-5 Z A 0.105ff
C3-6 Z B 0.109ff
C5-6 A B 0.104ff
*
*
*
.ends NR2LL



.subckt FA1HS A B CI CO Z gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 22:39:06 2001
*** spice backannotate
XMN5 CO net168 gnd gnd ENHSGP_BS3JU W=0.585U L=0.130U 
+  AS=0.327P AD=0.199P PS=2.429U PD=1.265U 
XMN2 net200 B gnd gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AD=0.160P AS=0.168P PD=1.600U PS=1.246U 
XMN3 net168 CI net200 gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AD=0.060P AS=0.160P PD=0.400U PS=1.600U 
XMN4 net168 B net204 gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AS=0.027P AD=0.060P PS=0.180U PD=0.400U 
XMN1 net200 A gnd gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AS=0.142P AD=0.160P PS=1.365U PD=1.600U 
XMN0 net204 A gnd gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AS=0.142P AD=0.027P PS=1.365U PD=0.180U 
XMN10 net188 A gnd gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AD=0.146P AS=0.290P PD=1.570U PS=3.240U 
XMN8 net188 B gnd gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AS=0.112P AD=0.146P PS=1.060U PD=1.570U 
XMN11 net188 CI gnd gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AD=0.146P AS=0.112P PD=1.570U PS=1.060U 
XMN9 net184 net168 net188 gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AD=0.110P AS=0.146P PD=1.030U PS=1.570U 
XMN6 net184 CI net156 gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AS=0.032P AD=0.110P PS=0.210U PD=1.030U 
XMN12 net156 A net176 gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AS=0.032P AD=0.032P PS=0.210U PD=0.210U 
XMN7 net176 B gnd gnd ENHSGP_BS3JU W=0.300U L=0.130U 
+  AS=0.160P AD=0.032P PS=1.286U PD=0.210U 
XMN13 Z net184 gnd gnd ENHSGP_BS3JU W=0.585U L=0.130U 
+  AD=0.240P AS=0.312P PD=1.405U PS=2.509U 
XMP7 CO net168 vdd vdd EPHSGP_BS3JU W=1.050U L=0.130U 
+  AS=0.373P AD=0.357P PS=2.475U PD=1.730U 
XMP1 net135 B vdd vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AD=0.172P AS=0.224P PD=1.210U PS=1.485U 
XMP2 net168 CI net135 vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AD=0.120P AS=0.172P PD=0.380U PS=1.210U 
XMP6 net168 B net114 vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AS=0.057P AD=0.120P PS=0.180U PD=0.380U 
XMP5 net114 A vdd vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AS=0.214P AD=0.057P PS=1.310U PD=0.180U 
XMP4 net135 A vdd vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AS=0.276P AD=0.214P PS=2.395U PD=1.310U 
XMP11 net146 A vdd vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AD=0.177P AS=0.276P PD=1.280U PS=2.395U 
XMP8 net146 B vdd vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AS=0.276P AD=0.177P PS=2.395U PD=1.280U 
XMP13 net146 CI vdd vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AD=0.177P AS=0.276P PD=1.280U PS=2.395U 
XMP12 net184 net168 net146 vdd EPHSGP_BS3JU W=0.630U L=0.130U 
+  AD=0.121P AS=0.177P PD=0.390U PS=1.280U 
XMP9 net184 CI net122 vdd EPHSGP_BS3JU W=0.680U L=0.130U 
+  AS=0.061P AD=0.131P PS=0.180U PD=0.420U 
XMP14 net122 A net98 vdd EPHSGP_BS3JU W=0.680U L=0.130U 
+  AS=0.061P AD=0.061P PS=0.180U PD=0.180U 
XMP10 net98 B vdd vdd EPHSGP_BS3JU W=0.680U L=0.130U 
+  AS=0.254P AD=0.061P PS=1.560U PD=0.180U 
XMP15 Z net184 vdd vdd EPHSGP_BS3JU W=1.050U L=0.130U 
+  AD=0.326P AS=0.392P PD=1.770U PS=2.410U 
C1 vdd gnd 0.484ff
C2 gnd gnd 2.079ff
C3 CO gnd 0.104ff
C5 net168 gnd 0.303ff
C8 net184 gnd 0.204ff
C11 Z gnd 0.078ff
C12 net135 gnd 0.018ff
C14 net146 gnd 0.021ff
C17 B gnd 0.459ff
C18 CI gnd 0.625ff
C19 A gnd 0.670ff
C1-2 vdd gnd 0.654ff
C1-5 vdd net168 0.009ff
C1-8 vdd net184 0.004ff
C1-12 vdd net135 0.087ff
C1-14 vdd net146 0.093ff
C1-17 vdd B 0.097ff
C1-18 vdd CI 0.291ff
C1-19 vdd A 0.085ff
C2-3 gnd CO 0.170ff
C2-5 gnd net168 0.388ff
C2-8 gnd net184 0.319ff
C2-11 gnd Z 0.104ff
C2-12 gnd net135 0.048ff
C2-14 gnd net146 0.052ff
C2-17 gnd B 0.391ff
C2-18 gnd CI 0.097ff
C2-19 gnd A 0.370ff
C3-5 CO net168 0.167ff
C3-17 CO B 0.006ff
C5-8 net168 net184 0.008ff
C5-12 net168 net135 0.012ff
C5-14 net168 net146 0.001ff
C5-17 net168 B 0.340ff
C5-18 net168 CI 0.291ff
C5-19 net168 A 0.088ff
C8-11 net184 Z 0.188ff
C8-17 net184 B 0.244ff
C8-18 net184 CI 0.025ff
C8-19 net184 A 0.051ff
C12-17 net135 B 0.003ff
C12-18 net135 CI 0.074ff
C12-19 net135 A 0.012ff
C14-17 net146 B 0.057ff
C14-18 net146 CI 0.020ff
C14-19 net146 A 0.003ff
C17-18 B CI 0.406ff
C17-19 B A 0.558ff
C18-19 CI A 0.173ff
*
*
*
.ends FA1HS
	

.subckt FD1QLL CP D Q gnd vdd
*** Version 5.500
*** Create time, Fri Jul 13 22:41:02 2001
*** spice backannotate
XMN2 net0176 D gnd gnd ENLLGP_BS3JU W=0.240U L=0.130U 
+  AS=0.099P AD=0.264P PS=0.684U PD=2.200U 
XMN0 CPN CP gnd gnd ENLLGP_BS3JU W=0.600U L=0.130U 
+  AS=0.246P AD=0.204P PS=1.711U PD=1.280U 
XMN1 CPI CPN gnd gnd ENLLGP_BS3JU W=0.300U L=0.130U 
+  AD=0.102P AS=0.123P PD=0.980U PS=0.855U 
XMN15 MN CPN net0176 gnd ENLLGP_BS3JU W=0.300U L=0.130U 
+  AD=0.111P AS=0.111P PD=1.040U PS=1.040U 
XMN8 M MN gnd gnd ENLLGP_BS3JU W=0.150U L=0.130U 
+  AS=0.065P AD=0.101P PS=0.514U PD=1.190U 
XMN9 net151 M gnd gnd ENLLGP_BS3JU W=0.540U L=0.130U 
+  AD=0.103P AS=0.234P PD=0.380U PS=1.851U 
XMN7 net040 M gnd gnd ENLLGP_BS3JU W=0.150U L=0.130U 
+  AD=0.014P AS=0.065P PD=0.180U PS=0.514U 
XMN6 MN CPI net040 gnd ENLLGP_BS3JU W=0.150U L=0.130U 
+  AD=0.101P AS=0.014P PD=1.190U PS=0.180U 
XMN10 SN CPI net151 gnd ENLLGP_BS3JU W=0.540U L=0.130U 
+  AD=0.155P AS=0.103P PD=0.994U PS=0.380U 
XMN13 SN CPN net0149 gnd ENLLGP_BS3JU W=0.150U L=0.130U 
+  AS=0.014P AD=0.043P PS=0.180U PD=0.276U 
XMN12 net0149 S gnd gnd ENLLGP_BS3JU W=0.150U L=0.130U 
+  AS=0.054P AD=0.014P PS=0.365U PD=0.180U 
XMN11 S SN gnd gnd ENLLGP_BS3JU W=0.230U L=0.130U 
+  AS=0.082P AD=0.157P PS=0.560U PD=1.450U 
XMN14 Q SN gnd gnd ENLLGP_BS3JU W=0.590U L=0.130U 
+  AD=0.182P AS=0.211P PD=1.270U PS=1.435U 
XMP3 net0218 D vdd vdd EPLLGP_BS3JU W=0.700U L=0.130U 
+  AS=0.333P AD=0.238P PS=1.488U PD=1.380U 
XMP0 CPN CP vdd vdd EPLLGP_BS3JU W=0.600U L=0.130U 
+  AS=0.285P AD=0.204P PS=1.276U PD=1.280U 
XMP1 CPI CPN vdd vdd EPLLGP_BS3JU W=0.600U L=0.130U 
+  AD=0.207P AS=0.285P PD=1.290U PS=1.276U 
XMP15 MN CPI net0218 vdd EPLLGP_BS3JU W=0.630U L=0.130U 
+  AD=0.198P AS=0.206P PD=1.310U PS=1.310U 
XMP8 M MN vdd vdd EPLLGP_BS3JU W=0.300U L=0.130U 
+  AS=0.152P AD=0.102P PS=0.993U PD=0.980U 
XMP9 net151 M vdd vdd EPLLGP_BS3JU W=0.750U L=0.130U 
+  AD=0.142P AS=0.381P PD=0.380U PS=2.481U 
XMP6 net075 M vdd vdd EPLLGP_BS3JU W=0.150U L=0.130U 
+  AD=0.014P AS=0.076P PD=0.180U PS=0.496U 
XMP10 SN CPN net151 vdd EPLLGP_BS3JU W=0.750U L=0.130U 
+  AD=0.207P AS=0.142P PD=1.183U PS=0.380U 
XMP7 MN CPN net075 vdd EPLLGP_BS3JU W=0.150U L=0.130U 
+  AD=0.101P AS=0.014P PD=1.190U PS=0.180U 
XMP12 SN CPI net0196 vdd EPLLGP_BS3JU W=0.150U L=0.130U 
+  AS=0.030P AD=0.041P PS=0.405U PD=0.237U 
XMP13 net0196 S vdd vdd EPLLGP_BS3JU W=0.150U L=0.130U 
+  AS=0.050P AD=0.030P PS=0.294U PD=0.405U 
XMP11 S SN vdd vdd EPLLGP_BS3JU W=0.280U L=0.130U 
+  AS=0.094P AD=0.159P PS=0.549U PD=1.390U 
XMP14 Q SN vdd vdd EPLLGP_BS3JU W=1.050U L=0.130U 
+  AD=0.305P AS=0.352P PD=1.730U PS=2.057U 
C1 vdd gnd 0.450ff
C2 net0176 gnd 0.052ff
C3 CPN gnd 0.614ff
C4 gnd gnd 2.037ff
C5 CPI gnd 0.252ff
C6 MN gnd 0.192ff
C7 M gnd 0.153ff
C8 net151 gnd 0.021ff
C10 SN gnd 0.340ff
C12 S gnd 0.146ff
C13 Q gnd 0.083ff
C14 net0218 gnd 0.049ff
C17 D gnd 0.267ff
C18 CP gnd 0.090ff
C1-3 vdd CPN 0.186ff
C1-4 vdd gnd 0.599ff
C1-5 vdd CPI 0.021ff
C1-6 vdd MN 0.076ff
C1-7 vdd M 0.007ff
C1-10 vdd SN 0.098ff
C1-12 vdd S 0.035ff
C1-14 vdd net0218 0.126ff
C1-17 vdd D 0.035ff
C1-18 vdd CP 0.001ff
C2-3 net0176 CPN 0.040ff
C2-4 net0176 gnd 0.216ff
C2-5 net0176 CPI 0.007ff
C2-6 net0176 MN 0.012ff
C2-17 net0176 D 0.039ff
C2-18 net0176 CP 0.010ff
C3-4 CPN gnd 0.317ff
C3-5 CPN CPI 0.262ff
C3-6 CPN MN 0.074ff
C3-7 CPN M 0.106ff
C3-8 CPN net151 0.011ff
C3-10 CPN SN 0.033ff
C3-12 CPN S 0.052ff
C3-14 CPN net0218 0.017ff
C3-17 CPN D 0.030ff
C3-18 CPN CP 0.190ff
C4-5 gnd CPI 0.189ff
C4-6 gnd MN 0.296ff
C4-7 gnd M 0.115ff
C4-8 gnd net151 0.049ff
C4-10 gnd SN 0.208ff
C4-12 gnd S 0.204ff
C4-13 gnd Q 0.148ff
C4-14 gnd net0218 0.091ff
C4-17 gnd D 0.130ff
C4-18 gnd CP 0.069ff
C5-6 CPI MN 0.189ff
C5-7 CPI M 0.182ff
C5-8 CPI net151 0.027ff
C5-10 CPI SN 0.089ff
C5-12 CPI S 0.065ff
C5-14 CPI net0218 0.013ff
C5-18 CPI CP 0.025ff
C6-7 MN M 0.213ff
C6-8 MN net151 0.023ff
C6-10 MN SN 0.018ff
C6-12 MN S 0.036ff
C6-14 MN net0218 0.005ff
C7-8 M net151 0.054ff
C8-10 net151 SN 0.077ff
C10-12 SN S 0.210ff
C10-13 SN Q 0.067ff
C12-13 S Q 0.059ff
C14-17 net0218 D 0.019ff
C14-18 net0218 CP 0.034ff
C17-18 D CP 0.095ff
*
*
*
.ends FD1QLL
