
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N5_M2_1 is

   port( S : in std_logic_vector (1 downto 0);  Q : in std_logic_vector (19 
         downto 0);  Y : out std_logic_vector (4 downto 0));

end mux_N5_M2_1;

architecture SYN_behav of mux_N5_M2_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => Y(4));
   U3 : AOI22_X1 port map( A1 => Q(4), A2 => n3, B1 => Q(14), B2 => n4, ZN => 
                           n2);
   U4 : AOI22_X1 port map( A1 => Q(19), A2 => n5, B1 => Q(9), B2 => n6, ZN => 
                           n1);
   U5 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => Q(3), A2 => n3, B1 => Q(13), B2 => n4, ZN => 
                           n8);
   U7 : AOI22_X1 port map( A1 => Q(18), A2 => n5, B1 => Q(8), B2 => n6, ZN => 
                           n7);
   U8 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => Q(2), A2 => n3, B1 => Q(12), B2 => n4, ZN => 
                           n10);
   U10 : AOI22_X1 port map( A1 => Q(17), A2 => n5, B1 => Q(7), B2 => n6, ZN => 
                           n9);
   U11 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => Q(1), A2 => n3, B1 => Q(11), B2 => n4, ZN => 
                           n12);
   U13 : AOI22_X1 port map( A1 => Q(16), A2 => n5, B1 => Q(6), B2 => n6, ZN => 
                           n11);
   U14 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => Y(0));
   U15 : AOI22_X1 port map( A1 => Q(0), A2 => n3, B1 => Q(10), B2 => n4, ZN => 
                           n14);
   U16 : NOR3_X1 port map( A1 => n5, A2 => n6, A3 => n4, ZN => n3);
   U17 : NOR2_X1 port map( A1 => n15, A2 => S(0), ZN => n4);
   U18 : AOI22_X1 port map( A1 => Q(15), A2 => n5, B1 => Q(5), B2 => n6, ZN => 
                           n13);
   U19 : NOR2_X1 port map( A1 => n16, A2 => S(1), ZN => n6);
   U20 : NOR2_X1 port map( A1 => n15, A2 => n16, ZN => n5);
   U21 : INV_X1 port map( A => S(0), ZN => n16);
   U22 : INV_X1 port map( A => S(1), ZN => n15);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity address_generator_N16_1 is

   port( clk, rst, enable : in std_logic;  done, working : out std_logic;  addr
         : out std_logic_vector (15 downto 0));

end address_generator_N16_1;

architecture SYN_struct of address_generator_N16_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal done_port, addr_14_port, addr_13_port, addr_12_port, addr_11_port, 
      addr_10_port, addr_9_port, addr_8_port, addr_7_port, addr_6_port, 
      addr_5_port, addr_4_port, addr_3_port, addr_2_port, addr_1_port, 
      addr_0_port, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
      N19, N20, N21, n2, n3, n4, n5, n6_port, n7_port, n8_port, n9_port, 
      n10_port, n11_port, n12_port, n13_port, n14_port, n15_port, n16_port, 
      n17_port, n18_port, working_port, n20_port : std_logic;

begin
   done <= done_port;
   working <= working_port;
   addr <= ( done_port, addr_14_port, addr_13_port, addr_12_port, addr_11_port,
      addr_10_port, addr_9_port, addr_8_port, addr_7_port, addr_6_port, 
      addr_5_port, addr_4_port, addr_3_port, addr_2_port, addr_1_port, 
      addr_0_port );
   
   curr_addr_reg_0_inst : DFF_X1 port map( D => N6, CK => clk, Q => addr_0_port
                           , QN => working_port);
   curr_addr_reg_1_inst : DFF_X1 port map( D => N7, CK => clk, Q => addr_1_port
                           , QN => n6_port);
   curr_addr_reg_2_inst : DFF_X1 port map( D => N8, CK => clk, Q => addr_2_port
                           , QN => n5);
   curr_addr_reg_3_inst : DFF_X1 port map( D => N9, CK => clk, Q => addr_3_port
                           , QN => n18_port);
   curr_addr_reg_4_inst : DFF_X1 port map( D => N10, CK => clk, Q => 
                           addr_4_port, QN => n17_port);
   curr_addr_reg_5_inst : DFF_X1 port map( D => N11, CK => clk, Q => 
                           addr_5_port, QN => n16_port);
   curr_addr_reg_6_inst : DFF_X1 port map( D => N12, CK => clk, Q => 
                           addr_6_port, QN => n15_port);
   curr_addr_reg_7_inst : DFF_X1 port map( D => N13, CK => clk, Q => 
                           addr_7_port, QN => n14_port);
   curr_addr_reg_8_inst : DFF_X1 port map( D => N14, CK => clk, Q => 
                           addr_8_port, QN => n13_port);
   curr_addr_reg_9_inst : DFF_X1 port map( D => N15, CK => clk, Q => 
                           addr_9_port, QN => n12_port);
   curr_addr_reg_10_inst : DFF_X1 port map( D => N16, CK => clk, Q => 
                           addr_10_port, QN => n11_port);
   curr_addr_reg_11_inst : DFF_X1 port map( D => N17, CK => clk, Q => 
                           addr_11_port, QN => n10_port);
   curr_addr_reg_12_inst : DFF_X1 port map( D => N18, CK => clk, Q => 
                           addr_12_port, QN => n9_port);
   curr_addr_reg_13_inst : DFF_X1 port map( D => N19, CK => clk, Q => 
                           addr_13_port, QN => n8_port);
   curr_addr_reg_14_inst : DFF_X1 port map( D => N20, CK => clk, Q => 
                           addr_14_port, QN => n7_port);
   curr_addr_reg_15_inst : DFF_X1 port map( D => N21, CK => clk, Q => done_port
                           , QN => n20_port);
   U3 : NOR2_X1 port map( A1 => n5, A2 => n2, ZN => N9);
   U4 : NOR2_X1 port map( A1 => n6_port, A2 => n2, ZN => N8);
   U5 : NOR2_X1 port map( A1 => working_port, A2 => n2, ZN => N7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n20_port, ZN => N6);
   U7 : NOR2_X1 port map( A1 => n7_port, A2 => n2, ZN => N21);
   U8 : NOR2_X1 port map( A1 => n8_port, A2 => n2, ZN => N20);
   U9 : NOR2_X1 port map( A1 => n9_port, A2 => n2, ZN => N19);
   U10 : NOR2_X1 port map( A1 => n10_port, A2 => n2, ZN => N18);
   U11 : NOR2_X1 port map( A1 => n11_port, A2 => n2, ZN => N17);
   U12 : NOR2_X1 port map( A1 => n12_port, A2 => n2, ZN => N16);
   U13 : NOR2_X1 port map( A1 => n13_port, A2 => n2, ZN => N15);
   U14 : NOR2_X1 port map( A1 => n14_port, A2 => n2, ZN => N14);
   U15 : NOR2_X1 port map( A1 => n15_port, A2 => n2, ZN => N13);
   U16 : NOR2_X1 port map( A1 => n16_port, A2 => n2, ZN => N12);
   U17 : NOR2_X1 port map( A1 => n17_port, A2 => n2, ZN => N11);
   U18 : NOR2_X1 port map( A1 => n18_port, A2 => n2, ZN => N10);
   U19 : INV_X1 port map( A => n3, ZN => n2);
   U20 : NOR2_X1 port map( A1 => rst, A2 => n4, ZN => n3);
   U21 : AOI21_X1 port map( B1 => working_port, B2 => n20_port, A => enable, ZN
                           => n4);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity equal_check_N5_1 is

   port( A, B : in std_logic_vector (4 downto 0);  EQUAL : out std_logic);

end equal_check_N5_1;

architecture SYN_behav of equal_check_N5_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => n1, A2 => n2, A3 => n3, ZN => EQUAL);
   U2 : XOR2_X1 port map( A => B(4), B => A(4), Z => n3);
   U3 : XOR2_X1 port map( A => B(2), B => A(2), Z => n2);
   U4 : NAND3_X1 port map( A1 => n4, A2 => n5, A3 => n6, ZN => n1);
   U5 : XNOR2_X1 port map( A => B(0), B => A(0), ZN => n6);
   U6 : XNOR2_X1 port map( A => B(1), B => A(1), ZN => n5);
   U7 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_39 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_39;

architecture SYN_behav of mux_N32_M1_39 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_38 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_38;

architecture SYN_behav of mux_N32_M1_38 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_37 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_37;

architecture SYN_behav of mux_N32_M1_37 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_36 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_36;

architecture SYN_behav of mux_N32_M1_36 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_35 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_35;

architecture SYN_behav of mux_N32_M1_35 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_34 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_34;

architecture SYN_behav of mux_N32_M1_34 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_33 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_33;

architecture SYN_behav of mux_N32_M1_33 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_32 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_32;

architecture SYN_behav of mux_N32_M1_32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_31 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_31;

architecture SYN_behav of mux_N32_M1_31 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_30 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_30;

architecture SYN_behav of mux_N32_M1_30 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_29 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_29;

architecture SYN_behav of mux_N32_M1_29 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_28 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_28;

architecture SYN_behav of mux_N32_M1_28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_27 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_27;

architecture SYN_behav of mux_N32_M1_27 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_26 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_26;

architecture SYN_behav of mux_N32_M1_26 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_25 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_25;

architecture SYN_behav of mux_N32_M1_25 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_24 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_24;

architecture SYN_behav of mux_N32_M1_24 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_23 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_23;

architecture SYN_behav of mux_N32_M1_23 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_22 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_22;

architecture SYN_behav of mux_N32_M1_22 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_21 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_21;

architecture SYN_behav of mux_N32_M1_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_20 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_20;

architecture SYN_behav of mux_N32_M1_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_19 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_19;

architecture SYN_behav of mux_N32_M1_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_18 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_18;

architecture SYN_behav of mux_N32_M1_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_17 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_17;

architecture SYN_behav of mux_N32_M1_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_16 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_16;

architecture SYN_behav of mux_N32_M1_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_15 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_15;

architecture SYN_behav of mux_N32_M1_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_14 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_14;

architecture SYN_behav of mux_N32_M1_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_13 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_13;

architecture SYN_behav of mux_N32_M1_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_12 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_12;

architecture SYN_behav of mux_N32_M1_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_11 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_11;

architecture SYN_behav of mux_N32_M1_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_10 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_10;

architecture SYN_behav of mux_N32_M1_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_9 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_9;

architecture SYN_behav of mux_N32_M1_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_8 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_8;

architecture SYN_behav of mux_N32_M1_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_7 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_7;

architecture SYN_behav of mux_N32_M1_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_6 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_6;

architecture SYN_behav of mux_N32_M1_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_5 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_5;

architecture SYN_behav of mux_N32_M1_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_4 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_4;

architecture SYN_behav of mux_N32_M1_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_3 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_3;

architecture SYN_behav of mux_N32_M1_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_2 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_2;

architecture SYN_behav of mux_N32_M1_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_1 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_1;

architecture SYN_behav of mux_N32_M1_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_89 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_89;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_88 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_88;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_87 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_87;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_86 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_86;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_85 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_85;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_84 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_84;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_83 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_83;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_82 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_82;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_81 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_81;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_80 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_80;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_79 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_79;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_78 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_78;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_77 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_77;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_76 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_76;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_75 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_75;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_74 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_74;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_73 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_73;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_72 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_72;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_71 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_71;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_70 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_70;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_69 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_69;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_68 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_68;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_67 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_67;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_66 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_66;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_65 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_65;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_64 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_64;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_63 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_63;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_62 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_62;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_61 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_61;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_60 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_60;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_59 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_59;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_58 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_58;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_57 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_57;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_56 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_56;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_55 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_55;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_54 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_54;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_53 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_53;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_52 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_52;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_51 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_51;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_50 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_50;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_49 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_49;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_48 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_48;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_47 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_47;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_46 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_46;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_45 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_45;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_44 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_44;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_43 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_43;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_42 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_42;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_41 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_41;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_40 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_40;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_39 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_39;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_38 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_38;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_37 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_37;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_36 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_36;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_35 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_35;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_34 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_34;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_33 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_33;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_32 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_32;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_31 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_31;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_30 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_30;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_29 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_29;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_28 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_28;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_27 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_27;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_26 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_26;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_25 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_25;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_24 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_24;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_23 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_23;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_22 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_22;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_21 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_21;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_20 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_20;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_19 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_19;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_18 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_18;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_17 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_17;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_16 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_16;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_15 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_15;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_14 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_14;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_13 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_13;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_12 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_12;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_11 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_11;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_10 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_10;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_9 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_9;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_8 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_8;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_7 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_7;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_6 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_6;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_5 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_5;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_4 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_4;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_3 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_3;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_2 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_2;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(31), QN => n68)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(30), QN => n67)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(29), QN => n66)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(28), QN => n65)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(27), QN => n64)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(26), QN => n63)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(25), QN => n62)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(24), QN => n61)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(23), QN => n60)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(22), QN => n59)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(21), QN => n58)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(20), QN => n57)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(19), QN => n56)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(18), QN => n55)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(17), QN => n54)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(16), QN => n53)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(15), QN => n52)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(14), QN => n51)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(13), QN => n50)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(12), QN => n49)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(11), QN => n48)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(10), QN => n47)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(9), QN => n46);
   Q_reg_8_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(8), QN => n45);
   Q_reg_7_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(7), QN => n44);
   Q_reg_6_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(6), QN => n43);
   Q_reg_5_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(5), QN => n42);
   Q_reg_4_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(4), QN => n41);
   Q_reg_3_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(3), QN => n40);
   Q_reg_2_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(2), QN => n39);
   Q_reg_1_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(1), QN => n38);
   Q_reg_0_inst : DFF_X1 port map( D => n100, CK => Clk, Q => Q(0), QN => n37);
   U3 : AND2_X1 port map( A1 => n3, A2 => n36, ZN => n1);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n3);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n46, A2 => n3, B1 => n2, B2 => n4, ZN => n69);
   U7 : INV_X1 port map( A => D(9), ZN => n4);
   U8 : OAI22_X1 port map( A1 => n45, A2 => n3, B1 => n2, B2 => n5, ZN => n70);
   U9 : INV_X1 port map( A => D(8), ZN => n5);
   U10 : OAI22_X1 port map( A1 => n44, A2 => n3, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U11 : INV_X1 port map( A => D(7), ZN => n6);
   U12 : OAI22_X1 port map( A1 => n43, A2 => n3, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U13 : INV_X1 port map( A => D(6), ZN => n7);
   U14 : OAI22_X1 port map( A1 => n42, A2 => n3, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U15 : INV_X1 port map( A => D(5), ZN => n8);
   U16 : OAI22_X1 port map( A1 => n41, A2 => n3, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U17 : INV_X1 port map( A => D(4), ZN => n9);
   U18 : OAI22_X1 port map( A1 => n40, A2 => n3, B1 => n2, B2 => n10, ZN => n75
                           );
   U19 : INV_X1 port map( A => D(3), ZN => n10);
   U20 : OAI22_X1 port map( A1 => n68, A2 => n3, B1 => n2, B2 => n11, ZN => n76
                           );
   U21 : INV_X1 port map( A => D(31), ZN => n11);
   U22 : OAI22_X1 port map( A1 => n67, A2 => n3, B1 => n2, B2 => n12, ZN => n77
                           );
   U23 : INV_X1 port map( A => D(30), ZN => n12);
   U24 : OAI22_X1 port map( A1 => n39, A2 => n3, B1 => n2, B2 => n13, ZN => n78
                           );
   U25 : INV_X1 port map( A => D(2), ZN => n13);
   U26 : OAI22_X1 port map( A1 => n66, A2 => n3, B1 => n2, B2 => n14, ZN => n79
                           );
   U27 : INV_X1 port map( A => D(29), ZN => n14);
   U28 : OAI22_X1 port map( A1 => n65, A2 => n3, B1 => n2, B2 => n15, ZN => n80
                           );
   U29 : INV_X1 port map( A => D(28), ZN => n15);
   U30 : OAI22_X1 port map( A1 => n64, A2 => n3, B1 => n2, B2 => n16, ZN => n81
                           );
   U31 : INV_X1 port map( A => D(27), ZN => n16);
   U32 : OAI22_X1 port map( A1 => n63, A2 => n3, B1 => n2, B2 => n17, ZN => n82
                           );
   U33 : INV_X1 port map( A => D(26), ZN => n17);
   U34 : OAI22_X1 port map( A1 => n62, A2 => n3, B1 => n2, B2 => n18, ZN => n83
                           );
   U35 : INV_X1 port map( A => D(25), ZN => n18);
   U36 : OAI22_X1 port map( A1 => n61, A2 => n3, B1 => n2, B2 => n19, ZN => n84
                           );
   U37 : INV_X1 port map( A => D(24), ZN => n19);
   U38 : OAI22_X1 port map( A1 => n60, A2 => n3, B1 => n2, B2 => n20, ZN => n85
                           );
   U39 : INV_X1 port map( A => D(23), ZN => n20);
   U40 : OAI22_X1 port map( A1 => n59, A2 => n3, B1 => n2, B2 => n21, ZN => n86
                           );
   U41 : INV_X1 port map( A => D(22), ZN => n21);
   U42 : OAI22_X1 port map( A1 => n58, A2 => n3, B1 => n2, B2 => n22, ZN => n87
                           );
   U43 : INV_X1 port map( A => D(21), ZN => n22);
   U44 : OAI22_X1 port map( A1 => n57, A2 => n3, B1 => n2, B2 => n23, ZN => n88
                           );
   U45 : INV_X1 port map( A => D(20), ZN => n23);
   U46 : OAI22_X1 port map( A1 => n38, A2 => n3, B1 => n2, B2 => n24, ZN => n89
                           );
   U47 : INV_X1 port map( A => D(1), ZN => n24);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n3, B1 => n2, B2 => n25, ZN => n90
                           );
   U49 : INV_X1 port map( A => D(19), ZN => n25);
   U50 : OAI22_X1 port map( A1 => n55, A2 => n3, B1 => n2, B2 => n26, ZN => n91
                           );
   U51 : INV_X1 port map( A => D(18), ZN => n26);
   U52 : OAI22_X1 port map( A1 => n54, A2 => n3, B1 => n2, B2 => n27, ZN => n92
                           );
   U53 : INV_X1 port map( A => D(17), ZN => n27);
   U54 : OAI22_X1 port map( A1 => n53, A2 => n3, B1 => n2, B2 => n28, ZN => n93
                           );
   U55 : INV_X1 port map( A => D(16), ZN => n28);
   U56 : OAI22_X1 port map( A1 => n52, A2 => n3, B1 => n2, B2 => n29, ZN => n94
                           );
   U57 : INV_X1 port map( A => D(15), ZN => n29);
   U58 : OAI22_X1 port map( A1 => n51, A2 => n3, B1 => n2, B2 => n30, ZN => n95
                           );
   U59 : INV_X1 port map( A => D(14), ZN => n30);
   U60 : OAI22_X1 port map( A1 => n50, A2 => n3, B1 => n2, B2 => n31, ZN => n96
                           );
   U61 : INV_X1 port map( A => D(13), ZN => n31);
   U62 : OAI22_X1 port map( A1 => n49, A2 => n3, B1 => n2, B2 => n32, ZN => n97
                           );
   U63 : INV_X1 port map( A => D(12), ZN => n32);
   U64 : OAI22_X1 port map( A1 => n48, A2 => n3, B1 => n2, B2 => n33, ZN => n98
                           );
   U65 : INV_X1 port map( A => D(11), ZN => n33);
   U66 : OAI22_X1 port map( A1 => n47, A2 => n3, B1 => n2, B2 => n34, ZN => n99
                           );
   U67 : INV_X1 port map( A => D(10), ZN => n34);
   U68 : OAI22_X1 port map( A1 => n37, A2 => n3, B1 => n2, B2 => n35, ZN => 
                           n100);
   U69 : INV_X1 port map( A => D(0), ZN => n35);
   U70 : INV_X1 port map( A => Rst, ZN => n36);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_1 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_1;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(9), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(8), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(7), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(6), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(5), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(4), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(3), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(31), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(30), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(2), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(29), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(28), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(27), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(26), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(25), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(24), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(23), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(22), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(21), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(20), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(1), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(19), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(18), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(17), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(16), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(15), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(14), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(13), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(12), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(11), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(10), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M5_1 is

   port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector (1023 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end mux_N32_M5_1;

architecture SYN_behav of mux_N32_M5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689 : 
      std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n661, A2 => n666, ZN => n16);
   U3 : AND2_X2 port map( A1 => n661, A2 => n664, ZN => n14);
   U4 : AND2_X2 port map( A1 => n663, A2 => n665, ZN => n12);
   U5 : AND2_X2 port map( A1 => n661, A2 => n662, ZN => n10);
   U6 : AND2_X2 port map( A1 => n666, A2 => n672, ZN => n22);
   U7 : AND2_X2 port map( A1 => n680, A2 => n665, ZN => n34);
   U8 : AND2_X2 port map( A1 => n662, A2 => n673, ZN => n28);
   U9 : AND2_X2 port map( A1 => n681, A2 => n664, ZN => n40);
   U10 : AND2_X2 port map( A1 => n665, A2 => n672, ZN => n26);
   U11 : AND2_X2 port map( A1 => n675, A2 => n664, ZN => n38);
   U12 : AND2_X2 port map( A1 => n681, A2 => n666, ZN => n52);
   U13 : AND2_X2 port map( A1 => n663, A2 => n662, ZN => n15);
   U14 : AND2_X2 port map( A1 => n662, A2 => n675, ZN => n46);
   U15 : AND2_X2 port map( A1 => n665, A2 => n673, ZN => n24);
   U16 : AND2_X2 port map( A1 => n680, A2 => n664, ZN => n36);
   U17 : AND2_X2 port map( A1 => n663, A2 => n666, ZN => n11);
   U18 : AND2_X2 port map( A1 => n682, A2 => n666, ZN => n50);
   U19 : AND2_X2 port map( A1 => n680, A2 => n662, ZN => n48);
   U20 : AND2_X2 port map( A1 => n661, A2 => n665, ZN => n13);
   U21 : AND2_X2 port map( A1 => n663, A2 => n664, ZN => n9);
   U22 : AND2_X2 port map( A1 => n664, A2 => n673, ZN => n21);
   U23 : AND2_X2 port map( A1 => n662, A2 => n672, ZN => n33);
   U24 : AND2_X2 port map( A1 => n675, A2 => n666, ZN => n27);
   U25 : AND2_X2 port map( A1 => n682, A2 => n665, ZN => n39);
   U26 : AND2_X2 port map( A1 => n682, A2 => n664, ZN => n45);
   U27 : AND2_X2 port map( A1 => n666, A2 => n673, ZN => n23);
   U28 : AND2_X2 port map( A1 => n675, A2 => n665, ZN => n35);
   U29 : AND2_X2 port map( A1 => n681, A2 => n662, ZN => n51);
   U30 : AND2_X2 port map( A1 => n672, A2 => n664, ZN => n25);
   U31 : AND2_X2 port map( A1 => n680, A2 => n666, ZN => n37);
   U32 : AND2_X2 port map( A1 => n682, A2 => n662, ZN => n49);
   U33 : AND2_X2 port map( A1 => n681, A2 => n665, ZN => n47);
   U34 : OR4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => Y(9));
   U35 : NAND4_X1 port map( A1 => n5, A2 => n6, A3 => n7, A4 => n8, ZN => n4);
   U36 : AOI22_X1 port map( A1 => Q(105), A2 => n9, B1 => Q(201), B2 => n10, ZN
                           => n8);
   U37 : AOI22_X1 port map( A1 => Q(169), A2 => n11, B1 => Q(41), B2 => n12, ZN
                           => n7);
   U38 : AOI22_X1 port map( A1 => Q(9), A2 => n13, B1 => Q(73), B2 => n14, ZN 
                           => n6);
   U39 : AOI22_X1 port map( A1 => Q(233), A2 => n15, B1 => Q(137), B2 => n16, 
                           ZN => n5);
   U40 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           n3);
   U41 : AOI22_X1 port map( A1 => Q(329), A2 => n21, B1 => Q(425), B2 => n22, 
                           ZN => n20);
   U42 : AOI22_X1 port map( A1 => Q(393), A2 => n23, B1 => Q(265), B2 => n24, 
                           ZN => n19);
   U43 : AOI22_X1 port map( A1 => Q(361), A2 => n25, B1 => Q(297), B2 => n26, 
                           ZN => n18);
   U44 : AOI22_X1 port map( A1 => Q(649), A2 => n27, B1 => Q(457), B2 => n28, 
                           ZN => n17);
   U45 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           n2);
   U46 : AOI22_X1 port map( A1 => Q(489), A2 => n33, B1 => Q(553), B2 => n34, 
                           ZN => n32);
   U47 : AOI22_X1 port map( A1 => Q(521), A2 => n35, B1 => Q(617), B2 => n36, 
                           ZN => n31);
   U48 : AOI22_X1 port map( A1 => Q(681), A2 => n37, B1 => Q(585), B2 => n38, 
                           ZN => n30);
   U49 : AOI22_X1 port map( A1 => Q(777), A2 => n39, B1 => Q(873), B2 => n40, 
                           ZN => n29);
   U50 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           n1);
   U51 : AOI22_X1 port map( A1 => Q(841), A2 => n45, B1 => Q(713), B2 => n46, 
                           ZN => n44);
   U52 : AOI22_X1 port map( A1 => Q(809), A2 => n47, B1 => Q(745), B2 => n48, 
                           ZN => n43);
   U53 : AOI22_X1 port map( A1 => Q(969), A2 => n49, B1 => Q(905), B2 => n50, 
                           ZN => n42);
   U54 : AOI22_X1 port map( A1 => Q(1001), A2 => n51, B1 => Q(937), B2 => n52, 
                           ZN => n41);
   U55 : OR4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           Y(8));
   U56 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n56);
   U57 : AOI22_X1 port map( A1 => Q(104), A2 => n9, B1 => Q(200), B2 => n10, ZN
                           => n60);
   U58 : AOI22_X1 port map( A1 => Q(168), A2 => n11, B1 => Q(40), B2 => n12, ZN
                           => n59);
   U59 : AOI22_X1 port map( A1 => Q(8), A2 => n13, B1 => Q(72), B2 => n14, ZN 
                           => n58);
   U60 : AOI22_X1 port map( A1 => Q(232), A2 => n15, B1 => Q(136), B2 => n16, 
                           ZN => n57);
   U61 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           n55);
   U62 : AOI22_X1 port map( A1 => Q(328), A2 => n21, B1 => Q(424), B2 => n22, 
                           ZN => n64);
   U63 : AOI22_X1 port map( A1 => Q(392), A2 => n23, B1 => Q(264), B2 => n24, 
                           ZN => n63);
   U64 : AOI22_X1 port map( A1 => Q(360), A2 => n25, B1 => Q(296), B2 => n26, 
                           ZN => n62);
   U65 : AOI22_X1 port map( A1 => Q(648), A2 => n27, B1 => Q(456), B2 => n28, 
                           ZN => n61);
   U66 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           n54);
   U67 : AOI22_X1 port map( A1 => Q(488), A2 => n33, B1 => Q(552), B2 => n34, 
                           ZN => n68);
   U68 : AOI22_X1 port map( A1 => Q(520), A2 => n35, B1 => Q(616), B2 => n36, 
                           ZN => n67);
   U69 : AOI22_X1 port map( A1 => Q(680), A2 => n37, B1 => Q(584), B2 => n38, 
                           ZN => n66);
   U70 : AOI22_X1 port map( A1 => Q(776), A2 => n39, B1 => Q(872), B2 => n40, 
                           ZN => n65);
   U71 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n53);
   U72 : AOI22_X1 port map( A1 => Q(840), A2 => n45, B1 => Q(712), B2 => n46, 
                           ZN => n72);
   U73 : AOI22_X1 port map( A1 => Q(808), A2 => n47, B1 => Q(744), B2 => n48, 
                           ZN => n71);
   U74 : AOI22_X1 port map( A1 => Q(968), A2 => n49, B1 => Q(904), B2 => n50, 
                           ZN => n70);
   U75 : AOI22_X1 port map( A1 => Q(1000), A2 => n51, B1 => Q(936), B2 => n52, 
                           ZN => n69);
   U76 : OR4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           Y(7));
   U77 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           n76);
   U78 : AOI22_X1 port map( A1 => Q(103), A2 => n9, B1 => Q(199), B2 => n10, ZN
                           => n80);
   U79 : AOI22_X1 port map( A1 => Q(167), A2 => n11, B1 => Q(39), B2 => n12, ZN
                           => n79);
   U80 : AOI22_X1 port map( A1 => Q(7), A2 => n13, B1 => Q(71), B2 => n14, ZN 
                           => n78);
   U81 : AOI22_X1 port map( A1 => Q(231), A2 => n15, B1 => Q(135), B2 => n16, 
                           ZN => n77);
   U82 : NAND4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           n75);
   U83 : AOI22_X1 port map( A1 => Q(327), A2 => n21, B1 => Q(423), B2 => n22, 
                           ZN => n84);
   U84 : AOI22_X1 port map( A1 => Q(391), A2 => n23, B1 => Q(263), B2 => n24, 
                           ZN => n83);
   U85 : AOI22_X1 port map( A1 => Q(359), A2 => n25, B1 => Q(295), B2 => n26, 
                           ZN => n82);
   U86 : AOI22_X1 port map( A1 => Q(647), A2 => n27, B1 => Q(455), B2 => n28, 
                           ZN => n81);
   U87 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           n74);
   U88 : AOI22_X1 port map( A1 => Q(487), A2 => n33, B1 => Q(551), B2 => n34, 
                           ZN => n88);
   U89 : AOI22_X1 port map( A1 => Q(519), A2 => n35, B1 => Q(615), B2 => n36, 
                           ZN => n87);
   U90 : AOI22_X1 port map( A1 => Q(679), A2 => n37, B1 => Q(583), B2 => n38, 
                           ZN => n86);
   U91 : AOI22_X1 port map( A1 => Q(775), A2 => n39, B1 => Q(871), B2 => n40, 
                           ZN => n85);
   U92 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           n73);
   U93 : AOI22_X1 port map( A1 => Q(839), A2 => n45, B1 => Q(711), B2 => n46, 
                           ZN => n92);
   U94 : AOI22_X1 port map( A1 => Q(807), A2 => n47, B1 => Q(743), B2 => n48, 
                           ZN => n91);
   U95 : AOI22_X1 port map( A1 => Q(967), A2 => n49, B1 => Q(903), B2 => n50, 
                           ZN => n90);
   U96 : AOI22_X1 port map( A1 => Q(999), A2 => n51, B1 => Q(935), B2 => n52, 
                           ZN => n89);
   U97 : OR4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           Y(6));
   U98 : NAND4_X1 port map( A1 => n97, A2 => n98, A3 => n99, A4 => n100, ZN => 
                           n96);
   U99 : AOI22_X1 port map( A1 => Q(102), A2 => n9, B1 => Q(198), B2 => n10, ZN
                           => n100);
   U100 : AOI22_X1 port map( A1 => Q(166), A2 => n11, B1 => Q(38), B2 => n12, 
                           ZN => n99);
   U101 : AOI22_X1 port map( A1 => Q(6), A2 => n13, B1 => Q(70), B2 => n14, ZN 
                           => n98);
   U102 : AOI22_X1 port map( A1 => Q(230), A2 => n15, B1 => Q(134), B2 => n16, 
                           ZN => n97);
   U103 : NAND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN
                           => n95);
   U104 : AOI22_X1 port map( A1 => Q(326), A2 => n21, B1 => Q(422), B2 => n22, 
                           ZN => n104);
   U105 : AOI22_X1 port map( A1 => Q(390), A2 => n23, B1 => Q(262), B2 => n24, 
                           ZN => n103);
   U106 : AOI22_X1 port map( A1 => Q(358), A2 => n25, B1 => Q(294), B2 => n26, 
                           ZN => n102);
   U107 : AOI22_X1 port map( A1 => Q(646), A2 => n27, B1 => Q(454), B2 => n28, 
                           ZN => n101);
   U108 : NAND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN
                           => n94);
   U109 : AOI22_X1 port map( A1 => Q(486), A2 => n33, B1 => Q(550), B2 => n34, 
                           ZN => n108);
   U110 : AOI22_X1 port map( A1 => Q(518), A2 => n35, B1 => Q(614), B2 => n36, 
                           ZN => n107);
   U111 : AOI22_X1 port map( A1 => Q(678), A2 => n37, B1 => Q(582), B2 => n38, 
                           ZN => n106);
   U112 : AOI22_X1 port map( A1 => Q(774), A2 => n39, B1 => Q(870), B2 => n40, 
                           ZN => n105);
   U113 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => n93);
   U114 : AOI22_X1 port map( A1 => Q(838), A2 => n45, B1 => Q(710), B2 => n46, 
                           ZN => n112);
   U115 : AOI22_X1 port map( A1 => Q(806), A2 => n47, B1 => Q(742), B2 => n48, 
                           ZN => n111);
   U116 : AOI22_X1 port map( A1 => Q(966), A2 => n49, B1 => Q(902), B2 => n50, 
                           ZN => n110);
   U117 : AOI22_X1 port map( A1 => Q(998), A2 => n51, B1 => Q(934), B2 => n52, 
                           ZN => n109);
   U118 : OR4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN 
                           => Y(5));
   U119 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN
                           => n116);
   U120 : AOI22_X1 port map( A1 => Q(101), A2 => n9, B1 => Q(197), B2 => n10, 
                           ZN => n120);
   U121 : AOI22_X1 port map( A1 => Q(165), A2 => n11, B1 => Q(37), B2 => n12, 
                           ZN => n119);
   U122 : AOI22_X1 port map( A1 => Q(5), A2 => n13, B1 => Q(69), B2 => n14, ZN 
                           => n118);
   U123 : AOI22_X1 port map( A1 => Q(229), A2 => n15, B1 => Q(133), B2 => n16, 
                           ZN => n117);
   U124 : NAND4_X1 port map( A1 => n121, A2 => n122, A3 => n123, A4 => n124, ZN
                           => n115);
   U125 : AOI22_X1 port map( A1 => Q(325), A2 => n21, B1 => Q(421), B2 => n22, 
                           ZN => n124);
   U126 : AOI22_X1 port map( A1 => Q(389), A2 => n23, B1 => Q(261), B2 => n24, 
                           ZN => n123);
   U127 : AOI22_X1 port map( A1 => Q(357), A2 => n25, B1 => Q(293), B2 => n26, 
                           ZN => n122);
   U128 : AOI22_X1 port map( A1 => Q(645), A2 => n27, B1 => Q(453), B2 => n28, 
                           ZN => n121);
   U129 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => n114);
   U130 : AOI22_X1 port map( A1 => Q(485), A2 => n33, B1 => Q(549), B2 => n34, 
                           ZN => n128);
   U131 : AOI22_X1 port map( A1 => Q(517), A2 => n35, B1 => Q(613), B2 => n36, 
                           ZN => n127);
   U132 : AOI22_X1 port map( A1 => Q(677), A2 => n37, B1 => Q(581), B2 => n38, 
                           ZN => n126);
   U133 : AOI22_X1 port map( A1 => Q(773), A2 => n39, B1 => Q(869), B2 => n40, 
                           ZN => n125);
   U134 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => n113);
   U135 : AOI22_X1 port map( A1 => Q(837), A2 => n45, B1 => Q(709), B2 => n46, 
                           ZN => n132);
   U136 : AOI22_X1 port map( A1 => Q(805), A2 => n47, B1 => Q(741), B2 => n48, 
                           ZN => n131);
   U137 : AOI22_X1 port map( A1 => Q(965), A2 => n49, B1 => Q(901), B2 => n50, 
                           ZN => n130);
   U138 : AOI22_X1 port map( A1 => Q(997), A2 => n51, B1 => Q(933), B2 => n52, 
                           ZN => n129);
   U139 : OR4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN 
                           => Y(4));
   U140 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => n136);
   U141 : AOI22_X1 port map( A1 => Q(100), A2 => n9, B1 => Q(196), B2 => n10, 
                           ZN => n140);
   U142 : AOI22_X1 port map( A1 => Q(164), A2 => n11, B1 => Q(36), B2 => n12, 
                           ZN => n139);
   U143 : AOI22_X1 port map( A1 => Q(4), A2 => n13, B1 => Q(68), B2 => n14, ZN 
                           => n138);
   U144 : AOI22_X1 port map( A1 => Q(228), A2 => n15, B1 => Q(132), B2 => n16, 
                           ZN => n137);
   U145 : NAND4_X1 port map( A1 => n141, A2 => n142, A3 => n143, A4 => n144, ZN
                           => n135);
   U146 : AOI22_X1 port map( A1 => Q(324), A2 => n21, B1 => Q(420), B2 => n22, 
                           ZN => n144);
   U147 : AOI22_X1 port map( A1 => Q(388), A2 => n23, B1 => Q(260), B2 => n24, 
                           ZN => n143);
   U148 : AOI22_X1 port map( A1 => Q(356), A2 => n25, B1 => Q(292), B2 => n26, 
                           ZN => n142);
   U149 : AOI22_X1 port map( A1 => Q(644), A2 => n27, B1 => Q(452), B2 => n28, 
                           ZN => n141);
   U150 : NAND4_X1 port map( A1 => n145, A2 => n146, A3 => n147, A4 => n148, ZN
                           => n134);
   U151 : AOI22_X1 port map( A1 => Q(484), A2 => n33, B1 => Q(548), B2 => n34, 
                           ZN => n148);
   U152 : AOI22_X1 port map( A1 => Q(516), A2 => n35, B1 => Q(612), B2 => n36, 
                           ZN => n147);
   U153 : AOI22_X1 port map( A1 => Q(676), A2 => n37, B1 => Q(580), B2 => n38, 
                           ZN => n146);
   U154 : AOI22_X1 port map( A1 => Q(772), A2 => n39, B1 => Q(868), B2 => n40, 
                           ZN => n145);
   U155 : NAND4_X1 port map( A1 => n149, A2 => n150, A3 => n151, A4 => n152, ZN
                           => n133);
   U156 : AOI22_X1 port map( A1 => Q(836), A2 => n45, B1 => Q(708), B2 => n46, 
                           ZN => n152);
   U157 : AOI22_X1 port map( A1 => Q(804), A2 => n47, B1 => Q(740), B2 => n48, 
                           ZN => n151);
   U158 : AOI22_X1 port map( A1 => Q(964), A2 => n49, B1 => Q(900), B2 => n50, 
                           ZN => n150);
   U159 : AOI22_X1 port map( A1 => Q(996), A2 => n51, B1 => Q(932), B2 => n52, 
                           ZN => n149);
   U160 : OR4_X1 port map( A1 => n153, A2 => n154, A3 => n155, A4 => n156, ZN 
                           => Y(3));
   U161 : NAND4_X1 port map( A1 => n157, A2 => n158, A3 => n159, A4 => n160, ZN
                           => n156);
   U162 : AOI22_X1 port map( A1 => Q(99), A2 => n9, B1 => Q(195), B2 => n10, ZN
                           => n160);
   U163 : AOI22_X1 port map( A1 => Q(163), A2 => n11, B1 => Q(35), B2 => n12, 
                           ZN => n159);
   U164 : AOI22_X1 port map( A1 => Q(3), A2 => n13, B1 => Q(67), B2 => n14, ZN 
                           => n158);
   U165 : AOI22_X1 port map( A1 => Q(227), A2 => n15, B1 => Q(131), B2 => n16, 
                           ZN => n157);
   U166 : NAND4_X1 port map( A1 => n161, A2 => n162, A3 => n163, A4 => n164, ZN
                           => n155);
   U167 : AOI22_X1 port map( A1 => Q(323), A2 => n21, B1 => Q(419), B2 => n22, 
                           ZN => n164);
   U168 : AOI22_X1 port map( A1 => Q(387), A2 => n23, B1 => Q(259), B2 => n24, 
                           ZN => n163);
   U169 : AOI22_X1 port map( A1 => Q(355), A2 => n25, B1 => Q(291), B2 => n26, 
                           ZN => n162);
   U170 : AOI22_X1 port map( A1 => Q(643), A2 => n27, B1 => Q(451), B2 => n28, 
                           ZN => n161);
   U171 : NAND4_X1 port map( A1 => n165, A2 => n166, A3 => n167, A4 => n168, ZN
                           => n154);
   U172 : AOI22_X1 port map( A1 => Q(483), A2 => n33, B1 => Q(547), B2 => n34, 
                           ZN => n168);
   U173 : AOI22_X1 port map( A1 => Q(515), A2 => n35, B1 => Q(611), B2 => n36, 
                           ZN => n167);
   U174 : AOI22_X1 port map( A1 => Q(675), A2 => n37, B1 => Q(579), B2 => n38, 
                           ZN => n166);
   U175 : AOI22_X1 port map( A1 => Q(771), A2 => n39, B1 => Q(867), B2 => n40, 
                           ZN => n165);
   U176 : NAND4_X1 port map( A1 => n169, A2 => n170, A3 => n171, A4 => n172, ZN
                           => n153);
   U177 : AOI22_X1 port map( A1 => Q(835), A2 => n45, B1 => Q(707), B2 => n46, 
                           ZN => n172);
   U178 : AOI22_X1 port map( A1 => Q(803), A2 => n47, B1 => Q(739), B2 => n48, 
                           ZN => n171);
   U179 : AOI22_X1 port map( A1 => Q(963), A2 => n49, B1 => Q(899), B2 => n50, 
                           ZN => n170);
   U180 : AOI22_X1 port map( A1 => Q(995), A2 => n51, B1 => Q(931), B2 => n52, 
                           ZN => n169);
   U181 : OR4_X1 port map( A1 => n173, A2 => n174, A3 => n175, A4 => n176, ZN 
                           => Y(31));
   U182 : NAND4_X1 port map( A1 => n177, A2 => n178, A3 => n179, A4 => n180, ZN
                           => n176);
   U183 : AOI22_X1 port map( A1 => Q(127), A2 => n9, B1 => Q(223), B2 => n10, 
                           ZN => n180);
   U184 : AOI22_X1 port map( A1 => Q(191), A2 => n11, B1 => Q(63), B2 => n12, 
                           ZN => n179);
   U185 : AOI22_X1 port map( A1 => Q(31), A2 => n13, B1 => Q(95), B2 => n14, ZN
                           => n178);
   U186 : AOI22_X1 port map( A1 => Q(255), A2 => n15, B1 => Q(159), B2 => n16, 
                           ZN => n177);
   U187 : NAND4_X1 port map( A1 => n181, A2 => n182, A3 => n183, A4 => n184, ZN
                           => n175);
   U188 : AOI22_X1 port map( A1 => Q(351), A2 => n21, B1 => Q(447), B2 => n22, 
                           ZN => n184);
   U189 : AOI22_X1 port map( A1 => Q(415), A2 => n23, B1 => Q(287), B2 => n24, 
                           ZN => n183);
   U190 : AOI22_X1 port map( A1 => Q(383), A2 => n25, B1 => Q(319), B2 => n26, 
                           ZN => n182);
   U191 : AOI22_X1 port map( A1 => Q(671), A2 => n27, B1 => Q(479), B2 => n28, 
                           ZN => n181);
   U192 : NAND4_X1 port map( A1 => n185, A2 => n186, A3 => n187, A4 => n188, ZN
                           => n174);
   U193 : AOI22_X1 port map( A1 => Q(511), A2 => n33, B1 => Q(575), B2 => n34, 
                           ZN => n188);
   U194 : AOI22_X1 port map( A1 => Q(543), A2 => n35, B1 => Q(639), B2 => n36, 
                           ZN => n187);
   U195 : AOI22_X1 port map( A1 => Q(703), A2 => n37, B1 => Q(607), B2 => n38, 
                           ZN => n186);
   U196 : AOI22_X1 port map( A1 => Q(799), A2 => n39, B1 => Q(895), B2 => n40, 
                           ZN => n185);
   U197 : NAND4_X1 port map( A1 => n189, A2 => n190, A3 => n191, A4 => n192, ZN
                           => n173);
   U198 : AOI22_X1 port map( A1 => Q(863), A2 => n45, B1 => Q(735), B2 => n46, 
                           ZN => n192);
   U199 : AOI22_X1 port map( A1 => Q(831), A2 => n47, B1 => Q(767), B2 => n48, 
                           ZN => n191);
   U200 : AOI22_X1 port map( A1 => Q(991), A2 => n49, B1 => Q(927), B2 => n50, 
                           ZN => n190);
   U201 : AOI22_X1 port map( A1 => Q(1023), A2 => n51, B1 => Q(959), B2 => n52,
                           ZN => n189);
   U202 : OR4_X1 port map( A1 => n193, A2 => n194, A3 => n195, A4 => n196, ZN 
                           => Y(30));
   U203 : NAND4_X1 port map( A1 => n197, A2 => n198, A3 => n199, A4 => n200, ZN
                           => n196);
   U204 : AOI22_X1 port map( A1 => Q(126), A2 => n9, B1 => Q(222), B2 => n10, 
                           ZN => n200);
   U205 : AOI22_X1 port map( A1 => Q(190), A2 => n11, B1 => Q(62), B2 => n12, 
                           ZN => n199);
   U206 : AOI22_X1 port map( A1 => Q(30), A2 => n13, B1 => Q(94), B2 => n14, ZN
                           => n198);
   U207 : AOI22_X1 port map( A1 => Q(254), A2 => n15, B1 => Q(158), B2 => n16, 
                           ZN => n197);
   U208 : NAND4_X1 port map( A1 => n201, A2 => n202, A3 => n203, A4 => n204, ZN
                           => n195);
   U209 : AOI22_X1 port map( A1 => Q(350), A2 => n21, B1 => Q(446), B2 => n22, 
                           ZN => n204);
   U210 : AOI22_X1 port map( A1 => Q(414), A2 => n23, B1 => Q(286), B2 => n24, 
                           ZN => n203);
   U211 : AOI22_X1 port map( A1 => Q(382), A2 => n25, B1 => Q(318), B2 => n26, 
                           ZN => n202);
   U212 : AOI22_X1 port map( A1 => Q(670), A2 => n27, B1 => Q(478), B2 => n28, 
                           ZN => n201);
   U213 : NAND4_X1 port map( A1 => n205, A2 => n206, A3 => n207, A4 => n208, ZN
                           => n194);
   U214 : AOI22_X1 port map( A1 => Q(510), A2 => n33, B1 => Q(574), B2 => n34, 
                           ZN => n208);
   U215 : AOI22_X1 port map( A1 => Q(542), A2 => n35, B1 => Q(638), B2 => n36, 
                           ZN => n207);
   U216 : AOI22_X1 port map( A1 => Q(702), A2 => n37, B1 => Q(606), B2 => n38, 
                           ZN => n206);
   U217 : AOI22_X1 port map( A1 => Q(798), A2 => n39, B1 => Q(894), B2 => n40, 
                           ZN => n205);
   U218 : NAND4_X1 port map( A1 => n209, A2 => n210, A3 => n211, A4 => n212, ZN
                           => n193);
   U219 : AOI22_X1 port map( A1 => Q(862), A2 => n45, B1 => Q(734), B2 => n46, 
                           ZN => n212);
   U220 : AOI22_X1 port map( A1 => Q(830), A2 => n47, B1 => Q(766), B2 => n48, 
                           ZN => n211);
   U221 : AOI22_X1 port map( A1 => Q(990), A2 => n49, B1 => Q(926), B2 => n50, 
                           ZN => n210);
   U222 : AOI22_X1 port map( A1 => Q(1022), A2 => n51, B1 => Q(958), B2 => n52,
                           ZN => n209);
   U223 : OR4_X1 port map( A1 => n213, A2 => n214, A3 => n215, A4 => n216, ZN 
                           => Y(2));
   U224 : NAND4_X1 port map( A1 => n217, A2 => n218, A3 => n219, A4 => n220, ZN
                           => n216);
   U225 : AOI22_X1 port map( A1 => Q(98), A2 => n9, B1 => Q(194), B2 => n10, ZN
                           => n220);
   U226 : AOI22_X1 port map( A1 => Q(162), A2 => n11, B1 => Q(34), B2 => n12, 
                           ZN => n219);
   U227 : AOI22_X1 port map( A1 => Q(2), A2 => n13, B1 => Q(66), B2 => n14, ZN 
                           => n218);
   U228 : AOI22_X1 port map( A1 => Q(226), A2 => n15, B1 => Q(130), B2 => n16, 
                           ZN => n217);
   U229 : NAND4_X1 port map( A1 => n221, A2 => n222, A3 => n223, A4 => n224, ZN
                           => n215);
   U230 : AOI22_X1 port map( A1 => Q(322), A2 => n21, B1 => Q(418), B2 => n22, 
                           ZN => n224);
   U231 : AOI22_X1 port map( A1 => Q(386), A2 => n23, B1 => Q(258), B2 => n24, 
                           ZN => n223);
   U232 : AOI22_X1 port map( A1 => Q(354), A2 => n25, B1 => Q(290), B2 => n26, 
                           ZN => n222);
   U233 : AOI22_X1 port map( A1 => Q(642), A2 => n27, B1 => Q(450), B2 => n28, 
                           ZN => n221);
   U234 : NAND4_X1 port map( A1 => n225, A2 => n226, A3 => n227, A4 => n228, ZN
                           => n214);
   U235 : AOI22_X1 port map( A1 => Q(482), A2 => n33, B1 => Q(546), B2 => n34, 
                           ZN => n228);
   U236 : AOI22_X1 port map( A1 => Q(514), A2 => n35, B1 => Q(610), B2 => n36, 
                           ZN => n227);
   U237 : AOI22_X1 port map( A1 => Q(674), A2 => n37, B1 => Q(578), B2 => n38, 
                           ZN => n226);
   U238 : AOI22_X1 port map( A1 => Q(770), A2 => n39, B1 => Q(866), B2 => n40, 
                           ZN => n225);
   U239 : NAND4_X1 port map( A1 => n229, A2 => n230, A3 => n231, A4 => n232, ZN
                           => n213);
   U240 : AOI22_X1 port map( A1 => Q(834), A2 => n45, B1 => Q(706), B2 => n46, 
                           ZN => n232);
   U241 : AOI22_X1 port map( A1 => Q(802), A2 => n47, B1 => Q(738), B2 => n48, 
                           ZN => n231);
   U242 : AOI22_X1 port map( A1 => Q(962), A2 => n49, B1 => Q(898), B2 => n50, 
                           ZN => n230);
   U243 : AOI22_X1 port map( A1 => Q(994), A2 => n51, B1 => Q(930), B2 => n52, 
                           ZN => n229);
   U244 : OR4_X1 port map( A1 => n233, A2 => n234, A3 => n235, A4 => n236, ZN 
                           => Y(29));
   U245 : NAND4_X1 port map( A1 => n237, A2 => n238, A3 => n239, A4 => n240, ZN
                           => n236);
   U246 : AOI22_X1 port map( A1 => Q(125), A2 => n9, B1 => Q(221), B2 => n10, 
                           ZN => n240);
   U247 : AOI22_X1 port map( A1 => Q(189), A2 => n11, B1 => Q(61), B2 => n12, 
                           ZN => n239);
   U248 : AOI22_X1 port map( A1 => Q(29), A2 => n13, B1 => Q(93), B2 => n14, ZN
                           => n238);
   U249 : AOI22_X1 port map( A1 => Q(253), A2 => n15, B1 => Q(157), B2 => n16, 
                           ZN => n237);
   U250 : NAND4_X1 port map( A1 => n241, A2 => n242, A3 => n243, A4 => n244, ZN
                           => n235);
   U251 : AOI22_X1 port map( A1 => Q(349), A2 => n21, B1 => Q(445), B2 => n22, 
                           ZN => n244);
   U252 : AOI22_X1 port map( A1 => Q(413), A2 => n23, B1 => Q(285), B2 => n24, 
                           ZN => n243);
   U253 : AOI22_X1 port map( A1 => Q(381), A2 => n25, B1 => Q(317), B2 => n26, 
                           ZN => n242);
   U254 : AOI22_X1 port map( A1 => Q(669), A2 => n27, B1 => Q(477), B2 => n28, 
                           ZN => n241);
   U255 : NAND4_X1 port map( A1 => n245, A2 => n246, A3 => n247, A4 => n248, ZN
                           => n234);
   U256 : AOI22_X1 port map( A1 => Q(509), A2 => n33, B1 => Q(573), B2 => n34, 
                           ZN => n248);
   U257 : AOI22_X1 port map( A1 => Q(541), A2 => n35, B1 => Q(637), B2 => n36, 
                           ZN => n247);
   U258 : AOI22_X1 port map( A1 => Q(701), A2 => n37, B1 => Q(605), B2 => n38, 
                           ZN => n246);
   U259 : AOI22_X1 port map( A1 => Q(797), A2 => n39, B1 => Q(893), B2 => n40, 
                           ZN => n245);
   U260 : NAND4_X1 port map( A1 => n249, A2 => n250, A3 => n251, A4 => n252, ZN
                           => n233);
   U261 : AOI22_X1 port map( A1 => Q(861), A2 => n45, B1 => Q(733), B2 => n46, 
                           ZN => n252);
   U262 : AOI22_X1 port map( A1 => Q(829), A2 => n47, B1 => Q(765), B2 => n48, 
                           ZN => n251);
   U263 : AOI22_X1 port map( A1 => Q(989), A2 => n49, B1 => Q(925), B2 => n50, 
                           ZN => n250);
   U264 : AOI22_X1 port map( A1 => Q(1021), A2 => n51, B1 => Q(957), B2 => n52,
                           ZN => n249);
   U265 : OR4_X1 port map( A1 => n253, A2 => n254, A3 => n255, A4 => n256, ZN 
                           => Y(28));
   U266 : NAND4_X1 port map( A1 => n257, A2 => n258, A3 => n259, A4 => n260, ZN
                           => n256);
   U267 : AOI22_X1 port map( A1 => Q(124), A2 => n9, B1 => Q(220), B2 => n10, 
                           ZN => n260);
   U268 : AOI22_X1 port map( A1 => Q(188), A2 => n11, B1 => Q(60), B2 => n12, 
                           ZN => n259);
   U269 : AOI22_X1 port map( A1 => Q(28), A2 => n13, B1 => Q(92), B2 => n14, ZN
                           => n258);
   U270 : AOI22_X1 port map( A1 => Q(252), A2 => n15, B1 => Q(156), B2 => n16, 
                           ZN => n257);
   U271 : NAND4_X1 port map( A1 => n261, A2 => n262, A3 => n263, A4 => n264, ZN
                           => n255);
   U272 : AOI22_X1 port map( A1 => Q(348), A2 => n21, B1 => Q(444), B2 => n22, 
                           ZN => n264);
   U273 : AOI22_X1 port map( A1 => Q(412), A2 => n23, B1 => Q(284), B2 => n24, 
                           ZN => n263);
   U274 : AOI22_X1 port map( A1 => Q(380), A2 => n25, B1 => Q(316), B2 => n26, 
                           ZN => n262);
   U275 : AOI22_X1 port map( A1 => Q(668), A2 => n27, B1 => Q(476), B2 => n28, 
                           ZN => n261);
   U276 : NAND4_X1 port map( A1 => n265, A2 => n266, A3 => n267, A4 => n268, ZN
                           => n254);
   U277 : AOI22_X1 port map( A1 => Q(508), A2 => n33, B1 => Q(572), B2 => n34, 
                           ZN => n268);
   U278 : AOI22_X1 port map( A1 => Q(540), A2 => n35, B1 => Q(636), B2 => n36, 
                           ZN => n267);
   U279 : AOI22_X1 port map( A1 => Q(700), A2 => n37, B1 => Q(604), B2 => n38, 
                           ZN => n266);
   U280 : AOI22_X1 port map( A1 => Q(796), A2 => n39, B1 => Q(892), B2 => n40, 
                           ZN => n265);
   U281 : NAND4_X1 port map( A1 => n269, A2 => n270, A3 => n271, A4 => n272, ZN
                           => n253);
   U282 : AOI22_X1 port map( A1 => Q(860), A2 => n45, B1 => Q(732), B2 => n46, 
                           ZN => n272);
   U283 : AOI22_X1 port map( A1 => Q(828), A2 => n47, B1 => Q(764), B2 => n48, 
                           ZN => n271);
   U284 : AOI22_X1 port map( A1 => Q(988), A2 => n49, B1 => Q(924), B2 => n50, 
                           ZN => n270);
   U285 : AOI22_X1 port map( A1 => Q(1020), A2 => n51, B1 => Q(956), B2 => n52,
                           ZN => n269);
   U286 : OR4_X1 port map( A1 => n273, A2 => n274, A3 => n275, A4 => n276, ZN 
                           => Y(27));
   U287 : NAND4_X1 port map( A1 => n277, A2 => n278, A3 => n279, A4 => n280, ZN
                           => n276);
   U288 : AOI22_X1 port map( A1 => Q(123), A2 => n9, B1 => Q(219), B2 => n10, 
                           ZN => n280);
   U289 : AOI22_X1 port map( A1 => Q(187), A2 => n11, B1 => Q(59), B2 => n12, 
                           ZN => n279);
   U290 : AOI22_X1 port map( A1 => Q(27), A2 => n13, B1 => Q(91), B2 => n14, ZN
                           => n278);
   U291 : AOI22_X1 port map( A1 => Q(251), A2 => n15, B1 => Q(155), B2 => n16, 
                           ZN => n277);
   U292 : NAND4_X1 port map( A1 => n281, A2 => n282, A3 => n283, A4 => n284, ZN
                           => n275);
   U293 : AOI22_X1 port map( A1 => Q(347), A2 => n21, B1 => Q(443), B2 => n22, 
                           ZN => n284);
   U294 : AOI22_X1 port map( A1 => Q(411), A2 => n23, B1 => Q(283), B2 => n24, 
                           ZN => n283);
   U295 : AOI22_X1 port map( A1 => Q(379), A2 => n25, B1 => Q(315), B2 => n26, 
                           ZN => n282);
   U296 : AOI22_X1 port map( A1 => Q(667), A2 => n27, B1 => Q(475), B2 => n28, 
                           ZN => n281);
   U297 : NAND4_X1 port map( A1 => n285, A2 => n286, A3 => n287, A4 => n288, ZN
                           => n274);
   U298 : AOI22_X1 port map( A1 => Q(507), A2 => n33, B1 => Q(571), B2 => n34, 
                           ZN => n288);
   U299 : AOI22_X1 port map( A1 => Q(539), A2 => n35, B1 => Q(635), B2 => n36, 
                           ZN => n287);
   U300 : AOI22_X1 port map( A1 => Q(699), A2 => n37, B1 => Q(603), B2 => n38, 
                           ZN => n286);
   U301 : AOI22_X1 port map( A1 => Q(795), A2 => n39, B1 => Q(891), B2 => n40, 
                           ZN => n285);
   U302 : NAND4_X1 port map( A1 => n289, A2 => n290, A3 => n291, A4 => n292, ZN
                           => n273);
   U303 : AOI22_X1 port map( A1 => Q(859), A2 => n45, B1 => Q(731), B2 => n46, 
                           ZN => n292);
   U304 : AOI22_X1 port map( A1 => Q(827), A2 => n47, B1 => Q(763), B2 => n48, 
                           ZN => n291);
   U305 : AOI22_X1 port map( A1 => Q(987), A2 => n49, B1 => Q(923), B2 => n50, 
                           ZN => n290);
   U306 : AOI22_X1 port map( A1 => Q(1019), A2 => n51, B1 => Q(955), B2 => n52,
                           ZN => n289);
   U307 : OR4_X1 port map( A1 => n293, A2 => n294, A3 => n295, A4 => n296, ZN 
                           => Y(26));
   U308 : NAND4_X1 port map( A1 => n297, A2 => n298, A3 => n299, A4 => n300, ZN
                           => n296);
   U309 : AOI22_X1 port map( A1 => Q(122), A2 => n9, B1 => Q(218), B2 => n10, 
                           ZN => n300);
   U310 : AOI22_X1 port map( A1 => Q(186), A2 => n11, B1 => Q(58), B2 => n12, 
                           ZN => n299);
   U311 : AOI22_X1 port map( A1 => Q(26), A2 => n13, B1 => Q(90), B2 => n14, ZN
                           => n298);
   U312 : AOI22_X1 port map( A1 => Q(250), A2 => n15, B1 => Q(154), B2 => n16, 
                           ZN => n297);
   U313 : NAND4_X1 port map( A1 => n301, A2 => n302, A3 => n303, A4 => n304, ZN
                           => n295);
   U314 : AOI22_X1 port map( A1 => Q(346), A2 => n21, B1 => Q(442), B2 => n22, 
                           ZN => n304);
   U315 : AOI22_X1 port map( A1 => Q(410), A2 => n23, B1 => Q(282), B2 => n24, 
                           ZN => n303);
   U316 : AOI22_X1 port map( A1 => Q(378), A2 => n25, B1 => Q(314), B2 => n26, 
                           ZN => n302);
   U317 : AOI22_X1 port map( A1 => Q(666), A2 => n27, B1 => Q(474), B2 => n28, 
                           ZN => n301);
   U318 : NAND4_X1 port map( A1 => n305, A2 => n306, A3 => n307, A4 => n308, ZN
                           => n294);
   U319 : AOI22_X1 port map( A1 => Q(506), A2 => n33, B1 => Q(570), B2 => n34, 
                           ZN => n308);
   U320 : AOI22_X1 port map( A1 => Q(538), A2 => n35, B1 => Q(634), B2 => n36, 
                           ZN => n307);
   U321 : AOI22_X1 port map( A1 => Q(698), A2 => n37, B1 => Q(602), B2 => n38, 
                           ZN => n306);
   U322 : AOI22_X1 port map( A1 => Q(794), A2 => n39, B1 => Q(890), B2 => n40, 
                           ZN => n305);
   U323 : NAND4_X1 port map( A1 => n309, A2 => n310, A3 => n311, A4 => n312, ZN
                           => n293);
   U324 : AOI22_X1 port map( A1 => Q(858), A2 => n45, B1 => Q(730), B2 => n46, 
                           ZN => n312);
   U325 : AOI22_X1 port map( A1 => Q(826), A2 => n47, B1 => Q(762), B2 => n48, 
                           ZN => n311);
   U326 : AOI22_X1 port map( A1 => Q(986), A2 => n49, B1 => Q(922), B2 => n50, 
                           ZN => n310);
   U327 : AOI22_X1 port map( A1 => Q(1018), A2 => n51, B1 => Q(954), B2 => n52,
                           ZN => n309);
   U328 : OR4_X1 port map( A1 => n313, A2 => n314, A3 => n315, A4 => n316, ZN 
                           => Y(25));
   U329 : NAND4_X1 port map( A1 => n317, A2 => n318, A3 => n319, A4 => n320, ZN
                           => n316);
   U330 : AOI22_X1 port map( A1 => Q(121), A2 => n9, B1 => Q(217), B2 => n10, 
                           ZN => n320);
   U331 : AOI22_X1 port map( A1 => Q(185), A2 => n11, B1 => Q(57), B2 => n12, 
                           ZN => n319);
   U332 : AOI22_X1 port map( A1 => Q(25), A2 => n13, B1 => Q(89), B2 => n14, ZN
                           => n318);
   U333 : AOI22_X1 port map( A1 => Q(249), A2 => n15, B1 => Q(153), B2 => n16, 
                           ZN => n317);
   U334 : NAND4_X1 port map( A1 => n321, A2 => n322, A3 => n323, A4 => n324, ZN
                           => n315);
   U335 : AOI22_X1 port map( A1 => Q(345), A2 => n21, B1 => Q(441), B2 => n22, 
                           ZN => n324);
   U336 : AOI22_X1 port map( A1 => Q(409), A2 => n23, B1 => Q(281), B2 => n24, 
                           ZN => n323);
   U337 : AOI22_X1 port map( A1 => Q(377), A2 => n25, B1 => Q(313), B2 => n26, 
                           ZN => n322);
   U338 : AOI22_X1 port map( A1 => Q(665), A2 => n27, B1 => Q(473), B2 => n28, 
                           ZN => n321);
   U339 : NAND4_X1 port map( A1 => n325, A2 => n326, A3 => n327, A4 => n328, ZN
                           => n314);
   U340 : AOI22_X1 port map( A1 => Q(505), A2 => n33, B1 => Q(569), B2 => n34, 
                           ZN => n328);
   U341 : AOI22_X1 port map( A1 => Q(537), A2 => n35, B1 => Q(633), B2 => n36, 
                           ZN => n327);
   U342 : AOI22_X1 port map( A1 => Q(697), A2 => n37, B1 => Q(601), B2 => n38, 
                           ZN => n326);
   U343 : AOI22_X1 port map( A1 => Q(793), A2 => n39, B1 => Q(889), B2 => n40, 
                           ZN => n325);
   U344 : NAND4_X1 port map( A1 => n329, A2 => n330, A3 => n331, A4 => n332, ZN
                           => n313);
   U345 : AOI22_X1 port map( A1 => Q(857), A2 => n45, B1 => Q(729), B2 => n46, 
                           ZN => n332);
   U346 : AOI22_X1 port map( A1 => Q(825), A2 => n47, B1 => Q(761), B2 => n48, 
                           ZN => n331);
   U347 : AOI22_X1 port map( A1 => Q(985), A2 => n49, B1 => Q(921), B2 => n50, 
                           ZN => n330);
   U348 : AOI22_X1 port map( A1 => Q(1017), A2 => n51, B1 => Q(953), B2 => n52,
                           ZN => n329);
   U349 : OR4_X1 port map( A1 => n333, A2 => n334, A3 => n335, A4 => n336, ZN 
                           => Y(24));
   U350 : NAND4_X1 port map( A1 => n337, A2 => n338, A3 => n339, A4 => n340, ZN
                           => n336);
   U351 : AOI22_X1 port map( A1 => Q(120), A2 => n9, B1 => Q(216), B2 => n10, 
                           ZN => n340);
   U352 : AOI22_X1 port map( A1 => Q(184), A2 => n11, B1 => Q(56), B2 => n12, 
                           ZN => n339);
   U353 : AOI22_X1 port map( A1 => Q(24), A2 => n13, B1 => Q(88), B2 => n14, ZN
                           => n338);
   U354 : AOI22_X1 port map( A1 => Q(248), A2 => n15, B1 => Q(152), B2 => n16, 
                           ZN => n337);
   U355 : NAND4_X1 port map( A1 => n341, A2 => n342, A3 => n343, A4 => n344, ZN
                           => n335);
   U356 : AOI22_X1 port map( A1 => Q(344), A2 => n21, B1 => Q(440), B2 => n22, 
                           ZN => n344);
   U357 : AOI22_X1 port map( A1 => Q(408), A2 => n23, B1 => Q(280), B2 => n24, 
                           ZN => n343);
   U358 : AOI22_X1 port map( A1 => Q(376), A2 => n25, B1 => Q(312), B2 => n26, 
                           ZN => n342);
   U359 : AOI22_X1 port map( A1 => Q(664), A2 => n27, B1 => Q(472), B2 => n28, 
                           ZN => n341);
   U360 : NAND4_X1 port map( A1 => n345, A2 => n346, A3 => n347, A4 => n348, ZN
                           => n334);
   U361 : AOI22_X1 port map( A1 => Q(504), A2 => n33, B1 => Q(568), B2 => n34, 
                           ZN => n348);
   U362 : AOI22_X1 port map( A1 => Q(536), A2 => n35, B1 => Q(632), B2 => n36, 
                           ZN => n347);
   U363 : AOI22_X1 port map( A1 => Q(696), A2 => n37, B1 => Q(600), B2 => n38, 
                           ZN => n346);
   U364 : AOI22_X1 port map( A1 => Q(792), A2 => n39, B1 => Q(888), B2 => n40, 
                           ZN => n345);
   U365 : NAND4_X1 port map( A1 => n349, A2 => n350, A3 => n351, A4 => n352, ZN
                           => n333);
   U366 : AOI22_X1 port map( A1 => Q(856), A2 => n45, B1 => Q(728), B2 => n46, 
                           ZN => n352);
   U367 : AOI22_X1 port map( A1 => Q(824), A2 => n47, B1 => Q(760), B2 => n48, 
                           ZN => n351);
   U368 : AOI22_X1 port map( A1 => Q(984), A2 => n49, B1 => Q(920), B2 => n50, 
                           ZN => n350);
   U369 : AOI22_X1 port map( A1 => Q(1016), A2 => n51, B1 => Q(952), B2 => n52,
                           ZN => n349);
   U370 : OR4_X1 port map( A1 => n353, A2 => n354, A3 => n355, A4 => n356, ZN 
                           => Y(23));
   U371 : NAND4_X1 port map( A1 => n357, A2 => n358, A3 => n359, A4 => n360, ZN
                           => n356);
   U372 : AOI22_X1 port map( A1 => Q(119), A2 => n9, B1 => Q(215), B2 => n10, 
                           ZN => n360);
   U373 : AOI22_X1 port map( A1 => Q(183), A2 => n11, B1 => Q(55), B2 => n12, 
                           ZN => n359);
   U374 : AOI22_X1 port map( A1 => Q(23), A2 => n13, B1 => Q(87), B2 => n14, ZN
                           => n358);
   U375 : AOI22_X1 port map( A1 => Q(247), A2 => n15, B1 => Q(151), B2 => n16, 
                           ZN => n357);
   U376 : NAND4_X1 port map( A1 => n361, A2 => n362, A3 => n363, A4 => n364, ZN
                           => n355);
   U377 : AOI22_X1 port map( A1 => Q(343), A2 => n21, B1 => Q(439), B2 => n22, 
                           ZN => n364);
   U378 : AOI22_X1 port map( A1 => Q(407), A2 => n23, B1 => Q(279), B2 => n24, 
                           ZN => n363);
   U379 : AOI22_X1 port map( A1 => Q(375), A2 => n25, B1 => Q(311), B2 => n26, 
                           ZN => n362);
   U380 : AOI22_X1 port map( A1 => Q(663), A2 => n27, B1 => Q(471), B2 => n28, 
                           ZN => n361);
   U381 : NAND4_X1 port map( A1 => n365, A2 => n366, A3 => n367, A4 => n368, ZN
                           => n354);
   U382 : AOI22_X1 port map( A1 => Q(503), A2 => n33, B1 => Q(567), B2 => n34, 
                           ZN => n368);
   U383 : AOI22_X1 port map( A1 => Q(535), A2 => n35, B1 => Q(631), B2 => n36, 
                           ZN => n367);
   U384 : AOI22_X1 port map( A1 => Q(695), A2 => n37, B1 => Q(599), B2 => n38, 
                           ZN => n366);
   U385 : AOI22_X1 port map( A1 => Q(791), A2 => n39, B1 => Q(887), B2 => n40, 
                           ZN => n365);
   U386 : NAND4_X1 port map( A1 => n369, A2 => n370, A3 => n371, A4 => n372, ZN
                           => n353);
   U387 : AOI22_X1 port map( A1 => Q(855), A2 => n45, B1 => Q(727), B2 => n46, 
                           ZN => n372);
   U388 : AOI22_X1 port map( A1 => Q(823), A2 => n47, B1 => Q(759), B2 => n48, 
                           ZN => n371);
   U389 : AOI22_X1 port map( A1 => Q(983), A2 => n49, B1 => Q(919), B2 => n50, 
                           ZN => n370);
   U390 : AOI22_X1 port map( A1 => Q(1015), A2 => n51, B1 => Q(951), B2 => n52,
                           ZN => n369);
   U391 : OR4_X1 port map( A1 => n373, A2 => n374, A3 => n375, A4 => n376, ZN 
                           => Y(22));
   U392 : NAND4_X1 port map( A1 => n377, A2 => n378, A3 => n379, A4 => n380, ZN
                           => n376);
   U393 : AOI22_X1 port map( A1 => Q(118), A2 => n9, B1 => Q(214), B2 => n10, 
                           ZN => n380);
   U394 : AOI22_X1 port map( A1 => Q(182), A2 => n11, B1 => Q(54), B2 => n12, 
                           ZN => n379);
   U395 : AOI22_X1 port map( A1 => Q(22), A2 => n13, B1 => Q(86), B2 => n14, ZN
                           => n378);
   U396 : AOI22_X1 port map( A1 => Q(246), A2 => n15, B1 => Q(150), B2 => n16, 
                           ZN => n377);
   U397 : NAND4_X1 port map( A1 => n381, A2 => n382, A3 => n383, A4 => n384, ZN
                           => n375);
   U398 : AOI22_X1 port map( A1 => Q(342), A2 => n21, B1 => Q(438), B2 => n22, 
                           ZN => n384);
   U399 : AOI22_X1 port map( A1 => Q(406), A2 => n23, B1 => Q(278), B2 => n24, 
                           ZN => n383);
   U400 : AOI22_X1 port map( A1 => Q(374), A2 => n25, B1 => Q(310), B2 => n26, 
                           ZN => n382);
   U401 : AOI22_X1 port map( A1 => Q(662), A2 => n27, B1 => Q(470), B2 => n28, 
                           ZN => n381);
   U402 : NAND4_X1 port map( A1 => n385, A2 => n386, A3 => n387, A4 => n388, ZN
                           => n374);
   U403 : AOI22_X1 port map( A1 => Q(502), A2 => n33, B1 => Q(566), B2 => n34, 
                           ZN => n388);
   U404 : AOI22_X1 port map( A1 => Q(534), A2 => n35, B1 => Q(630), B2 => n36, 
                           ZN => n387);
   U405 : AOI22_X1 port map( A1 => Q(694), A2 => n37, B1 => Q(598), B2 => n38, 
                           ZN => n386);
   U406 : AOI22_X1 port map( A1 => Q(790), A2 => n39, B1 => Q(886), B2 => n40, 
                           ZN => n385);
   U407 : NAND4_X1 port map( A1 => n389, A2 => n390, A3 => n391, A4 => n392, ZN
                           => n373);
   U408 : AOI22_X1 port map( A1 => Q(854), A2 => n45, B1 => Q(726), B2 => n46, 
                           ZN => n392);
   U409 : AOI22_X1 port map( A1 => Q(822), A2 => n47, B1 => Q(758), B2 => n48, 
                           ZN => n391);
   U410 : AOI22_X1 port map( A1 => Q(982), A2 => n49, B1 => Q(918), B2 => n50, 
                           ZN => n390);
   U411 : AOI22_X1 port map( A1 => Q(1014), A2 => n51, B1 => Q(950), B2 => n52,
                           ZN => n389);
   U412 : OR4_X1 port map( A1 => n393, A2 => n394, A3 => n395, A4 => n396, ZN 
                           => Y(21));
   U413 : NAND4_X1 port map( A1 => n397, A2 => n398, A3 => n399, A4 => n400, ZN
                           => n396);
   U414 : AOI22_X1 port map( A1 => Q(117), A2 => n9, B1 => Q(213), B2 => n10, 
                           ZN => n400);
   U415 : AOI22_X1 port map( A1 => Q(181), A2 => n11, B1 => Q(53), B2 => n12, 
                           ZN => n399);
   U416 : AOI22_X1 port map( A1 => Q(21), A2 => n13, B1 => Q(85), B2 => n14, ZN
                           => n398);
   U417 : AOI22_X1 port map( A1 => Q(245), A2 => n15, B1 => Q(149), B2 => n16, 
                           ZN => n397);
   U418 : NAND4_X1 port map( A1 => n401, A2 => n402, A3 => n403, A4 => n404, ZN
                           => n395);
   U419 : AOI22_X1 port map( A1 => Q(341), A2 => n21, B1 => Q(437), B2 => n22, 
                           ZN => n404);
   U420 : AOI22_X1 port map( A1 => Q(405), A2 => n23, B1 => Q(277), B2 => n24, 
                           ZN => n403);
   U421 : AOI22_X1 port map( A1 => Q(373), A2 => n25, B1 => Q(309), B2 => n26, 
                           ZN => n402);
   U422 : AOI22_X1 port map( A1 => Q(661), A2 => n27, B1 => Q(469), B2 => n28, 
                           ZN => n401);
   U423 : NAND4_X1 port map( A1 => n405, A2 => n406, A3 => n407, A4 => n408, ZN
                           => n394);
   U424 : AOI22_X1 port map( A1 => Q(501), A2 => n33, B1 => Q(565), B2 => n34, 
                           ZN => n408);
   U425 : AOI22_X1 port map( A1 => Q(533), A2 => n35, B1 => Q(629), B2 => n36, 
                           ZN => n407);
   U426 : AOI22_X1 port map( A1 => Q(693), A2 => n37, B1 => Q(597), B2 => n38, 
                           ZN => n406);
   U427 : AOI22_X1 port map( A1 => Q(789), A2 => n39, B1 => Q(885), B2 => n40, 
                           ZN => n405);
   U428 : NAND4_X1 port map( A1 => n409, A2 => n410, A3 => n411, A4 => n412, ZN
                           => n393);
   U429 : AOI22_X1 port map( A1 => Q(853), A2 => n45, B1 => Q(725), B2 => n46, 
                           ZN => n412);
   U430 : AOI22_X1 port map( A1 => Q(821), A2 => n47, B1 => Q(757), B2 => n48, 
                           ZN => n411);
   U431 : AOI22_X1 port map( A1 => Q(981), A2 => n49, B1 => Q(917), B2 => n50, 
                           ZN => n410);
   U432 : AOI22_X1 port map( A1 => Q(1013), A2 => n51, B1 => Q(949), B2 => n52,
                           ZN => n409);
   U433 : OR4_X1 port map( A1 => n413, A2 => n414, A3 => n415, A4 => n416, ZN 
                           => Y(20));
   U434 : NAND4_X1 port map( A1 => n417, A2 => n418, A3 => n419, A4 => n420, ZN
                           => n416);
   U435 : AOI22_X1 port map( A1 => Q(116), A2 => n9, B1 => Q(212), B2 => n10, 
                           ZN => n420);
   U436 : AOI22_X1 port map( A1 => Q(180), A2 => n11, B1 => Q(52), B2 => n12, 
                           ZN => n419);
   U437 : AOI22_X1 port map( A1 => Q(20), A2 => n13, B1 => Q(84), B2 => n14, ZN
                           => n418);
   U438 : AOI22_X1 port map( A1 => Q(244), A2 => n15, B1 => Q(148), B2 => n16, 
                           ZN => n417);
   U439 : NAND4_X1 port map( A1 => n421, A2 => n422, A3 => n423, A4 => n424, ZN
                           => n415);
   U440 : AOI22_X1 port map( A1 => Q(340), A2 => n21, B1 => Q(436), B2 => n22, 
                           ZN => n424);
   U441 : AOI22_X1 port map( A1 => Q(404), A2 => n23, B1 => Q(276), B2 => n24, 
                           ZN => n423);
   U442 : AOI22_X1 port map( A1 => Q(372), A2 => n25, B1 => Q(308), B2 => n26, 
                           ZN => n422);
   U443 : AOI22_X1 port map( A1 => Q(660), A2 => n27, B1 => Q(468), B2 => n28, 
                           ZN => n421);
   U444 : NAND4_X1 port map( A1 => n425, A2 => n426, A3 => n427, A4 => n428, ZN
                           => n414);
   U445 : AOI22_X1 port map( A1 => Q(500), A2 => n33, B1 => Q(564), B2 => n34, 
                           ZN => n428);
   U446 : AOI22_X1 port map( A1 => Q(532), A2 => n35, B1 => Q(628), B2 => n36, 
                           ZN => n427);
   U447 : AOI22_X1 port map( A1 => Q(692), A2 => n37, B1 => Q(596), B2 => n38, 
                           ZN => n426);
   U448 : AOI22_X1 port map( A1 => Q(788), A2 => n39, B1 => Q(884), B2 => n40, 
                           ZN => n425);
   U449 : NAND4_X1 port map( A1 => n429, A2 => n430, A3 => n431, A4 => n432, ZN
                           => n413);
   U450 : AOI22_X1 port map( A1 => Q(852), A2 => n45, B1 => Q(724), B2 => n46, 
                           ZN => n432);
   U451 : AOI22_X1 port map( A1 => Q(820), A2 => n47, B1 => Q(756), B2 => n48, 
                           ZN => n431);
   U452 : AOI22_X1 port map( A1 => Q(980), A2 => n49, B1 => Q(916), B2 => n50, 
                           ZN => n430);
   U453 : AOI22_X1 port map( A1 => Q(1012), A2 => n51, B1 => Q(948), B2 => n52,
                           ZN => n429);
   U454 : OR4_X1 port map( A1 => n433, A2 => n434, A3 => n435, A4 => n436, ZN 
                           => Y(1));
   U455 : NAND4_X1 port map( A1 => n437, A2 => n438, A3 => n439, A4 => n440, ZN
                           => n436);
   U456 : AOI22_X1 port map( A1 => Q(97), A2 => n9, B1 => Q(193), B2 => n10, ZN
                           => n440);
   U457 : AOI22_X1 port map( A1 => Q(161), A2 => n11, B1 => Q(33), B2 => n12, 
                           ZN => n439);
   U458 : AOI22_X1 port map( A1 => Q(1), A2 => n13, B1 => Q(65), B2 => n14, ZN 
                           => n438);
   U459 : AOI22_X1 port map( A1 => Q(225), A2 => n15, B1 => Q(129), B2 => n16, 
                           ZN => n437);
   U460 : NAND4_X1 port map( A1 => n441, A2 => n442, A3 => n443, A4 => n444, ZN
                           => n435);
   U461 : AOI22_X1 port map( A1 => Q(321), A2 => n21, B1 => Q(417), B2 => n22, 
                           ZN => n444);
   U462 : AOI22_X1 port map( A1 => Q(385), A2 => n23, B1 => Q(257), B2 => n24, 
                           ZN => n443);
   U463 : AOI22_X1 port map( A1 => Q(353), A2 => n25, B1 => Q(289), B2 => n26, 
                           ZN => n442);
   U464 : AOI22_X1 port map( A1 => Q(641), A2 => n27, B1 => Q(449), B2 => n28, 
                           ZN => n441);
   U465 : NAND4_X1 port map( A1 => n445, A2 => n446, A3 => n447, A4 => n448, ZN
                           => n434);
   U466 : AOI22_X1 port map( A1 => Q(481), A2 => n33, B1 => Q(545), B2 => n34, 
                           ZN => n448);
   U467 : AOI22_X1 port map( A1 => Q(513), A2 => n35, B1 => Q(609), B2 => n36, 
                           ZN => n447);
   U468 : AOI22_X1 port map( A1 => Q(673), A2 => n37, B1 => Q(577), B2 => n38, 
                           ZN => n446);
   U469 : AOI22_X1 port map( A1 => Q(769), A2 => n39, B1 => Q(865), B2 => n40, 
                           ZN => n445);
   U470 : NAND4_X1 port map( A1 => n449, A2 => n450, A3 => n451, A4 => n452, ZN
                           => n433);
   U471 : AOI22_X1 port map( A1 => Q(833), A2 => n45, B1 => Q(705), B2 => n46, 
                           ZN => n452);
   U472 : AOI22_X1 port map( A1 => Q(801), A2 => n47, B1 => Q(737), B2 => n48, 
                           ZN => n451);
   U473 : AOI22_X1 port map( A1 => Q(961), A2 => n49, B1 => Q(897), B2 => n50, 
                           ZN => n450);
   U474 : AOI22_X1 port map( A1 => Q(993), A2 => n51, B1 => Q(929), B2 => n52, 
                           ZN => n449);
   U475 : OR4_X1 port map( A1 => n453, A2 => n454, A3 => n455, A4 => n456, ZN 
                           => Y(19));
   U476 : NAND4_X1 port map( A1 => n457, A2 => n458, A3 => n459, A4 => n460, ZN
                           => n456);
   U477 : AOI22_X1 port map( A1 => Q(115), A2 => n9, B1 => Q(211), B2 => n10, 
                           ZN => n460);
   U478 : AOI22_X1 port map( A1 => Q(179), A2 => n11, B1 => Q(51), B2 => n12, 
                           ZN => n459);
   U479 : AOI22_X1 port map( A1 => Q(19), A2 => n13, B1 => Q(83), B2 => n14, ZN
                           => n458);
   U480 : AOI22_X1 port map( A1 => Q(243), A2 => n15, B1 => Q(147), B2 => n16, 
                           ZN => n457);
   U481 : NAND4_X1 port map( A1 => n461, A2 => n462, A3 => n463, A4 => n464, ZN
                           => n455);
   U482 : AOI22_X1 port map( A1 => Q(339), A2 => n21, B1 => Q(435), B2 => n22, 
                           ZN => n464);
   U483 : AOI22_X1 port map( A1 => Q(403), A2 => n23, B1 => Q(275), B2 => n24, 
                           ZN => n463);
   U484 : AOI22_X1 port map( A1 => Q(371), A2 => n25, B1 => Q(307), B2 => n26, 
                           ZN => n462);
   U485 : AOI22_X1 port map( A1 => Q(659), A2 => n27, B1 => Q(467), B2 => n28, 
                           ZN => n461);
   U486 : NAND4_X1 port map( A1 => n465, A2 => n466, A3 => n467, A4 => n468, ZN
                           => n454);
   U487 : AOI22_X1 port map( A1 => Q(499), A2 => n33, B1 => Q(563), B2 => n34, 
                           ZN => n468);
   U488 : AOI22_X1 port map( A1 => Q(531), A2 => n35, B1 => Q(627), B2 => n36, 
                           ZN => n467);
   U489 : AOI22_X1 port map( A1 => Q(691), A2 => n37, B1 => Q(595), B2 => n38, 
                           ZN => n466);
   U490 : AOI22_X1 port map( A1 => Q(787), A2 => n39, B1 => Q(883), B2 => n40, 
                           ZN => n465);
   U491 : NAND4_X1 port map( A1 => n469, A2 => n470, A3 => n471, A4 => n472, ZN
                           => n453);
   U492 : AOI22_X1 port map( A1 => Q(851), A2 => n45, B1 => Q(723), B2 => n46, 
                           ZN => n472);
   U493 : AOI22_X1 port map( A1 => Q(819), A2 => n47, B1 => Q(755), B2 => n48, 
                           ZN => n471);
   U494 : AOI22_X1 port map( A1 => Q(979), A2 => n49, B1 => Q(915), B2 => n50, 
                           ZN => n470);
   U495 : AOI22_X1 port map( A1 => Q(1011), A2 => n51, B1 => Q(947), B2 => n52,
                           ZN => n469);
   U496 : OR4_X1 port map( A1 => n473, A2 => n474, A3 => n475, A4 => n476, ZN 
                           => Y(18));
   U497 : NAND4_X1 port map( A1 => n477, A2 => n478, A3 => n479, A4 => n480, ZN
                           => n476);
   U498 : AOI22_X1 port map( A1 => Q(114), A2 => n9, B1 => Q(210), B2 => n10, 
                           ZN => n480);
   U499 : AOI22_X1 port map( A1 => Q(178), A2 => n11, B1 => Q(50), B2 => n12, 
                           ZN => n479);
   U500 : AOI22_X1 port map( A1 => Q(18), A2 => n13, B1 => Q(82), B2 => n14, ZN
                           => n478);
   U501 : AOI22_X1 port map( A1 => Q(242), A2 => n15, B1 => Q(146), B2 => n16, 
                           ZN => n477);
   U502 : NAND4_X1 port map( A1 => n481, A2 => n482, A3 => n483, A4 => n484, ZN
                           => n475);
   U503 : AOI22_X1 port map( A1 => Q(338), A2 => n21, B1 => Q(434), B2 => n22, 
                           ZN => n484);
   U504 : AOI22_X1 port map( A1 => Q(402), A2 => n23, B1 => Q(274), B2 => n24, 
                           ZN => n483);
   U505 : AOI22_X1 port map( A1 => Q(370), A2 => n25, B1 => Q(306), B2 => n26, 
                           ZN => n482);
   U506 : AOI22_X1 port map( A1 => Q(658), A2 => n27, B1 => Q(466), B2 => n28, 
                           ZN => n481);
   U507 : NAND4_X1 port map( A1 => n485, A2 => n486, A3 => n487, A4 => n488, ZN
                           => n474);
   U508 : AOI22_X1 port map( A1 => Q(498), A2 => n33, B1 => Q(562), B2 => n34, 
                           ZN => n488);
   U509 : AOI22_X1 port map( A1 => Q(530), A2 => n35, B1 => Q(626), B2 => n36, 
                           ZN => n487);
   U510 : AOI22_X1 port map( A1 => Q(690), A2 => n37, B1 => Q(594), B2 => n38, 
                           ZN => n486);
   U511 : AOI22_X1 port map( A1 => Q(786), A2 => n39, B1 => Q(882), B2 => n40, 
                           ZN => n485);
   U512 : NAND4_X1 port map( A1 => n489, A2 => n490, A3 => n491, A4 => n492, ZN
                           => n473);
   U513 : AOI22_X1 port map( A1 => Q(850), A2 => n45, B1 => Q(722), B2 => n46, 
                           ZN => n492);
   U514 : AOI22_X1 port map( A1 => Q(818), A2 => n47, B1 => Q(754), B2 => n48, 
                           ZN => n491);
   U515 : AOI22_X1 port map( A1 => Q(978), A2 => n49, B1 => Q(914), B2 => n50, 
                           ZN => n490);
   U516 : AOI22_X1 port map( A1 => Q(1010), A2 => n51, B1 => Q(946), B2 => n52,
                           ZN => n489);
   U517 : OR4_X1 port map( A1 => n493, A2 => n494, A3 => n495, A4 => n496, ZN 
                           => Y(17));
   U518 : NAND4_X1 port map( A1 => n497, A2 => n498, A3 => n499, A4 => n500, ZN
                           => n496);
   U519 : AOI22_X1 port map( A1 => Q(113), A2 => n9, B1 => Q(209), B2 => n10, 
                           ZN => n500);
   U520 : AOI22_X1 port map( A1 => Q(177), A2 => n11, B1 => Q(49), B2 => n12, 
                           ZN => n499);
   U521 : AOI22_X1 port map( A1 => Q(17), A2 => n13, B1 => Q(81), B2 => n14, ZN
                           => n498);
   U522 : AOI22_X1 port map( A1 => Q(241), A2 => n15, B1 => Q(145), B2 => n16, 
                           ZN => n497);
   U523 : NAND4_X1 port map( A1 => n501, A2 => n502, A3 => n503, A4 => n504, ZN
                           => n495);
   U524 : AOI22_X1 port map( A1 => Q(337), A2 => n21, B1 => Q(433), B2 => n22, 
                           ZN => n504);
   U525 : AOI22_X1 port map( A1 => Q(401), A2 => n23, B1 => Q(273), B2 => n24, 
                           ZN => n503);
   U526 : AOI22_X1 port map( A1 => Q(369), A2 => n25, B1 => Q(305), B2 => n26, 
                           ZN => n502);
   U527 : AOI22_X1 port map( A1 => Q(657), A2 => n27, B1 => Q(465), B2 => n28, 
                           ZN => n501);
   U528 : NAND4_X1 port map( A1 => n505, A2 => n506, A3 => n507, A4 => n508, ZN
                           => n494);
   U529 : AOI22_X1 port map( A1 => Q(497), A2 => n33, B1 => Q(561), B2 => n34, 
                           ZN => n508);
   U530 : AOI22_X1 port map( A1 => Q(529), A2 => n35, B1 => Q(625), B2 => n36, 
                           ZN => n507);
   U531 : AOI22_X1 port map( A1 => Q(689), A2 => n37, B1 => Q(593), B2 => n38, 
                           ZN => n506);
   U532 : AOI22_X1 port map( A1 => Q(785), A2 => n39, B1 => Q(881), B2 => n40, 
                           ZN => n505);
   U533 : NAND4_X1 port map( A1 => n509, A2 => n510, A3 => n511, A4 => n512, ZN
                           => n493);
   U534 : AOI22_X1 port map( A1 => Q(849), A2 => n45, B1 => Q(721), B2 => n46, 
                           ZN => n512);
   U535 : AOI22_X1 port map( A1 => Q(817), A2 => n47, B1 => Q(753), B2 => n48, 
                           ZN => n511);
   U536 : AOI22_X1 port map( A1 => Q(977), A2 => n49, B1 => Q(913), B2 => n50, 
                           ZN => n510);
   U537 : AOI22_X1 port map( A1 => Q(1009), A2 => n51, B1 => Q(945), B2 => n52,
                           ZN => n509);
   U538 : OR4_X1 port map( A1 => n513, A2 => n514, A3 => n515, A4 => n516, ZN 
                           => Y(16));
   U539 : NAND4_X1 port map( A1 => n517, A2 => n518, A3 => n519, A4 => n520, ZN
                           => n516);
   U540 : AOI22_X1 port map( A1 => Q(112), A2 => n9, B1 => Q(208), B2 => n10, 
                           ZN => n520);
   U541 : AOI22_X1 port map( A1 => Q(176), A2 => n11, B1 => Q(48), B2 => n12, 
                           ZN => n519);
   U542 : AOI22_X1 port map( A1 => Q(16), A2 => n13, B1 => Q(80), B2 => n14, ZN
                           => n518);
   U543 : AOI22_X1 port map( A1 => Q(240), A2 => n15, B1 => Q(144), B2 => n16, 
                           ZN => n517);
   U544 : NAND4_X1 port map( A1 => n521, A2 => n522, A3 => n523, A4 => n524, ZN
                           => n515);
   U545 : AOI22_X1 port map( A1 => Q(336), A2 => n21, B1 => Q(432), B2 => n22, 
                           ZN => n524);
   U546 : AOI22_X1 port map( A1 => Q(400), A2 => n23, B1 => Q(272), B2 => n24, 
                           ZN => n523);
   U547 : AOI22_X1 port map( A1 => Q(368), A2 => n25, B1 => Q(304), B2 => n26, 
                           ZN => n522);
   U548 : AOI22_X1 port map( A1 => Q(656), A2 => n27, B1 => Q(464), B2 => n28, 
                           ZN => n521);
   U549 : NAND4_X1 port map( A1 => n525, A2 => n526, A3 => n527, A4 => n528, ZN
                           => n514);
   U550 : AOI22_X1 port map( A1 => Q(496), A2 => n33, B1 => Q(560), B2 => n34, 
                           ZN => n528);
   U551 : AOI22_X1 port map( A1 => Q(528), A2 => n35, B1 => Q(624), B2 => n36, 
                           ZN => n527);
   U552 : AOI22_X1 port map( A1 => Q(688), A2 => n37, B1 => Q(592), B2 => n38, 
                           ZN => n526);
   U553 : AOI22_X1 port map( A1 => Q(784), A2 => n39, B1 => Q(880), B2 => n40, 
                           ZN => n525);
   U554 : NAND4_X1 port map( A1 => n529, A2 => n530, A3 => n531, A4 => n532, ZN
                           => n513);
   U555 : AOI22_X1 port map( A1 => Q(848), A2 => n45, B1 => Q(720), B2 => n46, 
                           ZN => n532);
   U556 : AOI22_X1 port map( A1 => Q(816), A2 => n47, B1 => Q(752), B2 => n48, 
                           ZN => n531);
   U557 : AOI22_X1 port map( A1 => Q(976), A2 => n49, B1 => Q(912), B2 => n50, 
                           ZN => n530);
   U558 : AOI22_X1 port map( A1 => Q(1008), A2 => n51, B1 => Q(944), B2 => n52,
                           ZN => n529);
   U559 : OR4_X1 port map( A1 => n533, A2 => n534, A3 => n535, A4 => n536, ZN 
                           => Y(15));
   U560 : NAND4_X1 port map( A1 => n537, A2 => n538, A3 => n539, A4 => n540, ZN
                           => n536);
   U561 : AOI22_X1 port map( A1 => Q(111), A2 => n9, B1 => Q(207), B2 => n10, 
                           ZN => n540);
   U562 : AOI22_X1 port map( A1 => Q(175), A2 => n11, B1 => Q(47), B2 => n12, 
                           ZN => n539);
   U563 : AOI22_X1 port map( A1 => Q(15), A2 => n13, B1 => Q(79), B2 => n14, ZN
                           => n538);
   U564 : AOI22_X1 port map( A1 => Q(239), A2 => n15, B1 => Q(143), B2 => n16, 
                           ZN => n537);
   U565 : NAND4_X1 port map( A1 => n541, A2 => n542, A3 => n543, A4 => n544, ZN
                           => n535);
   U566 : AOI22_X1 port map( A1 => Q(335), A2 => n21, B1 => Q(431), B2 => n22, 
                           ZN => n544);
   U567 : AOI22_X1 port map( A1 => Q(399), A2 => n23, B1 => Q(271), B2 => n24, 
                           ZN => n543);
   U568 : AOI22_X1 port map( A1 => Q(367), A2 => n25, B1 => Q(303), B2 => n26, 
                           ZN => n542);
   U569 : AOI22_X1 port map( A1 => Q(655), A2 => n27, B1 => Q(463), B2 => n28, 
                           ZN => n541);
   U570 : NAND4_X1 port map( A1 => n545, A2 => n546, A3 => n547, A4 => n548, ZN
                           => n534);
   U571 : AOI22_X1 port map( A1 => Q(495), A2 => n33, B1 => Q(559), B2 => n34, 
                           ZN => n548);
   U572 : AOI22_X1 port map( A1 => Q(527), A2 => n35, B1 => Q(623), B2 => n36, 
                           ZN => n547);
   U573 : AOI22_X1 port map( A1 => Q(687), A2 => n37, B1 => Q(591), B2 => n38, 
                           ZN => n546);
   U574 : AOI22_X1 port map( A1 => Q(783), A2 => n39, B1 => Q(879), B2 => n40, 
                           ZN => n545);
   U575 : NAND4_X1 port map( A1 => n549, A2 => n550, A3 => n551, A4 => n552, ZN
                           => n533);
   U576 : AOI22_X1 port map( A1 => Q(847), A2 => n45, B1 => Q(719), B2 => n46, 
                           ZN => n552);
   U577 : AOI22_X1 port map( A1 => Q(815), A2 => n47, B1 => Q(751), B2 => n48, 
                           ZN => n551);
   U578 : AOI22_X1 port map( A1 => Q(975), A2 => n49, B1 => Q(911), B2 => n50, 
                           ZN => n550);
   U579 : AOI22_X1 port map( A1 => Q(1007), A2 => n51, B1 => Q(943), B2 => n52,
                           ZN => n549);
   U580 : OR4_X1 port map( A1 => n553, A2 => n554, A3 => n555, A4 => n556, ZN 
                           => Y(14));
   U581 : NAND4_X1 port map( A1 => n557, A2 => n558, A3 => n559, A4 => n560, ZN
                           => n556);
   U582 : AOI22_X1 port map( A1 => Q(110), A2 => n9, B1 => Q(206), B2 => n10, 
                           ZN => n560);
   U583 : AOI22_X1 port map( A1 => Q(174), A2 => n11, B1 => Q(46), B2 => n12, 
                           ZN => n559);
   U584 : AOI22_X1 port map( A1 => Q(14), A2 => n13, B1 => Q(78), B2 => n14, ZN
                           => n558);
   U585 : AOI22_X1 port map( A1 => Q(238), A2 => n15, B1 => Q(142), B2 => n16, 
                           ZN => n557);
   U586 : NAND4_X1 port map( A1 => n561, A2 => n562, A3 => n563, A4 => n564, ZN
                           => n555);
   U587 : AOI22_X1 port map( A1 => Q(334), A2 => n21, B1 => Q(430), B2 => n22, 
                           ZN => n564);
   U588 : AOI22_X1 port map( A1 => Q(398), A2 => n23, B1 => Q(270), B2 => n24, 
                           ZN => n563);
   U589 : AOI22_X1 port map( A1 => Q(366), A2 => n25, B1 => Q(302), B2 => n26, 
                           ZN => n562);
   U590 : AOI22_X1 port map( A1 => Q(654), A2 => n27, B1 => Q(462), B2 => n28, 
                           ZN => n561);
   U591 : NAND4_X1 port map( A1 => n565, A2 => n566, A3 => n567, A4 => n568, ZN
                           => n554);
   U592 : AOI22_X1 port map( A1 => Q(494), A2 => n33, B1 => Q(558), B2 => n34, 
                           ZN => n568);
   U593 : AOI22_X1 port map( A1 => Q(526), A2 => n35, B1 => Q(622), B2 => n36, 
                           ZN => n567);
   U594 : AOI22_X1 port map( A1 => Q(686), A2 => n37, B1 => Q(590), B2 => n38, 
                           ZN => n566);
   U595 : AOI22_X1 port map( A1 => Q(782), A2 => n39, B1 => Q(878), B2 => n40, 
                           ZN => n565);
   U596 : NAND4_X1 port map( A1 => n569, A2 => n570, A3 => n571, A4 => n572, ZN
                           => n553);
   U597 : AOI22_X1 port map( A1 => Q(846), A2 => n45, B1 => Q(718), B2 => n46, 
                           ZN => n572);
   U598 : AOI22_X1 port map( A1 => Q(814), A2 => n47, B1 => Q(750), B2 => n48, 
                           ZN => n571);
   U599 : AOI22_X1 port map( A1 => Q(974), A2 => n49, B1 => Q(910), B2 => n50, 
                           ZN => n570);
   U600 : AOI22_X1 port map( A1 => Q(1006), A2 => n51, B1 => Q(942), B2 => n52,
                           ZN => n569);
   U601 : OR4_X1 port map( A1 => n573, A2 => n574, A3 => n575, A4 => n576, ZN 
                           => Y(13));
   U602 : NAND4_X1 port map( A1 => n577, A2 => n578, A3 => n579, A4 => n580, ZN
                           => n576);
   U603 : AOI22_X1 port map( A1 => Q(109), A2 => n9, B1 => Q(205), B2 => n10, 
                           ZN => n580);
   U604 : AOI22_X1 port map( A1 => Q(173), A2 => n11, B1 => Q(45), B2 => n12, 
                           ZN => n579);
   U605 : AOI22_X1 port map( A1 => Q(13), A2 => n13, B1 => Q(77), B2 => n14, ZN
                           => n578);
   U606 : AOI22_X1 port map( A1 => Q(237), A2 => n15, B1 => Q(141), B2 => n16, 
                           ZN => n577);
   U607 : NAND4_X1 port map( A1 => n581, A2 => n582, A3 => n583, A4 => n584, ZN
                           => n575);
   U608 : AOI22_X1 port map( A1 => Q(333), A2 => n21, B1 => Q(429), B2 => n22, 
                           ZN => n584);
   U609 : AOI22_X1 port map( A1 => Q(397), A2 => n23, B1 => Q(269), B2 => n24, 
                           ZN => n583);
   U610 : AOI22_X1 port map( A1 => Q(365), A2 => n25, B1 => Q(301), B2 => n26, 
                           ZN => n582);
   U611 : AOI22_X1 port map( A1 => Q(653), A2 => n27, B1 => Q(461), B2 => n28, 
                           ZN => n581);
   U612 : NAND4_X1 port map( A1 => n585, A2 => n586, A3 => n587, A4 => n588, ZN
                           => n574);
   U613 : AOI22_X1 port map( A1 => Q(493), A2 => n33, B1 => Q(557), B2 => n34, 
                           ZN => n588);
   U614 : AOI22_X1 port map( A1 => Q(525), A2 => n35, B1 => Q(621), B2 => n36, 
                           ZN => n587);
   U615 : AOI22_X1 port map( A1 => Q(685), A2 => n37, B1 => Q(589), B2 => n38, 
                           ZN => n586);
   U616 : AOI22_X1 port map( A1 => Q(781), A2 => n39, B1 => Q(877), B2 => n40, 
                           ZN => n585);
   U617 : NAND4_X1 port map( A1 => n589, A2 => n590, A3 => n591, A4 => n592, ZN
                           => n573);
   U618 : AOI22_X1 port map( A1 => Q(845), A2 => n45, B1 => Q(717), B2 => n46, 
                           ZN => n592);
   U619 : AOI22_X1 port map( A1 => Q(813), A2 => n47, B1 => Q(749), B2 => n48, 
                           ZN => n591);
   U620 : AOI22_X1 port map( A1 => Q(973), A2 => n49, B1 => Q(909), B2 => n50, 
                           ZN => n590);
   U621 : AOI22_X1 port map( A1 => Q(1005), A2 => n51, B1 => Q(941), B2 => n52,
                           ZN => n589);
   U622 : OR4_X1 port map( A1 => n593, A2 => n594, A3 => n595, A4 => n596, ZN 
                           => Y(12));
   U623 : NAND4_X1 port map( A1 => n597, A2 => n598, A3 => n599, A4 => n600, ZN
                           => n596);
   U624 : AOI22_X1 port map( A1 => Q(108), A2 => n9, B1 => Q(204), B2 => n10, 
                           ZN => n600);
   U625 : AOI22_X1 port map( A1 => Q(172), A2 => n11, B1 => Q(44), B2 => n12, 
                           ZN => n599);
   U626 : AOI22_X1 port map( A1 => Q(12), A2 => n13, B1 => Q(76), B2 => n14, ZN
                           => n598);
   U627 : AOI22_X1 port map( A1 => Q(236), A2 => n15, B1 => Q(140), B2 => n16, 
                           ZN => n597);
   U628 : NAND4_X1 port map( A1 => n601, A2 => n602, A3 => n603, A4 => n604, ZN
                           => n595);
   U629 : AOI22_X1 port map( A1 => Q(332), A2 => n21, B1 => Q(428), B2 => n22, 
                           ZN => n604);
   U630 : AOI22_X1 port map( A1 => Q(396), A2 => n23, B1 => Q(268), B2 => n24, 
                           ZN => n603);
   U631 : AOI22_X1 port map( A1 => Q(364), A2 => n25, B1 => Q(300), B2 => n26, 
                           ZN => n602);
   U632 : AOI22_X1 port map( A1 => Q(652), A2 => n27, B1 => Q(460), B2 => n28, 
                           ZN => n601);
   U633 : NAND4_X1 port map( A1 => n605, A2 => n606, A3 => n607, A4 => n608, ZN
                           => n594);
   U634 : AOI22_X1 port map( A1 => Q(492), A2 => n33, B1 => Q(556), B2 => n34, 
                           ZN => n608);
   U635 : AOI22_X1 port map( A1 => Q(524), A2 => n35, B1 => Q(620), B2 => n36, 
                           ZN => n607);
   U636 : AOI22_X1 port map( A1 => Q(684), A2 => n37, B1 => Q(588), B2 => n38, 
                           ZN => n606);
   U637 : AOI22_X1 port map( A1 => Q(780), A2 => n39, B1 => Q(876), B2 => n40, 
                           ZN => n605);
   U638 : NAND4_X1 port map( A1 => n609, A2 => n610, A3 => n611, A4 => n612, ZN
                           => n593);
   U639 : AOI22_X1 port map( A1 => Q(844), A2 => n45, B1 => Q(716), B2 => n46, 
                           ZN => n612);
   U640 : AOI22_X1 port map( A1 => Q(812), A2 => n47, B1 => Q(748), B2 => n48, 
                           ZN => n611);
   U641 : AOI22_X1 port map( A1 => Q(972), A2 => n49, B1 => Q(908), B2 => n50, 
                           ZN => n610);
   U642 : AOI22_X1 port map( A1 => Q(1004), A2 => n51, B1 => Q(940), B2 => n52,
                           ZN => n609);
   U643 : OR4_X1 port map( A1 => n613, A2 => n614, A3 => n615, A4 => n616, ZN 
                           => Y(11));
   U644 : NAND4_X1 port map( A1 => n617, A2 => n618, A3 => n619, A4 => n620, ZN
                           => n616);
   U645 : AOI22_X1 port map( A1 => Q(107), A2 => n9, B1 => Q(203), B2 => n10, 
                           ZN => n620);
   U646 : AOI22_X1 port map( A1 => Q(171), A2 => n11, B1 => Q(43), B2 => n12, 
                           ZN => n619);
   U647 : AOI22_X1 port map( A1 => Q(11), A2 => n13, B1 => Q(75), B2 => n14, ZN
                           => n618);
   U648 : AOI22_X1 port map( A1 => Q(235), A2 => n15, B1 => Q(139), B2 => n16, 
                           ZN => n617);
   U649 : NAND4_X1 port map( A1 => n621, A2 => n622, A3 => n623, A4 => n624, ZN
                           => n615);
   U650 : AOI22_X1 port map( A1 => Q(331), A2 => n21, B1 => Q(427), B2 => n22, 
                           ZN => n624);
   U651 : AOI22_X1 port map( A1 => Q(395), A2 => n23, B1 => Q(267), B2 => n24, 
                           ZN => n623);
   U652 : AOI22_X1 port map( A1 => Q(363), A2 => n25, B1 => Q(299), B2 => n26, 
                           ZN => n622);
   U653 : AOI22_X1 port map( A1 => Q(651), A2 => n27, B1 => Q(459), B2 => n28, 
                           ZN => n621);
   U654 : NAND4_X1 port map( A1 => n625, A2 => n626, A3 => n627, A4 => n628, ZN
                           => n614);
   U655 : AOI22_X1 port map( A1 => Q(491), A2 => n33, B1 => Q(555), B2 => n34, 
                           ZN => n628);
   U656 : AOI22_X1 port map( A1 => Q(523), A2 => n35, B1 => Q(619), B2 => n36, 
                           ZN => n627);
   U657 : AOI22_X1 port map( A1 => Q(683), A2 => n37, B1 => Q(587), B2 => n38, 
                           ZN => n626);
   U658 : AOI22_X1 port map( A1 => Q(779), A2 => n39, B1 => Q(875), B2 => n40, 
                           ZN => n625);
   U659 : NAND4_X1 port map( A1 => n629, A2 => n630, A3 => n631, A4 => n632, ZN
                           => n613);
   U660 : AOI22_X1 port map( A1 => Q(843), A2 => n45, B1 => Q(715), B2 => n46, 
                           ZN => n632);
   U661 : AOI22_X1 port map( A1 => Q(811), A2 => n47, B1 => Q(747), B2 => n48, 
                           ZN => n631);
   U662 : AOI22_X1 port map( A1 => Q(971), A2 => n49, B1 => Q(907), B2 => n50, 
                           ZN => n630);
   U663 : AOI22_X1 port map( A1 => Q(1003), A2 => n51, B1 => Q(939), B2 => n52,
                           ZN => n629);
   U664 : OR4_X1 port map( A1 => n633, A2 => n634, A3 => n635, A4 => n636, ZN 
                           => Y(10));
   U665 : NAND4_X1 port map( A1 => n637, A2 => n638, A3 => n639, A4 => n640, ZN
                           => n636);
   U666 : AOI22_X1 port map( A1 => Q(106), A2 => n9, B1 => Q(202), B2 => n10, 
                           ZN => n640);
   U667 : AOI22_X1 port map( A1 => Q(170), A2 => n11, B1 => Q(42), B2 => n12, 
                           ZN => n639);
   U668 : AOI22_X1 port map( A1 => Q(10), A2 => n13, B1 => Q(74), B2 => n14, ZN
                           => n638);
   U669 : AOI22_X1 port map( A1 => Q(234), A2 => n15, B1 => Q(138), B2 => n16, 
                           ZN => n637);
   U670 : NAND4_X1 port map( A1 => n641, A2 => n642, A3 => n643, A4 => n644, ZN
                           => n635);
   U671 : AOI22_X1 port map( A1 => Q(330), A2 => n21, B1 => Q(426), B2 => n22, 
                           ZN => n644);
   U672 : AOI22_X1 port map( A1 => Q(394), A2 => n23, B1 => Q(266), B2 => n24, 
                           ZN => n643);
   U673 : AOI22_X1 port map( A1 => Q(362), A2 => n25, B1 => Q(298), B2 => n26, 
                           ZN => n642);
   U674 : AOI22_X1 port map( A1 => Q(650), A2 => n27, B1 => Q(458), B2 => n28, 
                           ZN => n641);
   U675 : NAND4_X1 port map( A1 => n645, A2 => n646, A3 => n647, A4 => n648, ZN
                           => n634);
   U676 : AOI22_X1 port map( A1 => Q(490), A2 => n33, B1 => Q(554), B2 => n34, 
                           ZN => n648);
   U677 : AOI22_X1 port map( A1 => Q(522), A2 => n35, B1 => Q(618), B2 => n36, 
                           ZN => n647);
   U678 : AOI22_X1 port map( A1 => Q(682), A2 => n37, B1 => Q(586), B2 => n38, 
                           ZN => n646);
   U679 : AOI22_X1 port map( A1 => Q(778), A2 => n39, B1 => Q(874), B2 => n40, 
                           ZN => n645);
   U680 : NAND4_X1 port map( A1 => n649, A2 => n650, A3 => n651, A4 => n652, ZN
                           => n633);
   U681 : AOI22_X1 port map( A1 => Q(842), A2 => n45, B1 => Q(714), B2 => n46, 
                           ZN => n652);
   U682 : AOI22_X1 port map( A1 => Q(810), A2 => n47, B1 => Q(746), B2 => n48, 
                           ZN => n651);
   U683 : AOI22_X1 port map( A1 => Q(970), A2 => n49, B1 => Q(906), B2 => n50, 
                           ZN => n650);
   U684 : AOI22_X1 port map( A1 => Q(1002), A2 => n51, B1 => Q(938), B2 => n52,
                           ZN => n649);
   U685 : OR4_X1 port map( A1 => n653, A2 => n654, A3 => n655, A4 => n656, ZN 
                           => Y(0));
   U686 : NAND4_X1 port map( A1 => n657, A2 => n658, A3 => n659, A4 => n660, ZN
                           => n656);
   U687 : AOI22_X1 port map( A1 => Q(96), A2 => n9, B1 => Q(192), B2 => n10, ZN
                           => n660);
   U688 : AOI22_X1 port map( A1 => Q(160), A2 => n11, B1 => Q(32), B2 => n12, 
                           ZN => n659);
   U689 : AOI22_X1 port map( A1 => Q(0), A2 => n13, B1 => Q(64), B2 => n14, ZN 
                           => n658);
   U690 : AOI22_X1 port map( A1 => Q(224), A2 => n15, B1 => Q(128), B2 => n16, 
                           ZN => n657);
   U691 : NOR3_X1 port map( A1 => S(3), A2 => S(4), A3 => S(0), ZN => n661);
   U692 : NOR3_X1 port map( A1 => S(3), A2 => S(4), A3 => n667, ZN => n663);
   U693 : NAND4_X1 port map( A1 => n668, A2 => n669, A3 => n670, A4 => n671, ZN
                           => n655);
   U694 : AOI22_X1 port map( A1 => Q(320), A2 => n21, B1 => Q(416), B2 => n22, 
                           ZN => n671);
   U695 : AOI22_X1 port map( A1 => Q(384), A2 => n23, B1 => Q(256), B2 => n24, 
                           ZN => n670);
   U696 : AOI22_X1 port map( A1 => Q(352), A2 => n25, B1 => Q(288), B2 => n26, 
                           ZN => n669);
   U697 : AOI22_X1 port map( A1 => Q(640), A2 => n27, B1 => Q(448), B2 => n28, 
                           ZN => n668);
   U698 : NOR3_X1 port map( A1 => S(0), A2 => S(4), A3 => n674, ZN => n673);
   U699 : NAND4_X1 port map( A1 => n676, A2 => n677, A3 => n678, A4 => n679, ZN
                           => n654);
   U700 : AOI22_X1 port map( A1 => Q(480), A2 => n33, B1 => Q(544), B2 => n34, 
                           ZN => n679);
   U701 : NOR3_X1 port map( A1 => n674, A2 => S(4), A3 => n667, ZN => n672);
   U702 : AOI22_X1 port map( A1 => Q(512), A2 => n35, B1 => Q(608), B2 => n36, 
                           ZN => n678);
   U703 : AOI22_X1 port map( A1 => Q(672), A2 => n37, B1 => Q(576), B2 => n38, 
                           ZN => n677);
   U704 : AOI22_X1 port map( A1 => Q(768), A2 => n39, B1 => Q(864), B2 => n40, 
                           ZN => n676);
   U705 : NAND4_X1 port map( A1 => n683, A2 => n684, A3 => n685, A4 => n686, ZN
                           => n653);
   U706 : AOI22_X1 port map( A1 => Q(832), A2 => n45, B1 => Q(704), B2 => n46, 
                           ZN => n686);
   U707 : NOR3_X1 port map( A1 => S(0), A2 => S(3), A3 => n687, ZN => n675);
   U708 : NOR2_X1 port map( A1 => n688, A2 => S(2), ZN => n664);
   U709 : AOI22_X1 port map( A1 => Q(800), A2 => n47, B1 => Q(736), B2 => n48, 
                           ZN => n685);
   U710 : NOR3_X1 port map( A1 => n667, A2 => S(3), A3 => n687, ZN => n680);
   U711 : NOR2_X1 port map( A1 => S(1), A2 => S(2), ZN => n665);
   U712 : AOI22_X1 port map( A1 => Q(960), A2 => n49, B1 => Q(896), B2 => n50, 
                           ZN => n684);
   U713 : NOR3_X1 port map( A1 => n674, A2 => S(0), A3 => n687, ZN => n682);
   U714 : AOI22_X1 port map( A1 => Q(992), A2 => n51, B1 => Q(928), B2 => n52, 
                           ZN => n683);
   U715 : NOR2_X1 port map( A1 => n689, A2 => S(1), ZN => n666);
   U716 : NOR2_X1 port map( A1 => n689, A2 => n688, ZN => n662);
   U717 : INV_X1 port map( A => S(1), ZN => n688);
   U718 : INV_X1 port map( A => S(2), ZN => n689);
   U719 : NOR3_X1 port map( A1 => n667, A2 => n674, A3 => n687, ZN => n681);
   U720 : INV_X1 port map( A => S(4), ZN => n687);
   U721 : INV_X1 port map( A => S(3), ZN => n674);
   U722 : INV_X1 port map( A => S(0), ZN => n667);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N5_RSTVAL1_1 is

   port( D : in std_logic_vector (4 downto 0);  Q : out std_logic_vector (4 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N5_RSTVAL1_1;

architecture SYN_Behavioural of reg_generic_N5_RSTVAL1_1 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1, n2, n3, n4, n5,
      n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n18, n_1000 : 
      std_logic;

begin
   Q <= ( Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_4_inst : DFF_X1 port map( D => n17, CK => Clk, Q => Q_4_port, QN => 
                           n12);
   Q_reg_3_inst : DFF_X1 port map( D => n16, CK => Clk, Q => Q_3_port, QN => 
                           n11);
   Q_reg_2_inst : DFF_X1 port map( D => n15, CK => Clk, Q => Q_2_port, QN => 
                           n10);
   Q_reg_1_inst : DFF_X1 port map( D => n13, CK => Clk, Q => Q_1_port, QN => n9
                           );
   Q_reg_0_inst : DFF_X1 port map( D => n18, CK => Clk, Q => Q_0_port, QN => 
                           n_1000);
   U3 : OAI22_X1 port map( A1 => n9, A2 => n1, B1 => n2, B2 => n3, ZN => n13);
   U4 : INV_X1 port map( A => D(1), ZN => n3);
   U5 : OAI22_X1 port map( A1 => n10, A2 => n1, B1 => n2, B2 => n4, ZN => n15);
   U6 : INV_X1 port map( A => D(2), ZN => n4);
   U7 : OAI22_X1 port map( A1 => n11, A2 => n1, B1 => n2, B2 => n5, ZN => n16);
   U8 : INV_X1 port map( A => D(3), ZN => n5);
   U9 : OAI22_X1 port map( A1 => n12, A2 => n1, B1 => n2, B2 => n6, ZN => n17);
   U10 : INV_X1 port map( A => D(4), ZN => n6);
   U11 : OR2_X1 port map( A1 => n7, A2 => Rst, ZN => n2);
   U12 : MUX2_X1 port map( A => Q_0_port, B => n8, S => n1, Z => n18);
   U13 : INV_X1 port map( A => n7, ZN => n1);
   U14 : NOR2_X1 port map( A1 => Rst, A2 => Enable, ZN => n7);
   U15 : OR2_X1 port map( A1 => D(0), A2 => Rst, ZN => n8);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity nwin_calc_F5_1 is

   port( c_win : in std_logic_vector (4 downto 0);  sel : in std_logic_vector 
         (1 downto 0);  n_win : out std_logic_vector (4 downto 0));

end nwin_calc_F5_1;

architecture SYN_struct of nwin_calc_F5_1 is

   component mux_N5_M2_1
      port( S : in std_logic_vector (1 downto 0);  Q : in std_logic_vector (19 
            downto 0);  Y : out std_logic_vector (4 downto 0));
   end component;

begin
   
   MUX_SEL : mux_N5_M2_1 port map( S(1) => sel(1), S(0) => sel(0), Q(19) => 
                           c_win(4), Q(18) => c_win(3), Q(17) => c_win(2), 
                           Q(16) => c_win(1), Q(15) => c_win(0), Q(14) => 
                           c_win(0), Q(13) => c_win(4), Q(12) => c_win(3), 
                           Q(11) => c_win(2), Q(10) => c_win(1), Q(9) => 
                           c_win(3), Q(8) => c_win(2), Q(7) => c_win(1), Q(6) 
                           => c_win(0), Q(5) => c_win(4), Q(4) => c_win(4), 
                           Q(3) => c_win(3), Q(2) => c_win(2), Q(1) => c_win(1)
                           , Q(0) => c_win(0), Y(4) => n_win(4), Y(3) => 
                           n_win(3), Y(2) => n_win(2), Y(1) => n_win(1), Y(0) 
                           => n_win(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N5_M2_0 is

   port( S : in std_logic_vector (1 downto 0);  Q : in std_logic_vector (19 
         downto 0);  Y : out std_logic_vector (4 downto 0));

end mux_N5_M2_0;

architecture SYN_behav of mux_N5_M2_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => Y(4));
   U3 : AOI22_X1 port map( A1 => Q(4), A2 => n3, B1 => Q(14), B2 => n4, ZN => 
                           n2);
   U4 : AOI22_X1 port map( A1 => Q(19), A2 => n5, B1 => Q(9), B2 => n6, ZN => 
                           n1);
   U5 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Y(3));
   U6 : AOI22_X1 port map( A1 => Q(3), A2 => n3, B1 => Q(13), B2 => n4, ZN => 
                           n8);
   U7 : AOI22_X1 port map( A1 => Q(18), A2 => n5, B1 => Q(8), B2 => n6, ZN => 
                           n7);
   U8 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => Y(2));
   U9 : AOI22_X1 port map( A1 => Q(2), A2 => n3, B1 => Q(12), B2 => n4, ZN => 
                           n10);
   U10 : AOI22_X1 port map( A1 => Q(17), A2 => n5, B1 => Q(7), B2 => n6, ZN => 
                           n9);
   U11 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => Y(1));
   U12 : AOI22_X1 port map( A1 => Q(1), A2 => n3, B1 => Q(11), B2 => n4, ZN => 
                           n12);
   U13 : AOI22_X1 port map( A1 => Q(16), A2 => n5, B1 => Q(6), B2 => n6, ZN => 
                           n11);
   U14 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => Y(0));
   U15 : AOI22_X1 port map( A1 => Q(0), A2 => n3, B1 => Q(10), B2 => n4, ZN => 
                           n14);
   U16 : NOR3_X1 port map( A1 => n5, A2 => n6, A3 => n4, ZN => n3);
   U17 : NOR2_X1 port map( A1 => n15, A2 => S(0), ZN => n4);
   U18 : AOI22_X1 port map( A1 => Q(15), A2 => n5, B1 => Q(5), B2 => n6, ZN => 
                           n13);
   U19 : NOR2_X1 port map( A1 => n16, A2 => S(1), ZN => n6);
   U20 : NOR2_X1 port map( A1 => n15, A2 => n16, ZN => n5);
   U21 : INV_X1 port map( A => S(0), ZN => n16);
   U22 : INV_X1 port map( A => S(1), ZN => n15);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M4 is

   port( S : in std_logic_vector (3 downto 0);  Q : in std_logic_vector (511 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end mux_N32_M4;

architecture SYN_behav of mux_N32_M4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348 : std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n333, A2 => n338, ZN => n14);
   U3 : AND2_X2 port map( A1 => n335, A2 => n334, ZN => n12);
   U4 : AND2_X2 port map( A1 => n344, A2 => n334, ZN => n26);
   U5 : AND2_X2 port map( A1 => n337, A2 => n345, ZN => n24);
   U6 : AND2_X2 port map( A1 => n333, A2 => n336, ZN => n13);
   U7 : AND2_X2 port map( A1 => n335, A2 => n337, ZN => n10);
   U8 : AND2_X2 port map( A1 => n338, A2 => n345, ZN => n22);
   U9 : AND2_X2 port map( A1 => n336, A2 => n344, ZN => n25);
   U10 : AND2_X2 port map( A1 => n333, A2 => n334, ZN => n8);
   U11 : AND2_X2 port map( A1 => n344, A2 => n337, ZN => n20);
   U12 : AND2_X2 port map( A1 => n335, A2 => n338, ZN => n11);
   U13 : AND2_X2 port map( A1 => n336, A2 => n345, ZN => n23);
   U14 : AND2_X2 port map( A1 => n333, A2 => n337, ZN => n9);
   U15 : AND2_X2 port map( A1 => n335, A2 => n336, ZN => n7);
   U16 : AND2_X2 port map( A1 => n338, A2 => n344, ZN => n21);
   U17 : AND2_X2 port map( A1 => n345, A2 => n334, ZN => n19);
   U18 : OR2_X1 port map( A1 => n1, A2 => n2, ZN => Y(9));
   U19 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U20 : AOI22_X1 port map( A1 => Q(105), A2 => n7, B1 => Q(201), B2 => n8, ZN 
                           => n6);
   U21 : AOI22_X1 port map( A1 => Q(169), A2 => n9, B1 => Q(41), B2 => n10, ZN 
                           => n5);
   U22 : AOI22_X1 port map( A1 => Q(9), A2 => n11, B1 => Q(73), B2 => n12, ZN 
                           => n4);
   U23 : AOI22_X1 port map( A1 => Q(233), A2 => n13, B1 => Q(137), B2 => n14, 
                           ZN => n3);
   U24 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           n1);
   U25 : AOI22_X1 port map( A1 => Q(329), A2 => n19, B1 => Q(425), B2 => n20, 
                           ZN => n18);
   U26 : AOI22_X1 port map( A1 => Q(393), A2 => n21, B1 => Q(265), B2 => n22, 
                           ZN => n17);
   U27 : AOI22_X1 port map( A1 => Q(361), A2 => n23, B1 => Q(297), B2 => n24, 
                           ZN => n16);
   U28 : AOI22_X1 port map( A1 => Q(489), A2 => n25, B1 => Q(457), B2 => n26, 
                           ZN => n15);
   U29 : OR2_X1 port map( A1 => n27, A2 => n28, ZN => Y(8));
   U30 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           n28);
   U31 : AOI22_X1 port map( A1 => Q(104), A2 => n7, B1 => Q(200), B2 => n8, ZN 
                           => n32);
   U32 : AOI22_X1 port map( A1 => Q(168), A2 => n9, B1 => Q(40), B2 => n10, ZN 
                           => n31);
   U33 : AOI22_X1 port map( A1 => Q(8), A2 => n11, B1 => Q(72), B2 => n12, ZN 
                           => n30);
   U34 : AOI22_X1 port map( A1 => Q(232), A2 => n13, B1 => Q(136), B2 => n14, 
                           ZN => n29);
   U35 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           n27);
   U36 : AOI22_X1 port map( A1 => Q(328), A2 => n19, B1 => Q(424), B2 => n20, 
                           ZN => n36);
   U37 : AOI22_X1 port map( A1 => Q(392), A2 => n21, B1 => Q(264), B2 => n22, 
                           ZN => n35);
   U38 : AOI22_X1 port map( A1 => Q(360), A2 => n23, B1 => Q(296), B2 => n24, 
                           ZN => n34);
   U39 : AOI22_X1 port map( A1 => Q(488), A2 => n25, B1 => Q(456), B2 => n26, 
                           ZN => n33);
   U40 : OR2_X1 port map( A1 => n37, A2 => n38, ZN => Y(7));
   U41 : NAND4_X1 port map( A1 => n39, A2 => n40, A3 => n41, A4 => n42, ZN => 
                           n38);
   U42 : AOI22_X1 port map( A1 => Q(103), A2 => n7, B1 => Q(199), B2 => n8, ZN 
                           => n42);
   U43 : AOI22_X1 port map( A1 => Q(167), A2 => n9, B1 => Q(39), B2 => n10, ZN 
                           => n41);
   U44 : AOI22_X1 port map( A1 => Q(7), A2 => n11, B1 => Q(71), B2 => n12, ZN 
                           => n40);
   U45 : AOI22_X1 port map( A1 => Q(231), A2 => n13, B1 => Q(135), B2 => n14, 
                           ZN => n39);
   U46 : NAND4_X1 port map( A1 => n43, A2 => n44, A3 => n45, A4 => n46, ZN => 
                           n37);
   U47 : AOI22_X1 port map( A1 => Q(327), A2 => n19, B1 => Q(423), B2 => n20, 
                           ZN => n46);
   U48 : AOI22_X1 port map( A1 => Q(391), A2 => n21, B1 => Q(263), B2 => n22, 
                           ZN => n45);
   U49 : AOI22_X1 port map( A1 => Q(359), A2 => n23, B1 => Q(295), B2 => n24, 
                           ZN => n44);
   U50 : AOI22_X1 port map( A1 => Q(487), A2 => n25, B1 => Q(455), B2 => n26, 
                           ZN => n43);
   U51 : OR2_X1 port map( A1 => n47, A2 => n48, ZN => Y(6));
   U52 : NAND4_X1 port map( A1 => n49, A2 => n50, A3 => n51, A4 => n52, ZN => 
                           n48);
   U53 : AOI22_X1 port map( A1 => Q(102), A2 => n7, B1 => Q(198), B2 => n8, ZN 
                           => n52);
   U54 : AOI22_X1 port map( A1 => Q(166), A2 => n9, B1 => Q(38), B2 => n10, ZN 
                           => n51);
   U55 : AOI22_X1 port map( A1 => Q(6), A2 => n11, B1 => Q(70), B2 => n12, ZN 
                           => n50);
   U56 : AOI22_X1 port map( A1 => Q(230), A2 => n13, B1 => Q(134), B2 => n14, 
                           ZN => n49);
   U57 : NAND4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           n47);
   U58 : AOI22_X1 port map( A1 => Q(326), A2 => n19, B1 => Q(422), B2 => n20, 
                           ZN => n56);
   U59 : AOI22_X1 port map( A1 => Q(390), A2 => n21, B1 => Q(262), B2 => n22, 
                           ZN => n55);
   U60 : AOI22_X1 port map( A1 => Q(358), A2 => n23, B1 => Q(294), B2 => n24, 
                           ZN => n54);
   U61 : AOI22_X1 port map( A1 => Q(486), A2 => n25, B1 => Q(454), B2 => n26, 
                           ZN => n53);
   U62 : OR2_X1 port map( A1 => n57, A2 => n58, ZN => Y(5));
   U63 : NAND4_X1 port map( A1 => n59, A2 => n60, A3 => n61, A4 => n62, ZN => 
                           n58);
   U64 : AOI22_X1 port map( A1 => Q(101), A2 => n7, B1 => Q(197), B2 => n8, ZN 
                           => n62);
   U65 : AOI22_X1 port map( A1 => Q(165), A2 => n9, B1 => Q(37), B2 => n10, ZN 
                           => n61);
   U66 : AOI22_X1 port map( A1 => Q(5), A2 => n11, B1 => Q(69), B2 => n12, ZN 
                           => n60);
   U67 : AOI22_X1 port map( A1 => Q(229), A2 => n13, B1 => Q(133), B2 => n14, 
                           ZN => n59);
   U68 : NAND4_X1 port map( A1 => n63, A2 => n64, A3 => n65, A4 => n66, ZN => 
                           n57);
   U69 : AOI22_X1 port map( A1 => Q(325), A2 => n19, B1 => Q(421), B2 => n20, 
                           ZN => n66);
   U70 : AOI22_X1 port map( A1 => Q(389), A2 => n21, B1 => Q(261), B2 => n22, 
                           ZN => n65);
   U71 : AOI22_X1 port map( A1 => Q(357), A2 => n23, B1 => Q(293), B2 => n24, 
                           ZN => n64);
   U72 : AOI22_X1 port map( A1 => Q(485), A2 => n25, B1 => Q(453), B2 => n26, 
                           ZN => n63);
   U73 : OR2_X1 port map( A1 => n67, A2 => n68, ZN => Y(4));
   U74 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n68);
   U75 : AOI22_X1 port map( A1 => Q(100), A2 => n7, B1 => Q(196), B2 => n8, ZN 
                           => n72);
   U76 : AOI22_X1 port map( A1 => Q(164), A2 => n9, B1 => Q(36), B2 => n10, ZN 
                           => n71);
   U77 : AOI22_X1 port map( A1 => Q(4), A2 => n11, B1 => Q(68), B2 => n12, ZN 
                           => n70);
   U78 : AOI22_X1 port map( A1 => Q(228), A2 => n13, B1 => Q(132), B2 => n14, 
                           ZN => n69);
   U79 : NAND4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           n67);
   U80 : AOI22_X1 port map( A1 => Q(324), A2 => n19, B1 => Q(420), B2 => n20, 
                           ZN => n76);
   U81 : AOI22_X1 port map( A1 => Q(388), A2 => n21, B1 => Q(260), B2 => n22, 
                           ZN => n75);
   U82 : AOI22_X1 port map( A1 => Q(356), A2 => n23, B1 => Q(292), B2 => n24, 
                           ZN => n74);
   U83 : AOI22_X1 port map( A1 => Q(484), A2 => n25, B1 => Q(452), B2 => n26, 
                           ZN => n73);
   U84 : OR2_X1 port map( A1 => n77, A2 => n78, ZN => Y(3));
   U85 : NAND4_X1 port map( A1 => n79, A2 => n80, A3 => n81, A4 => n82, ZN => 
                           n78);
   U86 : AOI22_X1 port map( A1 => Q(99), A2 => n7, B1 => Q(195), B2 => n8, ZN 
                           => n82);
   U87 : AOI22_X1 port map( A1 => Q(163), A2 => n9, B1 => Q(35), B2 => n10, ZN 
                           => n81);
   U88 : AOI22_X1 port map( A1 => Q(3), A2 => n11, B1 => Q(67), B2 => n12, ZN 
                           => n80);
   U89 : AOI22_X1 port map( A1 => Q(227), A2 => n13, B1 => Q(131), B2 => n14, 
                           ZN => n79);
   U90 : NAND4_X1 port map( A1 => n83, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           n77);
   U91 : AOI22_X1 port map( A1 => Q(323), A2 => n19, B1 => Q(419), B2 => n20, 
                           ZN => n86);
   U92 : AOI22_X1 port map( A1 => Q(387), A2 => n21, B1 => Q(259), B2 => n22, 
                           ZN => n85);
   U93 : AOI22_X1 port map( A1 => Q(355), A2 => n23, B1 => Q(291), B2 => n24, 
                           ZN => n84);
   U94 : AOI22_X1 port map( A1 => Q(483), A2 => n25, B1 => Q(451), B2 => n26, 
                           ZN => n83);
   U95 : OR2_X1 port map( A1 => n87, A2 => n88, ZN => Y(31));
   U96 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           n88);
   U97 : AOI22_X1 port map( A1 => Q(127), A2 => n7, B1 => Q(223), B2 => n8, ZN 
                           => n92);
   U98 : AOI22_X1 port map( A1 => Q(191), A2 => n9, B1 => Q(63), B2 => n10, ZN 
                           => n91);
   U99 : AOI22_X1 port map( A1 => Q(31), A2 => n11, B1 => Q(95), B2 => n12, ZN 
                           => n90);
   U100 : AOI22_X1 port map( A1 => Q(255), A2 => n13, B1 => Q(159), B2 => n14, 
                           ZN => n89);
   U101 : NAND4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           n87);
   U102 : AOI22_X1 port map( A1 => Q(351), A2 => n19, B1 => Q(447), B2 => n20, 
                           ZN => n96);
   U103 : AOI22_X1 port map( A1 => Q(415), A2 => n21, B1 => Q(287), B2 => n22, 
                           ZN => n95);
   U104 : AOI22_X1 port map( A1 => Q(383), A2 => n23, B1 => Q(319), B2 => n24, 
                           ZN => n94);
   U105 : AOI22_X1 port map( A1 => Q(511), A2 => n25, B1 => Q(479), B2 => n26, 
                           ZN => n93);
   U106 : OR2_X1 port map( A1 => n97, A2 => n98, ZN => Y(30));
   U107 : NAND4_X1 port map( A1 => n99, A2 => n100, A3 => n101, A4 => n102, ZN 
                           => n98);
   U108 : AOI22_X1 port map( A1 => Q(126), A2 => n7, B1 => Q(222), B2 => n8, ZN
                           => n102);
   U109 : AOI22_X1 port map( A1 => Q(190), A2 => n9, B1 => Q(62), B2 => n10, ZN
                           => n101);
   U110 : AOI22_X1 port map( A1 => Q(30), A2 => n11, B1 => Q(94), B2 => n12, ZN
                           => n100);
   U111 : AOI22_X1 port map( A1 => Q(254), A2 => n13, B1 => Q(158), B2 => n14, 
                           ZN => n99);
   U112 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN
                           => n97);
   U113 : AOI22_X1 port map( A1 => Q(350), A2 => n19, B1 => Q(446), B2 => n20, 
                           ZN => n106);
   U114 : AOI22_X1 port map( A1 => Q(414), A2 => n21, B1 => Q(286), B2 => n22, 
                           ZN => n105);
   U115 : AOI22_X1 port map( A1 => Q(382), A2 => n23, B1 => Q(318), B2 => n24, 
                           ZN => n104);
   U116 : AOI22_X1 port map( A1 => Q(510), A2 => n25, B1 => Q(478), B2 => n26, 
                           ZN => n103);
   U117 : OR2_X1 port map( A1 => n107, A2 => n108, ZN => Y(2));
   U118 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => n108);
   U119 : AOI22_X1 port map( A1 => Q(98), A2 => n7, B1 => Q(194), B2 => n8, ZN 
                           => n112);
   U120 : AOI22_X1 port map( A1 => Q(162), A2 => n9, B1 => Q(34), B2 => n10, ZN
                           => n111);
   U121 : AOI22_X1 port map( A1 => Q(2), A2 => n11, B1 => Q(66), B2 => n12, ZN 
                           => n110);
   U122 : AOI22_X1 port map( A1 => Q(226), A2 => n13, B1 => Q(130), B2 => n14, 
                           ZN => n109);
   U123 : NAND4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN
                           => n107);
   U124 : AOI22_X1 port map( A1 => Q(322), A2 => n19, B1 => Q(418), B2 => n20, 
                           ZN => n116);
   U125 : AOI22_X1 port map( A1 => Q(386), A2 => n21, B1 => Q(258), B2 => n22, 
                           ZN => n115);
   U126 : AOI22_X1 port map( A1 => Q(354), A2 => n23, B1 => Q(290), B2 => n24, 
                           ZN => n114);
   U127 : AOI22_X1 port map( A1 => Q(482), A2 => n25, B1 => Q(450), B2 => n26, 
                           ZN => n113);
   U128 : OR2_X1 port map( A1 => n117, A2 => n118, ZN => Y(29));
   U129 : NAND4_X1 port map( A1 => n119, A2 => n120, A3 => n121, A4 => n122, ZN
                           => n118);
   U130 : AOI22_X1 port map( A1 => Q(125), A2 => n7, B1 => Q(221), B2 => n8, ZN
                           => n122);
   U131 : AOI22_X1 port map( A1 => Q(189), A2 => n9, B1 => Q(61), B2 => n10, ZN
                           => n121);
   U132 : AOI22_X1 port map( A1 => Q(29), A2 => n11, B1 => Q(93), B2 => n12, ZN
                           => n120);
   U133 : AOI22_X1 port map( A1 => Q(253), A2 => n13, B1 => Q(157), B2 => n14, 
                           ZN => n119);
   U134 : NAND4_X1 port map( A1 => n123, A2 => n124, A3 => n125, A4 => n126, ZN
                           => n117);
   U135 : AOI22_X1 port map( A1 => Q(349), A2 => n19, B1 => Q(445), B2 => n20, 
                           ZN => n126);
   U136 : AOI22_X1 port map( A1 => Q(413), A2 => n21, B1 => Q(285), B2 => n22, 
                           ZN => n125);
   U137 : AOI22_X1 port map( A1 => Q(381), A2 => n23, B1 => Q(317), B2 => n24, 
                           ZN => n124);
   U138 : AOI22_X1 port map( A1 => Q(509), A2 => n25, B1 => Q(477), B2 => n26, 
                           ZN => n123);
   U139 : OR2_X1 port map( A1 => n127, A2 => n128, ZN => Y(28));
   U140 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => n128);
   U141 : AOI22_X1 port map( A1 => Q(124), A2 => n7, B1 => Q(220), B2 => n8, ZN
                           => n132);
   U142 : AOI22_X1 port map( A1 => Q(188), A2 => n9, B1 => Q(60), B2 => n10, ZN
                           => n131);
   U143 : AOI22_X1 port map( A1 => Q(28), A2 => n11, B1 => Q(92), B2 => n12, ZN
                           => n130);
   U144 : AOI22_X1 port map( A1 => Q(252), A2 => n13, B1 => Q(156), B2 => n14, 
                           ZN => n129);
   U145 : NAND4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN
                           => n127);
   U146 : AOI22_X1 port map( A1 => Q(348), A2 => n19, B1 => Q(444), B2 => n20, 
                           ZN => n136);
   U147 : AOI22_X1 port map( A1 => Q(412), A2 => n21, B1 => Q(284), B2 => n22, 
                           ZN => n135);
   U148 : AOI22_X1 port map( A1 => Q(380), A2 => n23, B1 => Q(316), B2 => n24, 
                           ZN => n134);
   U149 : AOI22_X1 port map( A1 => Q(508), A2 => n25, B1 => Q(476), B2 => n26, 
                           ZN => n133);
   U150 : OR2_X1 port map( A1 => n137, A2 => n138, ZN => Y(27));
   U151 : NAND4_X1 port map( A1 => n139, A2 => n140, A3 => n141, A4 => n142, ZN
                           => n138);
   U152 : AOI22_X1 port map( A1 => Q(123), A2 => n7, B1 => Q(219), B2 => n8, ZN
                           => n142);
   U153 : AOI22_X1 port map( A1 => Q(187), A2 => n9, B1 => Q(59), B2 => n10, ZN
                           => n141);
   U154 : AOI22_X1 port map( A1 => Q(27), A2 => n11, B1 => Q(91), B2 => n12, ZN
                           => n140);
   U155 : AOI22_X1 port map( A1 => Q(251), A2 => n13, B1 => Q(155), B2 => n14, 
                           ZN => n139);
   U156 : NAND4_X1 port map( A1 => n143, A2 => n144, A3 => n145, A4 => n146, ZN
                           => n137);
   U157 : AOI22_X1 port map( A1 => Q(347), A2 => n19, B1 => Q(443), B2 => n20, 
                           ZN => n146);
   U158 : AOI22_X1 port map( A1 => Q(411), A2 => n21, B1 => Q(283), B2 => n22, 
                           ZN => n145);
   U159 : AOI22_X1 port map( A1 => Q(379), A2 => n23, B1 => Q(315), B2 => n24, 
                           ZN => n144);
   U160 : AOI22_X1 port map( A1 => Q(507), A2 => n25, B1 => Q(475), B2 => n26, 
                           ZN => n143);
   U161 : OR2_X1 port map( A1 => n147, A2 => n148, ZN => Y(26));
   U162 : NAND4_X1 port map( A1 => n149, A2 => n150, A3 => n151, A4 => n152, ZN
                           => n148);
   U163 : AOI22_X1 port map( A1 => Q(122), A2 => n7, B1 => Q(218), B2 => n8, ZN
                           => n152);
   U164 : AOI22_X1 port map( A1 => Q(186), A2 => n9, B1 => Q(58), B2 => n10, ZN
                           => n151);
   U165 : AOI22_X1 port map( A1 => Q(26), A2 => n11, B1 => Q(90), B2 => n12, ZN
                           => n150);
   U166 : AOI22_X1 port map( A1 => Q(250), A2 => n13, B1 => Q(154), B2 => n14, 
                           ZN => n149);
   U167 : NAND4_X1 port map( A1 => n153, A2 => n154, A3 => n155, A4 => n156, ZN
                           => n147);
   U168 : AOI22_X1 port map( A1 => Q(346), A2 => n19, B1 => Q(442), B2 => n20, 
                           ZN => n156);
   U169 : AOI22_X1 port map( A1 => Q(410), A2 => n21, B1 => Q(282), B2 => n22, 
                           ZN => n155);
   U170 : AOI22_X1 port map( A1 => Q(378), A2 => n23, B1 => Q(314), B2 => n24, 
                           ZN => n154);
   U171 : AOI22_X1 port map( A1 => Q(506), A2 => n25, B1 => Q(474), B2 => n26, 
                           ZN => n153);
   U172 : OR2_X1 port map( A1 => n157, A2 => n158, ZN => Y(25));
   U173 : NAND4_X1 port map( A1 => n159, A2 => n160, A3 => n161, A4 => n162, ZN
                           => n158);
   U174 : AOI22_X1 port map( A1 => Q(121), A2 => n7, B1 => Q(217), B2 => n8, ZN
                           => n162);
   U175 : AOI22_X1 port map( A1 => Q(185), A2 => n9, B1 => Q(57), B2 => n10, ZN
                           => n161);
   U176 : AOI22_X1 port map( A1 => Q(25), A2 => n11, B1 => Q(89), B2 => n12, ZN
                           => n160);
   U177 : AOI22_X1 port map( A1 => Q(249), A2 => n13, B1 => Q(153), B2 => n14, 
                           ZN => n159);
   U178 : NAND4_X1 port map( A1 => n163, A2 => n164, A3 => n165, A4 => n166, ZN
                           => n157);
   U179 : AOI22_X1 port map( A1 => Q(345), A2 => n19, B1 => Q(441), B2 => n20, 
                           ZN => n166);
   U180 : AOI22_X1 port map( A1 => Q(409), A2 => n21, B1 => Q(281), B2 => n22, 
                           ZN => n165);
   U181 : AOI22_X1 port map( A1 => Q(377), A2 => n23, B1 => Q(313), B2 => n24, 
                           ZN => n164);
   U182 : AOI22_X1 port map( A1 => Q(505), A2 => n25, B1 => Q(473), B2 => n26, 
                           ZN => n163);
   U183 : OR2_X1 port map( A1 => n167, A2 => n168, ZN => Y(24));
   U184 : NAND4_X1 port map( A1 => n169, A2 => n170, A3 => n171, A4 => n172, ZN
                           => n168);
   U185 : AOI22_X1 port map( A1 => Q(120), A2 => n7, B1 => Q(216), B2 => n8, ZN
                           => n172);
   U186 : AOI22_X1 port map( A1 => Q(184), A2 => n9, B1 => Q(56), B2 => n10, ZN
                           => n171);
   U187 : AOI22_X1 port map( A1 => Q(24), A2 => n11, B1 => Q(88), B2 => n12, ZN
                           => n170);
   U188 : AOI22_X1 port map( A1 => Q(248), A2 => n13, B1 => Q(152), B2 => n14, 
                           ZN => n169);
   U189 : NAND4_X1 port map( A1 => n173, A2 => n174, A3 => n175, A4 => n176, ZN
                           => n167);
   U190 : AOI22_X1 port map( A1 => Q(344), A2 => n19, B1 => Q(440), B2 => n20, 
                           ZN => n176);
   U191 : AOI22_X1 port map( A1 => Q(408), A2 => n21, B1 => Q(280), B2 => n22, 
                           ZN => n175);
   U192 : AOI22_X1 port map( A1 => Q(376), A2 => n23, B1 => Q(312), B2 => n24, 
                           ZN => n174);
   U193 : AOI22_X1 port map( A1 => Q(504), A2 => n25, B1 => Q(472), B2 => n26, 
                           ZN => n173);
   U194 : OR2_X1 port map( A1 => n177, A2 => n178, ZN => Y(23));
   U195 : NAND4_X1 port map( A1 => n179, A2 => n180, A3 => n181, A4 => n182, ZN
                           => n178);
   U196 : AOI22_X1 port map( A1 => Q(119), A2 => n7, B1 => Q(215), B2 => n8, ZN
                           => n182);
   U197 : AOI22_X1 port map( A1 => Q(183), A2 => n9, B1 => Q(55), B2 => n10, ZN
                           => n181);
   U198 : AOI22_X1 port map( A1 => Q(23), A2 => n11, B1 => Q(87), B2 => n12, ZN
                           => n180);
   U199 : AOI22_X1 port map( A1 => Q(247), A2 => n13, B1 => Q(151), B2 => n14, 
                           ZN => n179);
   U200 : NAND4_X1 port map( A1 => n183, A2 => n184, A3 => n185, A4 => n186, ZN
                           => n177);
   U201 : AOI22_X1 port map( A1 => Q(343), A2 => n19, B1 => Q(439), B2 => n20, 
                           ZN => n186);
   U202 : AOI22_X1 port map( A1 => Q(407), A2 => n21, B1 => Q(279), B2 => n22, 
                           ZN => n185);
   U203 : AOI22_X1 port map( A1 => Q(375), A2 => n23, B1 => Q(311), B2 => n24, 
                           ZN => n184);
   U204 : AOI22_X1 port map( A1 => Q(503), A2 => n25, B1 => Q(471), B2 => n26, 
                           ZN => n183);
   U205 : OR2_X1 port map( A1 => n187, A2 => n188, ZN => Y(22));
   U206 : NAND4_X1 port map( A1 => n189, A2 => n190, A3 => n191, A4 => n192, ZN
                           => n188);
   U207 : AOI22_X1 port map( A1 => Q(118), A2 => n7, B1 => Q(214), B2 => n8, ZN
                           => n192);
   U208 : AOI22_X1 port map( A1 => Q(182), A2 => n9, B1 => Q(54), B2 => n10, ZN
                           => n191);
   U209 : AOI22_X1 port map( A1 => Q(22), A2 => n11, B1 => Q(86), B2 => n12, ZN
                           => n190);
   U210 : AOI22_X1 port map( A1 => Q(246), A2 => n13, B1 => Q(150), B2 => n14, 
                           ZN => n189);
   U211 : NAND4_X1 port map( A1 => n193, A2 => n194, A3 => n195, A4 => n196, ZN
                           => n187);
   U212 : AOI22_X1 port map( A1 => Q(342), A2 => n19, B1 => Q(438), B2 => n20, 
                           ZN => n196);
   U213 : AOI22_X1 port map( A1 => Q(406), A2 => n21, B1 => Q(278), B2 => n22, 
                           ZN => n195);
   U214 : AOI22_X1 port map( A1 => Q(374), A2 => n23, B1 => Q(310), B2 => n24, 
                           ZN => n194);
   U215 : AOI22_X1 port map( A1 => Q(502), A2 => n25, B1 => Q(470), B2 => n26, 
                           ZN => n193);
   U216 : OR2_X1 port map( A1 => n197, A2 => n198, ZN => Y(21));
   U217 : NAND4_X1 port map( A1 => n199, A2 => n200, A3 => n201, A4 => n202, ZN
                           => n198);
   U218 : AOI22_X1 port map( A1 => Q(117), A2 => n7, B1 => Q(213), B2 => n8, ZN
                           => n202);
   U219 : AOI22_X1 port map( A1 => Q(181), A2 => n9, B1 => Q(53), B2 => n10, ZN
                           => n201);
   U220 : AOI22_X1 port map( A1 => Q(21), A2 => n11, B1 => Q(85), B2 => n12, ZN
                           => n200);
   U221 : AOI22_X1 port map( A1 => Q(245), A2 => n13, B1 => Q(149), B2 => n14, 
                           ZN => n199);
   U222 : NAND4_X1 port map( A1 => n203, A2 => n204, A3 => n205, A4 => n206, ZN
                           => n197);
   U223 : AOI22_X1 port map( A1 => Q(341), A2 => n19, B1 => Q(437), B2 => n20, 
                           ZN => n206);
   U224 : AOI22_X1 port map( A1 => Q(405), A2 => n21, B1 => Q(277), B2 => n22, 
                           ZN => n205);
   U225 : AOI22_X1 port map( A1 => Q(373), A2 => n23, B1 => Q(309), B2 => n24, 
                           ZN => n204);
   U226 : AOI22_X1 port map( A1 => Q(501), A2 => n25, B1 => Q(469), B2 => n26, 
                           ZN => n203);
   U227 : OR2_X1 port map( A1 => n207, A2 => n208, ZN => Y(20));
   U228 : NAND4_X1 port map( A1 => n209, A2 => n210, A3 => n211, A4 => n212, ZN
                           => n208);
   U229 : AOI22_X1 port map( A1 => Q(116), A2 => n7, B1 => Q(212), B2 => n8, ZN
                           => n212);
   U230 : AOI22_X1 port map( A1 => Q(180), A2 => n9, B1 => Q(52), B2 => n10, ZN
                           => n211);
   U231 : AOI22_X1 port map( A1 => Q(20), A2 => n11, B1 => Q(84), B2 => n12, ZN
                           => n210);
   U232 : AOI22_X1 port map( A1 => Q(244), A2 => n13, B1 => Q(148), B2 => n14, 
                           ZN => n209);
   U233 : NAND4_X1 port map( A1 => n213, A2 => n214, A3 => n215, A4 => n216, ZN
                           => n207);
   U234 : AOI22_X1 port map( A1 => Q(340), A2 => n19, B1 => Q(436), B2 => n20, 
                           ZN => n216);
   U235 : AOI22_X1 port map( A1 => Q(404), A2 => n21, B1 => Q(276), B2 => n22, 
                           ZN => n215);
   U236 : AOI22_X1 port map( A1 => Q(372), A2 => n23, B1 => Q(308), B2 => n24, 
                           ZN => n214);
   U237 : AOI22_X1 port map( A1 => Q(500), A2 => n25, B1 => Q(468), B2 => n26, 
                           ZN => n213);
   U238 : OR2_X1 port map( A1 => n217, A2 => n218, ZN => Y(1));
   U239 : NAND4_X1 port map( A1 => n219, A2 => n220, A3 => n221, A4 => n222, ZN
                           => n218);
   U240 : AOI22_X1 port map( A1 => Q(97), A2 => n7, B1 => Q(193), B2 => n8, ZN 
                           => n222);
   U241 : AOI22_X1 port map( A1 => Q(161), A2 => n9, B1 => Q(33), B2 => n10, ZN
                           => n221);
   U242 : AOI22_X1 port map( A1 => Q(1), A2 => n11, B1 => Q(65), B2 => n12, ZN 
                           => n220);
   U243 : AOI22_X1 port map( A1 => Q(225), A2 => n13, B1 => Q(129), B2 => n14, 
                           ZN => n219);
   U244 : NAND4_X1 port map( A1 => n223, A2 => n224, A3 => n225, A4 => n226, ZN
                           => n217);
   U245 : AOI22_X1 port map( A1 => Q(321), A2 => n19, B1 => Q(417), B2 => n20, 
                           ZN => n226);
   U246 : AOI22_X1 port map( A1 => Q(385), A2 => n21, B1 => Q(257), B2 => n22, 
                           ZN => n225);
   U247 : AOI22_X1 port map( A1 => Q(353), A2 => n23, B1 => Q(289), B2 => n24, 
                           ZN => n224);
   U248 : AOI22_X1 port map( A1 => Q(481), A2 => n25, B1 => Q(449), B2 => n26, 
                           ZN => n223);
   U249 : OR2_X1 port map( A1 => n227, A2 => n228, ZN => Y(19));
   U250 : NAND4_X1 port map( A1 => n229, A2 => n230, A3 => n231, A4 => n232, ZN
                           => n228);
   U251 : AOI22_X1 port map( A1 => Q(115), A2 => n7, B1 => Q(211), B2 => n8, ZN
                           => n232);
   U252 : AOI22_X1 port map( A1 => Q(179), A2 => n9, B1 => Q(51), B2 => n10, ZN
                           => n231);
   U253 : AOI22_X1 port map( A1 => Q(19), A2 => n11, B1 => Q(83), B2 => n12, ZN
                           => n230);
   U254 : AOI22_X1 port map( A1 => Q(243), A2 => n13, B1 => Q(147), B2 => n14, 
                           ZN => n229);
   U255 : NAND4_X1 port map( A1 => n233, A2 => n234, A3 => n235, A4 => n236, ZN
                           => n227);
   U256 : AOI22_X1 port map( A1 => Q(339), A2 => n19, B1 => Q(435), B2 => n20, 
                           ZN => n236);
   U257 : AOI22_X1 port map( A1 => Q(403), A2 => n21, B1 => Q(275), B2 => n22, 
                           ZN => n235);
   U258 : AOI22_X1 port map( A1 => Q(371), A2 => n23, B1 => Q(307), B2 => n24, 
                           ZN => n234);
   U259 : AOI22_X1 port map( A1 => Q(499), A2 => n25, B1 => Q(467), B2 => n26, 
                           ZN => n233);
   U260 : OR2_X1 port map( A1 => n237, A2 => n238, ZN => Y(18));
   U261 : NAND4_X1 port map( A1 => n239, A2 => n240, A3 => n241, A4 => n242, ZN
                           => n238);
   U262 : AOI22_X1 port map( A1 => Q(114), A2 => n7, B1 => Q(210), B2 => n8, ZN
                           => n242);
   U263 : AOI22_X1 port map( A1 => Q(178), A2 => n9, B1 => Q(50), B2 => n10, ZN
                           => n241);
   U264 : AOI22_X1 port map( A1 => Q(18), A2 => n11, B1 => Q(82), B2 => n12, ZN
                           => n240);
   U265 : AOI22_X1 port map( A1 => Q(242), A2 => n13, B1 => Q(146), B2 => n14, 
                           ZN => n239);
   U266 : NAND4_X1 port map( A1 => n243, A2 => n244, A3 => n245, A4 => n246, ZN
                           => n237);
   U267 : AOI22_X1 port map( A1 => Q(338), A2 => n19, B1 => Q(434), B2 => n20, 
                           ZN => n246);
   U268 : AOI22_X1 port map( A1 => Q(402), A2 => n21, B1 => Q(274), B2 => n22, 
                           ZN => n245);
   U269 : AOI22_X1 port map( A1 => Q(370), A2 => n23, B1 => Q(306), B2 => n24, 
                           ZN => n244);
   U270 : AOI22_X1 port map( A1 => Q(498), A2 => n25, B1 => Q(466), B2 => n26, 
                           ZN => n243);
   U271 : OR2_X1 port map( A1 => n247, A2 => n248, ZN => Y(17));
   U272 : NAND4_X1 port map( A1 => n249, A2 => n250, A3 => n251, A4 => n252, ZN
                           => n248);
   U273 : AOI22_X1 port map( A1 => Q(113), A2 => n7, B1 => Q(209), B2 => n8, ZN
                           => n252);
   U274 : AOI22_X1 port map( A1 => Q(177), A2 => n9, B1 => Q(49), B2 => n10, ZN
                           => n251);
   U275 : AOI22_X1 port map( A1 => Q(17), A2 => n11, B1 => Q(81), B2 => n12, ZN
                           => n250);
   U276 : AOI22_X1 port map( A1 => Q(241), A2 => n13, B1 => Q(145), B2 => n14, 
                           ZN => n249);
   U277 : NAND4_X1 port map( A1 => n253, A2 => n254, A3 => n255, A4 => n256, ZN
                           => n247);
   U278 : AOI22_X1 port map( A1 => Q(337), A2 => n19, B1 => Q(433), B2 => n20, 
                           ZN => n256);
   U279 : AOI22_X1 port map( A1 => Q(401), A2 => n21, B1 => Q(273), B2 => n22, 
                           ZN => n255);
   U280 : AOI22_X1 port map( A1 => Q(369), A2 => n23, B1 => Q(305), B2 => n24, 
                           ZN => n254);
   U281 : AOI22_X1 port map( A1 => Q(497), A2 => n25, B1 => Q(465), B2 => n26, 
                           ZN => n253);
   U282 : OR2_X1 port map( A1 => n257, A2 => n258, ZN => Y(16));
   U283 : NAND4_X1 port map( A1 => n259, A2 => n260, A3 => n261, A4 => n262, ZN
                           => n258);
   U284 : AOI22_X1 port map( A1 => Q(112), A2 => n7, B1 => Q(208), B2 => n8, ZN
                           => n262);
   U285 : AOI22_X1 port map( A1 => Q(176), A2 => n9, B1 => Q(48), B2 => n10, ZN
                           => n261);
   U286 : AOI22_X1 port map( A1 => Q(16), A2 => n11, B1 => Q(80), B2 => n12, ZN
                           => n260);
   U287 : AOI22_X1 port map( A1 => Q(240), A2 => n13, B1 => Q(144), B2 => n14, 
                           ZN => n259);
   U288 : NAND4_X1 port map( A1 => n263, A2 => n264, A3 => n265, A4 => n266, ZN
                           => n257);
   U289 : AOI22_X1 port map( A1 => Q(336), A2 => n19, B1 => Q(432), B2 => n20, 
                           ZN => n266);
   U290 : AOI22_X1 port map( A1 => Q(400), A2 => n21, B1 => Q(272), B2 => n22, 
                           ZN => n265);
   U291 : AOI22_X1 port map( A1 => Q(368), A2 => n23, B1 => Q(304), B2 => n24, 
                           ZN => n264);
   U292 : AOI22_X1 port map( A1 => Q(496), A2 => n25, B1 => Q(464), B2 => n26, 
                           ZN => n263);
   U293 : OR2_X1 port map( A1 => n267, A2 => n268, ZN => Y(15));
   U294 : NAND4_X1 port map( A1 => n269, A2 => n270, A3 => n271, A4 => n272, ZN
                           => n268);
   U295 : AOI22_X1 port map( A1 => Q(111), A2 => n7, B1 => Q(207), B2 => n8, ZN
                           => n272);
   U296 : AOI22_X1 port map( A1 => Q(175), A2 => n9, B1 => Q(47), B2 => n10, ZN
                           => n271);
   U297 : AOI22_X1 port map( A1 => Q(15), A2 => n11, B1 => Q(79), B2 => n12, ZN
                           => n270);
   U298 : AOI22_X1 port map( A1 => Q(239), A2 => n13, B1 => Q(143), B2 => n14, 
                           ZN => n269);
   U299 : NAND4_X1 port map( A1 => n273, A2 => n274, A3 => n275, A4 => n276, ZN
                           => n267);
   U300 : AOI22_X1 port map( A1 => Q(335), A2 => n19, B1 => Q(431), B2 => n20, 
                           ZN => n276);
   U301 : AOI22_X1 port map( A1 => Q(399), A2 => n21, B1 => Q(271), B2 => n22, 
                           ZN => n275);
   U302 : AOI22_X1 port map( A1 => Q(367), A2 => n23, B1 => Q(303), B2 => n24, 
                           ZN => n274);
   U303 : AOI22_X1 port map( A1 => Q(495), A2 => n25, B1 => Q(463), B2 => n26, 
                           ZN => n273);
   U304 : OR2_X1 port map( A1 => n277, A2 => n278, ZN => Y(14));
   U305 : NAND4_X1 port map( A1 => n279, A2 => n280, A3 => n281, A4 => n282, ZN
                           => n278);
   U306 : AOI22_X1 port map( A1 => Q(110), A2 => n7, B1 => Q(206), B2 => n8, ZN
                           => n282);
   U307 : AOI22_X1 port map( A1 => Q(174), A2 => n9, B1 => Q(46), B2 => n10, ZN
                           => n281);
   U308 : AOI22_X1 port map( A1 => Q(14), A2 => n11, B1 => Q(78), B2 => n12, ZN
                           => n280);
   U309 : AOI22_X1 port map( A1 => Q(238), A2 => n13, B1 => Q(142), B2 => n14, 
                           ZN => n279);
   U310 : NAND4_X1 port map( A1 => n283, A2 => n284, A3 => n285, A4 => n286, ZN
                           => n277);
   U311 : AOI22_X1 port map( A1 => Q(334), A2 => n19, B1 => Q(430), B2 => n20, 
                           ZN => n286);
   U312 : AOI22_X1 port map( A1 => Q(398), A2 => n21, B1 => Q(270), B2 => n22, 
                           ZN => n285);
   U313 : AOI22_X1 port map( A1 => Q(366), A2 => n23, B1 => Q(302), B2 => n24, 
                           ZN => n284);
   U314 : AOI22_X1 port map( A1 => Q(494), A2 => n25, B1 => Q(462), B2 => n26, 
                           ZN => n283);
   U315 : OR2_X1 port map( A1 => n287, A2 => n288, ZN => Y(13));
   U316 : NAND4_X1 port map( A1 => n289, A2 => n290, A3 => n291, A4 => n292, ZN
                           => n288);
   U317 : AOI22_X1 port map( A1 => Q(109), A2 => n7, B1 => Q(205), B2 => n8, ZN
                           => n292);
   U318 : AOI22_X1 port map( A1 => Q(173), A2 => n9, B1 => Q(45), B2 => n10, ZN
                           => n291);
   U319 : AOI22_X1 port map( A1 => Q(13), A2 => n11, B1 => Q(77), B2 => n12, ZN
                           => n290);
   U320 : AOI22_X1 port map( A1 => Q(237), A2 => n13, B1 => Q(141), B2 => n14, 
                           ZN => n289);
   U321 : NAND4_X1 port map( A1 => n293, A2 => n294, A3 => n295, A4 => n296, ZN
                           => n287);
   U322 : AOI22_X1 port map( A1 => Q(333), A2 => n19, B1 => Q(429), B2 => n20, 
                           ZN => n296);
   U323 : AOI22_X1 port map( A1 => Q(397), A2 => n21, B1 => Q(269), B2 => n22, 
                           ZN => n295);
   U324 : AOI22_X1 port map( A1 => Q(365), A2 => n23, B1 => Q(301), B2 => n24, 
                           ZN => n294);
   U325 : AOI22_X1 port map( A1 => Q(493), A2 => n25, B1 => Q(461), B2 => n26, 
                           ZN => n293);
   U326 : OR2_X1 port map( A1 => n297, A2 => n298, ZN => Y(12));
   U327 : NAND4_X1 port map( A1 => n299, A2 => n300, A3 => n301, A4 => n302, ZN
                           => n298);
   U328 : AOI22_X1 port map( A1 => Q(108), A2 => n7, B1 => Q(204), B2 => n8, ZN
                           => n302);
   U329 : AOI22_X1 port map( A1 => Q(172), A2 => n9, B1 => Q(44), B2 => n10, ZN
                           => n301);
   U330 : AOI22_X1 port map( A1 => Q(12), A2 => n11, B1 => Q(76), B2 => n12, ZN
                           => n300);
   U331 : AOI22_X1 port map( A1 => Q(236), A2 => n13, B1 => Q(140), B2 => n14, 
                           ZN => n299);
   U332 : NAND4_X1 port map( A1 => n303, A2 => n304, A3 => n305, A4 => n306, ZN
                           => n297);
   U333 : AOI22_X1 port map( A1 => Q(332), A2 => n19, B1 => Q(428), B2 => n20, 
                           ZN => n306);
   U334 : AOI22_X1 port map( A1 => Q(396), A2 => n21, B1 => Q(268), B2 => n22, 
                           ZN => n305);
   U335 : AOI22_X1 port map( A1 => Q(364), A2 => n23, B1 => Q(300), B2 => n24, 
                           ZN => n304);
   U336 : AOI22_X1 port map( A1 => Q(492), A2 => n25, B1 => Q(460), B2 => n26, 
                           ZN => n303);
   U337 : OR2_X1 port map( A1 => n307, A2 => n308, ZN => Y(11));
   U338 : NAND4_X1 port map( A1 => n309, A2 => n310, A3 => n311, A4 => n312, ZN
                           => n308);
   U339 : AOI22_X1 port map( A1 => Q(107), A2 => n7, B1 => Q(203), B2 => n8, ZN
                           => n312);
   U340 : AOI22_X1 port map( A1 => Q(171), A2 => n9, B1 => Q(43), B2 => n10, ZN
                           => n311);
   U341 : AOI22_X1 port map( A1 => Q(11), A2 => n11, B1 => Q(75), B2 => n12, ZN
                           => n310);
   U342 : AOI22_X1 port map( A1 => Q(235), A2 => n13, B1 => Q(139), B2 => n14, 
                           ZN => n309);
   U343 : NAND4_X1 port map( A1 => n313, A2 => n314, A3 => n315, A4 => n316, ZN
                           => n307);
   U344 : AOI22_X1 port map( A1 => Q(331), A2 => n19, B1 => Q(427), B2 => n20, 
                           ZN => n316);
   U345 : AOI22_X1 port map( A1 => Q(395), A2 => n21, B1 => Q(267), B2 => n22, 
                           ZN => n315);
   U346 : AOI22_X1 port map( A1 => Q(363), A2 => n23, B1 => Q(299), B2 => n24, 
                           ZN => n314);
   U347 : AOI22_X1 port map( A1 => Q(491), A2 => n25, B1 => Q(459), B2 => n26, 
                           ZN => n313);
   U348 : OR2_X1 port map( A1 => n317, A2 => n318, ZN => Y(10));
   U349 : NAND4_X1 port map( A1 => n319, A2 => n320, A3 => n321, A4 => n322, ZN
                           => n318);
   U350 : AOI22_X1 port map( A1 => Q(106), A2 => n7, B1 => Q(202), B2 => n8, ZN
                           => n322);
   U351 : AOI22_X1 port map( A1 => Q(170), A2 => n9, B1 => Q(42), B2 => n10, ZN
                           => n321);
   U352 : AOI22_X1 port map( A1 => Q(10), A2 => n11, B1 => Q(74), B2 => n12, ZN
                           => n320);
   U353 : AOI22_X1 port map( A1 => Q(234), A2 => n13, B1 => Q(138), B2 => n14, 
                           ZN => n319);
   U354 : NAND4_X1 port map( A1 => n323, A2 => n324, A3 => n325, A4 => n326, ZN
                           => n317);
   U355 : AOI22_X1 port map( A1 => Q(330), A2 => n19, B1 => Q(426), B2 => n20, 
                           ZN => n326);
   U356 : AOI22_X1 port map( A1 => Q(394), A2 => n21, B1 => Q(266), B2 => n22, 
                           ZN => n325);
   U357 : AOI22_X1 port map( A1 => Q(362), A2 => n23, B1 => Q(298), B2 => n24, 
                           ZN => n324);
   U358 : AOI22_X1 port map( A1 => Q(490), A2 => n25, B1 => Q(458), B2 => n26, 
                           ZN => n323);
   U359 : OR2_X1 port map( A1 => n327, A2 => n328, ZN => Y(0));
   U360 : NAND4_X1 port map( A1 => n329, A2 => n330, A3 => n331, A4 => n332, ZN
                           => n328);
   U361 : AOI22_X1 port map( A1 => Q(96), A2 => n7, B1 => Q(192), B2 => n8, ZN 
                           => n332);
   U362 : AOI22_X1 port map( A1 => Q(160), A2 => n9, B1 => Q(32), B2 => n10, ZN
                           => n331);
   U363 : AOI22_X1 port map( A1 => Q(0), A2 => n11, B1 => Q(64), B2 => n12, ZN 
                           => n330);
   U364 : NOR2_X1 port map( A1 => S(2), A2 => S(3), ZN => n335);
   U365 : AOI22_X1 port map( A1 => Q(224), A2 => n13, B1 => Q(128), B2 => n14, 
                           ZN => n329);
   U366 : NOR2_X1 port map( A1 => n339, A2 => S(3), ZN => n333);
   U367 : NAND4_X1 port map( A1 => n340, A2 => n341, A3 => n342, A4 => n343, ZN
                           => n327);
   U368 : AOI22_X1 port map( A1 => Q(320), A2 => n19, B1 => Q(416), B2 => n20, 
                           ZN => n343);
   U369 : AOI22_X1 port map( A1 => Q(384), A2 => n21, B1 => Q(256), B2 => n22, 
                           ZN => n342);
   U370 : NOR2_X1 port map( A1 => S(0), A2 => S(1), ZN => n338);
   U371 : AOI22_X1 port map( A1 => Q(352), A2 => n23, B1 => Q(288), B2 => n24, 
                           ZN => n341);
   U372 : NOR2_X1 port map( A1 => n346, A2 => S(1), ZN => n337);
   U373 : NOR2_X1 port map( A1 => n347, A2 => S(2), ZN => n345);
   U374 : AOI22_X1 port map( A1 => Q(480), A2 => n25, B1 => Q(448), B2 => n26, 
                           ZN => n340);
   U375 : NOR2_X1 port map( A1 => n348, A2 => S(0), ZN => n334);
   U376 : NOR2_X1 port map( A1 => n339, A2 => n347, ZN => n344);
   U377 : INV_X1 port map( A => S(3), ZN => n347);
   U378 : INV_X1 port map( A => S(2), ZN => n339);
   U379 : NOR2_X1 port map( A1 => n346, A2 => n348, ZN => n336);
   U380 : INV_X1 port map( A => S(1), ZN => n348);
   U381 : INV_X1 port map( A => S(0), ZN => n346);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity addr_encoder_N4 is

   port( Q : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (3 
         downto 0));

end addr_encoder_N4;

architecture SYN_behav of addr_encoder_N4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31 : std_logic;

begin
   
   U3 : NOR3_X1 port map( A1 => n1, A2 => n2, A3 => n3, ZN => Y(3));
   U4 : INV_X1 port map( A => n4, ZN => n3);
   U5 : NOR3_X1 port map( A1 => n5, A2 => n6, A3 => n7, ZN => n2);
   U6 : INV_X1 port map( A => n8, ZN => n6);
   U7 : AOI21_X1 port map( B1 => n4, B2 => n9, A => n1, ZN => Y(2));
   U8 : OR4_X1 port map( A1 => Q(0), A2 => Q(1), A3 => Q(2), A4 => Q(3), ZN => 
                           n1);
   U9 : OAI21_X1 port map( B1 => n7, B2 => n5, A => n8, ZN => n9);
   U10 : NOR4_X1 port map( A1 => Q(10), A2 => Q(11), A3 => Q(8), A4 => Q(9), ZN
                           => n8);
   U11 : INV_X1 port map( A => n10, ZN => n5);
   U12 : NOR4_X1 port map( A1 => Q(4), A2 => Q(5), A3 => Q(6), A4 => Q(7), ZN 
                           => n4);
   U13 : AOI211_X1 port map( C1 => n11, C2 => n12, A => Q(1), B => Q(0), ZN => 
                           Y(1));
   U14 : OAI211_X1 port map( C1 => n13, C2 => n14, A => n15, B => n16, ZN => 
                           n12);
   U15 : INV_X1 port map( A => Q(5), ZN => n16);
   U16 : INV_X1 port map( A => Q(4), ZN => n15);
   U17 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => n14);
   U18 : NOR3_X1 port map( A1 => n19, A2 => Q(9), A3 => Q(8), ZN => n13);
   U19 : AOI211_X1 port map( C1 => n10, C2 => n7, A => Q(11), B => Q(10), ZN =>
                           n19);
   U20 : OR2_X1 port map( A1 => Q(15), A2 => Q(14), ZN => n7);
   U21 : NOR2_X1 port map( A1 => Q(12), A2 => Q(13), ZN => n10);
   U22 : NOR2_X1 port map( A1 => Q(3), A2 => Q(2), ZN => n11);
   U23 : NOR2_X1 port map( A1 => Q(0), A2 => n20, ZN => Y(0));
   U24 : AOI21_X1 port map( B1 => n21, B2 => n22, A => Q(1), ZN => n20);
   U25 : INV_X1 port map( A => Q(2), ZN => n22);
   U26 : OAI21_X1 port map( B1 => Q(4), B2 => n23, A => n24, ZN => n21);
   U27 : INV_X1 port map( A => Q(3), ZN => n24);
   U28 : AOI21_X1 port map( B1 => n25, B2 => n17, A => Q(5), ZN => n23);
   U29 : INV_X1 port map( A => Q(6), ZN => n17);
   U30 : OAI21_X1 port map( B1 => Q(8), B2 => n26, A => n18, ZN => n25);
   U31 : INV_X1 port map( A => Q(7), ZN => n18);
   U32 : AOI21_X1 port map( B1 => n27, B2 => n28, A => Q(9), ZN => n26);
   U33 : INV_X1 port map( A => Q(10), ZN => n28);
   U34 : OAI21_X1 port map( B1 => Q(12), B2 => n29, A => n30, ZN => n27);
   U35 : INV_X1 port map( A => Q(11), ZN => n30);
   U36 : AOI21_X1 port map( B1 => Q(15), B2 => n31, A => Q(13), ZN => n29);
   U37 : INV_X1 port map( A => Q(14), ZN => n31);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity address_generator_N16_0 is

   port( clk, rst, enable : in std_logic;  done, working : out std_logic;  addr
         : out std_logic_vector (15 downto 0));

end address_generator_N16_0;

architecture SYN_struct of address_generator_N16_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal done_port, addr_14_port, addr_13_port, addr_12_port, addr_11_port, 
      addr_10_port, addr_9_port, addr_8_port, addr_7_port, addr_6_port, 
      addr_5_port, addr_4_port, addr_3_port, addr_2_port, addr_1_port, 
      addr_0_port, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
      N19, N20, N21, n1, working_port, n2, n3, n4, n5, n6_port, n7_port, 
      n8_port, n9_port, n10_port, n11_port, n12_port, n13_port, n14_port, 
      n15_port, n16_port, n17_port, n18_port : std_logic;

begin
   done <= done_port;
   working <= working_port;
   addr <= ( done_port, addr_14_port, addr_13_port, addr_12_port, addr_11_port,
      addr_10_port, addr_9_port, addr_8_port, addr_7_port, addr_6_port, 
      addr_5_port, addr_4_port, addr_3_port, addr_2_port, addr_1_port, 
      addr_0_port );
   
   curr_addr_reg_0_inst : DFF_X1 port map( D => N6, CK => clk, Q => addr_0_port
                           , QN => working_port);
   curr_addr_reg_1_inst : DFF_X1 port map( D => N7, CK => clk, Q => addr_1_port
                           , QN => n6_port);
   curr_addr_reg_2_inst : DFF_X1 port map( D => N8, CK => clk, Q => addr_2_port
                           , QN => n5);
   curr_addr_reg_3_inst : DFF_X1 port map( D => N9, CK => clk, Q => addr_3_port
                           , QN => n18_port);
   curr_addr_reg_4_inst : DFF_X1 port map( D => N10, CK => clk, Q => 
                           addr_4_port, QN => n17_port);
   curr_addr_reg_5_inst : DFF_X1 port map( D => N11, CK => clk, Q => 
                           addr_5_port, QN => n16_port);
   curr_addr_reg_6_inst : DFF_X1 port map( D => N12, CK => clk, Q => 
                           addr_6_port, QN => n15_port);
   curr_addr_reg_7_inst : DFF_X1 port map( D => N13, CK => clk, Q => 
                           addr_7_port, QN => n14_port);
   curr_addr_reg_8_inst : DFF_X1 port map( D => N14, CK => clk, Q => 
                           addr_8_port, QN => n13_port);
   curr_addr_reg_9_inst : DFF_X1 port map( D => N15, CK => clk, Q => 
                           addr_9_port, QN => n12_port);
   curr_addr_reg_10_inst : DFF_X1 port map( D => N16, CK => clk, Q => 
                           addr_10_port, QN => n11_port);
   curr_addr_reg_11_inst : DFF_X1 port map( D => N17, CK => clk, Q => 
                           addr_11_port, QN => n10_port);
   curr_addr_reg_12_inst : DFF_X1 port map( D => N18, CK => clk, Q => 
                           addr_12_port, QN => n9_port);
   curr_addr_reg_13_inst : DFF_X1 port map( D => N19, CK => clk, Q => 
                           addr_13_port, QN => n8_port);
   curr_addr_reg_14_inst : DFF_X1 port map( D => N20, CK => clk, Q => 
                           addr_14_port, QN => n7_port);
   curr_addr_reg_15_inst : DFF_X1 port map( D => N21, CK => clk, Q => done_port
                           , QN => n1);
   U3 : NOR2_X1 port map( A1 => n5, A2 => n2, ZN => N9);
   U4 : NOR2_X1 port map( A1 => n6_port, A2 => n2, ZN => N8);
   U5 : NOR2_X1 port map( A1 => working_port, A2 => n2, ZN => N7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => N6);
   U7 : NOR2_X1 port map( A1 => n7_port, A2 => n2, ZN => N21);
   U8 : NOR2_X1 port map( A1 => n8_port, A2 => n2, ZN => N20);
   U9 : NOR2_X1 port map( A1 => n9_port, A2 => n2, ZN => N19);
   U10 : NOR2_X1 port map( A1 => n10_port, A2 => n2, ZN => N18);
   U11 : NOR2_X1 port map( A1 => n11_port, A2 => n2, ZN => N17);
   U12 : NOR2_X1 port map( A1 => n12_port, A2 => n2, ZN => N16);
   U13 : NOR2_X1 port map( A1 => n13_port, A2 => n2, ZN => N15);
   U14 : NOR2_X1 port map( A1 => n14_port, A2 => n2, ZN => N14);
   U15 : NOR2_X1 port map( A1 => n15_port, A2 => n2, ZN => N13);
   U16 : NOR2_X1 port map( A1 => n16_port, A2 => n2, ZN => N12);
   U17 : NOR2_X1 port map( A1 => n17_port, A2 => n2, ZN => N11);
   U18 : NOR2_X1 port map( A1 => n18_port, A2 => n2, ZN => N10);
   U19 : INV_X1 port map( A => n3, ZN => n2);
   U20 : NOR2_X1 port map( A1 => rst, A2 => n4, ZN => n3);
   U21 : AOI21_X1 port map( B1 => working_port, B2 => n1, A => enable, ZN => n4
                           );

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity in_loc_selblock_NBIT_DATA32_N8_F5 is

   port( regs : in std_logic_vector (2559 downto 0);  win : in std_logic_vector
         (4 downto 0);  curr_proc_regs : out std_logic_vector (511 downto 0));

end in_loc_selblock_NBIT_DATA32_N8_F5;

architecture SYN_behav of in_loc_selblock_NBIT_DATA32_N8_F5 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292 : 
      std_logic;

begin
   
   U2 : BUF_X1 port map( A => n264, Z => n98);
   U3 : BUF_X1 port map( A => n264, Z => n99);
   U4 : BUF_X1 port map( A => n264, Z => n97);
   U5 : BUF_X1 port map( A => n264, Z => n102);
   U6 : BUF_X1 port map( A => n264, Z => n100);
   U7 : BUF_X1 port map( A => n264, Z => n96);
   U8 : BUF_X1 port map( A => n264, Z => n101);
   U9 : BUF_X1 port map( A => n264, Z => n103);
   U10 : BUF_X1 port map( A => n263, Z => n46);
   U11 : BUF_X1 port map( A => n263, Z => n47);
   U12 : BUF_X1 port map( A => n263, Z => n45);
   U13 : BUF_X1 port map( A => n263, Z => n50);
   U14 : BUF_X1 port map( A => n263, Z => n48);
   U15 : BUF_X1 port map( A => n263, Z => n44);
   U16 : BUF_X1 port map( A => n263, Z => n49);
   U17 : BUF_X1 port map( A => n263, Z => n51);
   U18 : BUF_X1 port map( A => n265, Z => n150);
   U19 : BUF_X1 port map( A => n265, Z => n151);
   U20 : BUF_X1 port map( A => n265, Z => n149);
   U21 : BUF_X1 port map( A => n265, Z => n154);
   U22 : BUF_X1 port map( A => n265, Z => n152);
   U23 : BUF_X1 port map( A => n265, Z => n148);
   U24 : BUF_X1 port map( A => n265, Z => n153);
   U25 : BUF_X1 port map( A => n265, Z => n155);
   U26 : BUF_X1 port map( A => n266, Z => n202);
   U27 : BUF_X1 port map( A => n266, Z => n203);
   U28 : BUF_X1 port map( A => n266, Z => n201);
   U29 : BUF_X1 port map( A => n266, Z => n206);
   U30 : BUF_X1 port map( A => n266, Z => n204);
   U31 : BUF_X1 port map( A => n266, Z => n200);
   U32 : BUF_X1 port map( A => n266, Z => n205);
   U33 : BUF_X1 port map( A => n266, Z => n207);
   U34 : BUF_X1 port map( A => n264, Z => n104);
   U35 : BUF_X1 port map( A => n263, Z => n52);
   U36 : BUF_X1 port map( A => n265, Z => n156);
   U37 : BUF_X1 port map( A => n266, Z => n208);
   U38 : BUF_X1 port map( A => win(4), Z => n252);
   U39 : BUF_X1 port map( A => win(4), Z => n253);
   U40 : BUF_X1 port map( A => win(4), Z => n255);
   U41 : BUF_X1 port map( A => win(4), Z => n256);
   U42 : BUF_X1 port map( A => win(4), Z => n258);
   U43 : BUF_X1 port map( A => win(4), Z => n254);
   U44 : BUF_X1 port map( A => win(4), Z => n259);
   U45 : BUF_X1 port map( A => win(4), Z => n257);
   U46 : BUF_X1 port map( A => win(4), Z => n260);
   U47 : CLKBUF_X1 port map( A => n52, Z => n1);
   U48 : CLKBUF_X1 port map( A => n52, Z => n2);
   U49 : CLKBUF_X1 port map( A => n52, Z => n3);
   U50 : CLKBUF_X1 port map( A => n51, Z => n4);
   U51 : CLKBUF_X1 port map( A => n51, Z => n5);
   U52 : CLKBUF_X1 port map( A => n51, Z => n6);
   U53 : CLKBUF_X1 port map( A => n51, Z => n7);
   U54 : CLKBUF_X1 port map( A => n51, Z => n8);
   U55 : CLKBUF_X1 port map( A => n50, Z => n9);
   U56 : CLKBUF_X1 port map( A => n50, Z => n10);
   U57 : CLKBUF_X1 port map( A => n50, Z => n11);
   U58 : CLKBUF_X1 port map( A => n50, Z => n12);
   U59 : CLKBUF_X1 port map( A => n50, Z => n13);
   U60 : CLKBUF_X1 port map( A => n49, Z => n14);
   U61 : CLKBUF_X1 port map( A => n49, Z => n15);
   U62 : CLKBUF_X1 port map( A => n49, Z => n16);
   U63 : CLKBUF_X1 port map( A => n49, Z => n17);
   U64 : CLKBUF_X1 port map( A => n49, Z => n18);
   U65 : CLKBUF_X1 port map( A => n48, Z => n19);
   U66 : CLKBUF_X1 port map( A => n48, Z => n20);
   U67 : CLKBUF_X1 port map( A => n48, Z => n21);
   U68 : CLKBUF_X1 port map( A => n48, Z => n22);
   U69 : CLKBUF_X1 port map( A => n48, Z => n23);
   U70 : CLKBUF_X1 port map( A => n47, Z => n24);
   U71 : CLKBUF_X1 port map( A => n47, Z => n25);
   U72 : CLKBUF_X1 port map( A => n47, Z => n26);
   U73 : CLKBUF_X1 port map( A => n47, Z => n27);
   U74 : CLKBUF_X1 port map( A => n47, Z => n28);
   U75 : CLKBUF_X1 port map( A => n46, Z => n29);
   U76 : CLKBUF_X1 port map( A => n46, Z => n30);
   U77 : CLKBUF_X1 port map( A => n46, Z => n31);
   U78 : CLKBUF_X1 port map( A => n46, Z => n32);
   U79 : CLKBUF_X1 port map( A => n46, Z => n33);
   U80 : CLKBUF_X1 port map( A => n45, Z => n34);
   U81 : CLKBUF_X1 port map( A => n45, Z => n35);
   U82 : CLKBUF_X1 port map( A => n45, Z => n36);
   U83 : CLKBUF_X1 port map( A => n45, Z => n37);
   U84 : CLKBUF_X1 port map( A => n45, Z => n38);
   U85 : CLKBUF_X1 port map( A => n44, Z => n39);
   U86 : CLKBUF_X1 port map( A => n44, Z => n40);
   U87 : CLKBUF_X1 port map( A => n44, Z => n41);
   U88 : CLKBUF_X1 port map( A => n44, Z => n42);
   U89 : CLKBUF_X1 port map( A => n44, Z => n43);
   U90 : CLKBUF_X1 port map( A => n104, Z => n53);
   U91 : CLKBUF_X1 port map( A => n104, Z => n54);
   U92 : CLKBUF_X1 port map( A => n104, Z => n55);
   U93 : CLKBUF_X1 port map( A => n103, Z => n56);
   U94 : CLKBUF_X1 port map( A => n103, Z => n57);
   U95 : CLKBUF_X1 port map( A => n103, Z => n58);
   U96 : CLKBUF_X1 port map( A => n103, Z => n59);
   U97 : CLKBUF_X1 port map( A => n103, Z => n60);
   U98 : CLKBUF_X1 port map( A => n102, Z => n61);
   U99 : CLKBUF_X1 port map( A => n102, Z => n62);
   U100 : CLKBUF_X1 port map( A => n102, Z => n63);
   U101 : CLKBUF_X1 port map( A => n102, Z => n64);
   U102 : CLKBUF_X1 port map( A => n102, Z => n65);
   U103 : CLKBUF_X1 port map( A => n101, Z => n66);
   U104 : CLKBUF_X1 port map( A => n101, Z => n67);
   U105 : CLKBUF_X1 port map( A => n101, Z => n68);
   U106 : CLKBUF_X1 port map( A => n101, Z => n69);
   U107 : CLKBUF_X1 port map( A => n101, Z => n70);
   U108 : CLKBUF_X1 port map( A => n100, Z => n71);
   U109 : CLKBUF_X1 port map( A => n100, Z => n72);
   U110 : CLKBUF_X1 port map( A => n100, Z => n73);
   U111 : CLKBUF_X1 port map( A => n100, Z => n74);
   U112 : CLKBUF_X1 port map( A => n100, Z => n75);
   U113 : CLKBUF_X1 port map( A => n99, Z => n76);
   U114 : CLKBUF_X1 port map( A => n99, Z => n77);
   U115 : CLKBUF_X1 port map( A => n99, Z => n78);
   U116 : CLKBUF_X1 port map( A => n99, Z => n79);
   U117 : CLKBUF_X1 port map( A => n99, Z => n80);
   U118 : CLKBUF_X1 port map( A => n98, Z => n81);
   U119 : CLKBUF_X1 port map( A => n98, Z => n82);
   U120 : CLKBUF_X1 port map( A => n98, Z => n83);
   U121 : CLKBUF_X1 port map( A => n98, Z => n84);
   U122 : CLKBUF_X1 port map( A => n98, Z => n85);
   U123 : CLKBUF_X1 port map( A => n97, Z => n86);
   U124 : CLKBUF_X1 port map( A => n97, Z => n87);
   U125 : CLKBUF_X1 port map( A => n97, Z => n88);
   U126 : CLKBUF_X1 port map( A => n97, Z => n89);
   U127 : CLKBUF_X1 port map( A => n97, Z => n90);
   U128 : CLKBUF_X1 port map( A => n96, Z => n91);
   U129 : CLKBUF_X1 port map( A => n96, Z => n92);
   U130 : CLKBUF_X1 port map( A => n96, Z => n93);
   U131 : CLKBUF_X1 port map( A => n96, Z => n94);
   U132 : CLKBUF_X1 port map( A => n96, Z => n95);
   U133 : CLKBUF_X1 port map( A => n156, Z => n105);
   U134 : CLKBUF_X1 port map( A => n156, Z => n106);
   U135 : CLKBUF_X1 port map( A => n156, Z => n107);
   U136 : CLKBUF_X1 port map( A => n155, Z => n108);
   U137 : CLKBUF_X1 port map( A => n155, Z => n109);
   U138 : CLKBUF_X1 port map( A => n155, Z => n110);
   U139 : CLKBUF_X1 port map( A => n155, Z => n111);
   U140 : CLKBUF_X1 port map( A => n155, Z => n112);
   U141 : CLKBUF_X1 port map( A => n154, Z => n113);
   U142 : CLKBUF_X1 port map( A => n154, Z => n114);
   U143 : CLKBUF_X1 port map( A => n154, Z => n115);
   U144 : CLKBUF_X1 port map( A => n154, Z => n116);
   U145 : CLKBUF_X1 port map( A => n154, Z => n117);
   U146 : CLKBUF_X1 port map( A => n153, Z => n118);
   U147 : CLKBUF_X1 port map( A => n153, Z => n119);
   U148 : CLKBUF_X1 port map( A => n153, Z => n120);
   U149 : CLKBUF_X1 port map( A => n153, Z => n121);
   U150 : CLKBUF_X1 port map( A => n153, Z => n122);
   U151 : CLKBUF_X1 port map( A => n152, Z => n123);
   U152 : CLKBUF_X1 port map( A => n152, Z => n124);
   U153 : CLKBUF_X1 port map( A => n152, Z => n125);
   U154 : CLKBUF_X1 port map( A => n152, Z => n126);
   U155 : CLKBUF_X1 port map( A => n152, Z => n127);
   U156 : CLKBUF_X1 port map( A => n151, Z => n128);
   U157 : CLKBUF_X1 port map( A => n151, Z => n129);
   U158 : CLKBUF_X1 port map( A => n151, Z => n130);
   U159 : CLKBUF_X1 port map( A => n151, Z => n131);
   U160 : CLKBUF_X1 port map( A => n151, Z => n132);
   U161 : CLKBUF_X1 port map( A => n150, Z => n133);
   U162 : CLKBUF_X1 port map( A => n150, Z => n134);
   U163 : CLKBUF_X1 port map( A => n150, Z => n135);
   U164 : CLKBUF_X1 port map( A => n150, Z => n136);
   U165 : CLKBUF_X1 port map( A => n150, Z => n137);
   U166 : CLKBUF_X1 port map( A => n149, Z => n138);
   U167 : CLKBUF_X1 port map( A => n149, Z => n139);
   U168 : CLKBUF_X1 port map( A => n149, Z => n140);
   U169 : CLKBUF_X1 port map( A => n149, Z => n141);
   U170 : CLKBUF_X1 port map( A => n149, Z => n142);
   U171 : CLKBUF_X1 port map( A => n148, Z => n143);
   U172 : CLKBUF_X1 port map( A => n148, Z => n144);
   U173 : CLKBUF_X1 port map( A => n148, Z => n145);
   U174 : CLKBUF_X1 port map( A => n148, Z => n146);
   U175 : CLKBUF_X1 port map( A => n148, Z => n147);
   U176 : CLKBUF_X1 port map( A => n208, Z => n157);
   U177 : CLKBUF_X1 port map( A => n208, Z => n158);
   U178 : CLKBUF_X1 port map( A => n208, Z => n159);
   U179 : CLKBUF_X1 port map( A => n207, Z => n160);
   U180 : CLKBUF_X1 port map( A => n207, Z => n161);
   U181 : CLKBUF_X1 port map( A => n207, Z => n162);
   U182 : CLKBUF_X1 port map( A => n207, Z => n163);
   U183 : CLKBUF_X1 port map( A => n207, Z => n164);
   U184 : CLKBUF_X1 port map( A => n206, Z => n165);
   U185 : CLKBUF_X1 port map( A => n206, Z => n166);
   U186 : CLKBUF_X1 port map( A => n206, Z => n167);
   U187 : CLKBUF_X1 port map( A => n206, Z => n168);
   U188 : CLKBUF_X1 port map( A => n206, Z => n169);
   U189 : CLKBUF_X1 port map( A => n205, Z => n170);
   U190 : CLKBUF_X1 port map( A => n205, Z => n171);
   U191 : CLKBUF_X1 port map( A => n205, Z => n172);
   U192 : CLKBUF_X1 port map( A => n205, Z => n173);
   U193 : CLKBUF_X1 port map( A => n205, Z => n174);
   U194 : CLKBUF_X1 port map( A => n204, Z => n175);
   U195 : CLKBUF_X1 port map( A => n204, Z => n176);
   U196 : CLKBUF_X1 port map( A => n204, Z => n177);
   U197 : CLKBUF_X1 port map( A => n204, Z => n178);
   U198 : CLKBUF_X1 port map( A => n204, Z => n179);
   U199 : CLKBUF_X1 port map( A => n203, Z => n180);
   U200 : CLKBUF_X1 port map( A => n203, Z => n181);
   U201 : CLKBUF_X1 port map( A => n203, Z => n182);
   U202 : CLKBUF_X1 port map( A => n203, Z => n183);
   U203 : CLKBUF_X1 port map( A => n203, Z => n184);
   U204 : CLKBUF_X1 port map( A => n202, Z => n185);
   U205 : CLKBUF_X1 port map( A => n202, Z => n186);
   U206 : CLKBUF_X1 port map( A => n202, Z => n187);
   U207 : CLKBUF_X1 port map( A => n202, Z => n188);
   U208 : CLKBUF_X1 port map( A => n202, Z => n189);
   U209 : CLKBUF_X1 port map( A => n201, Z => n190);
   U210 : CLKBUF_X1 port map( A => n201, Z => n191);
   U211 : CLKBUF_X1 port map( A => n201, Z => n192);
   U212 : CLKBUF_X1 port map( A => n201, Z => n193);
   U213 : CLKBUF_X1 port map( A => n201, Z => n194);
   U214 : CLKBUF_X1 port map( A => n200, Z => n195);
   U215 : CLKBUF_X1 port map( A => n200, Z => n196);
   U216 : CLKBUF_X1 port map( A => n200, Z => n197);
   U217 : CLKBUF_X1 port map( A => n200, Z => n198);
   U218 : CLKBUF_X1 port map( A => n200, Z => n199);
   U219 : CLKBUF_X1 port map( A => n260, Z => n209);
   U220 : CLKBUF_X1 port map( A => n260, Z => n210);
   U221 : CLKBUF_X1 port map( A => n260, Z => n211);
   U222 : CLKBUF_X1 port map( A => n259, Z => n212);
   U223 : CLKBUF_X1 port map( A => n259, Z => n213);
   U224 : CLKBUF_X1 port map( A => n259, Z => n214);
   U225 : CLKBUF_X1 port map( A => n259, Z => n215);
   U226 : CLKBUF_X1 port map( A => n259, Z => n216);
   U227 : CLKBUF_X1 port map( A => n258, Z => n217);
   U228 : CLKBUF_X1 port map( A => n258, Z => n218);
   U229 : CLKBUF_X1 port map( A => n258, Z => n219);
   U230 : CLKBUF_X1 port map( A => n258, Z => n220);
   U231 : CLKBUF_X1 port map( A => n258, Z => n221);
   U232 : CLKBUF_X1 port map( A => n257, Z => n222);
   U233 : CLKBUF_X1 port map( A => n257, Z => n223);
   U234 : CLKBUF_X1 port map( A => n257, Z => n224);
   U235 : CLKBUF_X1 port map( A => n257, Z => n225);
   U236 : CLKBUF_X1 port map( A => n257, Z => n226);
   U237 : CLKBUF_X1 port map( A => n256, Z => n227);
   U238 : CLKBUF_X1 port map( A => n256, Z => n228);
   U239 : CLKBUF_X1 port map( A => n256, Z => n229);
   U240 : CLKBUF_X1 port map( A => n256, Z => n230);
   U241 : CLKBUF_X1 port map( A => n256, Z => n231);
   U242 : CLKBUF_X1 port map( A => n255, Z => n232);
   U243 : CLKBUF_X1 port map( A => n255, Z => n233);
   U244 : CLKBUF_X1 port map( A => n255, Z => n234);
   U245 : CLKBUF_X1 port map( A => n255, Z => n235);
   U246 : CLKBUF_X1 port map( A => n255, Z => n236);
   U247 : CLKBUF_X1 port map( A => n254, Z => n237);
   U248 : CLKBUF_X1 port map( A => n254, Z => n238);
   U249 : CLKBUF_X1 port map( A => n254, Z => n239);
   U250 : CLKBUF_X1 port map( A => n254, Z => n240);
   U251 : CLKBUF_X1 port map( A => n254, Z => n241);
   U252 : CLKBUF_X1 port map( A => n253, Z => n242);
   U253 : CLKBUF_X1 port map( A => n253, Z => n243);
   U254 : CLKBUF_X1 port map( A => n253, Z => n244);
   U255 : CLKBUF_X1 port map( A => n253, Z => n245);
   U256 : CLKBUF_X1 port map( A => n253, Z => n246);
   U257 : CLKBUF_X1 port map( A => n252, Z => n247);
   U258 : CLKBUF_X1 port map( A => n252, Z => n248);
   U259 : CLKBUF_X1 port map( A => n252, Z => n249);
   U260 : CLKBUF_X1 port map( A => n252, Z => n250);
   U261 : CLKBUF_X1 port map( A => n252, Z => n251);
   U262 : NAND2_X1 port map( A1 => n261, A2 => n262, ZN => curr_proc_regs(9));
   U263 : AOI222_X1 port map( A1 => regs(9), A2 => n43, B1 => regs(1545), B2 =>
                           n95, C1 => regs(521), C2 => n147, ZN => n262);
   U264 : AOI22_X1 port map( A1 => regs(1033), A2 => n199, B1 => n251, B2 => 
                           regs(2057), ZN => n261);
   U265 : NAND2_X1 port map( A1 => n267, A2 => n268, ZN => curr_proc_regs(99));
   U266 : AOI222_X1 port map( A1 => regs(99), A2 => n43, B1 => regs(1635), B2 
                           => n95, C1 => regs(611), C2 => n147, ZN => n268);
   U267 : AOI22_X1 port map( A1 => regs(1123), A2 => n199, B1 => regs(2147), B2
                           => n240, ZN => n267);
   U268 : NAND2_X1 port map( A1 => n269, A2 => n270, ZN => curr_proc_regs(98));
   U269 : AOI222_X1 port map( A1 => regs(98), A2 => n43, B1 => regs(1634), B2 
                           => n95, C1 => regs(610), C2 => n147, ZN => n270);
   U270 : AOI22_X1 port map( A1 => regs(1122), A2 => n199, B1 => regs(2146), B2
                           => n240, ZN => n269);
   U271 : NAND2_X1 port map( A1 => n271, A2 => n272, ZN => curr_proc_regs(97));
   U272 : AOI222_X1 port map( A1 => regs(97), A2 => n43, B1 => regs(1633), B2 
                           => n95, C1 => regs(609), C2 => n147, ZN => n272);
   U273 : AOI22_X1 port map( A1 => regs(1121), A2 => n199, B1 => regs(2145), B2
                           => n240, ZN => n271);
   U274 : NAND2_X1 port map( A1 => n273, A2 => n274, ZN => curr_proc_regs(96));
   U275 : AOI222_X1 port map( A1 => regs(96), A2 => n43, B1 => regs(1632), B2 
                           => n95, C1 => regs(608), C2 => n147, ZN => n274);
   U276 : AOI22_X1 port map( A1 => regs(1120), A2 => n199, B1 => regs(2144), B2
                           => n240, ZN => n273);
   U277 : NAND2_X1 port map( A1 => n275, A2 => n276, ZN => curr_proc_regs(95));
   U278 : AOI222_X1 port map( A1 => regs(95), A2 => n43, B1 => regs(1631), B2 
                           => n95, C1 => regs(607), C2 => n147, ZN => n276);
   U279 : AOI22_X1 port map( A1 => regs(1119), A2 => n199, B1 => regs(2143), B2
                           => n240, ZN => n275);
   U280 : NAND2_X1 port map( A1 => n277, A2 => n278, ZN => curr_proc_regs(94));
   U281 : AOI222_X1 port map( A1 => regs(94), A2 => n43, B1 => regs(1630), B2 
                           => n95, C1 => regs(606), C2 => n147, ZN => n278);
   U282 : AOI22_X1 port map( A1 => regs(1118), A2 => n199, B1 => regs(2142), B2
                           => n240, ZN => n277);
   U283 : NAND2_X1 port map( A1 => n279, A2 => n280, ZN => curr_proc_regs(93));
   U284 : AOI222_X1 port map( A1 => regs(93), A2 => n43, B1 => regs(1629), B2 
                           => n95, C1 => regs(605), C2 => n147, ZN => n280);
   U285 : AOI22_X1 port map( A1 => regs(1117), A2 => n199, B1 => regs(2141), B2
                           => n240, ZN => n279);
   U286 : NAND2_X1 port map( A1 => n281, A2 => n282, ZN => curr_proc_regs(92));
   U287 : AOI222_X1 port map( A1 => regs(92), A2 => n42, B1 => regs(1628), B2 
                           => n94, C1 => regs(604), C2 => n146, ZN => n282);
   U288 : AOI22_X1 port map( A1 => regs(1116), A2 => n198, B1 => regs(2140), B2
                           => n240, ZN => n281);
   U289 : NAND2_X1 port map( A1 => n283, A2 => n284, ZN => curr_proc_regs(91));
   U290 : AOI222_X1 port map( A1 => regs(91), A2 => n42, B1 => regs(1627), B2 
                           => n94, C1 => regs(603), C2 => n146, ZN => n284);
   U291 : AOI22_X1 port map( A1 => regs(1115), A2 => n198, B1 => regs(2139), B2
                           => n240, ZN => n283);
   U292 : NAND2_X1 port map( A1 => n285, A2 => n286, ZN => curr_proc_regs(90));
   U293 : AOI222_X1 port map( A1 => regs(90), A2 => n42, B1 => regs(1626), B2 
                           => n94, C1 => regs(602), C2 => n146, ZN => n286);
   U294 : AOI22_X1 port map( A1 => regs(1114), A2 => n198, B1 => regs(2138), B2
                           => n240, ZN => n285);
   U295 : NAND2_X1 port map( A1 => n287, A2 => n288, ZN => curr_proc_regs(8));
   U296 : AOI222_X1 port map( A1 => regs(8), A2 => n42, B1 => regs(1544), B2 =>
                           n94, C1 => regs(520), C2 => n146, ZN => n288);
   U297 : AOI22_X1 port map( A1 => regs(1032), A2 => n198, B1 => regs(2056), B2
                           => n240, ZN => n287);
   U298 : NAND2_X1 port map( A1 => n289, A2 => n290, ZN => curr_proc_regs(89));
   U299 : AOI222_X1 port map( A1 => regs(89), A2 => n42, B1 => regs(1625), B2 
                           => n94, C1 => regs(601), C2 => n146, ZN => n290);
   U300 : AOI22_X1 port map( A1 => regs(1113), A2 => n198, B1 => regs(2137), B2
                           => n240, ZN => n289);
   U301 : NAND2_X1 port map( A1 => n291, A2 => n292, ZN => curr_proc_regs(88));
   U302 : AOI222_X1 port map( A1 => regs(88), A2 => n42, B1 => regs(1624), B2 
                           => n94, C1 => regs(600), C2 => n146, ZN => n292);
   U303 : AOI22_X1 port map( A1 => regs(1112), A2 => n198, B1 => regs(2136), B2
                           => n239, ZN => n291);
   U304 : NAND2_X1 port map( A1 => n293, A2 => n294, ZN => curr_proc_regs(87));
   U305 : AOI222_X1 port map( A1 => regs(87), A2 => n42, B1 => regs(1623), B2 
                           => n94, C1 => regs(599), C2 => n146, ZN => n294);
   U306 : AOI22_X1 port map( A1 => regs(1111), A2 => n198, B1 => regs(2135), B2
                           => n239, ZN => n293);
   U307 : NAND2_X1 port map( A1 => n295, A2 => n296, ZN => curr_proc_regs(86));
   U308 : AOI222_X1 port map( A1 => regs(86), A2 => n42, B1 => regs(1622), B2 
                           => n94, C1 => regs(598), C2 => n146, ZN => n296);
   U309 : AOI22_X1 port map( A1 => regs(1110), A2 => n198, B1 => regs(2134), B2
                           => n239, ZN => n295);
   U310 : NAND2_X1 port map( A1 => n297, A2 => n298, ZN => curr_proc_regs(85));
   U311 : AOI222_X1 port map( A1 => regs(85), A2 => n42, B1 => regs(1621), B2 
                           => n94, C1 => regs(597), C2 => n146, ZN => n298);
   U312 : AOI22_X1 port map( A1 => regs(1109), A2 => n198, B1 => regs(2133), B2
                           => n239, ZN => n297);
   U313 : NAND2_X1 port map( A1 => n299, A2 => n300, ZN => curr_proc_regs(84));
   U314 : AOI222_X1 port map( A1 => regs(84), A2 => n42, B1 => regs(1620), B2 
                           => n94, C1 => regs(596), C2 => n146, ZN => n300);
   U315 : AOI22_X1 port map( A1 => regs(1108), A2 => n198, B1 => regs(2132), B2
                           => n239, ZN => n299);
   U316 : NAND2_X1 port map( A1 => n301, A2 => n302, ZN => curr_proc_regs(83));
   U317 : AOI222_X1 port map( A1 => regs(83), A2 => n42, B1 => regs(1619), B2 
                           => n94, C1 => regs(595), C2 => n146, ZN => n302);
   U318 : AOI22_X1 port map( A1 => regs(1107), A2 => n198, B1 => regs(2131), B2
                           => n239, ZN => n301);
   U319 : NAND2_X1 port map( A1 => n303, A2 => n304, ZN => curr_proc_regs(82));
   U320 : AOI222_X1 port map( A1 => regs(82), A2 => n42, B1 => regs(1618), B2 
                           => n94, C1 => regs(594), C2 => n146, ZN => n304);
   U321 : AOI22_X1 port map( A1 => regs(1106), A2 => n198, B1 => regs(2130), B2
                           => n239, ZN => n303);
   U322 : NAND2_X1 port map( A1 => n305, A2 => n306, ZN => curr_proc_regs(81));
   U323 : AOI222_X1 port map( A1 => regs(81), A2 => n41, B1 => regs(1617), B2 
                           => n93, C1 => regs(593), C2 => n145, ZN => n306);
   U324 : AOI22_X1 port map( A1 => regs(1105), A2 => n197, B1 => regs(2129), B2
                           => n239, ZN => n305);
   U325 : NAND2_X1 port map( A1 => n307, A2 => n308, ZN => curr_proc_regs(80));
   U326 : AOI222_X1 port map( A1 => regs(80), A2 => n41, B1 => regs(1616), B2 
                           => n93, C1 => regs(592), C2 => n145, ZN => n308);
   U327 : AOI22_X1 port map( A1 => regs(1104), A2 => n197, B1 => regs(2128), B2
                           => n239, ZN => n307);
   U328 : NAND2_X1 port map( A1 => n309, A2 => n310, ZN => curr_proc_regs(7));
   U329 : AOI222_X1 port map( A1 => regs(7), A2 => n41, B1 => regs(1543), B2 =>
                           n93, C1 => regs(519), C2 => n145, ZN => n310);
   U330 : AOI22_X1 port map( A1 => regs(1031), A2 => n197, B1 => regs(2055), B2
                           => n239, ZN => n309);
   U331 : NAND2_X1 port map( A1 => n311, A2 => n312, ZN => curr_proc_regs(79));
   U332 : AOI222_X1 port map( A1 => regs(79), A2 => n41, B1 => regs(1615), B2 
                           => n93, C1 => regs(591), C2 => n145, ZN => n312);
   U333 : AOI22_X1 port map( A1 => regs(1103), A2 => n197, B1 => regs(2127), B2
                           => n239, ZN => n311);
   U334 : NAND2_X1 port map( A1 => n313, A2 => n314, ZN => curr_proc_regs(78));
   U335 : AOI222_X1 port map( A1 => regs(78), A2 => n41, B1 => regs(1614), B2 
                           => n93, C1 => regs(590), C2 => n145, ZN => n314);
   U336 : AOI22_X1 port map( A1 => regs(1102), A2 => n197, B1 => regs(2126), B2
                           => n239, ZN => n313);
   U337 : NAND2_X1 port map( A1 => n315, A2 => n316, ZN => curr_proc_regs(77));
   U338 : AOI222_X1 port map( A1 => regs(77), A2 => n41, B1 => regs(1613), B2 
                           => n93, C1 => regs(589), C2 => n145, ZN => n316);
   U339 : AOI22_X1 port map( A1 => regs(1101), A2 => n197, B1 => regs(2125), B2
                           => n238, ZN => n315);
   U340 : NAND2_X1 port map( A1 => n317, A2 => n318, ZN => curr_proc_regs(76));
   U341 : AOI222_X1 port map( A1 => regs(76), A2 => n41, B1 => regs(1612), B2 
                           => n93, C1 => regs(588), C2 => n145, ZN => n318);
   U342 : AOI22_X1 port map( A1 => regs(1100), A2 => n197, B1 => regs(2124), B2
                           => n238, ZN => n317);
   U343 : NAND2_X1 port map( A1 => n319, A2 => n320, ZN => curr_proc_regs(75));
   U344 : AOI222_X1 port map( A1 => regs(75), A2 => n41, B1 => regs(1611), B2 
                           => n93, C1 => regs(587), C2 => n145, ZN => n320);
   U345 : AOI22_X1 port map( A1 => regs(1099), A2 => n197, B1 => regs(2123), B2
                           => n238, ZN => n319);
   U346 : NAND2_X1 port map( A1 => n321, A2 => n322, ZN => curr_proc_regs(74));
   U347 : AOI222_X1 port map( A1 => regs(74), A2 => n41, B1 => regs(1610), B2 
                           => n93, C1 => regs(586), C2 => n145, ZN => n322);
   U348 : AOI22_X1 port map( A1 => regs(1098), A2 => n197, B1 => regs(2122), B2
                           => n238, ZN => n321);
   U349 : NAND2_X1 port map( A1 => n323, A2 => n324, ZN => curr_proc_regs(73));
   U350 : AOI222_X1 port map( A1 => regs(73), A2 => n41, B1 => regs(1609), B2 
                           => n93, C1 => regs(585), C2 => n145, ZN => n324);
   U351 : AOI22_X1 port map( A1 => regs(1097), A2 => n197, B1 => regs(2121), B2
                           => n238, ZN => n323);
   U352 : NAND2_X1 port map( A1 => n325, A2 => n326, ZN => curr_proc_regs(72));
   U353 : AOI222_X1 port map( A1 => regs(72), A2 => n41, B1 => regs(1608), B2 
                           => n93, C1 => regs(584), C2 => n145, ZN => n326);
   U354 : AOI22_X1 port map( A1 => regs(1096), A2 => n197, B1 => regs(2120), B2
                           => n238, ZN => n325);
   U355 : NAND2_X1 port map( A1 => n327, A2 => n328, ZN => curr_proc_regs(71));
   U356 : AOI222_X1 port map( A1 => regs(71), A2 => n41, B1 => regs(1607), B2 
                           => n93, C1 => regs(583), C2 => n145, ZN => n328);
   U357 : AOI22_X1 port map( A1 => regs(1095), A2 => n197, B1 => regs(2119), B2
                           => n238, ZN => n327);
   U358 : NAND2_X1 port map( A1 => n329, A2 => n330, ZN => curr_proc_regs(70));
   U359 : AOI222_X1 port map( A1 => regs(70), A2 => n40, B1 => regs(1606), B2 
                           => n92, C1 => regs(582), C2 => n144, ZN => n330);
   U360 : AOI22_X1 port map( A1 => regs(1094), A2 => n196, B1 => regs(2118), B2
                           => n238, ZN => n329);
   U361 : NAND2_X1 port map( A1 => n331, A2 => n332, ZN => curr_proc_regs(6));
   U362 : AOI222_X1 port map( A1 => regs(6), A2 => n40, B1 => regs(1542), B2 =>
                           n92, C1 => regs(518), C2 => n144, ZN => n332);
   U363 : AOI22_X1 port map( A1 => regs(1030), A2 => n196, B1 => regs(2054), B2
                           => n238, ZN => n331);
   U364 : NAND2_X1 port map( A1 => n333, A2 => n334, ZN => curr_proc_regs(69));
   U365 : AOI222_X1 port map( A1 => regs(69), A2 => n40, B1 => regs(1605), B2 
                           => n92, C1 => regs(581), C2 => n144, ZN => n334);
   U366 : AOI22_X1 port map( A1 => regs(1093), A2 => n196, B1 => regs(2117), B2
                           => n238, ZN => n333);
   U367 : NAND2_X1 port map( A1 => n335, A2 => n336, ZN => curr_proc_regs(68));
   U368 : AOI222_X1 port map( A1 => regs(68), A2 => n40, B1 => regs(1604), B2 
                           => n92, C1 => regs(580), C2 => n144, ZN => n336);
   U369 : AOI22_X1 port map( A1 => regs(1092), A2 => n196, B1 => regs(2116), B2
                           => n238, ZN => n335);
   U370 : NAND2_X1 port map( A1 => n337, A2 => n338, ZN => curr_proc_regs(67));
   U371 : AOI222_X1 port map( A1 => regs(67), A2 => n40, B1 => regs(1603), B2 
                           => n92, C1 => regs(579), C2 => n144, ZN => n338);
   U372 : AOI22_X1 port map( A1 => regs(1091), A2 => n196, B1 => regs(2115), B2
                           => n238, ZN => n337);
   U373 : NAND2_X1 port map( A1 => n339, A2 => n340, ZN => curr_proc_regs(66));
   U374 : AOI222_X1 port map( A1 => regs(66), A2 => n40, B1 => regs(1602), B2 
                           => n92, C1 => regs(578), C2 => n144, ZN => n340);
   U375 : AOI22_X1 port map( A1 => regs(1090), A2 => n196, B1 => regs(2114), B2
                           => n237, ZN => n339);
   U376 : NAND2_X1 port map( A1 => n341, A2 => n342, ZN => curr_proc_regs(65));
   U377 : AOI222_X1 port map( A1 => regs(65), A2 => n40, B1 => regs(1601), B2 
                           => n92, C1 => regs(577), C2 => n144, ZN => n342);
   U378 : AOI22_X1 port map( A1 => regs(1089), A2 => n196, B1 => regs(2113), B2
                           => n237, ZN => n341);
   U379 : NAND2_X1 port map( A1 => n343, A2 => n344, ZN => curr_proc_regs(64));
   U380 : AOI222_X1 port map( A1 => regs(64), A2 => n40, B1 => regs(1600), B2 
                           => n92, C1 => regs(576), C2 => n144, ZN => n344);
   U381 : AOI22_X1 port map( A1 => regs(1088), A2 => n196, B1 => regs(2112), B2
                           => n237, ZN => n343);
   U382 : NAND2_X1 port map( A1 => n345, A2 => n346, ZN => curr_proc_regs(63));
   U383 : AOI222_X1 port map( A1 => regs(63), A2 => n40, B1 => regs(1599), B2 
                           => n92, C1 => regs(575), C2 => n144, ZN => n346);
   U384 : AOI22_X1 port map( A1 => regs(1087), A2 => n196, B1 => regs(2111), B2
                           => n237, ZN => n345);
   U385 : NAND2_X1 port map( A1 => n347, A2 => n348, ZN => curr_proc_regs(62));
   U386 : AOI222_X1 port map( A1 => regs(62), A2 => n40, B1 => regs(1598), B2 
                           => n92, C1 => regs(574), C2 => n144, ZN => n348);
   U387 : AOI22_X1 port map( A1 => regs(1086), A2 => n196, B1 => regs(2110), B2
                           => n237, ZN => n347);
   U388 : NAND2_X1 port map( A1 => n349, A2 => n350, ZN => curr_proc_regs(61));
   U389 : AOI222_X1 port map( A1 => regs(61), A2 => n40, B1 => regs(1597), B2 
                           => n92, C1 => regs(573), C2 => n144, ZN => n350);
   U390 : AOI22_X1 port map( A1 => regs(1085), A2 => n196, B1 => regs(2109), B2
                           => n237, ZN => n349);
   U391 : NAND2_X1 port map( A1 => n351, A2 => n352, ZN => curr_proc_regs(60));
   U392 : AOI222_X1 port map( A1 => regs(60), A2 => n40, B1 => regs(1596), B2 
                           => n92, C1 => regs(572), C2 => n144, ZN => n352);
   U393 : AOI22_X1 port map( A1 => regs(1084), A2 => n196, B1 => regs(2108), B2
                           => n237, ZN => n351);
   U394 : NAND2_X1 port map( A1 => n353, A2 => n354, ZN => curr_proc_regs(5));
   U395 : AOI222_X1 port map( A1 => regs(5), A2 => n39, B1 => regs(1541), B2 =>
                           n91, C1 => regs(517), C2 => n143, ZN => n354);
   U396 : AOI22_X1 port map( A1 => regs(1029), A2 => n195, B1 => regs(2053), B2
                           => n237, ZN => n353);
   U397 : NAND2_X1 port map( A1 => n355, A2 => n356, ZN => curr_proc_regs(59));
   U398 : AOI222_X1 port map( A1 => regs(59), A2 => n39, B1 => regs(1595), B2 
                           => n91, C1 => regs(571), C2 => n143, ZN => n356);
   U399 : AOI22_X1 port map( A1 => regs(1083), A2 => n195, B1 => regs(2107), B2
                           => n237, ZN => n355);
   U400 : NAND2_X1 port map( A1 => n357, A2 => n358, ZN => curr_proc_regs(58));
   U401 : AOI222_X1 port map( A1 => regs(58), A2 => n39, B1 => regs(1594), B2 
                           => n91, C1 => regs(570), C2 => n143, ZN => n358);
   U402 : AOI22_X1 port map( A1 => regs(1082), A2 => n195, B1 => regs(2106), B2
                           => n237, ZN => n357);
   U403 : NAND2_X1 port map( A1 => n359, A2 => n360, ZN => curr_proc_regs(57));
   U404 : AOI222_X1 port map( A1 => regs(57), A2 => n39, B1 => regs(1593), B2 
                           => n91, C1 => regs(569), C2 => n143, ZN => n360);
   U405 : AOI22_X1 port map( A1 => regs(1081), A2 => n195, B1 => regs(2105), B2
                           => n237, ZN => n359);
   U406 : NAND2_X1 port map( A1 => n361, A2 => n362, ZN => curr_proc_regs(56));
   U407 : AOI222_X1 port map( A1 => regs(56), A2 => n39, B1 => regs(1592), B2 
                           => n91, C1 => regs(568), C2 => n143, ZN => n362);
   U408 : AOI22_X1 port map( A1 => regs(1080), A2 => n195, B1 => regs(2104), B2
                           => n237, ZN => n361);
   U409 : NAND2_X1 port map( A1 => n363, A2 => n364, ZN => curr_proc_regs(55));
   U410 : AOI222_X1 port map( A1 => regs(55), A2 => n39, B1 => regs(1591), B2 
                           => n91, C1 => regs(567), C2 => n143, ZN => n364);
   U411 : AOI22_X1 port map( A1 => regs(1079), A2 => n195, B1 => regs(2103), B2
                           => n236, ZN => n363);
   U412 : NAND2_X1 port map( A1 => n365, A2 => n366, ZN => curr_proc_regs(54));
   U413 : AOI222_X1 port map( A1 => regs(54), A2 => n39, B1 => regs(1590), B2 
                           => n91, C1 => regs(566), C2 => n143, ZN => n366);
   U414 : AOI22_X1 port map( A1 => regs(1078), A2 => n195, B1 => regs(2102), B2
                           => n236, ZN => n365);
   U415 : NAND2_X1 port map( A1 => n367, A2 => n368, ZN => curr_proc_regs(53));
   U416 : AOI222_X1 port map( A1 => regs(53), A2 => n39, B1 => regs(1589), B2 
                           => n91, C1 => regs(565), C2 => n143, ZN => n368);
   U417 : AOI22_X1 port map( A1 => regs(1077), A2 => n195, B1 => regs(2101), B2
                           => n236, ZN => n367);
   U418 : NAND2_X1 port map( A1 => n369, A2 => n370, ZN => curr_proc_regs(52));
   U419 : AOI222_X1 port map( A1 => regs(52), A2 => n39, B1 => regs(1588), B2 
                           => n91, C1 => regs(564), C2 => n143, ZN => n370);
   U420 : AOI22_X1 port map( A1 => regs(1076), A2 => n195, B1 => regs(2100), B2
                           => n236, ZN => n369);
   U421 : NAND2_X1 port map( A1 => n371, A2 => n372, ZN => curr_proc_regs(51));
   U422 : AOI222_X1 port map( A1 => regs(51), A2 => n39, B1 => regs(1587), B2 
                           => n91, C1 => regs(563), C2 => n143, ZN => n372);
   U423 : AOI22_X1 port map( A1 => regs(1075), A2 => n195, B1 => regs(2099), B2
                           => n236, ZN => n371);
   U424 : NAND2_X1 port map( A1 => n373, A2 => n374, ZN => curr_proc_regs(511))
                           ;
   U425 : AOI222_X1 port map( A1 => regs(511), A2 => n39, B1 => regs(2047), B2 
                           => n91, C1 => regs(1023), C2 => n143, ZN => n374);
   U426 : AOI22_X1 port map( A1 => regs(1535), A2 => n195, B1 => regs(2559), B2
                           => n236, ZN => n373);
   U427 : NAND2_X1 port map( A1 => n375, A2 => n376, ZN => curr_proc_regs(510))
                           ;
   U428 : AOI222_X1 port map( A1 => regs(510), A2 => n39, B1 => regs(2046), B2 
                           => n91, C1 => regs(1022), C2 => n143, ZN => n376);
   U429 : AOI22_X1 port map( A1 => regs(1534), A2 => n195, B1 => regs(2558), B2
                           => n236, ZN => n375);
   U430 : NAND2_X1 port map( A1 => n377, A2 => n378, ZN => curr_proc_regs(50));
   U431 : AOI222_X1 port map( A1 => regs(50), A2 => n38, B1 => regs(1586), B2 
                           => n90, C1 => regs(562), C2 => n142, ZN => n378);
   U432 : AOI22_X1 port map( A1 => regs(1074), A2 => n194, B1 => regs(2098), B2
                           => n236, ZN => n377);
   U433 : NAND2_X1 port map( A1 => n379, A2 => n380, ZN => curr_proc_regs(509))
                           ;
   U434 : AOI222_X1 port map( A1 => regs(509), A2 => n38, B1 => regs(2045), B2 
                           => n90, C1 => regs(1021), C2 => n142, ZN => n380);
   U435 : AOI22_X1 port map( A1 => regs(1533), A2 => n194, B1 => regs(2557), B2
                           => n236, ZN => n379);
   U436 : NAND2_X1 port map( A1 => n381, A2 => n382, ZN => curr_proc_regs(508))
                           ;
   U437 : AOI222_X1 port map( A1 => regs(508), A2 => n38, B1 => regs(2044), B2 
                           => n90, C1 => regs(1020), C2 => n142, ZN => n382);
   U438 : AOI22_X1 port map( A1 => regs(1532), A2 => n194, B1 => regs(2556), B2
                           => n236, ZN => n381);
   U439 : NAND2_X1 port map( A1 => n383, A2 => n384, ZN => curr_proc_regs(507))
                           ;
   U440 : AOI222_X1 port map( A1 => regs(507), A2 => n38, B1 => regs(2043), B2 
                           => n90, C1 => regs(1019), C2 => n142, ZN => n384);
   U441 : AOI22_X1 port map( A1 => regs(1531), A2 => n194, B1 => regs(2555), B2
                           => n236, ZN => n383);
   U442 : NAND2_X1 port map( A1 => n385, A2 => n386, ZN => curr_proc_regs(506))
                           ;
   U443 : AOI222_X1 port map( A1 => regs(506), A2 => n38, B1 => regs(2042), B2 
                           => n90, C1 => regs(1018), C2 => n142, ZN => n386);
   U444 : AOI22_X1 port map( A1 => regs(1530), A2 => n194, B1 => regs(2554), B2
                           => n236, ZN => n385);
   U445 : NAND2_X1 port map( A1 => n387, A2 => n388, ZN => curr_proc_regs(505))
                           ;
   U446 : AOI222_X1 port map( A1 => regs(505), A2 => n38, B1 => regs(2041), B2 
                           => n90, C1 => regs(1017), C2 => n142, ZN => n388);
   U447 : AOI22_X1 port map( A1 => regs(1529), A2 => n194, B1 => regs(2553), B2
                           => n235, ZN => n387);
   U448 : NAND2_X1 port map( A1 => n389, A2 => n390, ZN => curr_proc_regs(504))
                           ;
   U449 : AOI222_X1 port map( A1 => regs(504), A2 => n38, B1 => regs(2040), B2 
                           => n90, C1 => regs(1016), C2 => n142, ZN => n390);
   U450 : AOI22_X1 port map( A1 => regs(1528), A2 => n194, B1 => regs(2552), B2
                           => n235, ZN => n389);
   U451 : NAND2_X1 port map( A1 => n391, A2 => n392, ZN => curr_proc_regs(503))
                           ;
   U452 : AOI222_X1 port map( A1 => regs(503), A2 => n38, B1 => regs(2039), B2 
                           => n90, C1 => regs(1015), C2 => n142, ZN => n392);
   U453 : AOI22_X1 port map( A1 => regs(1527), A2 => n194, B1 => regs(2551), B2
                           => n235, ZN => n391);
   U454 : NAND2_X1 port map( A1 => n393, A2 => n394, ZN => curr_proc_regs(502))
                           ;
   U455 : AOI222_X1 port map( A1 => regs(502), A2 => n38, B1 => regs(2038), B2 
                           => n90, C1 => regs(1014), C2 => n142, ZN => n394);
   U456 : AOI22_X1 port map( A1 => regs(1526), A2 => n194, B1 => regs(2550), B2
                           => n241, ZN => n393);
   U457 : NAND2_X1 port map( A1 => n395, A2 => n396, ZN => curr_proc_regs(501))
                           ;
   U458 : AOI222_X1 port map( A1 => regs(501), A2 => n38, B1 => regs(2037), B2 
                           => n90, C1 => regs(1013), C2 => n142, ZN => n396);
   U459 : AOI22_X1 port map( A1 => regs(1525), A2 => n194, B1 => regs(2549), B2
                           => n235, ZN => n395);
   U460 : NAND2_X1 port map( A1 => n397, A2 => n398, ZN => curr_proc_regs(500))
                           ;
   U461 : AOI222_X1 port map( A1 => regs(500), A2 => n38, B1 => regs(2036), B2 
                           => n90, C1 => regs(1012), C2 => n142, ZN => n398);
   U462 : AOI22_X1 port map( A1 => regs(1524), A2 => n194, B1 => regs(2548), B2
                           => n235, ZN => n397);
   U463 : NAND2_X1 port map( A1 => n399, A2 => n400, ZN => curr_proc_regs(4));
   U464 : AOI222_X1 port map( A1 => regs(4), A2 => n38, B1 => regs(1540), B2 =>
                           n90, C1 => regs(516), C2 => n142, ZN => n400);
   U465 : AOI22_X1 port map( A1 => regs(1028), A2 => n194, B1 => regs(2052), B2
                           => n235, ZN => n399);
   U466 : NAND2_X1 port map( A1 => n401, A2 => n402, ZN => curr_proc_regs(49));
   U467 : AOI222_X1 port map( A1 => regs(49), A2 => n37, B1 => regs(1585), B2 
                           => n89, C1 => regs(561), C2 => n141, ZN => n402);
   U468 : AOI22_X1 port map( A1 => regs(1073), A2 => n193, B1 => regs(2097), B2
                           => n235, ZN => n401);
   U469 : NAND2_X1 port map( A1 => n403, A2 => n404, ZN => curr_proc_regs(499))
                           ;
   U470 : AOI222_X1 port map( A1 => regs(499), A2 => n37, B1 => regs(2035), B2 
                           => n89, C1 => regs(1011), C2 => n141, ZN => n404);
   U471 : AOI22_X1 port map( A1 => regs(1523), A2 => n193, B1 => regs(2547), B2
                           => n235, ZN => n403);
   U472 : NAND2_X1 port map( A1 => n405, A2 => n406, ZN => curr_proc_regs(498))
                           ;
   U473 : AOI222_X1 port map( A1 => regs(498), A2 => n37, B1 => regs(2034), B2 
                           => n89, C1 => regs(1010), C2 => n141, ZN => n406);
   U474 : AOI22_X1 port map( A1 => regs(1522), A2 => n193, B1 => regs(2546), B2
                           => n235, ZN => n405);
   U475 : NAND2_X1 port map( A1 => n407, A2 => n408, ZN => curr_proc_regs(497))
                           ;
   U476 : AOI222_X1 port map( A1 => regs(497), A2 => n37, B1 => regs(2033), B2 
                           => n89, C1 => regs(1009), C2 => n141, ZN => n408);
   U477 : AOI22_X1 port map( A1 => regs(1521), A2 => n193, B1 => regs(2545), B2
                           => n235, ZN => n407);
   U478 : NAND2_X1 port map( A1 => n409, A2 => n410, ZN => curr_proc_regs(496))
                           ;
   U479 : AOI222_X1 port map( A1 => regs(496), A2 => n37, B1 => regs(2032), B2 
                           => n89, C1 => regs(1008), C2 => n141, ZN => n410);
   U480 : AOI22_X1 port map( A1 => regs(1520), A2 => n193, B1 => regs(2544), B2
                           => n235, ZN => n409);
   U481 : NAND2_X1 port map( A1 => n411, A2 => n412, ZN => curr_proc_regs(495))
                           ;
   U482 : AOI222_X1 port map( A1 => regs(495), A2 => n37, B1 => regs(2031), B2 
                           => n89, C1 => regs(1007), C2 => n141, ZN => n412);
   U483 : AOI22_X1 port map( A1 => regs(1519), A2 => n193, B1 => regs(2543), B2
                           => n234, ZN => n411);
   U484 : NAND2_X1 port map( A1 => n413, A2 => n414, ZN => curr_proc_regs(494))
                           ;
   U485 : AOI222_X1 port map( A1 => regs(494), A2 => n37, B1 => regs(2030), B2 
                           => n89, C1 => regs(1006), C2 => n141, ZN => n414);
   U486 : AOI22_X1 port map( A1 => regs(1518), A2 => n193, B1 => regs(2542), B2
                           => n234, ZN => n413);
   U487 : NAND2_X1 port map( A1 => n415, A2 => n416, ZN => curr_proc_regs(493))
                           ;
   U488 : AOI222_X1 port map( A1 => regs(493), A2 => n37, B1 => regs(2029), B2 
                           => n89, C1 => regs(1005), C2 => n141, ZN => n416);
   U489 : AOI22_X1 port map( A1 => regs(1517), A2 => n193, B1 => regs(2541), B2
                           => n234, ZN => n415);
   U490 : NAND2_X1 port map( A1 => n417, A2 => n418, ZN => curr_proc_regs(492))
                           ;
   U491 : AOI222_X1 port map( A1 => regs(492), A2 => n37, B1 => regs(2028), B2 
                           => n89, C1 => regs(1004), C2 => n141, ZN => n418);
   U492 : AOI22_X1 port map( A1 => regs(1516), A2 => n193, B1 => regs(2540), B2
                           => n234, ZN => n417);
   U493 : NAND2_X1 port map( A1 => n419, A2 => n420, ZN => curr_proc_regs(491))
                           ;
   U494 : AOI222_X1 port map( A1 => regs(491), A2 => n37, B1 => regs(2027), B2 
                           => n89, C1 => regs(1003), C2 => n141, ZN => n420);
   U495 : AOI22_X1 port map( A1 => regs(1515), A2 => n193, B1 => regs(2539), B2
                           => n234, ZN => n419);
   U496 : NAND2_X1 port map( A1 => n421, A2 => n422, ZN => curr_proc_regs(490))
                           ;
   U497 : AOI222_X1 port map( A1 => regs(490), A2 => n37, B1 => regs(2026), B2 
                           => n89, C1 => regs(1002), C2 => n141, ZN => n422);
   U498 : AOI22_X1 port map( A1 => regs(1514), A2 => n193, B1 => regs(2538), B2
                           => n234, ZN => n421);
   U499 : NAND2_X1 port map( A1 => n423, A2 => n424, ZN => curr_proc_regs(48));
   U500 : AOI222_X1 port map( A1 => regs(48), A2 => n37, B1 => regs(1584), B2 
                           => n89, C1 => regs(560), C2 => n141, ZN => n424);
   U501 : AOI22_X1 port map( A1 => regs(1072), A2 => n193, B1 => regs(2096), B2
                           => n234, ZN => n423);
   U502 : NAND2_X1 port map( A1 => n425, A2 => n426, ZN => curr_proc_regs(489))
                           ;
   U503 : AOI222_X1 port map( A1 => regs(489), A2 => n36, B1 => regs(2025), B2 
                           => n88, C1 => regs(1001), C2 => n140, ZN => n426);
   U504 : AOI22_X1 port map( A1 => regs(1513), A2 => n192, B1 => regs(2537), B2
                           => n234, ZN => n425);
   U505 : NAND2_X1 port map( A1 => n427, A2 => n428, ZN => curr_proc_regs(488))
                           ;
   U506 : AOI222_X1 port map( A1 => regs(488), A2 => n36, B1 => regs(2024), B2 
                           => n88, C1 => regs(1000), C2 => n140, ZN => n428);
   U507 : AOI22_X1 port map( A1 => regs(1512), A2 => n192, B1 => regs(2536), B2
                           => n234, ZN => n427);
   U508 : NAND2_X1 port map( A1 => n429, A2 => n430, ZN => curr_proc_regs(487))
                           ;
   U509 : AOI222_X1 port map( A1 => regs(487), A2 => n36, B1 => regs(2023), B2 
                           => n88, C1 => regs(999), C2 => n140, ZN => n430);
   U510 : AOI22_X1 port map( A1 => regs(1511), A2 => n192, B1 => regs(2535), B2
                           => n234, ZN => n429);
   U511 : NAND2_X1 port map( A1 => n431, A2 => n432, ZN => curr_proc_regs(486))
                           ;
   U512 : AOI222_X1 port map( A1 => regs(486), A2 => n36, B1 => regs(2022), B2 
                           => n88, C1 => regs(998), C2 => n140, ZN => n432);
   U513 : AOI22_X1 port map( A1 => regs(1510), A2 => n192, B1 => regs(2534), B2
                           => n234, ZN => n431);
   U514 : NAND2_X1 port map( A1 => n433, A2 => n434, ZN => curr_proc_regs(485))
                           ;
   U515 : AOI222_X1 port map( A1 => regs(485), A2 => n36, B1 => regs(2021), B2 
                           => n88, C1 => regs(997), C2 => n140, ZN => n434);
   U516 : AOI22_X1 port map( A1 => regs(1509), A2 => n192, B1 => regs(2533), B2
                           => n234, ZN => n433);
   U517 : NAND2_X1 port map( A1 => n435, A2 => n436, ZN => curr_proc_regs(484))
                           ;
   U518 : AOI222_X1 port map( A1 => regs(484), A2 => n36, B1 => regs(2020), B2 
                           => n88, C1 => regs(996), C2 => n140, ZN => n436);
   U519 : AOI22_X1 port map( A1 => regs(1508), A2 => n192, B1 => regs(2532), B2
                           => n233, ZN => n435);
   U520 : NAND2_X1 port map( A1 => n437, A2 => n438, ZN => curr_proc_regs(483))
                           ;
   U521 : AOI222_X1 port map( A1 => regs(483), A2 => n36, B1 => regs(2019), B2 
                           => n88, C1 => regs(995), C2 => n140, ZN => n438);
   U522 : AOI22_X1 port map( A1 => regs(1507), A2 => n192, B1 => regs(2531), B2
                           => n233, ZN => n437);
   U523 : NAND2_X1 port map( A1 => n439, A2 => n440, ZN => curr_proc_regs(482))
                           ;
   U524 : AOI222_X1 port map( A1 => regs(482), A2 => n36, B1 => regs(2018), B2 
                           => n88, C1 => regs(994), C2 => n140, ZN => n440);
   U525 : AOI22_X1 port map( A1 => regs(1506), A2 => n192, B1 => regs(2530), B2
                           => n233, ZN => n439);
   U526 : NAND2_X1 port map( A1 => n441, A2 => n442, ZN => curr_proc_regs(481))
                           ;
   U527 : AOI222_X1 port map( A1 => regs(481), A2 => n36, B1 => regs(2017), B2 
                           => n88, C1 => regs(993), C2 => n140, ZN => n442);
   U528 : AOI22_X1 port map( A1 => regs(1505), A2 => n192, B1 => regs(2529), B2
                           => n233, ZN => n441);
   U529 : NAND2_X1 port map( A1 => n443, A2 => n444, ZN => curr_proc_regs(480))
                           ;
   U530 : AOI222_X1 port map( A1 => regs(480), A2 => n36, B1 => regs(2016), B2 
                           => n88, C1 => regs(992), C2 => n140, ZN => n444);
   U531 : AOI22_X1 port map( A1 => regs(1504), A2 => n192, B1 => regs(2528), B2
                           => n233, ZN => n443);
   U532 : NAND2_X1 port map( A1 => n445, A2 => n446, ZN => curr_proc_regs(47));
   U533 : AOI222_X1 port map( A1 => regs(47), A2 => n36, B1 => regs(1583), B2 
                           => n88, C1 => regs(559), C2 => n140, ZN => n446);
   U534 : AOI22_X1 port map( A1 => regs(1071), A2 => n192, B1 => regs(2095), B2
                           => n233, ZN => n445);
   U535 : NAND2_X1 port map( A1 => n447, A2 => n448, ZN => curr_proc_regs(479))
                           ;
   U536 : AOI222_X1 port map( A1 => regs(479), A2 => n36, B1 => regs(2015), B2 
                           => n88, C1 => regs(991), C2 => n140, ZN => n448);
   U537 : AOI22_X1 port map( A1 => regs(1503), A2 => n192, B1 => regs(2527), B2
                           => n233, ZN => n447);
   U538 : NAND2_X1 port map( A1 => n449, A2 => n450, ZN => curr_proc_regs(478))
                           ;
   U539 : AOI222_X1 port map( A1 => regs(478), A2 => n35, B1 => regs(2014), B2 
                           => n87, C1 => regs(990), C2 => n139, ZN => n450);
   U540 : AOI22_X1 port map( A1 => regs(1502), A2 => n191, B1 => regs(2526), B2
                           => n233, ZN => n449);
   U541 : NAND2_X1 port map( A1 => n451, A2 => n452, ZN => curr_proc_regs(477))
                           ;
   U542 : AOI222_X1 port map( A1 => regs(477), A2 => n35, B1 => regs(2013), B2 
                           => n87, C1 => regs(989), C2 => n139, ZN => n452);
   U543 : AOI22_X1 port map( A1 => regs(1501), A2 => n191, B1 => regs(2525), B2
                           => n233, ZN => n451);
   U544 : NAND2_X1 port map( A1 => n453, A2 => n454, ZN => curr_proc_regs(476))
                           ;
   U545 : AOI222_X1 port map( A1 => regs(476), A2 => n35, B1 => regs(2012), B2 
                           => n87, C1 => regs(988), C2 => n139, ZN => n454);
   U546 : AOI22_X1 port map( A1 => regs(1500), A2 => n191, B1 => regs(2524), B2
                           => n233, ZN => n453);
   U547 : NAND2_X1 port map( A1 => n455, A2 => n456, ZN => curr_proc_regs(475))
                           ;
   U548 : AOI222_X1 port map( A1 => regs(475), A2 => n35, B1 => regs(2011), B2 
                           => n87, C1 => regs(987), C2 => n139, ZN => n456);
   U549 : AOI22_X1 port map( A1 => regs(1499), A2 => n191, B1 => regs(2523), B2
                           => n233, ZN => n455);
   U550 : NAND2_X1 port map( A1 => n457, A2 => n458, ZN => curr_proc_regs(474))
                           ;
   U551 : AOI222_X1 port map( A1 => regs(474), A2 => n35, B1 => regs(2010), B2 
                           => n87, C1 => regs(986), C2 => n139, ZN => n458);
   U552 : AOI22_X1 port map( A1 => regs(1498), A2 => n191, B1 => regs(2522), B2
                           => n233, ZN => n457);
   U553 : NAND2_X1 port map( A1 => n459, A2 => n460, ZN => curr_proc_regs(473))
                           ;
   U554 : AOI222_X1 port map( A1 => regs(473), A2 => n35, B1 => regs(2009), B2 
                           => n87, C1 => regs(985), C2 => n139, ZN => n460);
   U555 : AOI22_X1 port map( A1 => regs(1497), A2 => n191, B1 => regs(2521), B2
                           => n232, ZN => n459);
   U556 : NAND2_X1 port map( A1 => n461, A2 => n462, ZN => curr_proc_regs(472))
                           ;
   U557 : AOI222_X1 port map( A1 => regs(472), A2 => n35, B1 => regs(2008), B2 
                           => n87, C1 => regs(984), C2 => n139, ZN => n462);
   U558 : AOI22_X1 port map( A1 => regs(1496), A2 => n191, B1 => regs(2520), B2
                           => n232, ZN => n461);
   U559 : NAND2_X1 port map( A1 => n463, A2 => n464, ZN => curr_proc_regs(471))
                           ;
   U560 : AOI222_X1 port map( A1 => regs(471), A2 => n35, B1 => regs(2007), B2 
                           => n87, C1 => regs(983), C2 => n139, ZN => n464);
   U561 : AOI22_X1 port map( A1 => regs(1495), A2 => n191, B1 => regs(2519), B2
                           => n232, ZN => n463);
   U562 : NAND2_X1 port map( A1 => n465, A2 => n466, ZN => curr_proc_regs(470))
                           ;
   U563 : AOI222_X1 port map( A1 => regs(470), A2 => n35, B1 => regs(2006), B2 
                           => n87, C1 => regs(982), C2 => n139, ZN => n466);
   U564 : AOI22_X1 port map( A1 => regs(1494), A2 => n191, B1 => regs(2518), B2
                           => n232, ZN => n465);
   U565 : NAND2_X1 port map( A1 => n467, A2 => n468, ZN => curr_proc_regs(46));
   U566 : AOI222_X1 port map( A1 => regs(46), A2 => n35, B1 => regs(1582), B2 
                           => n87, C1 => regs(558), C2 => n139, ZN => n468);
   U567 : AOI22_X1 port map( A1 => regs(1070), A2 => n191, B1 => regs(2094), B2
                           => n232, ZN => n467);
   U568 : NAND2_X1 port map( A1 => n469, A2 => n470, ZN => curr_proc_regs(469))
                           ;
   U569 : AOI222_X1 port map( A1 => regs(469), A2 => n35, B1 => regs(2005), B2 
                           => n87, C1 => regs(981), C2 => n139, ZN => n470);
   U570 : AOI22_X1 port map( A1 => regs(1493), A2 => n191, B1 => regs(2517), B2
                           => n232, ZN => n469);
   U571 : NAND2_X1 port map( A1 => n471, A2 => n472, ZN => curr_proc_regs(468))
                           ;
   U572 : AOI222_X1 port map( A1 => regs(468), A2 => n35, B1 => regs(2004), B2 
                           => n87, C1 => regs(980), C2 => n139, ZN => n472);
   U573 : AOI22_X1 port map( A1 => regs(1492), A2 => n191, B1 => regs(2516), B2
                           => n232, ZN => n471);
   U574 : NAND2_X1 port map( A1 => n473, A2 => n474, ZN => curr_proc_regs(467))
                           ;
   U575 : AOI222_X1 port map( A1 => regs(467), A2 => n34, B1 => regs(2003), B2 
                           => n86, C1 => regs(979), C2 => n138, ZN => n474);
   U576 : AOI22_X1 port map( A1 => regs(1491), A2 => n190, B1 => regs(2515), B2
                           => n232, ZN => n473);
   U577 : NAND2_X1 port map( A1 => n475, A2 => n476, ZN => curr_proc_regs(466))
                           ;
   U578 : AOI222_X1 port map( A1 => regs(466), A2 => n34, B1 => regs(2002), B2 
                           => n86, C1 => regs(978), C2 => n138, ZN => n476);
   U579 : AOI22_X1 port map( A1 => regs(1490), A2 => n190, B1 => regs(2514), B2
                           => n232, ZN => n475);
   U580 : NAND2_X1 port map( A1 => n477, A2 => n478, ZN => curr_proc_regs(465))
                           ;
   U581 : AOI222_X1 port map( A1 => regs(465), A2 => n34, B1 => regs(2001), B2 
                           => n86, C1 => regs(977), C2 => n138, ZN => n478);
   U582 : AOI22_X1 port map( A1 => regs(1489), A2 => n190, B1 => regs(2513), B2
                           => n232, ZN => n477);
   U583 : NAND2_X1 port map( A1 => n479, A2 => n480, ZN => curr_proc_regs(464))
                           ;
   U584 : AOI222_X1 port map( A1 => regs(464), A2 => n34, B1 => regs(2000), B2 
                           => n86, C1 => regs(976), C2 => n138, ZN => n480);
   U585 : AOI22_X1 port map( A1 => regs(1488), A2 => n190, B1 => regs(2512), B2
                           => n232, ZN => n479);
   U586 : NAND2_X1 port map( A1 => n481, A2 => n482, ZN => curr_proc_regs(463))
                           ;
   U587 : AOI222_X1 port map( A1 => regs(463), A2 => n34, B1 => regs(1999), B2 
                           => n86, C1 => regs(975), C2 => n138, ZN => n482);
   U588 : AOI22_X1 port map( A1 => regs(1487), A2 => n190, B1 => regs(2511), B2
                           => n232, ZN => n481);
   U589 : NAND2_X1 port map( A1 => n483, A2 => n484, ZN => curr_proc_regs(462))
                           ;
   U590 : AOI222_X1 port map( A1 => regs(462), A2 => n34, B1 => regs(1998), B2 
                           => n86, C1 => regs(974), C2 => n138, ZN => n484);
   U591 : AOI22_X1 port map( A1 => regs(1486), A2 => n190, B1 => regs(2510), B2
                           => n231, ZN => n483);
   U592 : NAND2_X1 port map( A1 => n485, A2 => n486, ZN => curr_proc_regs(461))
                           ;
   U593 : AOI222_X1 port map( A1 => regs(461), A2 => n34, B1 => regs(1997), B2 
                           => n86, C1 => regs(973), C2 => n138, ZN => n486);
   U594 : AOI22_X1 port map( A1 => regs(1485), A2 => n190, B1 => regs(2509), B2
                           => n231, ZN => n485);
   U595 : NAND2_X1 port map( A1 => n487, A2 => n488, ZN => curr_proc_regs(460))
                           ;
   U596 : AOI222_X1 port map( A1 => regs(460), A2 => n34, B1 => regs(1996), B2 
                           => n86, C1 => regs(972), C2 => n138, ZN => n488);
   U597 : AOI22_X1 port map( A1 => regs(1484), A2 => n190, B1 => regs(2508), B2
                           => n231, ZN => n487);
   U598 : NAND2_X1 port map( A1 => n489, A2 => n490, ZN => curr_proc_regs(45));
   U599 : AOI222_X1 port map( A1 => regs(45), A2 => n34, B1 => regs(1581), B2 
                           => n86, C1 => regs(557), C2 => n138, ZN => n490);
   U600 : AOI22_X1 port map( A1 => regs(1069), A2 => n190, B1 => regs(2093), B2
                           => n231, ZN => n489);
   U601 : NAND2_X1 port map( A1 => n491, A2 => n492, ZN => curr_proc_regs(459))
                           ;
   U602 : AOI222_X1 port map( A1 => regs(459), A2 => n34, B1 => regs(1995), B2 
                           => n86, C1 => regs(971), C2 => n138, ZN => n492);
   U603 : AOI22_X1 port map( A1 => regs(1483), A2 => n190, B1 => regs(2507), B2
                           => n231, ZN => n491);
   U604 : NAND2_X1 port map( A1 => n493, A2 => n494, ZN => curr_proc_regs(458))
                           ;
   U605 : AOI222_X1 port map( A1 => regs(458), A2 => n34, B1 => regs(1994), B2 
                           => n86, C1 => regs(970), C2 => n138, ZN => n494);
   U606 : AOI22_X1 port map( A1 => regs(1482), A2 => n190, B1 => regs(2506), B2
                           => n231, ZN => n493);
   U607 : NAND2_X1 port map( A1 => n495, A2 => n496, ZN => curr_proc_regs(457))
                           ;
   U608 : AOI222_X1 port map( A1 => regs(457), A2 => n34, B1 => regs(1993), B2 
                           => n86, C1 => regs(969), C2 => n138, ZN => n496);
   U609 : AOI22_X1 port map( A1 => regs(1481), A2 => n190, B1 => regs(2505), B2
                           => n231, ZN => n495);
   U610 : NAND2_X1 port map( A1 => n497, A2 => n498, ZN => curr_proc_regs(456))
                           ;
   U611 : AOI222_X1 port map( A1 => regs(456), A2 => n33, B1 => regs(1992), B2 
                           => n85, C1 => regs(968), C2 => n137, ZN => n498);
   U612 : AOI22_X1 port map( A1 => regs(1480), A2 => n189, B1 => regs(2504), B2
                           => n231, ZN => n497);
   U613 : NAND2_X1 port map( A1 => n499, A2 => n500, ZN => curr_proc_regs(455))
                           ;
   U614 : AOI222_X1 port map( A1 => regs(455), A2 => n33, B1 => regs(1991), B2 
                           => n85, C1 => regs(967), C2 => n137, ZN => n500);
   U615 : AOI22_X1 port map( A1 => regs(1479), A2 => n189, B1 => regs(2503), B2
                           => n231, ZN => n499);
   U616 : NAND2_X1 port map( A1 => n501, A2 => n502, ZN => curr_proc_regs(454))
                           ;
   U617 : AOI222_X1 port map( A1 => regs(454), A2 => n33, B1 => regs(1990), B2 
                           => n85, C1 => regs(966), C2 => n137, ZN => n502);
   U618 : AOI22_X1 port map( A1 => regs(1478), A2 => n189, B1 => regs(2502), B2
                           => n231, ZN => n501);
   U619 : NAND2_X1 port map( A1 => n503, A2 => n504, ZN => curr_proc_regs(453))
                           ;
   U620 : AOI222_X1 port map( A1 => regs(453), A2 => n33, B1 => regs(1989), B2 
                           => n85, C1 => regs(965), C2 => n137, ZN => n504);
   U621 : AOI22_X1 port map( A1 => regs(1477), A2 => n189, B1 => regs(2501), B2
                           => n231, ZN => n503);
   U622 : NAND2_X1 port map( A1 => n505, A2 => n506, ZN => curr_proc_regs(452))
                           ;
   U623 : AOI222_X1 port map( A1 => regs(452), A2 => n33, B1 => regs(1988), B2 
                           => n85, C1 => regs(964), C2 => n137, ZN => n506);
   U624 : AOI22_X1 port map( A1 => regs(1476), A2 => n189, B1 => regs(2500), B2
                           => n231, ZN => n505);
   U625 : NAND2_X1 port map( A1 => n507, A2 => n508, ZN => curr_proc_regs(451))
                           ;
   U626 : AOI222_X1 port map( A1 => regs(451), A2 => n33, B1 => regs(1987), B2 
                           => n85, C1 => regs(963), C2 => n137, ZN => n508);
   U627 : AOI22_X1 port map( A1 => regs(1475), A2 => n189, B1 => regs(2499), B2
                           => n230, ZN => n507);
   U628 : NAND2_X1 port map( A1 => n509, A2 => n510, ZN => curr_proc_regs(450))
                           ;
   U629 : AOI222_X1 port map( A1 => regs(450), A2 => n33, B1 => regs(1986), B2 
                           => n85, C1 => regs(962), C2 => n137, ZN => n510);
   U630 : AOI22_X1 port map( A1 => regs(1474), A2 => n189, B1 => regs(2498), B2
                           => n230, ZN => n509);
   U631 : NAND2_X1 port map( A1 => n511, A2 => n512, ZN => curr_proc_regs(44));
   U632 : AOI222_X1 port map( A1 => regs(44), A2 => n33, B1 => regs(1580), B2 
                           => n85, C1 => regs(556), C2 => n137, ZN => n512);
   U633 : AOI22_X1 port map( A1 => regs(1068), A2 => n189, B1 => regs(2092), B2
                           => n230, ZN => n511);
   U634 : NAND2_X1 port map( A1 => n513, A2 => n514, ZN => curr_proc_regs(449))
                           ;
   U635 : AOI222_X1 port map( A1 => regs(449), A2 => n33, B1 => regs(1985), B2 
                           => n85, C1 => regs(961), C2 => n137, ZN => n514);
   U636 : AOI22_X1 port map( A1 => regs(1473), A2 => n189, B1 => regs(2497), B2
                           => n230, ZN => n513);
   U637 : NAND2_X1 port map( A1 => n515, A2 => n516, ZN => curr_proc_regs(448))
                           ;
   U638 : AOI222_X1 port map( A1 => regs(448), A2 => n33, B1 => regs(1984), B2 
                           => n85, C1 => regs(960), C2 => n137, ZN => n516);
   U639 : AOI22_X1 port map( A1 => regs(1472), A2 => n189, B1 => regs(2496), B2
                           => n230, ZN => n515);
   U640 : NAND2_X1 port map( A1 => n517, A2 => n518, ZN => curr_proc_regs(447))
                           ;
   U641 : AOI222_X1 port map( A1 => regs(447), A2 => n33, B1 => regs(1983), B2 
                           => n85, C1 => regs(959), C2 => n137, ZN => n518);
   U642 : AOI22_X1 port map( A1 => regs(1471), A2 => n189, B1 => regs(2495), B2
                           => n230, ZN => n517);
   U643 : NAND2_X1 port map( A1 => n519, A2 => n520, ZN => curr_proc_regs(446))
                           ;
   U644 : AOI222_X1 port map( A1 => regs(446), A2 => n33, B1 => regs(1982), B2 
                           => n85, C1 => regs(958), C2 => n137, ZN => n520);
   U645 : AOI22_X1 port map( A1 => regs(1470), A2 => n189, B1 => regs(2494), B2
                           => n230, ZN => n519);
   U646 : NAND2_X1 port map( A1 => n521, A2 => n522, ZN => curr_proc_regs(445))
                           ;
   U647 : AOI222_X1 port map( A1 => regs(445), A2 => n32, B1 => regs(1981), B2 
                           => n84, C1 => regs(957), C2 => n136, ZN => n522);
   U648 : AOI22_X1 port map( A1 => regs(1469), A2 => n188, B1 => regs(2493), B2
                           => n235, ZN => n521);
   U649 : NAND2_X1 port map( A1 => n523, A2 => n524, ZN => curr_proc_regs(444))
                           ;
   U650 : AOI222_X1 port map( A1 => regs(444), A2 => n32, B1 => regs(1980), B2 
                           => n84, C1 => regs(956), C2 => n136, ZN => n524);
   U651 : AOI22_X1 port map( A1 => regs(1468), A2 => n188, B1 => regs(2492), B2
                           => n251, ZN => n523);
   U652 : NAND2_X1 port map( A1 => n525, A2 => n526, ZN => curr_proc_regs(443))
                           ;
   U653 : AOI222_X1 port map( A1 => regs(443), A2 => n32, B1 => regs(1979), B2 
                           => n84, C1 => regs(955), C2 => n136, ZN => n526);
   U654 : AOI22_X1 port map( A1 => regs(1467), A2 => n188, B1 => regs(2491), B2
                           => n251, ZN => n525);
   U655 : NAND2_X1 port map( A1 => n527, A2 => n528, ZN => curr_proc_regs(442))
                           ;
   U656 : AOI222_X1 port map( A1 => regs(442), A2 => n32, B1 => regs(1978), B2 
                           => n84, C1 => regs(954), C2 => n136, ZN => n528);
   U657 : AOI22_X1 port map( A1 => regs(1466), A2 => n188, B1 => regs(2490), B2
                           => n251, ZN => n527);
   U658 : NAND2_X1 port map( A1 => n529, A2 => n530, ZN => curr_proc_regs(441))
                           ;
   U659 : AOI222_X1 port map( A1 => regs(441), A2 => n32, B1 => regs(1977), B2 
                           => n84, C1 => regs(953), C2 => n136, ZN => n530);
   U660 : AOI22_X1 port map( A1 => regs(1465), A2 => n188, B1 => regs(2489), B2
                           => n251, ZN => n529);
   U661 : NAND2_X1 port map( A1 => n531, A2 => n532, ZN => curr_proc_regs(440))
                           ;
   U662 : AOI222_X1 port map( A1 => regs(440), A2 => n32, B1 => regs(1976), B2 
                           => n84, C1 => regs(952), C2 => n136, ZN => n532);
   U663 : AOI22_X1 port map( A1 => regs(1464), A2 => n188, B1 => regs(2488), B2
                           => n251, ZN => n531);
   U664 : NAND2_X1 port map( A1 => n533, A2 => n534, ZN => curr_proc_regs(43));
   U665 : AOI222_X1 port map( A1 => regs(43), A2 => n32, B1 => regs(1579), B2 
                           => n84, C1 => regs(555), C2 => n136, ZN => n534);
   U666 : AOI22_X1 port map( A1 => regs(1067), A2 => n188, B1 => regs(2091), B2
                           => n251, ZN => n533);
   U667 : NAND2_X1 port map( A1 => n535, A2 => n536, ZN => curr_proc_regs(439))
                           ;
   U668 : AOI222_X1 port map( A1 => regs(439), A2 => n32, B1 => regs(1975), B2 
                           => n84, C1 => regs(951), C2 => n136, ZN => n536);
   U669 : AOI22_X1 port map( A1 => regs(1463), A2 => n188, B1 => regs(2487), B2
                           => n251, ZN => n535);
   U670 : NAND2_X1 port map( A1 => n537, A2 => n538, ZN => curr_proc_regs(438))
                           ;
   U671 : AOI222_X1 port map( A1 => regs(438), A2 => n32, B1 => regs(1974), B2 
                           => n84, C1 => regs(950), C2 => n136, ZN => n538);
   U672 : AOI22_X1 port map( A1 => regs(1462), A2 => n188, B1 => regs(2486), B2
                           => n251, ZN => n537);
   U673 : NAND2_X1 port map( A1 => n539, A2 => n540, ZN => curr_proc_regs(437))
                           ;
   U674 : AOI222_X1 port map( A1 => regs(437), A2 => n32, B1 => regs(1973), B2 
                           => n84, C1 => regs(949), C2 => n136, ZN => n540);
   U675 : AOI22_X1 port map( A1 => regs(1461), A2 => n188, B1 => regs(2485), B2
                           => n250, ZN => n539);
   U676 : NAND2_X1 port map( A1 => n541, A2 => n542, ZN => curr_proc_regs(436))
                           ;
   U677 : AOI222_X1 port map( A1 => regs(436), A2 => n32, B1 => regs(1972), B2 
                           => n84, C1 => regs(948), C2 => n136, ZN => n542);
   U678 : AOI22_X1 port map( A1 => regs(1460), A2 => n188, B1 => regs(2484), B2
                           => n251, ZN => n541);
   U679 : NAND2_X1 port map( A1 => n543, A2 => n544, ZN => curr_proc_regs(435))
                           ;
   U680 : AOI222_X1 port map( A1 => regs(435), A2 => n32, B1 => regs(1971), B2 
                           => n84, C1 => regs(947), C2 => n136, ZN => n544);
   U681 : AOI22_X1 port map( A1 => regs(1459), A2 => n188, B1 => regs(2483), B2
                           => n250, ZN => n543);
   U682 : NAND2_X1 port map( A1 => n545, A2 => n546, ZN => curr_proc_regs(434))
                           ;
   U683 : AOI222_X1 port map( A1 => regs(434), A2 => n31, B1 => regs(1970), B2 
                           => n83, C1 => regs(946), C2 => n135, ZN => n546);
   U684 : AOI22_X1 port map( A1 => regs(1458), A2 => n187, B1 => regs(2482), B2
                           => n250, ZN => n545);
   U685 : NAND2_X1 port map( A1 => n547, A2 => n548, ZN => curr_proc_regs(433))
                           ;
   U686 : AOI222_X1 port map( A1 => regs(433), A2 => n31, B1 => regs(1969), B2 
                           => n83, C1 => regs(945), C2 => n135, ZN => n548);
   U687 : AOI22_X1 port map( A1 => regs(1457), A2 => n187, B1 => regs(2481), B2
                           => n250, ZN => n547);
   U688 : NAND2_X1 port map( A1 => n549, A2 => n550, ZN => curr_proc_regs(432))
                           ;
   U689 : AOI222_X1 port map( A1 => regs(432), A2 => n31, B1 => regs(1968), B2 
                           => n83, C1 => regs(944), C2 => n135, ZN => n550);
   U690 : AOI22_X1 port map( A1 => regs(1456), A2 => n187, B1 => regs(2480), B2
                           => n250, ZN => n549);
   U691 : NAND2_X1 port map( A1 => n551, A2 => n552, ZN => curr_proc_regs(431))
                           ;
   U692 : AOI222_X1 port map( A1 => regs(431), A2 => n31, B1 => regs(1967), B2 
                           => n83, C1 => regs(943), C2 => n135, ZN => n552);
   U693 : AOI22_X1 port map( A1 => regs(1455), A2 => n187, B1 => regs(2479), B2
                           => n250, ZN => n551);
   U694 : NAND2_X1 port map( A1 => n553, A2 => n554, ZN => curr_proc_regs(430))
                           ;
   U695 : AOI222_X1 port map( A1 => regs(430), A2 => n31, B1 => regs(1966), B2 
                           => n83, C1 => regs(942), C2 => n135, ZN => n554);
   U696 : AOI22_X1 port map( A1 => regs(1454), A2 => n187, B1 => regs(2478), B2
                           => n250, ZN => n553);
   U697 : NAND2_X1 port map( A1 => n555, A2 => n556, ZN => curr_proc_regs(42));
   U698 : AOI222_X1 port map( A1 => regs(42), A2 => n31, B1 => regs(1578), B2 
                           => n83, C1 => regs(554), C2 => n135, ZN => n556);
   U699 : AOI22_X1 port map( A1 => regs(1066), A2 => n187, B1 => regs(2090), B2
                           => n250, ZN => n555);
   U700 : NAND2_X1 port map( A1 => n557, A2 => n558, ZN => curr_proc_regs(429))
                           ;
   U701 : AOI222_X1 port map( A1 => regs(429), A2 => n31, B1 => regs(1965), B2 
                           => n83, C1 => regs(941), C2 => n135, ZN => n558);
   U702 : AOI22_X1 port map( A1 => regs(1453), A2 => n187, B1 => regs(2477), B2
                           => n250, ZN => n557);
   U703 : NAND2_X1 port map( A1 => n559, A2 => n560, ZN => curr_proc_regs(428))
                           ;
   U704 : AOI222_X1 port map( A1 => regs(428), A2 => n31, B1 => regs(1964), B2 
                           => n83, C1 => regs(940), C2 => n135, ZN => n560);
   U705 : AOI22_X1 port map( A1 => regs(1452), A2 => n187, B1 => regs(2476), B2
                           => n250, ZN => n559);
   U706 : NAND2_X1 port map( A1 => n561, A2 => n562, ZN => curr_proc_regs(427))
                           ;
   U707 : AOI222_X1 port map( A1 => regs(427), A2 => n31, B1 => regs(1963), B2 
                           => n83, C1 => regs(939), C2 => n135, ZN => n562);
   U708 : AOI22_X1 port map( A1 => regs(1451), A2 => n187, B1 => regs(2475), B2
                           => n250, ZN => n561);
   U709 : NAND2_X1 port map( A1 => n563, A2 => n564, ZN => curr_proc_regs(426))
                           ;
   U710 : AOI222_X1 port map( A1 => regs(426), A2 => n31, B1 => regs(1962), B2 
                           => n83, C1 => regs(938), C2 => n135, ZN => n564);
   U711 : AOI22_X1 port map( A1 => regs(1450), A2 => n187, B1 => regs(2474), B2
                           => n249, ZN => n563);
   U712 : NAND2_X1 port map( A1 => n565, A2 => n566, ZN => curr_proc_regs(425))
                           ;
   U713 : AOI222_X1 port map( A1 => regs(425), A2 => n31, B1 => regs(1961), B2 
                           => n83, C1 => regs(937), C2 => n135, ZN => n566);
   U714 : AOI22_X1 port map( A1 => regs(1449), A2 => n187, B1 => regs(2473), B2
                           => n250, ZN => n565);
   U715 : NAND2_X1 port map( A1 => n567, A2 => n568, ZN => curr_proc_regs(424))
                           ;
   U716 : AOI222_X1 port map( A1 => regs(424), A2 => n31, B1 => regs(1960), B2 
                           => n83, C1 => regs(936), C2 => n135, ZN => n568);
   U717 : AOI22_X1 port map( A1 => regs(1448), A2 => n187, B1 => regs(2472), B2
                           => n249, ZN => n567);
   U718 : NAND2_X1 port map( A1 => n569, A2 => n570, ZN => curr_proc_regs(423))
                           ;
   U719 : AOI222_X1 port map( A1 => regs(423), A2 => n30, B1 => regs(1959), B2 
                           => n82, C1 => regs(935), C2 => n134, ZN => n570);
   U720 : AOI22_X1 port map( A1 => regs(1447), A2 => n186, B1 => regs(2471), B2
                           => n249, ZN => n569);
   U721 : NAND2_X1 port map( A1 => n571, A2 => n572, ZN => curr_proc_regs(422))
                           ;
   U722 : AOI222_X1 port map( A1 => regs(422), A2 => n30, B1 => regs(1958), B2 
                           => n82, C1 => regs(934), C2 => n134, ZN => n572);
   U723 : AOI22_X1 port map( A1 => regs(1446), A2 => n186, B1 => regs(2470), B2
                           => n249, ZN => n571);
   U724 : NAND2_X1 port map( A1 => n573, A2 => n574, ZN => curr_proc_regs(421))
                           ;
   U725 : AOI222_X1 port map( A1 => regs(421), A2 => n30, B1 => regs(1957), B2 
                           => n82, C1 => regs(933), C2 => n134, ZN => n574);
   U726 : AOI22_X1 port map( A1 => regs(1445), A2 => n186, B1 => regs(2469), B2
                           => n249, ZN => n573);
   U727 : NAND2_X1 port map( A1 => n575, A2 => n576, ZN => curr_proc_regs(420))
                           ;
   U728 : AOI222_X1 port map( A1 => regs(420), A2 => n30, B1 => regs(1956), B2 
                           => n82, C1 => regs(932), C2 => n134, ZN => n576);
   U729 : AOI22_X1 port map( A1 => regs(1444), A2 => n186, B1 => regs(2468), B2
                           => n249, ZN => n575);
   U730 : NAND2_X1 port map( A1 => n577, A2 => n578, ZN => curr_proc_regs(41));
   U731 : AOI222_X1 port map( A1 => regs(41), A2 => n30, B1 => regs(1577), B2 
                           => n82, C1 => regs(553), C2 => n134, ZN => n578);
   U732 : AOI22_X1 port map( A1 => regs(1065), A2 => n186, B1 => regs(2089), B2
                           => n249, ZN => n577);
   U733 : NAND2_X1 port map( A1 => n579, A2 => n580, ZN => curr_proc_regs(419))
                           ;
   U734 : AOI222_X1 port map( A1 => regs(419), A2 => n30, B1 => regs(1955), B2 
                           => n82, C1 => regs(931), C2 => n134, ZN => n580);
   U735 : AOI22_X1 port map( A1 => regs(1443), A2 => n186, B1 => regs(2467), B2
                           => n249, ZN => n579);
   U736 : NAND2_X1 port map( A1 => n581, A2 => n582, ZN => curr_proc_regs(418))
                           ;
   U737 : AOI222_X1 port map( A1 => regs(418), A2 => n30, B1 => regs(1954), B2 
                           => n82, C1 => regs(930), C2 => n134, ZN => n582);
   U738 : AOI22_X1 port map( A1 => regs(1442), A2 => n186, B1 => regs(2466), B2
                           => n249, ZN => n581);
   U739 : NAND2_X1 port map( A1 => n583, A2 => n584, ZN => curr_proc_regs(417))
                           ;
   U740 : AOI222_X1 port map( A1 => regs(417), A2 => n30, B1 => regs(1953), B2 
                           => n82, C1 => regs(929), C2 => n134, ZN => n584);
   U741 : AOI22_X1 port map( A1 => regs(1441), A2 => n186, B1 => regs(2465), B2
                           => n249, ZN => n583);
   U742 : NAND2_X1 port map( A1 => n585, A2 => n586, ZN => curr_proc_regs(416))
                           ;
   U743 : AOI222_X1 port map( A1 => regs(416), A2 => n30, B1 => regs(1952), B2 
                           => n82, C1 => regs(928), C2 => n134, ZN => n586);
   U744 : AOI22_X1 port map( A1 => regs(1440), A2 => n186, B1 => regs(2464), B2
                           => n249, ZN => n585);
   U745 : NAND2_X1 port map( A1 => n587, A2 => n588, ZN => curr_proc_regs(415))
                           ;
   U746 : AOI222_X1 port map( A1 => regs(415), A2 => n30, B1 => regs(1951), B2 
                           => n82, C1 => regs(927), C2 => n134, ZN => n588);
   U747 : AOI22_X1 port map( A1 => regs(1439), A2 => n186, B1 => regs(2463), B2
                           => n248, ZN => n587);
   U748 : NAND2_X1 port map( A1 => n589, A2 => n590, ZN => curr_proc_regs(414))
                           ;
   U749 : AOI222_X1 port map( A1 => regs(414), A2 => n30, B1 => regs(1950), B2 
                           => n82, C1 => regs(926), C2 => n134, ZN => n590);
   U750 : AOI22_X1 port map( A1 => regs(1438), A2 => n186, B1 => regs(2462), B2
                           => n249, ZN => n589);
   U751 : NAND2_X1 port map( A1 => n591, A2 => n592, ZN => curr_proc_regs(413))
                           ;
   U752 : AOI222_X1 port map( A1 => regs(413), A2 => n30, B1 => regs(1949), B2 
                           => n82, C1 => regs(925), C2 => n134, ZN => n592);
   U753 : AOI22_X1 port map( A1 => regs(1437), A2 => n186, B1 => regs(2461), B2
                           => n248, ZN => n591);
   U754 : NAND2_X1 port map( A1 => n593, A2 => n594, ZN => curr_proc_regs(412))
                           ;
   U755 : AOI222_X1 port map( A1 => regs(412), A2 => n29, B1 => regs(1948), B2 
                           => n81, C1 => regs(924), C2 => n133, ZN => n594);
   U756 : AOI22_X1 port map( A1 => regs(1436), A2 => n185, B1 => regs(2460), B2
                           => n248, ZN => n593);
   U757 : NAND2_X1 port map( A1 => n595, A2 => n596, ZN => curr_proc_regs(411))
                           ;
   U758 : AOI222_X1 port map( A1 => regs(411), A2 => n29, B1 => regs(1947), B2 
                           => n81, C1 => regs(923), C2 => n133, ZN => n596);
   U759 : AOI22_X1 port map( A1 => regs(1435), A2 => n185, B1 => regs(2459), B2
                           => n248, ZN => n595);
   U760 : NAND2_X1 port map( A1 => n597, A2 => n598, ZN => curr_proc_regs(410))
                           ;
   U761 : AOI222_X1 port map( A1 => regs(410), A2 => n29, B1 => regs(1946), B2 
                           => n81, C1 => regs(922), C2 => n133, ZN => n598);
   U762 : AOI22_X1 port map( A1 => regs(1434), A2 => n185, B1 => regs(2458), B2
                           => n248, ZN => n597);
   U763 : NAND2_X1 port map( A1 => n599, A2 => n600, ZN => curr_proc_regs(40));
   U764 : AOI222_X1 port map( A1 => regs(40), A2 => n29, B1 => regs(1576), B2 
                           => n81, C1 => regs(552), C2 => n133, ZN => n600);
   U765 : AOI22_X1 port map( A1 => regs(1064), A2 => n185, B1 => regs(2088), B2
                           => n248, ZN => n599);
   U766 : NAND2_X1 port map( A1 => n601, A2 => n602, ZN => curr_proc_regs(409))
                           ;
   U767 : AOI222_X1 port map( A1 => regs(409), A2 => n29, B1 => regs(1945), B2 
                           => n81, C1 => regs(921), C2 => n133, ZN => n602);
   U768 : AOI22_X1 port map( A1 => regs(1433), A2 => n185, B1 => regs(2457), B2
                           => n248, ZN => n601);
   U769 : NAND2_X1 port map( A1 => n603, A2 => n604, ZN => curr_proc_regs(408))
                           ;
   U770 : AOI222_X1 port map( A1 => regs(408), A2 => n29, B1 => regs(1944), B2 
                           => n81, C1 => regs(920), C2 => n133, ZN => n604);
   U771 : AOI22_X1 port map( A1 => regs(1432), A2 => n185, B1 => regs(2456), B2
                           => n248, ZN => n603);
   U772 : NAND2_X1 port map( A1 => n605, A2 => n606, ZN => curr_proc_regs(407))
                           ;
   U773 : AOI222_X1 port map( A1 => regs(407), A2 => n29, B1 => regs(1943), B2 
                           => n81, C1 => regs(919), C2 => n133, ZN => n606);
   U774 : AOI22_X1 port map( A1 => regs(1431), A2 => n185, B1 => regs(2455), B2
                           => n248, ZN => n605);
   U775 : NAND2_X1 port map( A1 => n607, A2 => n608, ZN => curr_proc_regs(406))
                           ;
   U776 : AOI222_X1 port map( A1 => regs(406), A2 => n29, B1 => regs(1942), B2 
                           => n81, C1 => regs(918), C2 => n133, ZN => n608);
   U777 : AOI22_X1 port map( A1 => regs(1430), A2 => n185, B1 => regs(2454), B2
                           => n248, ZN => n607);
   U778 : NAND2_X1 port map( A1 => n609, A2 => n610, ZN => curr_proc_regs(405))
                           ;
   U779 : AOI222_X1 port map( A1 => regs(405), A2 => n29, B1 => regs(1941), B2 
                           => n81, C1 => regs(917), C2 => n133, ZN => n610);
   U780 : AOI22_X1 port map( A1 => regs(1429), A2 => n185, B1 => regs(2453), B2
                           => n248, ZN => n609);
   U781 : NAND2_X1 port map( A1 => n611, A2 => n612, ZN => curr_proc_regs(404))
                           ;
   U782 : AOI222_X1 port map( A1 => regs(404), A2 => n29, B1 => regs(1940), B2 
                           => n81, C1 => regs(916), C2 => n133, ZN => n612);
   U783 : AOI22_X1 port map( A1 => regs(1428), A2 => n185, B1 => regs(2452), B2
                           => n247, ZN => n611);
   U784 : NAND2_X1 port map( A1 => n613, A2 => n614, ZN => curr_proc_regs(403))
                           ;
   U785 : AOI222_X1 port map( A1 => regs(403), A2 => n29, B1 => regs(1939), B2 
                           => n81, C1 => regs(915), C2 => n133, ZN => n614);
   U786 : AOI22_X1 port map( A1 => regs(1427), A2 => n185, B1 => regs(2451), B2
                           => n248, ZN => n613);
   U787 : NAND2_X1 port map( A1 => n615, A2 => n616, ZN => curr_proc_regs(402))
                           ;
   U788 : AOI222_X1 port map( A1 => regs(402), A2 => n29, B1 => regs(1938), B2 
                           => n81, C1 => regs(914), C2 => n133, ZN => n616);
   U789 : AOI22_X1 port map( A1 => regs(1426), A2 => n185, B1 => regs(2450), B2
                           => n247, ZN => n615);
   U790 : NAND2_X1 port map( A1 => n617, A2 => n618, ZN => curr_proc_regs(401))
                           ;
   U791 : AOI222_X1 port map( A1 => regs(401), A2 => n28, B1 => regs(1937), B2 
                           => n80, C1 => regs(913), C2 => n132, ZN => n618);
   U792 : AOI22_X1 port map( A1 => regs(1425), A2 => n184, B1 => regs(2449), B2
                           => n247, ZN => n617);
   U793 : NAND2_X1 port map( A1 => n619, A2 => n620, ZN => curr_proc_regs(400))
                           ;
   U794 : AOI222_X1 port map( A1 => regs(400), A2 => n28, B1 => regs(1936), B2 
                           => n80, C1 => regs(912), C2 => n132, ZN => n620);
   U795 : AOI22_X1 port map( A1 => regs(1424), A2 => n184, B1 => regs(2448), B2
                           => n247, ZN => n619);
   U796 : NAND2_X1 port map( A1 => n621, A2 => n622, ZN => curr_proc_regs(3));
   U797 : AOI222_X1 port map( A1 => regs(3), A2 => n28, B1 => regs(1539), B2 =>
                           n80, C1 => regs(515), C2 => n132, ZN => n622);
   U798 : AOI22_X1 port map( A1 => regs(1027), A2 => n184, B1 => regs(2051), B2
                           => n247, ZN => n621);
   U799 : NAND2_X1 port map( A1 => n623, A2 => n624, ZN => curr_proc_regs(39));
   U800 : AOI222_X1 port map( A1 => regs(39), A2 => n28, B1 => regs(1575), B2 
                           => n80, C1 => regs(551), C2 => n132, ZN => n624);
   U801 : AOI22_X1 port map( A1 => regs(1063), A2 => n184, B1 => regs(2087), B2
                           => n247, ZN => n623);
   U802 : NAND2_X1 port map( A1 => n625, A2 => n626, ZN => curr_proc_regs(399))
                           ;
   U803 : AOI222_X1 port map( A1 => regs(399), A2 => n28, B1 => regs(1935), B2 
                           => n80, C1 => regs(911), C2 => n132, ZN => n626);
   U804 : AOI22_X1 port map( A1 => regs(1423), A2 => n184, B1 => regs(2447), B2
                           => n247, ZN => n625);
   U805 : NAND2_X1 port map( A1 => n627, A2 => n628, ZN => curr_proc_regs(398))
                           ;
   U806 : AOI222_X1 port map( A1 => regs(398), A2 => n28, B1 => regs(1934), B2 
                           => n80, C1 => regs(910), C2 => n132, ZN => n628);
   U807 : AOI22_X1 port map( A1 => regs(1422), A2 => n184, B1 => regs(2446), B2
                           => n247, ZN => n627);
   U808 : NAND2_X1 port map( A1 => n629, A2 => n630, ZN => curr_proc_regs(397))
                           ;
   U809 : AOI222_X1 port map( A1 => regs(397), A2 => n28, B1 => regs(1933), B2 
                           => n80, C1 => regs(909), C2 => n132, ZN => n630);
   U810 : AOI22_X1 port map( A1 => regs(1421), A2 => n184, B1 => regs(2445), B2
                           => n247, ZN => n629);
   U811 : NAND2_X1 port map( A1 => n631, A2 => n632, ZN => curr_proc_regs(396))
                           ;
   U812 : AOI222_X1 port map( A1 => regs(396), A2 => n28, B1 => regs(1932), B2 
                           => n80, C1 => regs(908), C2 => n132, ZN => n632);
   U813 : AOI22_X1 port map( A1 => regs(1420), A2 => n184, B1 => regs(2444), B2
                           => n247, ZN => n631);
   U814 : NAND2_X1 port map( A1 => n633, A2 => n634, ZN => curr_proc_regs(395))
                           ;
   U815 : AOI222_X1 port map( A1 => regs(395), A2 => n28, B1 => regs(1931), B2 
                           => n80, C1 => regs(907), C2 => n132, ZN => n634);
   U816 : AOI22_X1 port map( A1 => regs(1419), A2 => n184, B1 => regs(2443), B2
                           => n247, ZN => n633);
   U817 : NAND2_X1 port map( A1 => n635, A2 => n636, ZN => curr_proc_regs(394))
                           ;
   U818 : AOI222_X1 port map( A1 => regs(394), A2 => n28, B1 => regs(1930), B2 
                           => n80, C1 => regs(906), C2 => n132, ZN => n636);
   U819 : AOI22_X1 port map( A1 => regs(1418), A2 => n184, B1 => regs(2442), B2
                           => n246, ZN => n635);
   U820 : NAND2_X1 port map( A1 => n637, A2 => n638, ZN => curr_proc_regs(393))
                           ;
   U821 : AOI222_X1 port map( A1 => regs(393), A2 => n28, B1 => regs(1929), B2 
                           => n80, C1 => regs(905), C2 => n132, ZN => n638);
   U822 : AOI22_X1 port map( A1 => regs(1417), A2 => n184, B1 => regs(2441), B2
                           => n247, ZN => n637);
   U823 : NAND2_X1 port map( A1 => n639, A2 => n640, ZN => curr_proc_regs(392))
                           ;
   U824 : AOI222_X1 port map( A1 => regs(392), A2 => n28, B1 => regs(1928), B2 
                           => n80, C1 => regs(904), C2 => n132, ZN => n640);
   U825 : AOI22_X1 port map( A1 => regs(1416), A2 => n184, B1 => regs(2440), B2
                           => n246, ZN => n639);
   U826 : NAND2_X1 port map( A1 => n641, A2 => n642, ZN => curr_proc_regs(391))
                           ;
   U827 : AOI222_X1 port map( A1 => regs(391), A2 => n27, B1 => regs(1927), B2 
                           => n79, C1 => regs(903), C2 => n131, ZN => n642);
   U828 : AOI22_X1 port map( A1 => regs(1415), A2 => n183, B1 => regs(2439), B2
                           => n246, ZN => n641);
   U829 : NAND2_X1 port map( A1 => n643, A2 => n644, ZN => curr_proc_regs(390))
                           ;
   U830 : AOI222_X1 port map( A1 => regs(390), A2 => n27, B1 => regs(1926), B2 
                           => n79, C1 => regs(902), C2 => n131, ZN => n644);
   U831 : AOI22_X1 port map( A1 => regs(1414), A2 => n183, B1 => regs(2438), B2
                           => n246, ZN => n643);
   U832 : NAND2_X1 port map( A1 => n645, A2 => n646, ZN => curr_proc_regs(38));
   U833 : AOI222_X1 port map( A1 => regs(38), A2 => n27, B1 => regs(1574), B2 
                           => n79, C1 => regs(550), C2 => n131, ZN => n646);
   U834 : AOI22_X1 port map( A1 => regs(1062), A2 => n183, B1 => regs(2086), B2
                           => n246, ZN => n645);
   U835 : NAND2_X1 port map( A1 => n647, A2 => n648, ZN => curr_proc_regs(389))
                           ;
   U836 : AOI222_X1 port map( A1 => regs(389), A2 => n27, B1 => regs(1925), B2 
                           => n79, C1 => regs(901), C2 => n131, ZN => n648);
   U837 : AOI22_X1 port map( A1 => regs(1413), A2 => n183, B1 => regs(2437), B2
                           => n246, ZN => n647);
   U838 : NAND2_X1 port map( A1 => n649, A2 => n650, ZN => curr_proc_regs(388))
                           ;
   U839 : AOI222_X1 port map( A1 => regs(388), A2 => n27, B1 => regs(1924), B2 
                           => n79, C1 => regs(900), C2 => n131, ZN => n650);
   U840 : AOI22_X1 port map( A1 => regs(1412), A2 => n183, B1 => regs(2436), B2
                           => n246, ZN => n649);
   U841 : NAND2_X1 port map( A1 => n651, A2 => n652, ZN => curr_proc_regs(387))
                           ;
   U842 : AOI222_X1 port map( A1 => regs(387), A2 => n27, B1 => regs(1923), B2 
                           => n79, C1 => regs(899), C2 => n131, ZN => n652);
   U843 : AOI22_X1 port map( A1 => regs(1411), A2 => n183, B1 => regs(2435), B2
                           => n246, ZN => n651);
   U844 : NAND2_X1 port map( A1 => n653, A2 => n654, ZN => curr_proc_regs(386))
                           ;
   U845 : AOI222_X1 port map( A1 => regs(386), A2 => n27, B1 => regs(1922), B2 
                           => n79, C1 => regs(898), C2 => n131, ZN => n654);
   U846 : AOI22_X1 port map( A1 => regs(1410), A2 => n183, B1 => regs(2434), B2
                           => n246, ZN => n653);
   U847 : NAND2_X1 port map( A1 => n655, A2 => n656, ZN => curr_proc_regs(385))
                           ;
   U848 : AOI222_X1 port map( A1 => regs(385), A2 => n27, B1 => regs(1921), B2 
                           => n79, C1 => regs(897), C2 => n131, ZN => n656);
   U849 : AOI22_X1 port map( A1 => regs(1409), A2 => n183, B1 => regs(2433), B2
                           => n246, ZN => n655);
   U850 : NAND2_X1 port map( A1 => n657, A2 => n658, ZN => curr_proc_regs(384))
                           ;
   U851 : AOI222_X1 port map( A1 => regs(384), A2 => n27, B1 => regs(1920), B2 
                           => n79, C1 => regs(896), C2 => n131, ZN => n658);
   U852 : AOI22_X1 port map( A1 => regs(1408), A2 => n183, B1 => regs(2432), B2
                           => n246, ZN => n657);
   U853 : NAND2_X1 port map( A1 => n659, A2 => n660, ZN => curr_proc_regs(383))
                           ;
   U854 : AOI222_X1 port map( A1 => regs(383), A2 => n27, B1 => regs(1919), B2 
                           => n79, C1 => regs(895), C2 => n131, ZN => n660);
   U855 : AOI22_X1 port map( A1 => regs(1407), A2 => n183, B1 => regs(2431), B2
                           => n245, ZN => n659);
   U856 : NAND2_X1 port map( A1 => n661, A2 => n662, ZN => curr_proc_regs(382))
                           ;
   U857 : AOI222_X1 port map( A1 => regs(382), A2 => n27, B1 => regs(1918), B2 
                           => n79, C1 => regs(894), C2 => n131, ZN => n662);
   U858 : AOI22_X1 port map( A1 => regs(1406), A2 => n183, B1 => regs(2430), B2
                           => n245, ZN => n661);
   U859 : NAND2_X1 port map( A1 => n663, A2 => n664, ZN => curr_proc_regs(381))
                           ;
   U860 : AOI222_X1 port map( A1 => regs(381), A2 => n27, B1 => regs(1917), B2 
                           => n79, C1 => regs(893), C2 => n131, ZN => n664);
   U861 : AOI22_X1 port map( A1 => regs(1405), A2 => n183, B1 => regs(2429), B2
                           => n245, ZN => n663);
   U862 : NAND2_X1 port map( A1 => n665, A2 => n666, ZN => curr_proc_regs(380))
                           ;
   U863 : AOI222_X1 port map( A1 => regs(380), A2 => n26, B1 => regs(1916), B2 
                           => n78, C1 => regs(892), C2 => n130, ZN => n666);
   U864 : AOI22_X1 port map( A1 => regs(1404), A2 => n182, B1 => regs(2428), B2
                           => n245, ZN => n665);
   U865 : NAND2_X1 port map( A1 => n667, A2 => n668, ZN => curr_proc_regs(37));
   U866 : AOI222_X1 port map( A1 => regs(37), A2 => n26, B1 => regs(1573), B2 
                           => n78, C1 => regs(549), C2 => n130, ZN => n668);
   U867 : AOI22_X1 port map( A1 => regs(1061), A2 => n182, B1 => regs(2085), B2
                           => n245, ZN => n667);
   U868 : NAND2_X1 port map( A1 => n669, A2 => n670, ZN => curr_proc_regs(379))
                           ;
   U869 : AOI222_X1 port map( A1 => regs(379), A2 => n26, B1 => regs(1915), B2 
                           => n78, C1 => regs(891), C2 => n130, ZN => n670);
   U870 : AOI22_X1 port map( A1 => regs(1403), A2 => n182, B1 => regs(2427), B2
                           => n245, ZN => n669);
   U871 : NAND2_X1 port map( A1 => n671, A2 => n672, ZN => curr_proc_regs(378))
                           ;
   U872 : AOI222_X1 port map( A1 => regs(378), A2 => n26, B1 => regs(1914), B2 
                           => n78, C1 => regs(890), C2 => n130, ZN => n672);
   U873 : AOI22_X1 port map( A1 => regs(1402), A2 => n182, B1 => regs(2426), B2
                           => n245, ZN => n671);
   U874 : NAND2_X1 port map( A1 => n673, A2 => n674, ZN => curr_proc_regs(377))
                           ;
   U875 : AOI222_X1 port map( A1 => regs(377), A2 => n26, B1 => regs(1913), B2 
                           => n78, C1 => regs(889), C2 => n130, ZN => n674);
   U876 : AOI22_X1 port map( A1 => regs(1401), A2 => n182, B1 => regs(2425), B2
                           => n245, ZN => n673);
   U877 : NAND2_X1 port map( A1 => n675, A2 => n676, ZN => curr_proc_regs(376))
                           ;
   U878 : AOI222_X1 port map( A1 => regs(376), A2 => n26, B1 => regs(1912), B2 
                           => n78, C1 => regs(888), C2 => n130, ZN => n676);
   U879 : AOI22_X1 port map( A1 => regs(1400), A2 => n182, B1 => regs(2424), B2
                           => n245, ZN => n675);
   U880 : NAND2_X1 port map( A1 => n677, A2 => n678, ZN => curr_proc_regs(375))
                           ;
   U881 : AOI222_X1 port map( A1 => regs(375), A2 => n26, B1 => regs(1911), B2 
                           => n78, C1 => regs(887), C2 => n130, ZN => n678);
   U882 : AOI22_X1 port map( A1 => regs(1399), A2 => n182, B1 => regs(2423), B2
                           => n245, ZN => n677);
   U883 : NAND2_X1 port map( A1 => n679, A2 => n680, ZN => curr_proc_regs(374))
                           ;
   U884 : AOI222_X1 port map( A1 => regs(374), A2 => n26, B1 => regs(1910), B2 
                           => n78, C1 => regs(886), C2 => n130, ZN => n680);
   U885 : AOI22_X1 port map( A1 => regs(1398), A2 => n182, B1 => regs(2422), B2
                           => n245, ZN => n679);
   U886 : NAND2_X1 port map( A1 => n681, A2 => n682, ZN => curr_proc_regs(373))
                           ;
   U887 : AOI222_X1 port map( A1 => regs(373), A2 => n26, B1 => regs(1909), B2 
                           => n78, C1 => regs(885), C2 => n130, ZN => n682);
   U888 : AOI22_X1 port map( A1 => regs(1397), A2 => n182, B1 => regs(2421), B2
                           => n245, ZN => n681);
   U889 : NAND2_X1 port map( A1 => n683, A2 => n684, ZN => curr_proc_regs(372))
                           ;
   U890 : AOI222_X1 port map( A1 => regs(372), A2 => n26, B1 => regs(1908), B2 
                           => n78, C1 => regs(884), C2 => n130, ZN => n684);
   U891 : AOI22_X1 port map( A1 => regs(1396), A2 => n182, B1 => regs(2420), B2
                           => n244, ZN => n683);
   U892 : NAND2_X1 port map( A1 => n685, A2 => n686, ZN => curr_proc_regs(371))
                           ;
   U893 : AOI222_X1 port map( A1 => regs(371), A2 => n26, B1 => regs(1907), B2 
                           => n78, C1 => regs(883), C2 => n130, ZN => n686);
   U894 : AOI22_X1 port map( A1 => regs(1395), A2 => n182, B1 => regs(2419), B2
                           => n244, ZN => n685);
   U895 : NAND2_X1 port map( A1 => n687, A2 => n688, ZN => curr_proc_regs(370))
                           ;
   U896 : AOI222_X1 port map( A1 => regs(370), A2 => n26, B1 => regs(1906), B2 
                           => n78, C1 => regs(882), C2 => n130, ZN => n688);
   U897 : AOI22_X1 port map( A1 => regs(1394), A2 => n182, B1 => regs(2418), B2
                           => n244, ZN => n687);
   U898 : NAND2_X1 port map( A1 => n689, A2 => n690, ZN => curr_proc_regs(36));
   U899 : AOI222_X1 port map( A1 => regs(36), A2 => n25, B1 => regs(1572), B2 
                           => n77, C1 => regs(548), C2 => n129, ZN => n690);
   U900 : AOI22_X1 port map( A1 => regs(1060), A2 => n181, B1 => regs(2084), B2
                           => n244, ZN => n689);
   U901 : NAND2_X1 port map( A1 => n691, A2 => n692, ZN => curr_proc_regs(369))
                           ;
   U902 : AOI222_X1 port map( A1 => regs(369), A2 => n25, B1 => regs(1905), B2 
                           => n77, C1 => regs(881), C2 => n129, ZN => n692);
   U903 : AOI22_X1 port map( A1 => regs(1393), A2 => n181, B1 => regs(2417), B2
                           => n244, ZN => n691);
   U904 : NAND2_X1 port map( A1 => n693, A2 => n694, ZN => curr_proc_regs(368))
                           ;
   U905 : AOI222_X1 port map( A1 => regs(368), A2 => n25, B1 => regs(1904), B2 
                           => n77, C1 => regs(880), C2 => n129, ZN => n694);
   U906 : AOI22_X1 port map( A1 => regs(1392), A2 => n181, B1 => regs(2416), B2
                           => n244, ZN => n693);
   U907 : NAND2_X1 port map( A1 => n695, A2 => n696, ZN => curr_proc_regs(367))
                           ;
   U908 : AOI222_X1 port map( A1 => regs(367), A2 => n25, B1 => regs(1903), B2 
                           => n77, C1 => regs(879), C2 => n129, ZN => n696);
   U909 : AOI22_X1 port map( A1 => regs(1391), A2 => n181, B1 => regs(2415), B2
                           => n244, ZN => n695);
   U910 : NAND2_X1 port map( A1 => n697, A2 => n698, ZN => curr_proc_regs(366))
                           ;
   U911 : AOI222_X1 port map( A1 => regs(366), A2 => n25, B1 => regs(1902), B2 
                           => n77, C1 => regs(878), C2 => n129, ZN => n698);
   U912 : AOI22_X1 port map( A1 => regs(1390), A2 => n181, B1 => regs(2414), B2
                           => n244, ZN => n697);
   U913 : NAND2_X1 port map( A1 => n699, A2 => n700, ZN => curr_proc_regs(365))
                           ;
   U914 : AOI222_X1 port map( A1 => regs(365), A2 => n25, B1 => regs(1901), B2 
                           => n77, C1 => regs(877), C2 => n129, ZN => n700);
   U915 : AOI22_X1 port map( A1 => regs(1389), A2 => n181, B1 => regs(2413), B2
                           => n244, ZN => n699);
   U916 : NAND2_X1 port map( A1 => n701, A2 => n702, ZN => curr_proc_regs(364))
                           ;
   U917 : AOI222_X1 port map( A1 => regs(364), A2 => n25, B1 => regs(1900), B2 
                           => n77, C1 => regs(876), C2 => n129, ZN => n702);
   U918 : AOI22_X1 port map( A1 => regs(1388), A2 => n181, B1 => regs(2412), B2
                           => n244, ZN => n701);
   U919 : NAND2_X1 port map( A1 => n703, A2 => n704, ZN => curr_proc_regs(363))
                           ;
   U920 : AOI222_X1 port map( A1 => regs(363), A2 => n25, B1 => regs(1899), B2 
                           => n77, C1 => regs(875), C2 => n129, ZN => n704);
   U921 : AOI22_X1 port map( A1 => regs(1387), A2 => n181, B1 => regs(2411), B2
                           => n244, ZN => n703);
   U922 : NAND2_X1 port map( A1 => n705, A2 => n706, ZN => curr_proc_regs(362))
                           ;
   U923 : AOI222_X1 port map( A1 => regs(362), A2 => n25, B1 => regs(1898), B2 
                           => n77, C1 => regs(874), C2 => n129, ZN => n706);
   U924 : AOI22_X1 port map( A1 => regs(1386), A2 => n181, B1 => regs(2410), B2
                           => n244, ZN => n705);
   U925 : NAND2_X1 port map( A1 => n707, A2 => n708, ZN => curr_proc_regs(361))
                           ;
   U926 : AOI222_X1 port map( A1 => regs(361), A2 => n25, B1 => regs(1897), B2 
                           => n77, C1 => regs(873), C2 => n129, ZN => n708);
   U927 : AOI22_X1 port map( A1 => regs(1385), A2 => n181, B1 => regs(2409), B2
                           => n243, ZN => n707);
   U928 : NAND2_X1 port map( A1 => n709, A2 => n710, ZN => curr_proc_regs(360))
                           ;
   U929 : AOI222_X1 port map( A1 => regs(360), A2 => n25, B1 => regs(1896), B2 
                           => n77, C1 => regs(872), C2 => n129, ZN => n710);
   U930 : AOI22_X1 port map( A1 => regs(1384), A2 => n181, B1 => regs(2408), B2
                           => n243, ZN => n709);
   U931 : NAND2_X1 port map( A1 => n711, A2 => n712, ZN => curr_proc_regs(35));
   U932 : AOI222_X1 port map( A1 => regs(35), A2 => n25, B1 => regs(1571), B2 
                           => n77, C1 => regs(547), C2 => n129, ZN => n712);
   U933 : AOI22_X1 port map( A1 => regs(1059), A2 => n181, B1 => regs(2083), B2
                           => n243, ZN => n711);
   U934 : NAND2_X1 port map( A1 => n713, A2 => n714, ZN => curr_proc_regs(359))
                           ;
   U935 : AOI222_X1 port map( A1 => regs(359), A2 => n24, B1 => regs(1895), B2 
                           => n76, C1 => regs(871), C2 => n128, ZN => n714);
   U936 : AOI22_X1 port map( A1 => regs(1383), A2 => n180, B1 => regs(2407), B2
                           => n243, ZN => n713);
   U937 : NAND2_X1 port map( A1 => n715, A2 => n716, ZN => curr_proc_regs(358))
                           ;
   U938 : AOI222_X1 port map( A1 => regs(358), A2 => n24, B1 => regs(1894), B2 
                           => n76, C1 => regs(870), C2 => n128, ZN => n716);
   U939 : AOI22_X1 port map( A1 => regs(1382), A2 => n180, B1 => regs(2406), B2
                           => n243, ZN => n715);
   U940 : NAND2_X1 port map( A1 => n717, A2 => n718, ZN => curr_proc_regs(357))
                           ;
   U941 : AOI222_X1 port map( A1 => regs(357), A2 => n24, B1 => regs(1893), B2 
                           => n76, C1 => regs(869), C2 => n128, ZN => n718);
   U942 : AOI22_X1 port map( A1 => regs(1381), A2 => n180, B1 => regs(2405), B2
                           => n243, ZN => n717);
   U943 : NAND2_X1 port map( A1 => n719, A2 => n720, ZN => curr_proc_regs(356))
                           ;
   U944 : AOI222_X1 port map( A1 => regs(356), A2 => n24, B1 => regs(1892), B2 
                           => n76, C1 => regs(868), C2 => n128, ZN => n720);
   U945 : AOI22_X1 port map( A1 => regs(1380), A2 => n180, B1 => regs(2404), B2
                           => n243, ZN => n719);
   U946 : NAND2_X1 port map( A1 => n721, A2 => n722, ZN => curr_proc_regs(355))
                           ;
   U947 : AOI222_X1 port map( A1 => regs(355), A2 => n24, B1 => regs(1891), B2 
                           => n76, C1 => regs(867), C2 => n128, ZN => n722);
   U948 : AOI22_X1 port map( A1 => regs(1379), A2 => n180, B1 => regs(2403), B2
                           => n243, ZN => n721);
   U949 : NAND2_X1 port map( A1 => n723, A2 => n724, ZN => curr_proc_regs(354))
                           ;
   U950 : AOI222_X1 port map( A1 => regs(354), A2 => n24, B1 => regs(1890), B2 
                           => n76, C1 => regs(866), C2 => n128, ZN => n724);
   U951 : AOI22_X1 port map( A1 => regs(1378), A2 => n180, B1 => regs(2402), B2
                           => n243, ZN => n723);
   U952 : NAND2_X1 port map( A1 => n725, A2 => n726, ZN => curr_proc_regs(353))
                           ;
   U953 : AOI222_X1 port map( A1 => regs(353), A2 => n24, B1 => regs(1889), B2 
                           => n76, C1 => regs(865), C2 => n128, ZN => n726);
   U954 : AOI22_X1 port map( A1 => regs(1377), A2 => n180, B1 => regs(2401), B2
                           => n243, ZN => n725);
   U955 : NAND2_X1 port map( A1 => n727, A2 => n728, ZN => curr_proc_regs(352))
                           ;
   U956 : AOI222_X1 port map( A1 => regs(352), A2 => n24, B1 => regs(1888), B2 
                           => n76, C1 => regs(864), C2 => n128, ZN => n728);
   U957 : AOI22_X1 port map( A1 => regs(1376), A2 => n180, B1 => regs(2400), B2
                           => n243, ZN => n727);
   U958 : NAND2_X1 port map( A1 => n729, A2 => n730, ZN => curr_proc_regs(351))
                           ;
   U959 : AOI222_X1 port map( A1 => regs(351), A2 => n24, B1 => regs(1887), B2 
                           => n76, C1 => regs(863), C2 => n128, ZN => n730);
   U960 : AOI22_X1 port map( A1 => regs(1375), A2 => n180, B1 => regs(2399), B2
                           => n243, ZN => n729);
   U961 : NAND2_X1 port map( A1 => n731, A2 => n732, ZN => curr_proc_regs(350))
                           ;
   U962 : AOI222_X1 port map( A1 => regs(350), A2 => n24, B1 => regs(1886), B2 
                           => n76, C1 => regs(862), C2 => n128, ZN => n732);
   U963 : AOI22_X1 port map( A1 => regs(1374), A2 => n180, B1 => regs(2398), B2
                           => n242, ZN => n731);
   U964 : NAND2_X1 port map( A1 => n733, A2 => n734, ZN => curr_proc_regs(34));
   U965 : AOI222_X1 port map( A1 => regs(34), A2 => n24, B1 => regs(1570), B2 
                           => n76, C1 => regs(546), C2 => n128, ZN => n734);
   U966 : AOI22_X1 port map( A1 => regs(1058), A2 => n180, B1 => regs(2082), B2
                           => n242, ZN => n733);
   U967 : NAND2_X1 port map( A1 => n735, A2 => n736, ZN => curr_proc_regs(349))
                           ;
   U968 : AOI222_X1 port map( A1 => regs(349), A2 => n24, B1 => regs(1885), B2 
                           => n76, C1 => regs(861), C2 => n128, ZN => n736);
   U969 : AOI22_X1 port map( A1 => regs(1373), A2 => n180, B1 => regs(2397), B2
                           => n242, ZN => n735);
   U970 : NAND2_X1 port map( A1 => n737, A2 => n738, ZN => curr_proc_regs(348))
                           ;
   U971 : AOI222_X1 port map( A1 => regs(348), A2 => n23, B1 => regs(1884), B2 
                           => n75, C1 => regs(860), C2 => n127, ZN => n738);
   U972 : AOI22_X1 port map( A1 => regs(1372), A2 => n179, B1 => regs(2396), B2
                           => n242, ZN => n737);
   U973 : NAND2_X1 port map( A1 => n739, A2 => n740, ZN => curr_proc_regs(347))
                           ;
   U974 : AOI222_X1 port map( A1 => regs(347), A2 => n23, B1 => regs(1883), B2 
                           => n75, C1 => regs(859), C2 => n127, ZN => n740);
   U975 : AOI22_X1 port map( A1 => regs(1371), A2 => n179, B1 => regs(2395), B2
                           => n242, ZN => n739);
   U976 : NAND2_X1 port map( A1 => n741, A2 => n742, ZN => curr_proc_regs(346))
                           ;
   U977 : AOI222_X1 port map( A1 => regs(346), A2 => n23, B1 => regs(1882), B2 
                           => n75, C1 => regs(858), C2 => n127, ZN => n742);
   U978 : AOI22_X1 port map( A1 => regs(1370), A2 => n179, B1 => regs(2394), B2
                           => n242, ZN => n741);
   U979 : NAND2_X1 port map( A1 => n743, A2 => n744, ZN => curr_proc_regs(345))
                           ;
   U980 : AOI222_X1 port map( A1 => regs(345), A2 => n23, B1 => regs(1881), B2 
                           => n75, C1 => regs(857), C2 => n127, ZN => n744);
   U981 : AOI22_X1 port map( A1 => regs(1369), A2 => n179, B1 => regs(2393), B2
                           => n242, ZN => n743);
   U982 : NAND2_X1 port map( A1 => n745, A2 => n746, ZN => curr_proc_regs(344))
                           ;
   U983 : AOI222_X1 port map( A1 => regs(344), A2 => n23, B1 => regs(1880), B2 
                           => n75, C1 => regs(856), C2 => n127, ZN => n746);
   U984 : AOI22_X1 port map( A1 => regs(1368), A2 => n179, B1 => regs(2392), B2
                           => n242, ZN => n745);
   U985 : NAND2_X1 port map( A1 => n747, A2 => n748, ZN => curr_proc_regs(343))
                           ;
   U986 : AOI222_X1 port map( A1 => regs(343), A2 => n23, B1 => regs(1879), B2 
                           => n75, C1 => regs(855), C2 => n127, ZN => n748);
   U987 : AOI22_X1 port map( A1 => regs(1367), A2 => n179, B1 => regs(2391), B2
                           => n242, ZN => n747);
   U988 : NAND2_X1 port map( A1 => n749, A2 => n750, ZN => curr_proc_regs(342))
                           ;
   U989 : AOI222_X1 port map( A1 => regs(342), A2 => n23, B1 => regs(1878), B2 
                           => n75, C1 => regs(854), C2 => n127, ZN => n750);
   U990 : AOI22_X1 port map( A1 => regs(1366), A2 => n179, B1 => regs(2390), B2
                           => n242, ZN => n749);
   U991 : NAND2_X1 port map( A1 => n751, A2 => n752, ZN => curr_proc_regs(341))
                           ;
   U992 : AOI222_X1 port map( A1 => regs(341), A2 => n23, B1 => regs(1877), B2 
                           => n75, C1 => regs(853), C2 => n127, ZN => n752);
   U993 : AOI22_X1 port map( A1 => regs(1365), A2 => n179, B1 => regs(2389), B2
                           => n242, ZN => n751);
   U994 : NAND2_X1 port map( A1 => n753, A2 => n754, ZN => curr_proc_regs(340))
                           ;
   U995 : AOI222_X1 port map( A1 => regs(340), A2 => n23, B1 => regs(1876), B2 
                           => n75, C1 => regs(852), C2 => n127, ZN => n754);
   U996 : AOI22_X1 port map( A1 => regs(1364), A2 => n179, B1 => regs(2388), B2
                           => n242, ZN => n753);
   U997 : NAND2_X1 port map( A1 => n755, A2 => n756, ZN => curr_proc_regs(33));
   U998 : AOI222_X1 port map( A1 => regs(33), A2 => n23, B1 => regs(1569), B2 
                           => n75, C1 => regs(545), C2 => n127, ZN => n756);
   U999 : AOI22_X1 port map( A1 => regs(1057), A2 => n179, B1 => regs(2081), B2
                           => n241, ZN => n755);
   U1000 : NAND2_X1 port map( A1 => n757, A2 => n758, ZN => curr_proc_regs(339)
                           );
   U1001 : AOI222_X1 port map( A1 => regs(339), A2 => n23, B1 => regs(1875), B2
                           => n75, C1 => regs(851), C2 => n127, ZN => n758);
   U1002 : AOI22_X1 port map( A1 => regs(1363), A2 => n179, B1 => regs(2387), 
                           B2 => n241, ZN => n757);
   U1003 : NAND2_X1 port map( A1 => n759, A2 => n760, ZN => curr_proc_regs(338)
                           );
   U1004 : AOI222_X1 port map( A1 => regs(338), A2 => n23, B1 => regs(1874), B2
                           => n75, C1 => regs(850), C2 => n127, ZN => n760);
   U1005 : AOI22_X1 port map( A1 => regs(1362), A2 => n179, B1 => regs(2386), 
                           B2 => n241, ZN => n759);
   U1006 : NAND2_X1 port map( A1 => n761, A2 => n762, ZN => curr_proc_regs(337)
                           );
   U1007 : AOI222_X1 port map( A1 => regs(337), A2 => n22, B1 => regs(1873), B2
                           => n74, C1 => regs(849), C2 => n126, ZN => n762);
   U1008 : AOI22_X1 port map( A1 => regs(1361), A2 => n178, B1 => regs(2385), 
                           B2 => n241, ZN => n761);
   U1009 : NAND2_X1 port map( A1 => n763, A2 => n764, ZN => curr_proc_regs(336)
                           );
   U1010 : AOI222_X1 port map( A1 => regs(336), A2 => n22, B1 => regs(1872), B2
                           => n74, C1 => regs(848), C2 => n126, ZN => n764);
   U1011 : AOI22_X1 port map( A1 => regs(1360), A2 => n178, B1 => regs(2384), 
                           B2 => n241, ZN => n763);
   U1012 : NAND2_X1 port map( A1 => n765, A2 => n766, ZN => curr_proc_regs(335)
                           );
   U1013 : AOI222_X1 port map( A1 => regs(335), A2 => n22, B1 => regs(1871), B2
                           => n74, C1 => regs(847), C2 => n126, ZN => n766);
   U1014 : AOI22_X1 port map( A1 => regs(1359), A2 => n178, B1 => regs(2383), 
                           B2 => n241, ZN => n765);
   U1015 : NAND2_X1 port map( A1 => n767, A2 => n768, ZN => curr_proc_regs(334)
                           );
   U1016 : AOI222_X1 port map( A1 => regs(334), A2 => n22, B1 => regs(1870), B2
                           => n74, C1 => regs(846), C2 => n126, ZN => n768);
   U1017 : AOI22_X1 port map( A1 => regs(1358), A2 => n178, B1 => regs(2382), 
                           B2 => n241, ZN => n767);
   U1018 : NAND2_X1 port map( A1 => n769, A2 => n770, ZN => curr_proc_regs(333)
                           );
   U1019 : AOI222_X1 port map( A1 => regs(333), A2 => n22, B1 => regs(1869), B2
                           => n74, C1 => regs(845), C2 => n126, ZN => n770);
   U1020 : AOI22_X1 port map( A1 => regs(1357), A2 => n178, B1 => regs(2381), 
                           B2 => n241, ZN => n769);
   U1021 : NAND2_X1 port map( A1 => n771, A2 => n772, ZN => curr_proc_regs(332)
                           );
   U1022 : AOI222_X1 port map( A1 => regs(332), A2 => n22, B1 => regs(1868), B2
                           => n74, C1 => regs(844), C2 => n126, ZN => n772);
   U1023 : AOI22_X1 port map( A1 => regs(1356), A2 => n178, B1 => regs(2380), 
                           B2 => n241, ZN => n771);
   U1024 : NAND2_X1 port map( A1 => n773, A2 => n774, ZN => curr_proc_regs(331)
                           );
   U1025 : AOI222_X1 port map( A1 => regs(331), A2 => n22, B1 => regs(1867), B2
                           => n74, C1 => regs(843), C2 => n126, ZN => n774);
   U1026 : AOI22_X1 port map( A1 => regs(1355), A2 => n178, B1 => regs(2379), 
                           B2 => n241, ZN => n773);
   U1027 : NAND2_X1 port map( A1 => n775, A2 => n776, ZN => curr_proc_regs(330)
                           );
   U1028 : AOI222_X1 port map( A1 => regs(330), A2 => n22, B1 => regs(1866), B2
                           => n74, C1 => regs(842), C2 => n126, ZN => n776);
   U1029 : AOI22_X1 port map( A1 => regs(1354), A2 => n178, B1 => regs(2378), 
                           B2 => n241, ZN => n775);
   U1030 : NAND2_X1 port map( A1 => n777, A2 => n778, ZN => curr_proc_regs(32))
                           ;
   U1031 : AOI222_X1 port map( A1 => regs(32), A2 => n22, B1 => regs(1568), B2 
                           => n74, C1 => regs(544), C2 => n126, ZN => n778);
   U1032 : AOI22_X1 port map( A1 => regs(1056), A2 => n178, B1 => regs(2080), 
                           B2 => n246, ZN => n777);
   U1033 : NAND2_X1 port map( A1 => n779, A2 => n780, ZN => curr_proc_regs(329)
                           );
   U1034 : AOI222_X1 port map( A1 => regs(329), A2 => n22, B1 => regs(1865), B2
                           => n74, C1 => regs(841), C2 => n126, ZN => n780);
   U1035 : AOI22_X1 port map( A1 => regs(1353), A2 => n178, B1 => regs(2377), 
                           B2 => n219, ZN => n779);
   U1036 : NAND2_X1 port map( A1 => n781, A2 => n782, ZN => curr_proc_regs(328)
                           );
   U1037 : AOI222_X1 port map( A1 => regs(328), A2 => n22, B1 => regs(1864), B2
                           => n74, C1 => regs(840), C2 => n126, ZN => n782);
   U1038 : AOI22_X1 port map( A1 => regs(1352), A2 => n178, B1 => regs(2376), 
                           B2 => n219, ZN => n781);
   U1039 : NAND2_X1 port map( A1 => n783, A2 => n784, ZN => curr_proc_regs(327)
                           );
   U1040 : AOI222_X1 port map( A1 => regs(327), A2 => n22, B1 => regs(1863), B2
                           => n74, C1 => regs(839), C2 => n126, ZN => n784);
   U1041 : AOI22_X1 port map( A1 => regs(1351), A2 => n178, B1 => regs(2375), 
                           B2 => n219, ZN => n783);
   U1042 : NAND2_X1 port map( A1 => n785, A2 => n786, ZN => curr_proc_regs(326)
                           );
   U1043 : AOI222_X1 port map( A1 => regs(326), A2 => n21, B1 => regs(1862), B2
                           => n73, C1 => regs(838), C2 => n125, ZN => n786);
   U1044 : AOI22_X1 port map( A1 => regs(1350), A2 => n177, B1 => regs(2374), 
                           B2 => n219, ZN => n785);
   U1045 : NAND2_X1 port map( A1 => n787, A2 => n788, ZN => curr_proc_regs(325)
                           );
   U1046 : AOI222_X1 port map( A1 => regs(325), A2 => n21, B1 => regs(1861), B2
                           => n73, C1 => regs(837), C2 => n125, ZN => n788);
   U1047 : AOI22_X1 port map( A1 => regs(1349), A2 => n177, B1 => regs(2373), 
                           B2 => n219, ZN => n787);
   U1048 : NAND2_X1 port map( A1 => n789, A2 => n790, ZN => curr_proc_regs(324)
                           );
   U1049 : AOI222_X1 port map( A1 => regs(324), A2 => n21, B1 => regs(1860), B2
                           => n73, C1 => regs(836), C2 => n125, ZN => n790);
   U1050 : AOI22_X1 port map( A1 => regs(1348), A2 => n177, B1 => regs(2372), 
                           B2 => n219, ZN => n789);
   U1051 : NAND2_X1 port map( A1 => n791, A2 => n792, ZN => curr_proc_regs(323)
                           );
   U1052 : AOI222_X1 port map( A1 => regs(323), A2 => n21, B1 => regs(1859), B2
                           => n73, C1 => regs(835), C2 => n125, ZN => n792);
   U1053 : AOI22_X1 port map( A1 => regs(1347), A2 => n177, B1 => regs(2371), 
                           B2 => n219, ZN => n791);
   U1054 : NAND2_X1 port map( A1 => n793, A2 => n794, ZN => curr_proc_regs(322)
                           );
   U1055 : AOI222_X1 port map( A1 => regs(322), A2 => n21, B1 => regs(1858), B2
                           => n73, C1 => regs(834), C2 => n125, ZN => n794);
   U1056 : AOI22_X1 port map( A1 => regs(1346), A2 => n177, B1 => regs(2370), 
                           B2 => n219, ZN => n793);
   U1057 : NAND2_X1 port map( A1 => n795, A2 => n796, ZN => curr_proc_regs(321)
                           );
   U1058 : AOI222_X1 port map( A1 => regs(321), A2 => n21, B1 => regs(1857), B2
                           => n73, C1 => regs(833), C2 => n125, ZN => n796);
   U1059 : AOI22_X1 port map( A1 => regs(1345), A2 => n177, B1 => regs(2369), 
                           B2 => n219, ZN => n795);
   U1060 : NAND2_X1 port map( A1 => n797, A2 => n798, ZN => curr_proc_regs(320)
                           );
   U1061 : AOI222_X1 port map( A1 => regs(320), A2 => n21, B1 => regs(1856), B2
                           => n73, C1 => regs(832), C2 => n125, ZN => n798);
   U1062 : AOI22_X1 port map( A1 => regs(1344), A2 => n177, B1 => regs(2368), 
                           B2 => n219, ZN => n797);
   U1063 : NAND2_X1 port map( A1 => n799, A2 => n800, ZN => curr_proc_regs(31))
                           ;
   U1064 : AOI222_X1 port map( A1 => regs(31), A2 => n21, B1 => regs(1567), B2 
                           => n73, C1 => regs(543), C2 => n125, ZN => n800);
   U1065 : AOI22_X1 port map( A1 => regs(1055), A2 => n177, B1 => regs(2079), 
                           B2 => n218, ZN => n799);
   U1066 : NAND2_X1 port map( A1 => n801, A2 => n802, ZN => curr_proc_regs(319)
                           );
   U1067 : AOI222_X1 port map( A1 => regs(319), A2 => n21, B1 => regs(1855), B2
                           => n73, C1 => regs(831), C2 => n125, ZN => n802);
   U1068 : AOI22_X1 port map( A1 => regs(1343), A2 => n177, B1 => regs(2367), 
                           B2 => n218, ZN => n801);
   U1069 : NAND2_X1 port map( A1 => n803, A2 => n804, ZN => curr_proc_regs(318)
                           );
   U1070 : AOI222_X1 port map( A1 => regs(318), A2 => n21, B1 => regs(1854), B2
                           => n73, C1 => regs(830), C2 => n125, ZN => n804);
   U1071 : AOI22_X1 port map( A1 => regs(1342), A2 => n177, B1 => regs(2366), 
                           B2 => n218, ZN => n803);
   U1072 : NAND2_X1 port map( A1 => n805, A2 => n806, ZN => curr_proc_regs(317)
                           );
   U1073 : AOI222_X1 port map( A1 => regs(317), A2 => n21, B1 => regs(1853), B2
                           => n73, C1 => regs(829), C2 => n125, ZN => n806);
   U1074 : AOI22_X1 port map( A1 => regs(1341), A2 => n177, B1 => regs(2365), 
                           B2 => n218, ZN => n805);
   U1075 : NAND2_X1 port map( A1 => n807, A2 => n808, ZN => curr_proc_regs(316)
                           );
   U1076 : AOI222_X1 port map( A1 => regs(316), A2 => n21, B1 => regs(1852), B2
                           => n73, C1 => regs(828), C2 => n125, ZN => n808);
   U1077 : AOI22_X1 port map( A1 => regs(1340), A2 => n177, B1 => regs(2364), 
                           B2 => n218, ZN => n807);
   U1078 : NAND2_X1 port map( A1 => n809, A2 => n810, ZN => curr_proc_regs(315)
                           );
   U1079 : AOI222_X1 port map( A1 => regs(315), A2 => n20, B1 => regs(1851), B2
                           => n72, C1 => regs(827), C2 => n124, ZN => n810);
   U1080 : AOI22_X1 port map( A1 => regs(1339), A2 => n176, B1 => regs(2363), 
                           B2 => n218, ZN => n809);
   U1081 : NAND2_X1 port map( A1 => n811, A2 => n812, ZN => curr_proc_regs(314)
                           );
   U1082 : AOI222_X1 port map( A1 => regs(314), A2 => n20, B1 => regs(1850), B2
                           => n72, C1 => regs(826), C2 => n124, ZN => n812);
   U1083 : AOI22_X1 port map( A1 => regs(1338), A2 => n176, B1 => regs(2362), 
                           B2 => n218, ZN => n811);
   U1084 : NAND2_X1 port map( A1 => n813, A2 => n814, ZN => curr_proc_regs(313)
                           );
   U1085 : AOI222_X1 port map( A1 => regs(313), A2 => n20, B1 => regs(1849), B2
                           => n72, C1 => regs(825), C2 => n124, ZN => n814);
   U1086 : AOI22_X1 port map( A1 => regs(1337), A2 => n176, B1 => regs(2361), 
                           B2 => n218, ZN => n813);
   U1087 : NAND2_X1 port map( A1 => n815, A2 => n816, ZN => curr_proc_regs(312)
                           );
   U1088 : AOI222_X1 port map( A1 => regs(312), A2 => n20, B1 => regs(1848), B2
                           => n72, C1 => regs(824), C2 => n124, ZN => n816);
   U1089 : AOI22_X1 port map( A1 => regs(1336), A2 => n176, B1 => regs(2360), 
                           B2 => n218, ZN => n815);
   U1090 : NAND2_X1 port map( A1 => n817, A2 => n818, ZN => curr_proc_regs(311)
                           );
   U1091 : AOI222_X1 port map( A1 => regs(311), A2 => n20, B1 => regs(1847), B2
                           => n72, C1 => regs(823), C2 => n124, ZN => n818);
   U1092 : AOI22_X1 port map( A1 => regs(1335), A2 => n176, B1 => regs(2359), 
                           B2 => n218, ZN => n817);
   U1093 : NAND2_X1 port map( A1 => n819, A2 => n820, ZN => curr_proc_regs(310)
                           );
   U1094 : AOI222_X1 port map( A1 => regs(310), A2 => n20, B1 => regs(1846), B2
                           => n72, C1 => regs(822), C2 => n124, ZN => n820);
   U1095 : AOI22_X1 port map( A1 => regs(1334), A2 => n176, B1 => regs(2358), 
                           B2 => n218, ZN => n819);
   U1096 : NAND2_X1 port map( A1 => n821, A2 => n822, ZN => curr_proc_regs(30))
                           ;
   U1097 : AOI222_X1 port map( A1 => regs(30), A2 => n20, B1 => regs(1566), B2 
                           => n72, C1 => regs(542), C2 => n124, ZN => n822);
   U1098 : AOI22_X1 port map( A1 => regs(1054), A2 => n176, B1 => regs(2078), 
                           B2 => n218, ZN => n821);
   U1099 : NAND2_X1 port map( A1 => n823, A2 => n824, ZN => curr_proc_regs(309)
                           );
   U1100 : AOI222_X1 port map( A1 => regs(309), A2 => n20, B1 => regs(1845), B2
                           => n72, C1 => regs(821), C2 => n124, ZN => n824);
   U1101 : AOI22_X1 port map( A1 => regs(1333), A2 => n176, B1 => regs(2357), 
                           B2 => n217, ZN => n823);
   U1102 : NAND2_X1 port map( A1 => n825, A2 => n826, ZN => curr_proc_regs(308)
                           );
   U1103 : AOI222_X1 port map( A1 => regs(308), A2 => n20, B1 => regs(1844), B2
                           => n72, C1 => regs(820), C2 => n124, ZN => n826);
   U1104 : AOI22_X1 port map( A1 => regs(1332), A2 => n176, B1 => regs(2356), 
                           B2 => n217, ZN => n825);
   U1105 : NAND2_X1 port map( A1 => n827, A2 => n828, ZN => curr_proc_regs(307)
                           );
   U1106 : AOI222_X1 port map( A1 => regs(307), A2 => n20, B1 => regs(1843), B2
                           => n72, C1 => regs(819), C2 => n124, ZN => n828);
   U1107 : AOI22_X1 port map( A1 => regs(1331), A2 => n176, B1 => regs(2355), 
                           B2 => n217, ZN => n827);
   U1108 : NAND2_X1 port map( A1 => n829, A2 => n830, ZN => curr_proc_regs(306)
                           );
   U1109 : AOI222_X1 port map( A1 => regs(306), A2 => n20, B1 => regs(1842), B2
                           => n72, C1 => regs(818), C2 => n124, ZN => n830);
   U1110 : AOI22_X1 port map( A1 => regs(1330), A2 => n176, B1 => regs(2354), 
                           B2 => n217, ZN => n829);
   U1111 : NAND2_X1 port map( A1 => n831, A2 => n832, ZN => curr_proc_regs(305)
                           );
   U1112 : AOI222_X1 port map( A1 => regs(305), A2 => n20, B1 => regs(1841), B2
                           => n72, C1 => regs(817), C2 => n124, ZN => n832);
   U1113 : AOI22_X1 port map( A1 => regs(1329), A2 => n176, B1 => regs(2353), 
                           B2 => n217, ZN => n831);
   U1114 : NAND2_X1 port map( A1 => n833, A2 => n834, ZN => curr_proc_regs(304)
                           );
   U1115 : AOI222_X1 port map( A1 => regs(304), A2 => n19, B1 => regs(1840), B2
                           => n71, C1 => regs(816), C2 => n123, ZN => n834);
   U1116 : AOI22_X1 port map( A1 => regs(1328), A2 => n175, B1 => regs(2352), 
                           B2 => n217, ZN => n833);
   U1117 : NAND2_X1 port map( A1 => n835, A2 => n836, ZN => curr_proc_regs(303)
                           );
   U1118 : AOI222_X1 port map( A1 => regs(303), A2 => n19, B1 => regs(1839), B2
                           => n71, C1 => regs(815), C2 => n123, ZN => n836);
   U1119 : AOI22_X1 port map( A1 => regs(1327), A2 => n175, B1 => regs(2351), 
                           B2 => n217, ZN => n835);
   U1120 : NAND2_X1 port map( A1 => n837, A2 => n838, ZN => curr_proc_regs(302)
                           );
   U1121 : AOI222_X1 port map( A1 => regs(302), A2 => n19, B1 => regs(1838), B2
                           => n71, C1 => regs(814), C2 => n123, ZN => n838);
   U1122 : AOI22_X1 port map( A1 => regs(1326), A2 => n175, B1 => regs(2350), 
                           B2 => n217, ZN => n837);
   U1123 : NAND2_X1 port map( A1 => n839, A2 => n840, ZN => curr_proc_regs(301)
                           );
   U1124 : AOI222_X1 port map( A1 => regs(301), A2 => n19, B1 => regs(1837), B2
                           => n71, C1 => regs(813), C2 => n123, ZN => n840);
   U1125 : AOI22_X1 port map( A1 => regs(1325), A2 => n175, B1 => regs(2349), 
                           B2 => n217, ZN => n839);
   U1126 : NAND2_X1 port map( A1 => n841, A2 => n842, ZN => curr_proc_regs(300)
                           );
   U1127 : AOI222_X1 port map( A1 => regs(300), A2 => n19, B1 => regs(1836), B2
                           => n71, C1 => regs(812), C2 => n123, ZN => n842);
   U1128 : AOI22_X1 port map( A1 => regs(1324), A2 => n175, B1 => regs(2348), 
                           B2 => n217, ZN => n841);
   U1129 : NAND2_X1 port map( A1 => n843, A2 => n844, ZN => curr_proc_regs(2));
   U1130 : AOI222_X1 port map( A1 => regs(2), A2 => n19, B1 => regs(1538), B2 
                           => n71, C1 => regs(514), C2 => n123, ZN => n844);
   U1131 : AOI22_X1 port map( A1 => regs(1026), A2 => n175, B1 => regs(2050), 
                           B2 => n217, ZN => n843);
   U1132 : NAND2_X1 port map( A1 => n845, A2 => n846, ZN => curr_proc_regs(29))
                           ;
   U1133 : AOI222_X1 port map( A1 => regs(29), A2 => n19, B1 => regs(1565), B2 
                           => n71, C1 => regs(541), C2 => n123, ZN => n846);
   U1134 : AOI22_X1 port map( A1 => regs(1053), A2 => n175, B1 => regs(2077), 
                           B2 => n217, ZN => n845);
   U1135 : NAND2_X1 port map( A1 => n847, A2 => n848, ZN => curr_proc_regs(299)
                           );
   U1136 : AOI222_X1 port map( A1 => regs(299), A2 => n19, B1 => regs(1835), B2
                           => n71, C1 => regs(811), C2 => n123, ZN => n848);
   U1137 : AOI22_X1 port map( A1 => regs(1323), A2 => n175, B1 => regs(2347), 
                           B2 => n216, ZN => n847);
   U1138 : NAND2_X1 port map( A1 => n849, A2 => n850, ZN => curr_proc_regs(298)
                           );
   U1139 : AOI222_X1 port map( A1 => regs(298), A2 => n19, B1 => regs(1834), B2
                           => n71, C1 => regs(810), C2 => n123, ZN => n850);
   U1140 : AOI22_X1 port map( A1 => regs(1322), A2 => n175, B1 => regs(2346), 
                           B2 => n216, ZN => n849);
   U1141 : NAND2_X1 port map( A1 => n851, A2 => n852, ZN => curr_proc_regs(297)
                           );
   U1142 : AOI222_X1 port map( A1 => regs(297), A2 => n19, B1 => regs(1833), B2
                           => n71, C1 => regs(809), C2 => n123, ZN => n852);
   U1143 : AOI22_X1 port map( A1 => regs(1321), A2 => n175, B1 => regs(2345), 
                           B2 => n216, ZN => n851);
   U1144 : NAND2_X1 port map( A1 => n853, A2 => n854, ZN => curr_proc_regs(296)
                           );
   U1145 : AOI222_X1 port map( A1 => regs(296), A2 => n19, B1 => regs(1832), B2
                           => n71, C1 => regs(808), C2 => n123, ZN => n854);
   U1146 : AOI22_X1 port map( A1 => regs(1320), A2 => n175, B1 => regs(2344), 
                           B2 => n216, ZN => n853);
   U1147 : NAND2_X1 port map( A1 => n855, A2 => n856, ZN => curr_proc_regs(295)
                           );
   U1148 : AOI222_X1 port map( A1 => regs(295), A2 => n19, B1 => regs(1831), B2
                           => n71, C1 => regs(807), C2 => n123, ZN => n856);
   U1149 : AOI22_X1 port map( A1 => regs(1319), A2 => n175, B1 => regs(2343), 
                           B2 => n216, ZN => n855);
   U1150 : NAND2_X1 port map( A1 => n857, A2 => n858, ZN => curr_proc_regs(294)
                           );
   U1151 : AOI222_X1 port map( A1 => regs(294), A2 => n18, B1 => regs(1830), B2
                           => n70, C1 => regs(806), C2 => n122, ZN => n858);
   U1152 : AOI22_X1 port map( A1 => regs(1318), A2 => n174, B1 => regs(2342), 
                           B2 => n216, ZN => n857);
   U1153 : NAND2_X1 port map( A1 => n859, A2 => n860, ZN => curr_proc_regs(293)
                           );
   U1154 : AOI222_X1 port map( A1 => regs(293), A2 => n18, B1 => regs(1829), B2
                           => n70, C1 => regs(805), C2 => n122, ZN => n860);
   U1155 : AOI22_X1 port map( A1 => regs(1317), A2 => n174, B1 => regs(2341), 
                           B2 => n216, ZN => n859);
   U1156 : NAND2_X1 port map( A1 => n861, A2 => n862, ZN => curr_proc_regs(292)
                           );
   U1157 : AOI222_X1 port map( A1 => regs(292), A2 => n18, B1 => regs(1828), B2
                           => n70, C1 => regs(804), C2 => n122, ZN => n862);
   U1158 : AOI22_X1 port map( A1 => regs(1316), A2 => n174, B1 => regs(2340), 
                           B2 => n216, ZN => n861);
   U1159 : NAND2_X1 port map( A1 => n863, A2 => n864, ZN => curr_proc_regs(291)
                           );
   U1160 : AOI222_X1 port map( A1 => regs(291), A2 => n18, B1 => regs(1827), B2
                           => n70, C1 => regs(803), C2 => n122, ZN => n864);
   U1161 : AOI22_X1 port map( A1 => regs(1315), A2 => n174, B1 => regs(2339), 
                           B2 => n216, ZN => n863);
   U1162 : NAND2_X1 port map( A1 => n865, A2 => n866, ZN => curr_proc_regs(290)
                           );
   U1163 : AOI222_X1 port map( A1 => regs(290), A2 => n18, B1 => regs(1826), B2
                           => n70, C1 => regs(802), C2 => n122, ZN => n866);
   U1164 : AOI22_X1 port map( A1 => regs(1314), A2 => n174, B1 => regs(2338), 
                           B2 => n216, ZN => n865);
   U1165 : NAND2_X1 port map( A1 => n867, A2 => n868, ZN => curr_proc_regs(28))
                           ;
   U1166 : AOI222_X1 port map( A1 => regs(28), A2 => n18, B1 => regs(1564), B2 
                           => n70, C1 => regs(540), C2 => n122, ZN => n868);
   U1167 : AOI22_X1 port map( A1 => regs(1052), A2 => n174, B1 => regs(2076), 
                           B2 => n216, ZN => n867);
   U1168 : NAND2_X1 port map( A1 => n869, A2 => n870, ZN => curr_proc_regs(289)
                           );
   U1169 : AOI222_X1 port map( A1 => regs(289), A2 => n18, B1 => regs(1825), B2
                           => n70, C1 => regs(801), C2 => n122, ZN => n870);
   U1170 : AOI22_X1 port map( A1 => regs(1313), A2 => n174, B1 => regs(2337), 
                           B2 => n216, ZN => n869);
   U1171 : NAND2_X1 port map( A1 => n871, A2 => n872, ZN => curr_proc_regs(288)
                           );
   U1172 : AOI222_X1 port map( A1 => regs(288), A2 => n18, B1 => regs(1824), B2
                           => n70, C1 => regs(800), C2 => n122, ZN => n872);
   U1173 : AOI22_X1 port map( A1 => regs(1312), A2 => n174, B1 => regs(2336), 
                           B2 => n215, ZN => n871);
   U1174 : NAND2_X1 port map( A1 => n873, A2 => n874, ZN => curr_proc_regs(287)
                           );
   U1175 : AOI222_X1 port map( A1 => regs(287), A2 => n18, B1 => regs(1823), B2
                           => n70, C1 => regs(799), C2 => n122, ZN => n874);
   U1176 : AOI22_X1 port map( A1 => regs(1311), A2 => n174, B1 => regs(2335), 
                           B2 => n215, ZN => n873);
   U1177 : NAND2_X1 port map( A1 => n875, A2 => n876, ZN => curr_proc_regs(286)
                           );
   U1178 : AOI222_X1 port map( A1 => regs(286), A2 => n18, B1 => regs(1822), B2
                           => n70, C1 => regs(798), C2 => n122, ZN => n876);
   U1179 : AOI22_X1 port map( A1 => regs(1310), A2 => n174, B1 => regs(2334), 
                           B2 => n215, ZN => n875);
   U1180 : NAND2_X1 port map( A1 => n877, A2 => n878, ZN => curr_proc_regs(285)
                           );
   U1181 : AOI222_X1 port map( A1 => regs(285), A2 => n18, B1 => regs(1821), B2
                           => n70, C1 => regs(797), C2 => n122, ZN => n878);
   U1182 : AOI22_X1 port map( A1 => regs(1309), A2 => n174, B1 => regs(2333), 
                           B2 => n215, ZN => n877);
   U1183 : NAND2_X1 port map( A1 => n879, A2 => n880, ZN => curr_proc_regs(284)
                           );
   U1184 : AOI222_X1 port map( A1 => regs(284), A2 => n18, B1 => regs(1820), B2
                           => n70, C1 => regs(796), C2 => n122, ZN => n880);
   U1185 : AOI22_X1 port map( A1 => regs(1308), A2 => n174, B1 => regs(2332), 
                           B2 => n215, ZN => n879);
   U1186 : NAND2_X1 port map( A1 => n881, A2 => n882, ZN => curr_proc_regs(283)
                           );
   U1187 : AOI222_X1 port map( A1 => regs(283), A2 => n17, B1 => regs(1819), B2
                           => n69, C1 => regs(795), C2 => n121, ZN => n882);
   U1188 : AOI22_X1 port map( A1 => regs(1307), A2 => n173, B1 => regs(2331), 
                           B2 => n215, ZN => n881);
   U1189 : NAND2_X1 port map( A1 => n883, A2 => n884, ZN => curr_proc_regs(282)
                           );
   U1190 : AOI222_X1 port map( A1 => regs(282), A2 => n17, B1 => regs(1818), B2
                           => n69, C1 => regs(794), C2 => n121, ZN => n884);
   U1191 : AOI22_X1 port map( A1 => regs(1306), A2 => n173, B1 => regs(2330), 
                           B2 => n215, ZN => n883);
   U1192 : NAND2_X1 port map( A1 => n885, A2 => n886, ZN => curr_proc_regs(281)
                           );
   U1193 : AOI222_X1 port map( A1 => regs(281), A2 => n17, B1 => regs(1817), B2
                           => n69, C1 => regs(793), C2 => n121, ZN => n886);
   U1194 : AOI22_X1 port map( A1 => regs(1305), A2 => n173, B1 => regs(2329), 
                           B2 => n215, ZN => n885);
   U1195 : NAND2_X1 port map( A1 => n887, A2 => n888, ZN => curr_proc_regs(280)
                           );
   U1196 : AOI222_X1 port map( A1 => regs(280), A2 => n17, B1 => regs(1816), B2
                           => n69, C1 => regs(792), C2 => n121, ZN => n888);
   U1197 : AOI22_X1 port map( A1 => regs(1304), A2 => n173, B1 => regs(2328), 
                           B2 => n215, ZN => n887);
   U1198 : NAND2_X1 port map( A1 => n889, A2 => n890, ZN => curr_proc_regs(27))
                           ;
   U1199 : AOI222_X1 port map( A1 => regs(27), A2 => n17, B1 => regs(1563), B2 
                           => n69, C1 => regs(539), C2 => n121, ZN => n890);
   U1200 : AOI22_X1 port map( A1 => regs(1051), A2 => n173, B1 => regs(2075), 
                           B2 => n215, ZN => n889);
   U1201 : NAND2_X1 port map( A1 => n891, A2 => n892, ZN => curr_proc_regs(279)
                           );
   U1202 : AOI222_X1 port map( A1 => regs(279), A2 => n17, B1 => regs(1815), B2
                           => n69, C1 => regs(791), C2 => n121, ZN => n892);
   U1203 : AOI22_X1 port map( A1 => regs(1303), A2 => n173, B1 => regs(2327), 
                           B2 => n215, ZN => n891);
   U1204 : NAND2_X1 port map( A1 => n893, A2 => n894, ZN => curr_proc_regs(278)
                           );
   U1205 : AOI222_X1 port map( A1 => regs(278), A2 => n17, B1 => regs(1814), B2
                           => n69, C1 => regs(790), C2 => n121, ZN => n894);
   U1206 : AOI22_X1 port map( A1 => regs(1302), A2 => n173, B1 => regs(2326), 
                           B2 => n215, ZN => n893);
   U1207 : NAND2_X1 port map( A1 => n895, A2 => n896, ZN => curr_proc_regs(277)
                           );
   U1208 : AOI222_X1 port map( A1 => regs(277), A2 => n17, B1 => regs(1813), B2
                           => n69, C1 => regs(789), C2 => n121, ZN => n896);
   U1209 : AOI22_X1 port map( A1 => regs(1301), A2 => n173, B1 => regs(2325), 
                           B2 => n214, ZN => n895);
   U1210 : NAND2_X1 port map( A1 => n897, A2 => n898, ZN => curr_proc_regs(276)
                           );
   U1211 : AOI222_X1 port map( A1 => regs(276), A2 => n17, B1 => regs(1812), B2
                           => n69, C1 => regs(788), C2 => n121, ZN => n898);
   U1212 : AOI22_X1 port map( A1 => regs(1300), A2 => n173, B1 => regs(2324), 
                           B2 => n214, ZN => n897);
   U1213 : NAND2_X1 port map( A1 => n899, A2 => n900, ZN => curr_proc_regs(275)
                           );
   U1214 : AOI222_X1 port map( A1 => regs(275), A2 => n17, B1 => regs(1811), B2
                           => n69, C1 => regs(787), C2 => n121, ZN => n900);
   U1215 : AOI22_X1 port map( A1 => regs(1299), A2 => n173, B1 => regs(2323), 
                           B2 => n214, ZN => n899);
   U1216 : NAND2_X1 port map( A1 => n901, A2 => n902, ZN => curr_proc_regs(274)
                           );
   U1217 : AOI222_X1 port map( A1 => regs(274), A2 => n17, B1 => regs(1810), B2
                           => n69, C1 => regs(786), C2 => n121, ZN => n902);
   U1218 : AOI22_X1 port map( A1 => regs(1298), A2 => n173, B1 => regs(2322), 
                           B2 => n214, ZN => n901);
   U1219 : NAND2_X1 port map( A1 => n903, A2 => n904, ZN => curr_proc_regs(273)
                           );
   U1220 : AOI222_X1 port map( A1 => regs(273), A2 => n17, B1 => regs(1809), B2
                           => n69, C1 => regs(785), C2 => n121, ZN => n904);
   U1221 : AOI22_X1 port map( A1 => regs(1297), A2 => n173, B1 => regs(2321), 
                           B2 => n214, ZN => n903);
   U1222 : NAND2_X1 port map( A1 => n905, A2 => n906, ZN => curr_proc_regs(272)
                           );
   U1223 : AOI222_X1 port map( A1 => regs(272), A2 => n16, B1 => regs(1808), B2
                           => n68, C1 => regs(784), C2 => n120, ZN => n906);
   U1224 : AOI22_X1 port map( A1 => regs(1296), A2 => n172, B1 => regs(2320), 
                           B2 => n214, ZN => n905);
   U1225 : NAND2_X1 port map( A1 => n907, A2 => n908, ZN => curr_proc_regs(271)
                           );
   U1226 : AOI222_X1 port map( A1 => regs(271), A2 => n16, B1 => regs(1807), B2
                           => n68, C1 => regs(783), C2 => n120, ZN => n908);
   U1227 : AOI22_X1 port map( A1 => regs(1295), A2 => n172, B1 => regs(2319), 
                           B2 => n214, ZN => n907);
   U1228 : NAND2_X1 port map( A1 => n909, A2 => n910, ZN => curr_proc_regs(270)
                           );
   U1229 : AOI222_X1 port map( A1 => regs(270), A2 => n16, B1 => regs(1806), B2
                           => n68, C1 => regs(782), C2 => n120, ZN => n910);
   U1230 : AOI22_X1 port map( A1 => regs(1294), A2 => n172, B1 => regs(2318), 
                           B2 => n214, ZN => n909);
   U1231 : NAND2_X1 port map( A1 => n911, A2 => n912, ZN => curr_proc_regs(26))
                           ;
   U1232 : AOI222_X1 port map( A1 => regs(26), A2 => n16, B1 => regs(1562), B2 
                           => n68, C1 => regs(538), C2 => n120, ZN => n912);
   U1233 : AOI22_X1 port map( A1 => regs(1050), A2 => n172, B1 => regs(2074), 
                           B2 => n214, ZN => n911);
   U1234 : NAND2_X1 port map( A1 => n913, A2 => n914, ZN => curr_proc_regs(269)
                           );
   U1235 : AOI222_X1 port map( A1 => regs(269), A2 => n16, B1 => regs(1805), B2
                           => n68, C1 => regs(781), C2 => n120, ZN => n914);
   U1236 : AOI22_X1 port map( A1 => regs(1293), A2 => n172, B1 => regs(2317), 
                           B2 => n214, ZN => n913);
   U1237 : NAND2_X1 port map( A1 => n915, A2 => n916, ZN => curr_proc_regs(268)
                           );
   U1238 : AOI222_X1 port map( A1 => regs(268), A2 => n16, B1 => regs(1804), B2
                           => n68, C1 => regs(780), C2 => n120, ZN => n916);
   U1239 : AOI22_X1 port map( A1 => regs(1292), A2 => n172, B1 => regs(2316), 
                           B2 => n214, ZN => n915);
   U1240 : NAND2_X1 port map( A1 => n917, A2 => n918, ZN => curr_proc_regs(267)
                           );
   U1241 : AOI222_X1 port map( A1 => regs(267), A2 => n16, B1 => regs(1803), B2
                           => n68, C1 => regs(779), C2 => n120, ZN => n918);
   U1242 : AOI22_X1 port map( A1 => regs(1291), A2 => n172, B1 => regs(2315), 
                           B2 => n213, ZN => n917);
   U1243 : NAND2_X1 port map( A1 => n919, A2 => n920, ZN => curr_proc_regs(266)
                           );
   U1244 : AOI222_X1 port map( A1 => regs(266), A2 => n16, B1 => regs(1802), B2
                           => n68, C1 => regs(778), C2 => n120, ZN => n920);
   U1245 : AOI22_X1 port map( A1 => regs(1290), A2 => n172, B1 => regs(2314), 
                           B2 => n213, ZN => n919);
   U1246 : NAND2_X1 port map( A1 => n921, A2 => n922, ZN => curr_proc_regs(265)
                           );
   U1247 : AOI222_X1 port map( A1 => regs(265), A2 => n16, B1 => regs(1801), B2
                           => n68, C1 => regs(777), C2 => n120, ZN => n922);
   U1248 : AOI22_X1 port map( A1 => regs(1289), A2 => n172, B1 => regs(2313), 
                           B2 => n213, ZN => n921);
   U1249 : NAND2_X1 port map( A1 => n923, A2 => n924, ZN => curr_proc_regs(264)
                           );
   U1250 : AOI222_X1 port map( A1 => regs(264), A2 => n16, B1 => regs(1800), B2
                           => n68, C1 => regs(776), C2 => n120, ZN => n924);
   U1251 : AOI22_X1 port map( A1 => regs(1288), A2 => n172, B1 => regs(2312), 
                           B2 => n213, ZN => n923);
   U1252 : NAND2_X1 port map( A1 => n925, A2 => n926, ZN => curr_proc_regs(263)
                           );
   U1253 : AOI222_X1 port map( A1 => regs(263), A2 => n16, B1 => regs(1799), B2
                           => n68, C1 => regs(775), C2 => n120, ZN => n926);
   U1254 : AOI22_X1 port map( A1 => regs(1287), A2 => n172, B1 => regs(2311), 
                           B2 => n213, ZN => n925);
   U1255 : NAND2_X1 port map( A1 => n927, A2 => n928, ZN => curr_proc_regs(262)
                           );
   U1256 : AOI222_X1 port map( A1 => regs(262), A2 => n16, B1 => regs(1798), B2
                           => n68, C1 => regs(774), C2 => n120, ZN => n928);
   U1257 : AOI22_X1 port map( A1 => regs(1286), A2 => n172, B1 => regs(2310), 
                           B2 => n213, ZN => n927);
   U1258 : NAND2_X1 port map( A1 => n929, A2 => n930, ZN => curr_proc_regs(261)
                           );
   U1259 : AOI222_X1 port map( A1 => regs(261), A2 => n15, B1 => regs(1797), B2
                           => n67, C1 => regs(773), C2 => n119, ZN => n930);
   U1260 : AOI22_X1 port map( A1 => regs(1285), A2 => n171, B1 => regs(2309), 
                           B2 => n213, ZN => n929);
   U1261 : NAND2_X1 port map( A1 => n931, A2 => n932, ZN => curr_proc_regs(260)
                           );
   U1262 : AOI222_X1 port map( A1 => regs(260), A2 => n15, B1 => regs(1796), B2
                           => n67, C1 => regs(772), C2 => n119, ZN => n932);
   U1263 : AOI22_X1 port map( A1 => regs(1284), A2 => n171, B1 => regs(2308), 
                           B2 => n213, ZN => n931);
   U1264 : NAND2_X1 port map( A1 => n933, A2 => n934, ZN => curr_proc_regs(25))
                           ;
   U1265 : AOI222_X1 port map( A1 => regs(25), A2 => n15, B1 => regs(1561), B2 
                           => n67, C1 => regs(537), C2 => n119, ZN => n934);
   U1266 : AOI22_X1 port map( A1 => regs(1049), A2 => n171, B1 => regs(2073), 
                           B2 => n213, ZN => n933);
   U1267 : NAND2_X1 port map( A1 => n935, A2 => n936, ZN => curr_proc_regs(259)
                           );
   U1268 : AOI222_X1 port map( A1 => regs(259), A2 => n15, B1 => regs(1795), B2
                           => n67, C1 => regs(771), C2 => n119, ZN => n936);
   U1269 : AOI22_X1 port map( A1 => regs(1283), A2 => n171, B1 => regs(2307), 
                           B2 => n213, ZN => n935);
   U1270 : NAND2_X1 port map( A1 => n937, A2 => n938, ZN => curr_proc_regs(258)
                           );
   U1271 : AOI222_X1 port map( A1 => regs(258), A2 => n15, B1 => regs(1794), B2
                           => n67, C1 => regs(770), C2 => n119, ZN => n938);
   U1272 : AOI22_X1 port map( A1 => regs(1282), A2 => n171, B1 => regs(2306), 
                           B2 => n213, ZN => n937);
   U1273 : NAND2_X1 port map( A1 => n939, A2 => n940, ZN => curr_proc_regs(257)
                           );
   U1274 : AOI222_X1 port map( A1 => regs(257), A2 => n15, B1 => regs(1793), B2
                           => n67, C1 => regs(769), C2 => n119, ZN => n940);
   U1275 : AOI22_X1 port map( A1 => regs(1281), A2 => n171, B1 => regs(2305), 
                           B2 => n213, ZN => n939);
   U1276 : NAND2_X1 port map( A1 => n941, A2 => n942, ZN => curr_proc_regs(256)
                           );
   U1277 : AOI222_X1 port map( A1 => regs(256), A2 => n15, B1 => regs(1792), B2
                           => n67, C1 => regs(768), C2 => n119, ZN => n942);
   U1278 : AOI22_X1 port map( A1 => regs(1280), A2 => n171, B1 => regs(2304), 
                           B2 => n212, ZN => n941);
   U1279 : NAND2_X1 port map( A1 => n943, A2 => n944, ZN => curr_proc_regs(255)
                           );
   U1280 : AOI222_X1 port map( A1 => regs(255), A2 => n15, B1 => regs(1791), B2
                           => n67, C1 => regs(767), C2 => n119, ZN => n944);
   U1281 : AOI22_X1 port map( A1 => regs(1279), A2 => n171, B1 => regs(2303), 
                           B2 => n212, ZN => n943);
   U1282 : NAND2_X1 port map( A1 => n945, A2 => n946, ZN => curr_proc_regs(254)
                           );
   U1283 : AOI222_X1 port map( A1 => regs(254), A2 => n15, B1 => regs(1790), B2
                           => n67, C1 => regs(766), C2 => n119, ZN => n946);
   U1284 : AOI22_X1 port map( A1 => regs(1278), A2 => n171, B1 => regs(2302), 
                           B2 => n212, ZN => n945);
   U1285 : NAND2_X1 port map( A1 => n947, A2 => n948, ZN => curr_proc_regs(253)
                           );
   U1286 : AOI222_X1 port map( A1 => regs(253), A2 => n15, B1 => regs(1789), B2
                           => n67, C1 => regs(765), C2 => n119, ZN => n948);
   U1287 : AOI22_X1 port map( A1 => regs(1277), A2 => n171, B1 => regs(2301), 
                           B2 => n212, ZN => n947);
   U1288 : NAND2_X1 port map( A1 => n949, A2 => n950, ZN => curr_proc_regs(252)
                           );
   U1289 : AOI222_X1 port map( A1 => regs(252), A2 => n15, B1 => regs(1788), B2
                           => n67, C1 => regs(764), C2 => n119, ZN => n950);
   U1290 : AOI22_X1 port map( A1 => regs(1276), A2 => n171, B1 => regs(2300), 
                           B2 => n212, ZN => n949);
   U1291 : NAND2_X1 port map( A1 => n951, A2 => n952, ZN => curr_proc_regs(251)
                           );
   U1292 : AOI222_X1 port map( A1 => regs(251), A2 => n15, B1 => regs(1787), B2
                           => n67, C1 => regs(763), C2 => n119, ZN => n952);
   U1293 : AOI22_X1 port map( A1 => regs(1275), A2 => n171, B1 => regs(2299), 
                           B2 => n212, ZN => n951);
   U1294 : NAND2_X1 port map( A1 => n953, A2 => n954, ZN => curr_proc_regs(250)
                           );
   U1295 : AOI222_X1 port map( A1 => regs(250), A2 => n14, B1 => regs(1786), B2
                           => n66, C1 => regs(762), C2 => n118, ZN => n954);
   U1296 : AOI22_X1 port map( A1 => regs(1274), A2 => n170, B1 => regs(2298), 
                           B2 => n212, ZN => n953);
   U1297 : NAND2_X1 port map( A1 => n955, A2 => n956, ZN => curr_proc_regs(24))
                           ;
   U1298 : AOI222_X1 port map( A1 => regs(24), A2 => n14, B1 => regs(1560), B2 
                           => n66, C1 => regs(536), C2 => n118, ZN => n956);
   U1299 : AOI22_X1 port map( A1 => regs(1048), A2 => n170, B1 => regs(2072), 
                           B2 => n212, ZN => n955);
   U1300 : NAND2_X1 port map( A1 => n957, A2 => n958, ZN => curr_proc_regs(249)
                           );
   U1301 : AOI222_X1 port map( A1 => regs(249), A2 => n14, B1 => regs(1785), B2
                           => n66, C1 => regs(761), C2 => n118, ZN => n958);
   U1302 : AOI22_X1 port map( A1 => regs(1273), A2 => n170, B1 => regs(2297), 
                           B2 => n212, ZN => n957);
   U1303 : NAND2_X1 port map( A1 => n959, A2 => n960, ZN => curr_proc_regs(248)
                           );
   U1304 : AOI222_X1 port map( A1 => regs(248), A2 => n14, B1 => regs(1784), B2
                           => n66, C1 => regs(760), C2 => n118, ZN => n960);
   U1305 : AOI22_X1 port map( A1 => regs(1272), A2 => n170, B1 => regs(2296), 
                           B2 => n212, ZN => n959);
   U1306 : NAND2_X1 port map( A1 => n961, A2 => n962, ZN => curr_proc_regs(247)
                           );
   U1307 : AOI222_X1 port map( A1 => regs(247), A2 => n14, B1 => regs(1783), B2
                           => n66, C1 => regs(759), C2 => n118, ZN => n962);
   U1308 : AOI22_X1 port map( A1 => regs(1271), A2 => n170, B1 => regs(2295), 
                           B2 => n212, ZN => n961);
   U1309 : NAND2_X1 port map( A1 => n963, A2 => n964, ZN => curr_proc_regs(246)
                           );
   U1310 : AOI222_X1 port map( A1 => regs(246), A2 => n14, B1 => regs(1782), B2
                           => n66, C1 => regs(758), C2 => n118, ZN => n964);
   U1311 : AOI22_X1 port map( A1 => regs(1270), A2 => n170, B1 => regs(2294), 
                           B2 => n212, ZN => n963);
   U1312 : NAND2_X1 port map( A1 => n965, A2 => n966, ZN => curr_proc_regs(245)
                           );
   U1313 : AOI222_X1 port map( A1 => regs(245), A2 => n14, B1 => regs(1781), B2
                           => n66, C1 => regs(757), C2 => n118, ZN => n966);
   U1314 : AOI22_X1 port map( A1 => regs(1269), A2 => n170, B1 => regs(2293), 
                           B2 => n211, ZN => n965);
   U1315 : NAND2_X1 port map( A1 => n967, A2 => n968, ZN => curr_proc_regs(244)
                           );
   U1316 : AOI222_X1 port map( A1 => regs(244), A2 => n14, B1 => regs(1780), B2
                           => n66, C1 => regs(756), C2 => n118, ZN => n968);
   U1317 : AOI22_X1 port map( A1 => regs(1268), A2 => n170, B1 => regs(2292), 
                           B2 => n211, ZN => n967);
   U1318 : NAND2_X1 port map( A1 => n969, A2 => n970, ZN => curr_proc_regs(243)
                           );
   U1319 : AOI222_X1 port map( A1 => regs(243), A2 => n14, B1 => regs(1779), B2
                           => n66, C1 => regs(755), C2 => n118, ZN => n970);
   U1320 : AOI22_X1 port map( A1 => regs(1267), A2 => n170, B1 => regs(2291), 
                           B2 => n211, ZN => n969);
   U1321 : NAND2_X1 port map( A1 => n971, A2 => n972, ZN => curr_proc_regs(242)
                           );
   U1322 : AOI222_X1 port map( A1 => regs(242), A2 => n14, B1 => regs(1778), B2
                           => n66, C1 => regs(754), C2 => n118, ZN => n972);
   U1323 : AOI22_X1 port map( A1 => regs(1266), A2 => n170, B1 => regs(2290), 
                           B2 => n211, ZN => n971);
   U1324 : NAND2_X1 port map( A1 => n973, A2 => n974, ZN => curr_proc_regs(241)
                           );
   U1325 : AOI222_X1 port map( A1 => regs(241), A2 => n14, B1 => regs(1777), B2
                           => n66, C1 => regs(753), C2 => n118, ZN => n974);
   U1326 : AOI22_X1 port map( A1 => regs(1265), A2 => n170, B1 => regs(2289), 
                           B2 => n211, ZN => n973);
   U1327 : NAND2_X1 port map( A1 => n975, A2 => n976, ZN => curr_proc_regs(240)
                           );
   U1328 : AOI222_X1 port map( A1 => regs(240), A2 => n14, B1 => regs(1776), B2
                           => n66, C1 => regs(752), C2 => n118, ZN => n976);
   U1329 : AOI22_X1 port map( A1 => regs(1264), A2 => n170, B1 => regs(2288), 
                           B2 => n211, ZN => n975);
   U1330 : NAND2_X1 port map( A1 => n977, A2 => n978, ZN => curr_proc_regs(23))
                           ;
   U1331 : AOI222_X1 port map( A1 => regs(23), A2 => n13, B1 => regs(1559), B2 
                           => n65, C1 => regs(535), C2 => n117, ZN => n978);
   U1332 : AOI22_X1 port map( A1 => regs(1047), A2 => n169, B1 => regs(2071), 
                           B2 => n211, ZN => n977);
   U1333 : NAND2_X1 port map( A1 => n979, A2 => n980, ZN => curr_proc_regs(239)
                           );
   U1334 : AOI222_X1 port map( A1 => regs(239), A2 => n13, B1 => regs(1775), B2
                           => n65, C1 => regs(751), C2 => n117, ZN => n980);
   U1335 : AOI22_X1 port map( A1 => regs(1263), A2 => n169, B1 => regs(2287), 
                           B2 => n211, ZN => n979);
   U1336 : NAND2_X1 port map( A1 => n981, A2 => n982, ZN => curr_proc_regs(238)
                           );
   U1337 : AOI222_X1 port map( A1 => regs(238), A2 => n13, B1 => regs(1774), B2
                           => n65, C1 => regs(750), C2 => n117, ZN => n982);
   U1338 : AOI22_X1 port map( A1 => regs(1262), A2 => n169, B1 => regs(2286), 
                           B2 => n211, ZN => n981);
   U1339 : NAND2_X1 port map( A1 => n983, A2 => n984, ZN => curr_proc_regs(237)
                           );
   U1340 : AOI222_X1 port map( A1 => regs(237), A2 => n13, B1 => regs(1773), B2
                           => n65, C1 => regs(749), C2 => n117, ZN => n984);
   U1341 : AOI22_X1 port map( A1 => regs(1261), A2 => n169, B1 => regs(2285), 
                           B2 => n211, ZN => n983);
   U1342 : NAND2_X1 port map( A1 => n985, A2 => n986, ZN => curr_proc_regs(236)
                           );
   U1343 : AOI222_X1 port map( A1 => regs(236), A2 => n13, B1 => regs(1772), B2
                           => n65, C1 => regs(748), C2 => n117, ZN => n986);
   U1344 : AOI22_X1 port map( A1 => regs(1260), A2 => n169, B1 => regs(2284), 
                           B2 => n211, ZN => n985);
   U1345 : NAND2_X1 port map( A1 => n987, A2 => n988, ZN => curr_proc_regs(235)
                           );
   U1346 : AOI222_X1 port map( A1 => regs(235), A2 => n13, B1 => regs(1771), B2
                           => n65, C1 => regs(747), C2 => n117, ZN => n988);
   U1347 : AOI22_X1 port map( A1 => regs(1259), A2 => n169, B1 => regs(2283), 
                           B2 => n211, ZN => n987);
   U1348 : NAND2_X1 port map( A1 => n989, A2 => n990, ZN => curr_proc_regs(234)
                           );
   U1349 : AOI222_X1 port map( A1 => regs(234), A2 => n13, B1 => regs(1770), B2
                           => n65, C1 => regs(746), C2 => n117, ZN => n990);
   U1350 : AOI22_X1 port map( A1 => regs(1258), A2 => n169, B1 => regs(2282), 
                           B2 => n210, ZN => n989);
   U1351 : NAND2_X1 port map( A1 => n991, A2 => n992, ZN => curr_proc_regs(233)
                           );
   U1352 : AOI222_X1 port map( A1 => regs(233), A2 => n13, B1 => regs(1769), B2
                           => n65, C1 => regs(745), C2 => n117, ZN => n992);
   U1353 : AOI22_X1 port map( A1 => regs(1257), A2 => n169, B1 => regs(2281), 
                           B2 => n210, ZN => n991);
   U1354 : NAND2_X1 port map( A1 => n993, A2 => n994, ZN => curr_proc_regs(232)
                           );
   U1355 : AOI222_X1 port map( A1 => regs(232), A2 => n13, B1 => regs(1768), B2
                           => n65, C1 => regs(744), C2 => n117, ZN => n994);
   U1356 : AOI22_X1 port map( A1 => regs(1256), A2 => n169, B1 => regs(2280), 
                           B2 => n210, ZN => n993);
   U1357 : NAND2_X1 port map( A1 => n995, A2 => n996, ZN => curr_proc_regs(231)
                           );
   U1358 : AOI222_X1 port map( A1 => regs(231), A2 => n13, B1 => regs(1767), B2
                           => n65, C1 => regs(743), C2 => n117, ZN => n996);
   U1359 : AOI22_X1 port map( A1 => regs(1255), A2 => n169, B1 => regs(2279), 
                           B2 => n210, ZN => n995);
   U1360 : NAND2_X1 port map( A1 => n997, A2 => n998, ZN => curr_proc_regs(230)
                           );
   U1361 : AOI222_X1 port map( A1 => regs(230), A2 => n13, B1 => regs(1766), B2
                           => n65, C1 => regs(742), C2 => n117, ZN => n998);
   U1362 : AOI22_X1 port map( A1 => regs(1254), A2 => n169, B1 => regs(2278), 
                           B2 => n210, ZN => n997);
   U1363 : NAND2_X1 port map( A1 => n999, A2 => n1000, ZN => curr_proc_regs(22)
                           );
   U1364 : AOI222_X1 port map( A1 => regs(22), A2 => n13, B1 => regs(1558), B2 
                           => n65, C1 => regs(534), C2 => n117, ZN => n1000);
   U1365 : AOI22_X1 port map( A1 => regs(1046), A2 => n169, B1 => regs(2070), 
                           B2 => n210, ZN => n999);
   U1366 : NAND2_X1 port map( A1 => n1001, A2 => n1002, ZN => 
                           curr_proc_regs(229));
   U1367 : AOI222_X1 port map( A1 => regs(229), A2 => n12, B1 => regs(1765), B2
                           => n64, C1 => regs(741), C2 => n116, ZN => n1002);
   U1368 : AOI22_X1 port map( A1 => regs(1253), A2 => n168, B1 => regs(2277), 
                           B2 => n210, ZN => n1001);
   U1369 : NAND2_X1 port map( A1 => n1003, A2 => n1004, ZN => 
                           curr_proc_regs(228));
   U1370 : AOI222_X1 port map( A1 => regs(228), A2 => n12, B1 => regs(1764), B2
                           => n64, C1 => regs(740), C2 => n116, ZN => n1004);
   U1371 : AOI22_X1 port map( A1 => regs(1252), A2 => n168, B1 => regs(2276), 
                           B2 => n210, ZN => n1003);
   U1372 : NAND2_X1 port map( A1 => n1005, A2 => n1006, ZN => 
                           curr_proc_regs(227));
   U1373 : AOI222_X1 port map( A1 => regs(227), A2 => n12, B1 => regs(1763), B2
                           => n64, C1 => regs(739), C2 => n116, ZN => n1006);
   U1374 : AOI22_X1 port map( A1 => regs(1251), A2 => n168, B1 => regs(2275), 
                           B2 => n210, ZN => n1005);
   U1375 : NAND2_X1 port map( A1 => n1007, A2 => n1008, ZN => 
                           curr_proc_regs(226));
   U1376 : AOI222_X1 port map( A1 => regs(226), A2 => n12, B1 => regs(1762), B2
                           => n64, C1 => regs(738), C2 => n116, ZN => n1008);
   U1377 : AOI22_X1 port map( A1 => regs(1250), A2 => n168, B1 => regs(2274), 
                           B2 => n210, ZN => n1007);
   U1378 : NAND2_X1 port map( A1 => n1009, A2 => n1010, ZN => 
                           curr_proc_regs(225));
   U1379 : AOI222_X1 port map( A1 => regs(225), A2 => n12, B1 => regs(1761), B2
                           => n64, C1 => regs(737), C2 => n116, ZN => n1010);
   U1380 : AOI22_X1 port map( A1 => regs(1249), A2 => n168, B1 => regs(2273), 
                           B2 => n210, ZN => n1009);
   U1381 : NAND2_X1 port map( A1 => n1011, A2 => n1012, ZN => 
                           curr_proc_regs(224));
   U1382 : AOI222_X1 port map( A1 => regs(224), A2 => n12, B1 => regs(1760), B2
                           => n64, C1 => regs(736), C2 => n116, ZN => n1012);
   U1383 : AOI22_X1 port map( A1 => regs(1248), A2 => n168, B1 => regs(2272), 
                           B2 => n210, ZN => n1011);
   U1384 : NAND2_X1 port map( A1 => n1013, A2 => n1014, ZN => 
                           curr_proc_regs(223));
   U1385 : AOI222_X1 port map( A1 => regs(223), A2 => n12, B1 => regs(1759), B2
                           => n64, C1 => regs(735), C2 => n116, ZN => n1014);
   U1386 : AOI22_X1 port map( A1 => regs(1247), A2 => n168, B1 => regs(2271), 
                           B2 => n209, ZN => n1013);
   U1387 : NAND2_X1 port map( A1 => n1015, A2 => n1016, ZN => 
                           curr_proc_regs(222));
   U1388 : AOI222_X1 port map( A1 => regs(222), A2 => n12, B1 => regs(1758), B2
                           => n64, C1 => regs(734), C2 => n116, ZN => n1016);
   U1389 : AOI22_X1 port map( A1 => regs(1246), A2 => n168, B1 => regs(2270), 
                           B2 => n209, ZN => n1015);
   U1390 : NAND2_X1 port map( A1 => n1017, A2 => n1018, ZN => 
                           curr_proc_regs(221));
   U1391 : AOI222_X1 port map( A1 => regs(221), A2 => n12, B1 => regs(1757), B2
                           => n64, C1 => regs(733), C2 => n116, ZN => n1018);
   U1392 : AOI22_X1 port map( A1 => regs(1245), A2 => n168, B1 => regs(2269), 
                           B2 => n209, ZN => n1017);
   U1393 : NAND2_X1 port map( A1 => n1019, A2 => n1020, ZN => 
                           curr_proc_regs(220));
   U1394 : AOI222_X1 port map( A1 => regs(220), A2 => n12, B1 => regs(1756), B2
                           => n64, C1 => regs(732), C2 => n116, ZN => n1020);
   U1395 : AOI22_X1 port map( A1 => regs(1244), A2 => n168, B1 => regs(2268), 
                           B2 => n209, ZN => n1019);
   U1396 : NAND2_X1 port map( A1 => n1021, A2 => n1022, ZN => 
                           curr_proc_regs(21));
   U1397 : AOI222_X1 port map( A1 => regs(21), A2 => n12, B1 => regs(1557), B2 
                           => n64, C1 => regs(533), C2 => n116, ZN => n1022);
   U1398 : AOI22_X1 port map( A1 => regs(1045), A2 => n168, B1 => regs(2069), 
                           B2 => n209, ZN => n1021);
   U1399 : NAND2_X1 port map( A1 => n1023, A2 => n1024, ZN => 
                           curr_proc_regs(219));
   U1400 : AOI222_X1 port map( A1 => regs(219), A2 => n12, B1 => regs(1755), B2
                           => n64, C1 => regs(731), C2 => n116, ZN => n1024);
   U1401 : AOI22_X1 port map( A1 => regs(1243), A2 => n168, B1 => regs(2267), 
                           B2 => n209, ZN => n1023);
   U1402 : NAND2_X1 port map( A1 => n1025, A2 => n1026, ZN => 
                           curr_proc_regs(218));
   U1403 : AOI222_X1 port map( A1 => regs(218), A2 => n11, B1 => regs(1754), B2
                           => n63, C1 => regs(730), C2 => n115, ZN => n1026);
   U1404 : AOI22_X1 port map( A1 => regs(1242), A2 => n167, B1 => regs(2266), 
                           B2 => n209, ZN => n1025);
   U1405 : NAND2_X1 port map( A1 => n1027, A2 => n1028, ZN => 
                           curr_proc_regs(217));
   U1406 : AOI222_X1 port map( A1 => regs(217), A2 => n11, B1 => regs(1753), B2
                           => n63, C1 => regs(729), C2 => n115, ZN => n1028);
   U1407 : AOI22_X1 port map( A1 => regs(1241), A2 => n167, B1 => regs(2265), 
                           B2 => n209, ZN => n1027);
   U1408 : NAND2_X1 port map( A1 => n1029, A2 => n1030, ZN => 
                           curr_proc_regs(216));
   U1409 : AOI222_X1 port map( A1 => regs(216), A2 => n11, B1 => regs(1752), B2
                           => n63, C1 => regs(728), C2 => n115, ZN => n1030);
   U1410 : AOI22_X1 port map( A1 => regs(1240), A2 => n167, B1 => regs(2264), 
                           B2 => n209, ZN => n1029);
   U1411 : NAND2_X1 port map( A1 => n1031, A2 => n1032, ZN => 
                           curr_proc_regs(215));
   U1412 : AOI222_X1 port map( A1 => regs(215), A2 => n11, B1 => regs(1751), B2
                           => n63, C1 => regs(727), C2 => n115, ZN => n1032);
   U1413 : AOI22_X1 port map( A1 => regs(1239), A2 => n167, B1 => regs(2263), 
                           B2 => n214, ZN => n1031);
   U1414 : NAND2_X1 port map( A1 => n1033, A2 => n1034, ZN => 
                           curr_proc_regs(214));
   U1415 : AOI222_X1 port map( A1 => regs(214), A2 => n11, B1 => regs(1750), B2
                           => n63, C1 => regs(726), C2 => n115, ZN => n1034);
   U1416 : AOI22_X1 port map( A1 => regs(1238), A2 => n167, B1 => regs(2262), 
                           B2 => n230, ZN => n1033);
   U1417 : NAND2_X1 port map( A1 => n1035, A2 => n1036, ZN => 
                           curr_proc_regs(213));
   U1418 : AOI222_X1 port map( A1 => regs(213), A2 => n11, B1 => regs(1749), B2
                           => n63, C1 => regs(725), C2 => n115, ZN => n1036);
   U1419 : AOI22_X1 port map( A1 => regs(1237), A2 => n167, B1 => regs(2261), 
                           B2 => n230, ZN => n1035);
   U1420 : NAND2_X1 port map( A1 => n1037, A2 => n1038, ZN => 
                           curr_proc_regs(212));
   U1421 : AOI222_X1 port map( A1 => regs(212), A2 => n11, B1 => regs(1748), B2
                           => n63, C1 => regs(724), C2 => n115, ZN => n1038);
   U1422 : AOI22_X1 port map( A1 => regs(1236), A2 => n167, B1 => regs(2260), 
                           B2 => n230, ZN => n1037);
   U1423 : NAND2_X1 port map( A1 => n1039, A2 => n1040, ZN => 
                           curr_proc_regs(211));
   U1424 : AOI222_X1 port map( A1 => regs(211), A2 => n11, B1 => regs(1747), B2
                           => n63, C1 => regs(723), C2 => n115, ZN => n1040);
   U1425 : AOI22_X1 port map( A1 => regs(1235), A2 => n167, B1 => regs(2259), 
                           B2 => n230, ZN => n1039);
   U1426 : NAND2_X1 port map( A1 => n1041, A2 => n1042, ZN => 
                           curr_proc_regs(210));
   U1427 : AOI222_X1 port map( A1 => regs(210), A2 => n11, B1 => regs(1746), B2
                           => n63, C1 => regs(722), C2 => n115, ZN => n1042);
   U1428 : AOI22_X1 port map( A1 => regs(1234), A2 => n167, B1 => regs(2258), 
                           B2 => n230, ZN => n1041);
   U1429 : NAND2_X1 port map( A1 => n1043, A2 => n1044, ZN => 
                           curr_proc_regs(20));
   U1430 : AOI222_X1 port map( A1 => regs(20), A2 => n11, B1 => regs(1556), B2 
                           => n63, C1 => regs(532), C2 => n115, ZN => n1044);
   U1431 : AOI22_X1 port map( A1 => regs(1044), A2 => n167, B1 => regs(2068), 
                           B2 => n229, ZN => n1043);
   U1432 : NAND2_X1 port map( A1 => n1045, A2 => n1046, ZN => 
                           curr_proc_regs(209));
   U1433 : AOI222_X1 port map( A1 => regs(209), A2 => n11, B1 => regs(1745), B2
                           => n63, C1 => regs(721), C2 => n115, ZN => n1046);
   U1434 : AOI22_X1 port map( A1 => regs(1233), A2 => n167, B1 => regs(2257), 
                           B2 => n229, ZN => n1045);
   U1435 : NAND2_X1 port map( A1 => n1047, A2 => n1048, ZN => 
                           curr_proc_regs(208));
   U1436 : AOI222_X1 port map( A1 => regs(208), A2 => n11, B1 => regs(1744), B2
                           => n63, C1 => regs(720), C2 => n115, ZN => n1048);
   U1437 : AOI22_X1 port map( A1 => regs(1232), A2 => n167, B1 => regs(2256), 
                           B2 => n229, ZN => n1047);
   U1438 : NAND2_X1 port map( A1 => n1049, A2 => n1050, ZN => 
                           curr_proc_regs(207));
   U1439 : AOI222_X1 port map( A1 => regs(207), A2 => n10, B1 => regs(1743), B2
                           => n62, C1 => regs(719), C2 => n114, ZN => n1050);
   U1440 : AOI22_X1 port map( A1 => regs(1231), A2 => n166, B1 => regs(2255), 
                           B2 => n229, ZN => n1049);
   U1441 : NAND2_X1 port map( A1 => n1051, A2 => n1052, ZN => 
                           curr_proc_regs(206));
   U1442 : AOI222_X1 port map( A1 => regs(206), A2 => n10, B1 => regs(1742), B2
                           => n62, C1 => regs(718), C2 => n114, ZN => n1052);
   U1443 : AOI22_X1 port map( A1 => regs(1230), A2 => n166, B1 => regs(2254), 
                           B2 => n229, ZN => n1051);
   U1444 : NAND2_X1 port map( A1 => n1053, A2 => n1054, ZN => 
                           curr_proc_regs(205));
   U1445 : AOI222_X1 port map( A1 => regs(205), A2 => n10, B1 => regs(1741), B2
                           => n62, C1 => regs(717), C2 => n114, ZN => n1054);
   U1446 : AOI22_X1 port map( A1 => regs(1229), A2 => n166, B1 => regs(2253), 
                           B2 => n229, ZN => n1053);
   U1447 : NAND2_X1 port map( A1 => n1055, A2 => n1056, ZN => 
                           curr_proc_regs(204));
   U1448 : AOI222_X1 port map( A1 => regs(204), A2 => n10, B1 => regs(1740), B2
                           => n62, C1 => regs(716), C2 => n114, ZN => n1056);
   U1449 : AOI22_X1 port map( A1 => regs(1228), A2 => n166, B1 => regs(2252), 
                           B2 => n229, ZN => n1055);
   U1450 : NAND2_X1 port map( A1 => n1057, A2 => n1058, ZN => 
                           curr_proc_regs(203));
   U1451 : AOI222_X1 port map( A1 => regs(203), A2 => n10, B1 => regs(1739), B2
                           => n62, C1 => regs(715), C2 => n114, ZN => n1058);
   U1452 : AOI22_X1 port map( A1 => regs(1227), A2 => n166, B1 => regs(2251), 
                           B2 => n229, ZN => n1057);
   U1453 : NAND2_X1 port map( A1 => n1059, A2 => n1060, ZN => 
                           curr_proc_regs(202));
   U1454 : AOI222_X1 port map( A1 => regs(202), A2 => n10, B1 => regs(1738), B2
                           => n62, C1 => regs(714), C2 => n114, ZN => n1060);
   U1455 : AOI22_X1 port map( A1 => regs(1226), A2 => n166, B1 => regs(2250), 
                           B2 => n229, ZN => n1059);
   U1456 : NAND2_X1 port map( A1 => n1061, A2 => n1062, ZN => 
                           curr_proc_regs(201));
   U1457 : AOI222_X1 port map( A1 => regs(201), A2 => n10, B1 => regs(1737), B2
                           => n62, C1 => regs(713), C2 => n114, ZN => n1062);
   U1458 : AOI22_X1 port map( A1 => regs(1225), A2 => n166, B1 => regs(2249), 
                           B2 => n229, ZN => n1061);
   U1459 : NAND2_X1 port map( A1 => n1063, A2 => n1064, ZN => 
                           curr_proc_regs(200));
   U1460 : AOI222_X1 port map( A1 => regs(200), A2 => n10, B1 => regs(1736), B2
                           => n62, C1 => regs(712), C2 => n114, ZN => n1064);
   U1461 : AOI22_X1 port map( A1 => regs(1224), A2 => n166, B1 => regs(2248), 
                           B2 => n229, ZN => n1063);
   U1462 : NAND2_X1 port map( A1 => n1065, A2 => n1066, ZN => curr_proc_regs(1)
                           );
   U1463 : AOI222_X1 port map( A1 => regs(1), A2 => n10, B1 => regs(1537), B2 
                           => n62, C1 => regs(513), C2 => n114, ZN => n1066);
   U1464 : AOI22_X1 port map( A1 => regs(1025), A2 => n166, B1 => regs(2049), 
                           B2 => n229, ZN => n1065);
   U1465 : NAND2_X1 port map( A1 => n1067, A2 => n1068, ZN => 
                           curr_proc_regs(19));
   U1466 : AOI222_X1 port map( A1 => regs(19), A2 => n10, B1 => regs(1555), B2 
                           => n62, C1 => regs(531), C2 => n114, ZN => n1068);
   U1467 : AOI22_X1 port map( A1 => regs(1043), A2 => n166, B1 => regs(2067), 
                           B2 => n228, ZN => n1067);
   U1468 : NAND2_X1 port map( A1 => n1069, A2 => n1070, ZN => 
                           curr_proc_regs(199));
   U1469 : AOI222_X1 port map( A1 => regs(199), A2 => n10, B1 => regs(1735), B2
                           => n62, C1 => regs(711), C2 => n114, ZN => n1070);
   U1470 : AOI22_X1 port map( A1 => regs(1223), A2 => n166, B1 => regs(2247), 
                           B2 => n228, ZN => n1069);
   U1471 : NAND2_X1 port map( A1 => n1071, A2 => n1072, ZN => 
                           curr_proc_regs(198));
   U1472 : AOI222_X1 port map( A1 => regs(198), A2 => n10, B1 => regs(1734), B2
                           => n62, C1 => regs(710), C2 => n114, ZN => n1072);
   U1473 : AOI22_X1 port map( A1 => regs(1222), A2 => n166, B1 => regs(2246), 
                           B2 => n228, ZN => n1071);
   U1474 : NAND2_X1 port map( A1 => n1073, A2 => n1074, ZN => 
                           curr_proc_regs(197));
   U1475 : AOI222_X1 port map( A1 => regs(197), A2 => n9, B1 => regs(1733), B2 
                           => n61, C1 => regs(709), C2 => n113, ZN => n1074);
   U1476 : AOI22_X1 port map( A1 => regs(1221), A2 => n165, B1 => regs(2245), 
                           B2 => n228, ZN => n1073);
   U1477 : NAND2_X1 port map( A1 => n1075, A2 => n1076, ZN => 
                           curr_proc_regs(196));
   U1478 : AOI222_X1 port map( A1 => regs(196), A2 => n9, B1 => regs(1732), B2 
                           => n61, C1 => regs(708), C2 => n113, ZN => n1076);
   U1479 : AOI22_X1 port map( A1 => regs(1220), A2 => n165, B1 => regs(2244), 
                           B2 => n228, ZN => n1075);
   U1480 : NAND2_X1 port map( A1 => n1077, A2 => n1078, ZN => 
                           curr_proc_regs(195));
   U1481 : AOI222_X1 port map( A1 => regs(195), A2 => n9, B1 => regs(1731), B2 
                           => n61, C1 => regs(707), C2 => n113, ZN => n1078);
   U1482 : AOI22_X1 port map( A1 => regs(1219), A2 => n165, B1 => regs(2243), 
                           B2 => n228, ZN => n1077);
   U1483 : NAND2_X1 port map( A1 => n1079, A2 => n1080, ZN => 
                           curr_proc_regs(194));
   U1484 : AOI222_X1 port map( A1 => regs(194), A2 => n9, B1 => regs(1730), B2 
                           => n61, C1 => regs(706), C2 => n113, ZN => n1080);
   U1485 : AOI22_X1 port map( A1 => regs(1218), A2 => n165, B1 => regs(2242), 
                           B2 => n228, ZN => n1079);
   U1486 : NAND2_X1 port map( A1 => n1081, A2 => n1082, ZN => 
                           curr_proc_regs(193));
   U1487 : AOI222_X1 port map( A1 => regs(193), A2 => n9, B1 => regs(1729), B2 
                           => n61, C1 => regs(705), C2 => n113, ZN => n1082);
   U1488 : AOI22_X1 port map( A1 => regs(1217), A2 => n165, B1 => regs(2241), 
                           B2 => n228, ZN => n1081);
   U1489 : NAND2_X1 port map( A1 => n1083, A2 => n1084, ZN => 
                           curr_proc_regs(192));
   U1490 : AOI222_X1 port map( A1 => regs(192), A2 => n9, B1 => regs(1728), B2 
                           => n61, C1 => regs(704), C2 => n113, ZN => n1084);
   U1491 : AOI22_X1 port map( A1 => regs(1216), A2 => n165, B1 => regs(2240), 
                           B2 => n228, ZN => n1083);
   U1492 : NAND2_X1 port map( A1 => n1085, A2 => n1086, ZN => 
                           curr_proc_regs(191));
   U1493 : AOI222_X1 port map( A1 => regs(191), A2 => n9, B1 => regs(1727), B2 
                           => n61, C1 => regs(703), C2 => n113, ZN => n1086);
   U1494 : AOI22_X1 port map( A1 => regs(1215), A2 => n165, B1 => regs(2239), 
                           B2 => n228, ZN => n1085);
   U1495 : NAND2_X1 port map( A1 => n1087, A2 => n1088, ZN => 
                           curr_proc_regs(190));
   U1496 : AOI222_X1 port map( A1 => regs(190), A2 => n9, B1 => regs(1726), B2 
                           => n61, C1 => regs(702), C2 => n113, ZN => n1088);
   U1497 : AOI22_X1 port map( A1 => regs(1214), A2 => n165, B1 => regs(2238), 
                           B2 => n228, ZN => n1087);
   U1498 : NAND2_X1 port map( A1 => n1089, A2 => n1090, ZN => 
                           curr_proc_regs(18));
   U1499 : AOI222_X1 port map( A1 => regs(18), A2 => n9, B1 => regs(1554), B2 
                           => n61, C1 => regs(530), C2 => n113, ZN => n1090);
   U1500 : AOI22_X1 port map( A1 => regs(1042), A2 => n165, B1 => regs(2066), 
                           B2 => n228, ZN => n1089);
   U1501 : NAND2_X1 port map( A1 => n1091, A2 => n1092, ZN => 
                           curr_proc_regs(189));
   U1502 : AOI222_X1 port map( A1 => regs(189), A2 => n9, B1 => regs(1725), B2 
                           => n61, C1 => regs(701), C2 => n113, ZN => n1092);
   U1503 : AOI22_X1 port map( A1 => regs(1213), A2 => n165, B1 => regs(2237), 
                           B2 => n227, ZN => n1091);
   U1504 : NAND2_X1 port map( A1 => n1093, A2 => n1094, ZN => 
                           curr_proc_regs(188));
   U1505 : AOI222_X1 port map( A1 => regs(188), A2 => n9, B1 => regs(1724), B2 
                           => n61, C1 => regs(700), C2 => n113, ZN => n1094);
   U1506 : AOI22_X1 port map( A1 => regs(1212), A2 => n165, B1 => regs(2236), 
                           B2 => n227, ZN => n1093);
   U1507 : NAND2_X1 port map( A1 => n1095, A2 => n1096, ZN => 
                           curr_proc_regs(187));
   U1508 : AOI222_X1 port map( A1 => regs(187), A2 => n9, B1 => regs(1723), B2 
                           => n61, C1 => regs(699), C2 => n113, ZN => n1096);
   U1509 : AOI22_X1 port map( A1 => regs(1211), A2 => n165, B1 => regs(2235), 
                           B2 => n227, ZN => n1095);
   U1510 : NAND2_X1 port map( A1 => n1097, A2 => n1098, ZN => 
                           curr_proc_regs(186));
   U1511 : AOI222_X1 port map( A1 => regs(186), A2 => n8, B1 => regs(1722), B2 
                           => n60, C1 => regs(698), C2 => n112, ZN => n1098);
   U1512 : AOI22_X1 port map( A1 => regs(1210), A2 => n164, B1 => regs(2234), 
                           B2 => n227, ZN => n1097);
   U1513 : NAND2_X1 port map( A1 => n1099, A2 => n1100, ZN => 
                           curr_proc_regs(185));
   U1514 : AOI222_X1 port map( A1 => regs(185), A2 => n8, B1 => regs(1721), B2 
                           => n60, C1 => regs(697), C2 => n112, ZN => n1100);
   U1515 : AOI22_X1 port map( A1 => regs(1209), A2 => n164, B1 => regs(2233), 
                           B2 => n227, ZN => n1099);
   U1516 : NAND2_X1 port map( A1 => n1101, A2 => n1102, ZN => 
                           curr_proc_regs(184));
   U1517 : AOI222_X1 port map( A1 => regs(184), A2 => n8, B1 => regs(1720), B2 
                           => n60, C1 => regs(696), C2 => n112, ZN => n1102);
   U1518 : AOI22_X1 port map( A1 => regs(1208), A2 => n164, B1 => regs(2232), 
                           B2 => n227, ZN => n1101);
   U1519 : NAND2_X1 port map( A1 => n1103, A2 => n1104, ZN => 
                           curr_proc_regs(183));
   U1520 : AOI222_X1 port map( A1 => regs(183), A2 => n8, B1 => regs(1719), B2 
                           => n60, C1 => regs(695), C2 => n112, ZN => n1104);
   U1521 : AOI22_X1 port map( A1 => regs(1207), A2 => n164, B1 => regs(2231), 
                           B2 => n227, ZN => n1103);
   U1522 : NAND2_X1 port map( A1 => n1105, A2 => n1106, ZN => 
                           curr_proc_regs(182));
   U1523 : AOI222_X1 port map( A1 => regs(182), A2 => n8, B1 => regs(1718), B2 
                           => n60, C1 => regs(694), C2 => n112, ZN => n1106);
   U1524 : AOI22_X1 port map( A1 => regs(1206), A2 => n164, B1 => regs(2230), 
                           B2 => n227, ZN => n1105);
   U1525 : NAND2_X1 port map( A1 => n1107, A2 => n1108, ZN => 
                           curr_proc_regs(181));
   U1526 : AOI222_X1 port map( A1 => regs(181), A2 => n8, B1 => regs(1717), B2 
                           => n60, C1 => regs(693), C2 => n112, ZN => n1108);
   U1527 : AOI22_X1 port map( A1 => regs(1205), A2 => n164, B1 => regs(2229), 
                           B2 => n227, ZN => n1107);
   U1528 : NAND2_X1 port map( A1 => n1109, A2 => n1110, ZN => 
                           curr_proc_regs(180));
   U1529 : AOI222_X1 port map( A1 => regs(180), A2 => n8, B1 => regs(1716), B2 
                           => n60, C1 => regs(692), C2 => n112, ZN => n1110);
   U1530 : AOI22_X1 port map( A1 => regs(1204), A2 => n164, B1 => regs(2228), 
                           B2 => n227, ZN => n1109);
   U1531 : NAND2_X1 port map( A1 => n1111, A2 => n1112, ZN => 
                           curr_proc_regs(17));
   U1532 : AOI222_X1 port map( A1 => regs(17), A2 => n8, B1 => regs(1553), B2 
                           => n60, C1 => regs(529), C2 => n112, ZN => n1112);
   U1533 : AOI22_X1 port map( A1 => regs(1041), A2 => n164, B1 => regs(2065), 
                           B2 => n227, ZN => n1111);
   U1534 : NAND2_X1 port map( A1 => n1113, A2 => n1114, ZN => 
                           curr_proc_regs(179));
   U1535 : AOI222_X1 port map( A1 => regs(179), A2 => n8, B1 => regs(1715), B2 
                           => n60, C1 => regs(691), C2 => n112, ZN => n1114);
   U1536 : AOI22_X1 port map( A1 => regs(1203), A2 => n164, B1 => regs(2227), 
                           B2 => n227, ZN => n1113);
   U1537 : NAND2_X1 port map( A1 => n1115, A2 => n1116, ZN => 
                           curr_proc_regs(178));
   U1538 : AOI222_X1 port map( A1 => regs(178), A2 => n8, B1 => regs(1714), B2 
                           => n60, C1 => regs(690), C2 => n112, ZN => n1116);
   U1539 : AOI22_X1 port map( A1 => regs(1202), A2 => n164, B1 => regs(2226), 
                           B2 => n226, ZN => n1115);
   U1540 : NAND2_X1 port map( A1 => n1117, A2 => n1118, ZN => 
                           curr_proc_regs(177));
   U1541 : AOI222_X1 port map( A1 => regs(177), A2 => n8, B1 => regs(1713), B2 
                           => n60, C1 => regs(689), C2 => n112, ZN => n1118);
   U1542 : AOI22_X1 port map( A1 => regs(1201), A2 => n164, B1 => regs(2225), 
                           B2 => n226, ZN => n1117);
   U1543 : NAND2_X1 port map( A1 => n1119, A2 => n1120, ZN => 
                           curr_proc_regs(176));
   U1544 : AOI222_X1 port map( A1 => regs(176), A2 => n8, B1 => regs(1712), B2 
                           => n60, C1 => regs(688), C2 => n112, ZN => n1120);
   U1545 : AOI22_X1 port map( A1 => regs(1200), A2 => n164, B1 => regs(2224), 
                           B2 => n226, ZN => n1119);
   U1546 : NAND2_X1 port map( A1 => n1121, A2 => n1122, ZN => 
                           curr_proc_regs(175));
   U1547 : AOI222_X1 port map( A1 => regs(175), A2 => n7, B1 => regs(1711), B2 
                           => n59, C1 => regs(687), C2 => n111, ZN => n1122);
   U1548 : AOI22_X1 port map( A1 => regs(1199), A2 => n163, B1 => regs(2223), 
                           B2 => n226, ZN => n1121);
   U1549 : NAND2_X1 port map( A1 => n1123, A2 => n1124, ZN => 
                           curr_proc_regs(174));
   U1550 : AOI222_X1 port map( A1 => regs(174), A2 => n7, B1 => regs(1710), B2 
                           => n59, C1 => regs(686), C2 => n111, ZN => n1124);
   U1551 : AOI22_X1 port map( A1 => regs(1198), A2 => n163, B1 => regs(2222), 
                           B2 => n226, ZN => n1123);
   U1552 : NAND2_X1 port map( A1 => n1125, A2 => n1126, ZN => 
                           curr_proc_regs(173));
   U1553 : AOI222_X1 port map( A1 => regs(173), A2 => n7, B1 => regs(1709), B2 
                           => n59, C1 => regs(685), C2 => n111, ZN => n1126);
   U1554 : AOI22_X1 port map( A1 => regs(1197), A2 => n163, B1 => regs(2221), 
                           B2 => n226, ZN => n1125);
   U1555 : NAND2_X1 port map( A1 => n1127, A2 => n1128, ZN => 
                           curr_proc_regs(172));
   U1556 : AOI222_X1 port map( A1 => regs(172), A2 => n7, B1 => regs(1708), B2 
                           => n59, C1 => regs(684), C2 => n111, ZN => n1128);
   U1557 : AOI22_X1 port map( A1 => regs(1196), A2 => n163, B1 => regs(2220), 
                           B2 => n226, ZN => n1127);
   U1558 : NAND2_X1 port map( A1 => n1129, A2 => n1130, ZN => 
                           curr_proc_regs(171));
   U1559 : AOI222_X1 port map( A1 => regs(171), A2 => n7, B1 => regs(1707), B2 
                           => n59, C1 => regs(683), C2 => n111, ZN => n1130);
   U1560 : AOI22_X1 port map( A1 => regs(1195), A2 => n163, B1 => regs(2219), 
                           B2 => n226, ZN => n1129);
   U1561 : NAND2_X1 port map( A1 => n1131, A2 => n1132, ZN => 
                           curr_proc_regs(170));
   U1562 : AOI222_X1 port map( A1 => regs(170), A2 => n7, B1 => regs(1706), B2 
                           => n59, C1 => regs(682), C2 => n111, ZN => n1132);
   U1563 : AOI22_X1 port map( A1 => regs(1194), A2 => n163, B1 => regs(2218), 
                           B2 => n226, ZN => n1131);
   U1564 : NAND2_X1 port map( A1 => n1133, A2 => n1134, ZN => 
                           curr_proc_regs(16));
   U1565 : AOI222_X1 port map( A1 => regs(16), A2 => n7, B1 => regs(1552), B2 
                           => n59, C1 => regs(528), C2 => n111, ZN => n1134);
   U1566 : AOI22_X1 port map( A1 => regs(1040), A2 => n163, B1 => regs(2064), 
                           B2 => n226, ZN => n1133);
   U1567 : NAND2_X1 port map( A1 => n1135, A2 => n1136, ZN => 
                           curr_proc_regs(169));
   U1568 : AOI222_X1 port map( A1 => regs(169), A2 => n7, B1 => regs(1705), B2 
                           => n59, C1 => regs(681), C2 => n111, ZN => n1136);
   U1569 : AOI22_X1 port map( A1 => regs(1193), A2 => n163, B1 => regs(2217), 
                           B2 => n226, ZN => n1135);
   U1570 : NAND2_X1 port map( A1 => n1137, A2 => n1138, ZN => 
                           curr_proc_regs(168));
   U1571 : AOI222_X1 port map( A1 => regs(168), A2 => n7, B1 => regs(1704), B2 
                           => n59, C1 => regs(680), C2 => n111, ZN => n1138);
   U1572 : AOI22_X1 port map( A1 => regs(1192), A2 => n163, B1 => regs(2216), 
                           B2 => n226, ZN => n1137);
   U1573 : NAND2_X1 port map( A1 => n1139, A2 => n1140, ZN => 
                           curr_proc_regs(167));
   U1574 : AOI222_X1 port map( A1 => regs(167), A2 => n7, B1 => regs(1703), B2 
                           => n59, C1 => regs(679), C2 => n111, ZN => n1140);
   U1575 : AOI22_X1 port map( A1 => regs(1191), A2 => n163, B1 => regs(2215), 
                           B2 => n225, ZN => n1139);
   U1576 : NAND2_X1 port map( A1 => n1141, A2 => n1142, ZN => 
                           curr_proc_regs(166));
   U1577 : AOI222_X1 port map( A1 => regs(166), A2 => n7, B1 => regs(1702), B2 
                           => n59, C1 => regs(678), C2 => n111, ZN => n1142);
   U1578 : AOI22_X1 port map( A1 => regs(1190), A2 => n163, B1 => regs(2214), 
                           B2 => n225, ZN => n1141);
   U1579 : NAND2_X1 port map( A1 => n1143, A2 => n1144, ZN => 
                           curr_proc_regs(165));
   U1580 : AOI222_X1 port map( A1 => regs(165), A2 => n7, B1 => regs(1701), B2 
                           => n59, C1 => regs(677), C2 => n111, ZN => n1144);
   U1581 : AOI22_X1 port map( A1 => regs(1189), A2 => n163, B1 => regs(2213), 
                           B2 => n225, ZN => n1143);
   U1582 : NAND2_X1 port map( A1 => n1145, A2 => n1146, ZN => 
                           curr_proc_regs(164));
   U1583 : AOI222_X1 port map( A1 => regs(164), A2 => n6, B1 => regs(1700), B2 
                           => n58, C1 => regs(676), C2 => n110, ZN => n1146);
   U1584 : AOI22_X1 port map( A1 => regs(1188), A2 => n162, B1 => regs(2212), 
                           B2 => n225, ZN => n1145);
   U1585 : NAND2_X1 port map( A1 => n1147, A2 => n1148, ZN => 
                           curr_proc_regs(163));
   U1586 : AOI222_X1 port map( A1 => regs(163), A2 => n6, B1 => regs(1699), B2 
                           => n58, C1 => regs(675), C2 => n110, ZN => n1148);
   U1587 : AOI22_X1 port map( A1 => regs(1187), A2 => n162, B1 => regs(2211), 
                           B2 => n225, ZN => n1147);
   U1588 : NAND2_X1 port map( A1 => n1149, A2 => n1150, ZN => 
                           curr_proc_regs(162));
   U1589 : AOI222_X1 port map( A1 => regs(162), A2 => n6, B1 => regs(1698), B2 
                           => n58, C1 => regs(674), C2 => n110, ZN => n1150);
   U1590 : AOI22_X1 port map( A1 => regs(1186), A2 => n162, B1 => regs(2210), 
                           B2 => n225, ZN => n1149);
   U1591 : NAND2_X1 port map( A1 => n1151, A2 => n1152, ZN => 
                           curr_proc_regs(161));
   U1592 : AOI222_X1 port map( A1 => regs(161), A2 => n6, B1 => regs(1697), B2 
                           => n58, C1 => regs(673), C2 => n110, ZN => n1152);
   U1593 : AOI22_X1 port map( A1 => regs(1185), A2 => n162, B1 => regs(2209), 
                           B2 => n225, ZN => n1151);
   U1594 : NAND2_X1 port map( A1 => n1153, A2 => n1154, ZN => 
                           curr_proc_regs(160));
   U1595 : AOI222_X1 port map( A1 => regs(160), A2 => n6, B1 => regs(1696), B2 
                           => n58, C1 => regs(672), C2 => n110, ZN => n1154);
   U1596 : AOI22_X1 port map( A1 => regs(1184), A2 => n162, B1 => regs(2208), 
                           B2 => n225, ZN => n1153);
   U1597 : NAND2_X1 port map( A1 => n1155, A2 => n1156, ZN => 
                           curr_proc_regs(15));
   U1598 : AOI222_X1 port map( A1 => regs(15), A2 => n6, B1 => regs(1551), B2 
                           => n58, C1 => regs(527), C2 => n110, ZN => n1156);
   U1599 : AOI22_X1 port map( A1 => regs(1039), A2 => n162, B1 => regs(2063), 
                           B2 => n225, ZN => n1155);
   U1600 : NAND2_X1 port map( A1 => n1157, A2 => n1158, ZN => 
                           curr_proc_regs(159));
   U1601 : AOI222_X1 port map( A1 => regs(159), A2 => n6, B1 => regs(1695), B2 
                           => n58, C1 => regs(671), C2 => n110, ZN => n1158);
   U1602 : AOI22_X1 port map( A1 => regs(1183), A2 => n162, B1 => regs(2207), 
                           B2 => n225, ZN => n1157);
   U1603 : NAND2_X1 port map( A1 => n1159, A2 => n1160, ZN => 
                           curr_proc_regs(158));
   U1604 : AOI222_X1 port map( A1 => regs(158), A2 => n6, B1 => regs(1694), B2 
                           => n58, C1 => regs(670), C2 => n110, ZN => n1160);
   U1605 : AOI22_X1 port map( A1 => regs(1182), A2 => n162, B1 => regs(2206), 
                           B2 => n225, ZN => n1159);
   U1606 : NAND2_X1 port map( A1 => n1161, A2 => n1162, ZN => 
                           curr_proc_regs(157));
   U1607 : AOI222_X1 port map( A1 => regs(157), A2 => n6, B1 => regs(1693), B2 
                           => n58, C1 => regs(669), C2 => n110, ZN => n1162);
   U1608 : AOI22_X1 port map( A1 => regs(1181), A2 => n162, B1 => regs(2205), 
                           B2 => n224, ZN => n1161);
   U1609 : NAND2_X1 port map( A1 => n1163, A2 => n1164, ZN => 
                           curr_proc_regs(156));
   U1610 : AOI222_X1 port map( A1 => regs(156), A2 => n6, B1 => regs(1692), B2 
                           => n58, C1 => regs(668), C2 => n110, ZN => n1164);
   U1611 : AOI22_X1 port map( A1 => regs(1180), A2 => n162, B1 => regs(2204), 
                           B2 => n224, ZN => n1163);
   U1612 : NAND2_X1 port map( A1 => n1165, A2 => n1166, ZN => 
                           curr_proc_regs(155));
   U1613 : AOI222_X1 port map( A1 => regs(155), A2 => n6, B1 => regs(1691), B2 
                           => n58, C1 => regs(667), C2 => n110, ZN => n1166);
   U1614 : AOI22_X1 port map( A1 => regs(1179), A2 => n162, B1 => regs(2203), 
                           B2 => n224, ZN => n1165);
   U1615 : NAND2_X1 port map( A1 => n1167, A2 => n1168, ZN => 
                           curr_proc_regs(154));
   U1616 : AOI222_X1 port map( A1 => regs(154), A2 => n6, B1 => regs(1690), B2 
                           => n58, C1 => regs(666), C2 => n110, ZN => n1168);
   U1617 : AOI22_X1 port map( A1 => regs(1178), A2 => n162, B1 => regs(2202), 
                           B2 => n224, ZN => n1167);
   U1618 : NAND2_X1 port map( A1 => n1169, A2 => n1170, ZN => 
                           curr_proc_regs(153));
   U1619 : AOI222_X1 port map( A1 => regs(153), A2 => n5, B1 => regs(1689), B2 
                           => n57, C1 => regs(665), C2 => n109, ZN => n1170);
   U1620 : AOI22_X1 port map( A1 => regs(1177), A2 => n161, B1 => regs(2201), 
                           B2 => n224, ZN => n1169);
   U1621 : NAND2_X1 port map( A1 => n1171, A2 => n1172, ZN => 
                           curr_proc_regs(152));
   U1622 : AOI222_X1 port map( A1 => regs(152), A2 => n5, B1 => regs(1688), B2 
                           => n57, C1 => regs(664), C2 => n109, ZN => n1172);
   U1623 : AOI22_X1 port map( A1 => regs(1176), A2 => n161, B1 => regs(2200), 
                           B2 => n224, ZN => n1171);
   U1624 : NAND2_X1 port map( A1 => n1173, A2 => n1174, ZN => 
                           curr_proc_regs(151));
   U1625 : AOI222_X1 port map( A1 => regs(151), A2 => n5, B1 => regs(1687), B2 
                           => n57, C1 => regs(663), C2 => n109, ZN => n1174);
   U1626 : AOI22_X1 port map( A1 => regs(1175), A2 => n161, B1 => regs(2199), 
                           B2 => n224, ZN => n1173);
   U1627 : NAND2_X1 port map( A1 => n1175, A2 => n1176, ZN => 
                           curr_proc_regs(150));
   U1628 : AOI222_X1 port map( A1 => regs(150), A2 => n5, B1 => regs(1686), B2 
                           => n57, C1 => regs(662), C2 => n109, ZN => n1176);
   U1629 : AOI22_X1 port map( A1 => regs(1174), A2 => n161, B1 => regs(2198), 
                           B2 => n224, ZN => n1175);
   U1630 : NAND2_X1 port map( A1 => n1177, A2 => n1178, ZN => 
                           curr_proc_regs(14));
   U1631 : AOI222_X1 port map( A1 => regs(14), A2 => n5, B1 => regs(1550), B2 
                           => n57, C1 => regs(526), C2 => n109, ZN => n1178);
   U1632 : AOI22_X1 port map( A1 => regs(1038), A2 => n161, B1 => regs(2062), 
                           B2 => n224, ZN => n1177);
   U1633 : NAND2_X1 port map( A1 => n1179, A2 => n1180, ZN => 
                           curr_proc_regs(149));
   U1634 : AOI222_X1 port map( A1 => regs(149), A2 => n5, B1 => regs(1685), B2 
                           => n57, C1 => regs(661), C2 => n109, ZN => n1180);
   U1635 : AOI22_X1 port map( A1 => regs(1173), A2 => n161, B1 => regs(2197), 
                           B2 => n224, ZN => n1179);
   U1636 : NAND2_X1 port map( A1 => n1181, A2 => n1182, ZN => 
                           curr_proc_regs(148));
   U1637 : AOI222_X1 port map( A1 => regs(148), A2 => n5, B1 => regs(1684), B2 
                           => n57, C1 => regs(660), C2 => n109, ZN => n1182);
   U1638 : AOI22_X1 port map( A1 => regs(1172), A2 => n161, B1 => regs(2196), 
                           B2 => n224, ZN => n1181);
   U1639 : NAND2_X1 port map( A1 => n1183, A2 => n1184, ZN => 
                           curr_proc_regs(147));
   U1640 : AOI222_X1 port map( A1 => regs(147), A2 => n5, B1 => regs(1683), B2 
                           => n57, C1 => regs(659), C2 => n109, ZN => n1184);
   U1641 : AOI22_X1 port map( A1 => regs(1171), A2 => n161, B1 => regs(2195), 
                           B2 => n224, ZN => n1183);
   U1642 : NAND2_X1 port map( A1 => n1185, A2 => n1186, ZN => 
                           curr_proc_regs(146));
   U1643 : AOI222_X1 port map( A1 => regs(146), A2 => n5, B1 => regs(1682), B2 
                           => n57, C1 => regs(658), C2 => n109, ZN => n1186);
   U1644 : AOI22_X1 port map( A1 => regs(1170), A2 => n161, B1 => regs(2194), 
                           B2 => n223, ZN => n1185);
   U1645 : NAND2_X1 port map( A1 => n1187, A2 => n1188, ZN => 
                           curr_proc_regs(145));
   U1646 : AOI222_X1 port map( A1 => regs(145), A2 => n5, B1 => regs(1681), B2 
                           => n57, C1 => regs(657), C2 => n109, ZN => n1188);
   U1647 : AOI22_X1 port map( A1 => regs(1169), A2 => n161, B1 => regs(2193), 
                           B2 => n223, ZN => n1187);
   U1648 : NAND2_X1 port map( A1 => n1189, A2 => n1190, ZN => 
                           curr_proc_regs(144));
   U1649 : AOI222_X1 port map( A1 => regs(144), A2 => n5, B1 => regs(1680), B2 
                           => n57, C1 => regs(656), C2 => n109, ZN => n1190);
   U1650 : AOI22_X1 port map( A1 => regs(1168), A2 => n161, B1 => regs(2192), 
                           B2 => n223, ZN => n1189);
   U1651 : NAND2_X1 port map( A1 => n1191, A2 => n1192, ZN => 
                           curr_proc_regs(143));
   U1652 : AOI222_X1 port map( A1 => regs(143), A2 => n5, B1 => regs(1679), B2 
                           => n57, C1 => regs(655), C2 => n109, ZN => n1192);
   U1653 : AOI22_X1 port map( A1 => regs(1167), A2 => n161, B1 => regs(2191), 
                           B2 => n223, ZN => n1191);
   U1654 : NAND2_X1 port map( A1 => n1193, A2 => n1194, ZN => 
                           curr_proc_regs(142));
   U1655 : AOI222_X1 port map( A1 => regs(142), A2 => n4, B1 => regs(1678), B2 
                           => n56, C1 => regs(654), C2 => n108, ZN => n1194);
   U1656 : AOI22_X1 port map( A1 => regs(1166), A2 => n160, B1 => regs(2190), 
                           B2 => n223, ZN => n1193);
   U1657 : NAND2_X1 port map( A1 => n1195, A2 => n1196, ZN => 
                           curr_proc_regs(141));
   U1658 : AOI222_X1 port map( A1 => regs(141), A2 => n4, B1 => regs(1677), B2 
                           => n56, C1 => regs(653), C2 => n108, ZN => n1196);
   U1659 : AOI22_X1 port map( A1 => regs(1165), A2 => n160, B1 => regs(2189), 
                           B2 => n223, ZN => n1195);
   U1660 : NAND2_X1 port map( A1 => n1197, A2 => n1198, ZN => 
                           curr_proc_regs(140));
   U1661 : AOI222_X1 port map( A1 => regs(140), A2 => n4, B1 => regs(1676), B2 
                           => n56, C1 => regs(652), C2 => n108, ZN => n1198);
   U1662 : AOI22_X1 port map( A1 => regs(1164), A2 => n160, B1 => regs(2188), 
                           B2 => n223, ZN => n1197);
   U1663 : NAND2_X1 port map( A1 => n1199, A2 => n1200, ZN => 
                           curr_proc_regs(13));
   U1664 : AOI222_X1 port map( A1 => regs(13), A2 => n4, B1 => regs(1549), B2 
                           => n56, C1 => regs(525), C2 => n108, ZN => n1200);
   U1665 : AOI22_X1 port map( A1 => regs(1037), A2 => n160, B1 => regs(2061), 
                           B2 => n223, ZN => n1199);
   U1666 : NAND2_X1 port map( A1 => n1201, A2 => n1202, ZN => 
                           curr_proc_regs(139));
   U1667 : AOI222_X1 port map( A1 => regs(139), A2 => n4, B1 => regs(1675), B2 
                           => n56, C1 => regs(651), C2 => n108, ZN => n1202);
   U1668 : AOI22_X1 port map( A1 => regs(1163), A2 => n160, B1 => regs(2187), 
                           B2 => n223, ZN => n1201);
   U1669 : NAND2_X1 port map( A1 => n1203, A2 => n1204, ZN => 
                           curr_proc_regs(138));
   U1670 : AOI222_X1 port map( A1 => regs(138), A2 => n4, B1 => regs(1674), B2 
                           => n56, C1 => regs(650), C2 => n108, ZN => n1204);
   U1671 : AOI22_X1 port map( A1 => regs(1162), A2 => n160, B1 => regs(2186), 
                           B2 => n223, ZN => n1203);
   U1672 : NAND2_X1 port map( A1 => n1205, A2 => n1206, ZN => 
                           curr_proc_regs(137));
   U1673 : AOI222_X1 port map( A1 => regs(137), A2 => n4, B1 => regs(1673), B2 
                           => n56, C1 => regs(649), C2 => n108, ZN => n1206);
   U1674 : AOI22_X1 port map( A1 => regs(1161), A2 => n160, B1 => regs(2185), 
                           B2 => n223, ZN => n1205);
   U1675 : NAND2_X1 port map( A1 => n1207, A2 => n1208, ZN => 
                           curr_proc_regs(136));
   U1676 : AOI222_X1 port map( A1 => regs(136), A2 => n4, B1 => regs(1672), B2 
                           => n56, C1 => regs(648), C2 => n108, ZN => n1208);
   U1677 : AOI22_X1 port map( A1 => regs(1160), A2 => n160, B1 => regs(2184), 
                           B2 => n223, ZN => n1207);
   U1678 : NAND2_X1 port map( A1 => n1209, A2 => n1210, ZN => 
                           curr_proc_regs(135));
   U1679 : AOI222_X1 port map( A1 => regs(135), A2 => n4, B1 => regs(1671), B2 
                           => n56, C1 => regs(647), C2 => n108, ZN => n1210);
   U1680 : AOI22_X1 port map( A1 => regs(1159), A2 => n160, B1 => regs(2183), 
                           B2 => n222, ZN => n1209);
   U1681 : NAND2_X1 port map( A1 => n1211, A2 => n1212, ZN => 
                           curr_proc_regs(134));
   U1682 : AOI222_X1 port map( A1 => regs(134), A2 => n4, B1 => regs(1670), B2 
                           => n56, C1 => regs(646), C2 => n108, ZN => n1212);
   U1683 : AOI22_X1 port map( A1 => regs(1158), A2 => n160, B1 => regs(2182), 
                           B2 => n222, ZN => n1211);
   U1684 : NAND2_X1 port map( A1 => n1213, A2 => n1214, ZN => 
                           curr_proc_regs(133));
   U1685 : AOI222_X1 port map( A1 => regs(133), A2 => n4, B1 => regs(1669), B2 
                           => n56, C1 => regs(645), C2 => n108, ZN => n1214);
   U1686 : AOI22_X1 port map( A1 => regs(1157), A2 => n160, B1 => regs(2181), 
                           B2 => n222, ZN => n1213);
   U1687 : NAND2_X1 port map( A1 => n1215, A2 => n1216, ZN => 
                           curr_proc_regs(132));
   U1688 : AOI222_X1 port map( A1 => regs(132), A2 => n4, B1 => regs(1668), B2 
                           => n56, C1 => regs(644), C2 => n108, ZN => n1216);
   U1689 : AOI22_X1 port map( A1 => regs(1156), A2 => n160, B1 => regs(2180), 
                           B2 => n222, ZN => n1215);
   U1690 : NAND2_X1 port map( A1 => n1217, A2 => n1218, ZN => 
                           curr_proc_regs(131));
   U1691 : AOI222_X1 port map( A1 => regs(131), A2 => n3, B1 => regs(1667), B2 
                           => n55, C1 => regs(643), C2 => n107, ZN => n1218);
   U1692 : AOI22_X1 port map( A1 => regs(1155), A2 => n159, B1 => regs(2179), 
                           B2 => n222, ZN => n1217);
   U1693 : NAND2_X1 port map( A1 => n1219, A2 => n1220, ZN => 
                           curr_proc_regs(130));
   U1694 : AOI222_X1 port map( A1 => regs(130), A2 => n3, B1 => regs(1666), B2 
                           => n55, C1 => regs(642), C2 => n107, ZN => n1220);
   U1695 : AOI22_X1 port map( A1 => regs(1154), A2 => n159, B1 => regs(2178), 
                           B2 => n222, ZN => n1219);
   U1696 : NAND2_X1 port map( A1 => n1221, A2 => n1222, ZN => 
                           curr_proc_regs(12));
   U1697 : AOI222_X1 port map( A1 => regs(12), A2 => n3, B1 => regs(1548), B2 
                           => n55, C1 => regs(524), C2 => n107, ZN => n1222);
   U1698 : AOI22_X1 port map( A1 => regs(1036), A2 => n159, B1 => regs(2060), 
                           B2 => n222, ZN => n1221);
   U1699 : NAND2_X1 port map( A1 => n1223, A2 => n1224, ZN => 
                           curr_proc_regs(129));
   U1700 : AOI222_X1 port map( A1 => regs(129), A2 => n3, B1 => regs(1665), B2 
                           => n55, C1 => regs(641), C2 => n107, ZN => n1224);
   U1701 : AOI22_X1 port map( A1 => regs(1153), A2 => n159, B1 => regs(2177), 
                           B2 => n222, ZN => n1223);
   U1702 : NAND2_X1 port map( A1 => n1225, A2 => n1226, ZN => 
                           curr_proc_regs(128));
   U1703 : AOI222_X1 port map( A1 => regs(128), A2 => n3, B1 => regs(1664), B2 
                           => n55, C1 => regs(640), C2 => n107, ZN => n1226);
   U1704 : AOI22_X1 port map( A1 => regs(1152), A2 => n159, B1 => regs(2176), 
                           B2 => n222, ZN => n1225);
   U1705 : NAND2_X1 port map( A1 => n1227, A2 => n1228, ZN => 
                           curr_proc_regs(127));
   U1706 : AOI222_X1 port map( A1 => regs(127), A2 => n3, B1 => regs(1663), B2 
                           => n55, C1 => regs(639), C2 => n107, ZN => n1228);
   U1707 : AOI22_X1 port map( A1 => regs(1151), A2 => n159, B1 => regs(2175), 
                           B2 => n222, ZN => n1227);
   U1708 : NAND2_X1 port map( A1 => n1229, A2 => n1230, ZN => 
                           curr_proc_regs(126));
   U1709 : AOI222_X1 port map( A1 => regs(126), A2 => n3, B1 => regs(1662), B2 
                           => n55, C1 => regs(638), C2 => n107, ZN => n1230);
   U1710 : AOI22_X1 port map( A1 => regs(1150), A2 => n159, B1 => regs(2174), 
                           B2 => n222, ZN => n1229);
   U1711 : NAND2_X1 port map( A1 => n1231, A2 => n1232, ZN => 
                           curr_proc_regs(125));
   U1712 : AOI222_X1 port map( A1 => regs(125), A2 => n3, B1 => regs(1661), B2 
                           => n55, C1 => regs(637), C2 => n107, ZN => n1232);
   U1713 : AOI22_X1 port map( A1 => regs(1149), A2 => n159, B1 => regs(2173), 
                           B2 => n222, ZN => n1231);
   U1714 : NAND2_X1 port map( A1 => n1233, A2 => n1234, ZN => 
                           curr_proc_regs(124));
   U1715 : AOI222_X1 port map( A1 => regs(124), A2 => n3, B1 => regs(1660), B2 
                           => n55, C1 => regs(636), C2 => n107, ZN => n1234);
   U1716 : AOI22_X1 port map( A1 => regs(1148), A2 => n159, B1 => regs(2172), 
                           B2 => n221, ZN => n1233);
   U1717 : NAND2_X1 port map( A1 => n1235, A2 => n1236, ZN => 
                           curr_proc_regs(123));
   U1718 : AOI222_X1 port map( A1 => regs(123), A2 => n3, B1 => regs(1659), B2 
                           => n55, C1 => regs(635), C2 => n107, ZN => n1236);
   U1719 : AOI22_X1 port map( A1 => regs(1147), A2 => n159, B1 => regs(2171), 
                           B2 => n221, ZN => n1235);
   U1720 : NAND2_X1 port map( A1 => n1237, A2 => n1238, ZN => 
                           curr_proc_regs(122));
   U1721 : AOI222_X1 port map( A1 => regs(122), A2 => n3, B1 => regs(1658), B2 
                           => n55, C1 => regs(634), C2 => n107, ZN => n1238);
   U1722 : AOI22_X1 port map( A1 => regs(1146), A2 => n159, B1 => regs(2170), 
                           B2 => n221, ZN => n1237);
   U1723 : NAND2_X1 port map( A1 => n1239, A2 => n1240, ZN => 
                           curr_proc_regs(121));
   U1724 : AOI222_X1 port map( A1 => regs(121), A2 => n3, B1 => regs(1657), B2 
                           => n55, C1 => regs(633), C2 => n107, ZN => n1240);
   U1725 : AOI22_X1 port map( A1 => regs(1145), A2 => n159, B1 => regs(2169), 
                           B2 => n221, ZN => n1239);
   U1726 : NAND2_X1 port map( A1 => n1241, A2 => n1242, ZN => 
                           curr_proc_regs(120));
   U1727 : AOI222_X1 port map( A1 => regs(120), A2 => n2, B1 => regs(1656), B2 
                           => n54, C1 => regs(632), C2 => n106, ZN => n1242);
   U1728 : AOI22_X1 port map( A1 => regs(1144), A2 => n158, B1 => regs(2168), 
                           B2 => n221, ZN => n1241);
   U1729 : NAND2_X1 port map( A1 => n1243, A2 => n1244, ZN => 
                           curr_proc_regs(11));
   U1730 : AOI222_X1 port map( A1 => regs(11), A2 => n2, B1 => regs(1547), B2 
                           => n54, C1 => regs(523), C2 => n106, ZN => n1244);
   U1731 : AOI22_X1 port map( A1 => regs(1035), A2 => n158, B1 => regs(2059), 
                           B2 => n221, ZN => n1243);
   U1732 : NAND2_X1 port map( A1 => n1245, A2 => n1246, ZN => 
                           curr_proc_regs(119));
   U1733 : AOI222_X1 port map( A1 => regs(119), A2 => n2, B1 => regs(1655), B2 
                           => n54, C1 => regs(631), C2 => n106, ZN => n1246);
   U1734 : AOI22_X1 port map( A1 => regs(1143), A2 => n158, B1 => regs(2167), 
                           B2 => n221, ZN => n1245);
   U1735 : NAND2_X1 port map( A1 => n1247, A2 => n1248, ZN => 
                           curr_proc_regs(118));
   U1736 : AOI222_X1 port map( A1 => regs(118), A2 => n2, B1 => regs(1654), B2 
                           => n54, C1 => regs(630), C2 => n106, ZN => n1248);
   U1737 : AOI22_X1 port map( A1 => regs(1142), A2 => n158, B1 => regs(2166), 
                           B2 => n221, ZN => n1247);
   U1738 : NAND2_X1 port map( A1 => n1249, A2 => n1250, ZN => 
                           curr_proc_regs(117));
   U1739 : AOI222_X1 port map( A1 => regs(117), A2 => n2, B1 => regs(1653), B2 
                           => n54, C1 => regs(629), C2 => n106, ZN => n1250);
   U1740 : AOI22_X1 port map( A1 => regs(1141), A2 => n158, B1 => regs(2165), 
                           B2 => n221, ZN => n1249);
   U1741 : NAND2_X1 port map( A1 => n1251, A2 => n1252, ZN => 
                           curr_proc_regs(116));
   U1742 : AOI222_X1 port map( A1 => regs(116), A2 => n2, B1 => regs(1652), B2 
                           => n54, C1 => regs(628), C2 => n106, ZN => n1252);
   U1743 : AOI22_X1 port map( A1 => regs(1140), A2 => n158, B1 => regs(2164), 
                           B2 => n221, ZN => n1251);
   U1744 : NAND2_X1 port map( A1 => n1253, A2 => n1254, ZN => 
                           curr_proc_regs(115));
   U1745 : AOI222_X1 port map( A1 => regs(115), A2 => n2, B1 => regs(1651), B2 
                           => n54, C1 => regs(627), C2 => n106, ZN => n1254);
   U1746 : AOI22_X1 port map( A1 => regs(1139), A2 => n158, B1 => regs(2163), 
                           B2 => n221, ZN => n1253);
   U1747 : NAND2_X1 port map( A1 => n1255, A2 => n1256, ZN => 
                           curr_proc_regs(114));
   U1748 : AOI222_X1 port map( A1 => regs(114), A2 => n2, B1 => regs(1650), B2 
                           => n54, C1 => regs(626), C2 => n106, ZN => n1256);
   U1749 : AOI22_X1 port map( A1 => regs(1138), A2 => n158, B1 => regs(2162), 
                           B2 => n221, ZN => n1255);
   U1750 : NAND2_X1 port map( A1 => n1257, A2 => n1258, ZN => 
                           curr_proc_regs(113));
   U1751 : AOI222_X1 port map( A1 => regs(113), A2 => n2, B1 => regs(1649), B2 
                           => n54, C1 => regs(625), C2 => n106, ZN => n1258);
   U1752 : AOI22_X1 port map( A1 => regs(1137), A2 => n158, B1 => regs(2161), 
                           B2 => n220, ZN => n1257);
   U1753 : NAND2_X1 port map( A1 => n1259, A2 => n1260, ZN => 
                           curr_proc_regs(112));
   U1754 : AOI222_X1 port map( A1 => regs(112), A2 => n2, B1 => regs(1648), B2 
                           => n54, C1 => regs(624), C2 => n106, ZN => n1260);
   U1755 : AOI22_X1 port map( A1 => regs(1136), A2 => n158, B1 => regs(2160), 
                           B2 => n220, ZN => n1259);
   U1756 : NAND2_X1 port map( A1 => n1261, A2 => n1262, ZN => 
                           curr_proc_regs(111));
   U1757 : AOI222_X1 port map( A1 => regs(111), A2 => n2, B1 => regs(1647), B2 
                           => n54, C1 => regs(623), C2 => n106, ZN => n1262);
   U1758 : AOI22_X1 port map( A1 => regs(1135), A2 => n158, B1 => regs(2159), 
                           B2 => n220, ZN => n1261);
   U1759 : NAND2_X1 port map( A1 => n1263, A2 => n1264, ZN => 
                           curr_proc_regs(110));
   U1760 : AOI222_X1 port map( A1 => regs(110), A2 => n2, B1 => regs(1646), B2 
                           => n54, C1 => regs(622), C2 => n106, ZN => n1264);
   U1761 : AOI22_X1 port map( A1 => regs(1134), A2 => n158, B1 => regs(2158), 
                           B2 => n220, ZN => n1263);
   U1762 : NAND2_X1 port map( A1 => n1265, A2 => n1266, ZN => 
                           curr_proc_regs(10));
   U1763 : AOI222_X1 port map( A1 => regs(10), A2 => n1, B1 => regs(1546), B2 
                           => n53, C1 => regs(522), C2 => n105, ZN => n1266);
   U1764 : AOI22_X1 port map( A1 => regs(1034), A2 => n157, B1 => regs(2058), 
                           B2 => n220, ZN => n1265);
   U1765 : NAND2_X1 port map( A1 => n1267, A2 => n1268, ZN => 
                           curr_proc_regs(109));
   U1766 : AOI222_X1 port map( A1 => regs(109), A2 => n1, B1 => regs(1645), B2 
                           => n53, C1 => regs(621), C2 => n105, ZN => n1268);
   U1767 : AOI22_X1 port map( A1 => regs(1133), A2 => n157, B1 => regs(2157), 
                           B2 => n220, ZN => n1267);
   U1768 : NAND2_X1 port map( A1 => n1269, A2 => n1270, ZN => 
                           curr_proc_regs(108));
   U1769 : AOI222_X1 port map( A1 => regs(108), A2 => n1, B1 => regs(1644), B2 
                           => n53, C1 => regs(620), C2 => n105, ZN => n1270);
   U1770 : AOI22_X1 port map( A1 => regs(1132), A2 => n157, B1 => regs(2156), 
                           B2 => n220, ZN => n1269);
   U1771 : NAND2_X1 port map( A1 => n1271, A2 => n1272, ZN => 
                           curr_proc_regs(107));
   U1772 : AOI222_X1 port map( A1 => regs(107), A2 => n1, B1 => regs(1643), B2 
                           => n53, C1 => regs(619), C2 => n105, ZN => n1272);
   U1773 : AOI22_X1 port map( A1 => regs(1131), A2 => n157, B1 => regs(2155), 
                           B2 => n220, ZN => n1271);
   U1774 : NAND2_X1 port map( A1 => n1273, A2 => n1274, ZN => 
                           curr_proc_regs(106));
   U1775 : AOI222_X1 port map( A1 => regs(106), A2 => n1, B1 => regs(1642), B2 
                           => n53, C1 => regs(618), C2 => n105, ZN => n1274);
   U1776 : AOI22_X1 port map( A1 => regs(1130), A2 => n157, B1 => regs(2154), 
                           B2 => n220, ZN => n1273);
   U1777 : NAND2_X1 port map( A1 => n1275, A2 => n1276, ZN => 
                           curr_proc_regs(105));
   U1778 : AOI222_X1 port map( A1 => regs(105), A2 => n1, B1 => regs(1641), B2 
                           => n53, C1 => regs(617), C2 => n105, ZN => n1276);
   U1779 : AOI22_X1 port map( A1 => regs(1129), A2 => n157, B1 => regs(2153), 
                           B2 => n220, ZN => n1275);
   U1780 : NAND2_X1 port map( A1 => n1277, A2 => n1278, ZN => 
                           curr_proc_regs(104));
   U1781 : AOI222_X1 port map( A1 => regs(104), A2 => n1, B1 => regs(1640), B2 
                           => n53, C1 => regs(616), C2 => n105, ZN => n1278);
   U1782 : AOI22_X1 port map( A1 => regs(1128), A2 => n157, B1 => regs(2152), 
                           B2 => n220, ZN => n1277);
   U1783 : NAND2_X1 port map( A1 => n1279, A2 => n1280, ZN => 
                           curr_proc_regs(103));
   U1784 : AOI222_X1 port map( A1 => regs(103), A2 => n1, B1 => regs(1639), B2 
                           => n53, C1 => regs(615), C2 => n105, ZN => n1280);
   U1785 : AOI22_X1 port map( A1 => regs(1127), A2 => n157, B1 => regs(2151), 
                           B2 => n220, ZN => n1279);
   U1786 : NAND2_X1 port map( A1 => n1281, A2 => n1282, ZN => 
                           curr_proc_regs(102));
   U1787 : AOI222_X1 port map( A1 => regs(102), A2 => n1, B1 => regs(1638), B2 
                           => n53, C1 => regs(614), C2 => n105, ZN => n1282);
   U1788 : AOI22_X1 port map( A1 => regs(1126), A2 => n157, B1 => regs(2150), 
                           B2 => n219, ZN => n1281);
   U1789 : NAND2_X1 port map( A1 => n1283, A2 => n1284, ZN => 
                           curr_proc_regs(101));
   U1790 : AOI222_X1 port map( A1 => regs(101), A2 => n1, B1 => regs(1637), B2 
                           => n53, C1 => regs(613), C2 => n105, ZN => n1284);
   U1791 : AOI22_X1 port map( A1 => regs(1125), A2 => n157, B1 => regs(2149), 
                           B2 => n219, ZN => n1283);
   U1792 : NAND2_X1 port map( A1 => n1285, A2 => n1286, ZN => 
                           curr_proc_regs(100));
   U1793 : AOI222_X1 port map( A1 => regs(100), A2 => n1, B1 => regs(1636), B2 
                           => n53, C1 => regs(612), C2 => n105, ZN => n1286);
   U1794 : AOI22_X1 port map( A1 => regs(1124), A2 => n157, B1 => regs(2148), 
                           B2 => n225, ZN => n1285);
   U1795 : NAND2_X1 port map( A1 => n1287, A2 => n1288, ZN => curr_proc_regs(0)
                           );
   U1796 : AOI222_X1 port map( A1 => regs(0), A2 => n1, B1 => regs(1536), B2 =>
                           n53, C1 => regs(512), C2 => n105, ZN => n1288);
   U1797 : AND3_X1 port map( A1 => n1289, A2 => n1290, A3 => win(1), ZN => n265
                           );
   U1798 : NOR2_X1 port map( A1 => n1291, A2 => n209, ZN => n264);
   U1799 : INV_X1 port map( A => win(3), ZN => n1291);
   U1800 : AND4_X1 port map( A1 => win(0), A2 => n1289, A3 => n1292, A4 => 
                           n1290, ZN => n263);
   U1801 : INV_X1 port map( A => win(2), ZN => n1290);
   U1802 : INV_X1 port map( A => win(1), ZN => n1292);
   U1803 : AOI22_X1 port map( A1 => regs(1024), A2 => n157, B1 => regs(2048), 
                           B2 => n209, ZN => n1287);
   U1804 : AND2_X1 port map( A1 => win(2), A2 => n1289, ZN => n266);
   U1805 : NOR2_X1 port map( A1 => win(3), A2 => n209, ZN => n1289);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity equal_check_N5_0 is

   port( A, B : in std_logic_vector (4 downto 0);  EQUAL : out std_logic);

end equal_check_N5_0;

architecture SYN_behav of equal_check_N5_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NOR3_X1 port map( A1 => n1, A2 => n2, A3 => n3, ZN => EQUAL);
   U2 : XOR2_X1 port map( A => B(4), B => A(4), Z => n3);
   U3 : XOR2_X1 port map( A => B(2), B => A(2), Z => n2);
   U4 : NAND3_X1 port map( A1 => n4, A2 => n5, A3 => n6, ZN => n1);
   U5 : XNOR2_X1 port map( A => B(0), B => A(0), ZN => n6);
   U6 : XNOR2_X1 port map( A => B(1), B => A(1), ZN => n5);
   U7 : XNOR2_X1 port map( A => B(3), B => A(3), ZN => n4);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity connection_mtx_M8_N8_F5 is

   port( dec : in std_logic_vector (31 downto 0);  addr_pop : in 
         std_logic_vector (15 downto 0);  win, swp : in std_logic_vector (4 
         downto 0);  sel : out std_logic_vector (87 downto 0));

end connection_mtx_M8_N8_F5;

architecture SYN_struct of connection_mtx_M8_N8_F5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal sel_87_port, sel_86_port, sel_85_port, sel_84_port, sel_83_port, 
      sel_82_port, sel_81_port, sel_80_port, sel_79_port, sel_78_port, 
      sel_77_port, sel_76_port, sel_75_port, sel_74_port, sel_73_port, 
      sel_72_port, sel_71_port, sel_70_port, sel_69_port, sel_68_port, 
      sel_67_port, sel_66_port, sel_65_port, sel_64_port, sel_63_port, 
      sel_62_port, sel_61_port, sel_60_port, sel_59_port, sel_58_port, 
      sel_57_port, sel_56_port, sel_55_port, sel_54_port, sel_53_port, 
      sel_52_port, sel_51_port, sel_50_port, sel_49_port, sel_48_port, 
      sel_47_port, sel_46_port, sel_45_port, sel_44_port, sel_43_port, 
      sel_42_port, sel_41_port, sel_40_port, sel_39_port, sel_38_port, 
      sel_37_port, sel_36_port, sel_35_port, sel_34_port, sel_33_port, 
      sel_32_port, sel_31_port, sel_30_port, sel_29_port, sel_28_port, 
      sel_27_port, sel_26_port, sel_25_port, sel_24_port, sel_23_port, 
      sel_22_port, sel_21_port, sel_20_port, sel_19_port, sel_18_port, 
      sel_17_port, sel_16_port, sel_15_port, sel_14_port, sel_13_port, 
      sel_12_port, sel_11_port, sel_10_port, sel_9_port, sel_8_port, n1, n2, n3
      , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50 : std_logic;

begin
   sel <= ( sel_87_port, sel_86_port, sel_85_port, sel_84_port, sel_83_port, 
      sel_82_port, sel_81_port, sel_80_port, sel_79_port, sel_78_port, 
      sel_77_port, sel_76_port, sel_75_port, sel_74_port, sel_73_port, 
      sel_72_port, sel_71_port, sel_70_port, sel_69_port, sel_68_port, 
      sel_67_port, sel_66_port, sel_65_port, sel_64_port, sel_63_port, 
      sel_62_port, sel_61_port, sel_60_port, sel_59_port, sel_58_port, 
      sel_57_port, sel_56_port, sel_55_port, sel_54_port, sel_53_port, 
      sel_52_port, sel_51_port, sel_50_port, sel_49_port, sel_48_port, 
      sel_47_port, sel_46_port, sel_45_port, sel_44_port, sel_43_port, 
      sel_42_port, sel_41_port, sel_40_port, sel_39_port, sel_38_port, 
      sel_37_port, sel_36_port, sel_35_port, sel_34_port, sel_33_port, 
      sel_32_port, sel_31_port, sel_30_port, sel_29_port, sel_28_port, 
      sel_27_port, sel_26_port, sel_25_port, sel_24_port, sel_23_port, 
      sel_22_port, sel_21_port, sel_20_port, sel_19_port, sel_18_port, 
      sel_17_port, sel_16_port, sel_15_port, sel_14_port, sel_13_port, 
      sel_12_port, sel_11_port, sel_10_port, sel_9_port, sel_8_port, dec(7), 
      dec(6), dec(5), dec(4), dec(3), dec(2), dec(1), dec(0) );
   
   U1 : INV_X1 port map( A => swp(4), ZN => n1);
   U2 : INV_X1 port map( A => swp(3), ZN => n2);
   U3 : INV_X1 port map( A => swp(2), ZN => n3);
   U4 : INV_X1 port map( A => swp(1), ZN => n4);
   U5 : INV_X1 port map( A => swp(0), ZN => n5);
   U6 : OAI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n5, C1 => n9, 
                           C2 => n10, ZN => sel_9_port);
   U7 : OAI222_X1 port map( A1 => n7, A2 => n11, B1 => n5, B2 => n12, C1 => n10
                           , C2 => n13, ZN => sel_8_port);
   U8 : OAI22_X1 port map( A1 => n7, A2 => n14, B1 => n15, B2 => n1, ZN => 
                           sel_87_port);
   U9 : OAI22_X1 port map( A1 => n7, A2 => n16, B1 => n1, B2 => n17, ZN => 
                           sel_86_port);
   U10 : OAI22_X1 port map( A1 => n7, A2 => n18, B1 => n1, B2 => n19, ZN => 
                           sel_85_port);
   U11 : OAI22_X1 port map( A1 => n7, A2 => n20, B1 => n1, B2 => n21, ZN => 
                           sel_84_port);
   U12 : OAI22_X1 port map( A1 => n7, A2 => n22, B1 => n1, B2 => n23, ZN => 
                           sel_83_port);
   U13 : OAI22_X1 port map( A1 => n7, A2 => n24, B1 => n1, B2 => n25, ZN => 
                           sel_82_port);
   U14 : OAI22_X1 port map( A1 => n7, A2 => n26, B1 => n1, B2 => n27, ZN => 
                           sel_81_port);
   U15 : OAI22_X1 port map( A1 => n7, A2 => n28, B1 => n1, B2 => n29, ZN => 
                           sel_80_port);
   U16 : OAI222_X1 port map( A1 => n7, A2 => n30, B1 => n1, B2 => n31, C1 => 
                           n32, C2 => n33, ZN => sel_79_port);
   U17 : OAI222_X1 port map( A1 => n7, A2 => n34, B1 => n1, B2 => n35, C1 => 
                           n33, C2 => n36, ZN => sel_78_port);
   U18 : OAI222_X1 port map( A1 => n7, A2 => n37, B1 => n1, B2 => n38, C1 => 
                           n33, C2 => n39, ZN => sel_77_port);
   U19 : OAI222_X1 port map( A1 => n7, A2 => n40, B1 => n1, B2 => n41, C1 => 
                           n33, C2 => n42, ZN => sel_76_port);
   U20 : OAI222_X1 port map( A1 => n7, A2 => n43, B1 => n1, B2 => n44, C1 => 
                           n33, C2 => n45, ZN => sel_75_port);
   U21 : OAI222_X1 port map( A1 => n7, A2 => n46, B1 => n1, B2 => n47, C1 => 
                           n33, C2 => n48, ZN => sel_74_port);
   U22 : OAI222_X1 port map( A1 => n6, A2 => n33, B1 => n8, B2 => n1, C1 => n7,
                           C2 => n9, ZN => sel_73_port);
   U23 : OAI222_X1 port map( A1 => n11, A2 => n33, B1 => n12, B2 => n1, C1 => 
                           n7, C2 => n13, ZN => sel_72_port);
   U24 : OAI22_X1 port map( A1 => n14, A2 => n33, B1 => n15, B2 => n2, ZN => 
                           sel_71_port);
   U25 : OAI22_X1 port map( A1 => n16, A2 => n33, B1 => n17, B2 => n2, ZN => 
                           sel_70_port);
   U26 : OAI22_X1 port map( A1 => n18, A2 => n33, B1 => n19, B2 => n2, ZN => 
                           sel_69_port);
   U27 : OAI22_X1 port map( A1 => n20, A2 => n33, B1 => n21, B2 => n2, ZN => 
                           sel_68_port);
   U28 : OAI22_X1 port map( A1 => n22, A2 => n33, B1 => n23, B2 => n2, ZN => 
                           sel_67_port);
   U29 : OAI22_X1 port map( A1 => n24, A2 => n33, B1 => n25, B2 => n2, ZN => 
                           sel_66_port);
   U30 : OAI22_X1 port map( A1 => n26, A2 => n33, B1 => n27, B2 => n2, ZN => 
                           sel_65_port);
   U31 : OAI22_X1 port map( A1 => n28, A2 => n33, B1 => n29, B2 => n2, ZN => 
                           sel_64_port);
   U32 : OAI222_X1 port map( A1 => n30, A2 => n33, B1 => n31, B2 => n2, C1 => 
                           n32, C2 => n49, ZN => sel_63_port);
   U33 : OAI222_X1 port map( A1 => n33, A2 => n34, B1 => n35, B2 => n2, C1 => 
                           n36, C2 => n49, ZN => sel_62_port);
   U34 : OAI222_X1 port map( A1 => n33, A2 => n37, B1 => n38, B2 => n2, C1 => 
                           n39, C2 => n49, ZN => sel_61_port);
   U35 : OAI222_X1 port map( A1 => n33, A2 => n40, B1 => n41, B2 => n2, C1 => 
                           n42, C2 => n49, ZN => sel_60_port);
   U36 : OAI222_X1 port map( A1 => n33, A2 => n43, B1 => n44, B2 => n2, C1 => 
                           n45, C2 => n49, ZN => sel_59_port);
   U37 : OAI222_X1 port map( A1 => n33, A2 => n46, B1 => n47, B2 => n2, C1 => 
                           n48, C2 => n49, ZN => sel_58_port);
   U38 : OAI222_X1 port map( A1 => n6, A2 => n49, B1 => n8, B2 => n2, C1 => n9,
                           C2 => n33, ZN => sel_57_port);
   U39 : OAI222_X1 port map( A1 => n11, A2 => n49, B1 => n12, B2 => n2, C1 => 
                           n13, C2 => n33, ZN => sel_56_port);
   U40 : INV_X1 port map( A => win(3), ZN => n33);
   U41 : OAI22_X1 port map( A1 => n14, A2 => n49, B1 => n15, B2 => n3, ZN => 
                           sel_55_port);
   U42 : OAI22_X1 port map( A1 => n16, A2 => n49, B1 => n17, B2 => n3, ZN => 
                           sel_54_port);
   U43 : OAI22_X1 port map( A1 => n18, A2 => n49, B1 => n19, B2 => n3, ZN => 
                           sel_53_port);
   U44 : OAI22_X1 port map( A1 => n20, A2 => n49, B1 => n21, B2 => n3, ZN => 
                           sel_52_port);
   U45 : OAI22_X1 port map( A1 => n22, A2 => n49, B1 => n23, B2 => n3, ZN => 
                           sel_51_port);
   U46 : OAI22_X1 port map( A1 => n24, A2 => n49, B1 => n25, B2 => n3, ZN => 
                           sel_50_port);
   U47 : OAI22_X1 port map( A1 => n26, A2 => n49, B1 => n27, B2 => n3, ZN => 
                           sel_49_port);
   U48 : OAI22_X1 port map( A1 => n28, A2 => n49, B1 => n29, B2 => n3, ZN => 
                           sel_48_port);
   U49 : OAI222_X1 port map( A1 => n30, A2 => n49, B1 => n31, B2 => n3, C1 => 
                           n32, C2 => n50, ZN => sel_47_port);
   U50 : OAI222_X1 port map( A1 => n34, A2 => n49, B1 => n35, B2 => n3, C1 => 
                           n36, C2 => n50, ZN => sel_46_port);
   U51 : OAI222_X1 port map( A1 => n37, A2 => n49, B1 => n38, B2 => n3, C1 => 
                           n39, C2 => n50, ZN => sel_45_port);
   U52 : OAI222_X1 port map( A1 => n40, A2 => n49, B1 => n41, B2 => n3, C1 => 
                           n42, C2 => n50, ZN => sel_44_port);
   U53 : OAI222_X1 port map( A1 => n43, A2 => n49, B1 => n44, B2 => n3, C1 => 
                           n45, C2 => n50, ZN => sel_43_port);
   U54 : OAI222_X1 port map( A1 => n46, A2 => n49, B1 => n47, B2 => n3, C1 => 
                           n48, C2 => n50, ZN => sel_42_port);
   U55 : OAI222_X1 port map( A1 => n6, A2 => n50, B1 => n8, B2 => n3, C1 => n9,
                           C2 => n49, ZN => sel_41_port);
   U56 : OAI222_X1 port map( A1 => n11, A2 => n50, B1 => n12, B2 => n3, C1 => 
                           n13, C2 => n49, ZN => sel_40_port);
   U57 : INV_X1 port map( A => win(2), ZN => n49);
   U58 : OAI22_X1 port map( A1 => n14, A2 => n50, B1 => n15, B2 => n4, ZN => 
                           sel_39_port);
   U59 : OAI22_X1 port map( A1 => n16, A2 => n50, B1 => n17, B2 => n4, ZN => 
                           sel_38_port);
   U60 : OAI22_X1 port map( A1 => n18, A2 => n50, B1 => n19, B2 => n4, ZN => 
                           sel_37_port);
   U61 : OAI22_X1 port map( A1 => n20, A2 => n50, B1 => n21, B2 => n4, ZN => 
                           sel_36_port);
   U62 : OAI22_X1 port map( A1 => n22, A2 => n50, B1 => n23, B2 => n4, ZN => 
                           sel_35_port);
   U63 : OAI22_X1 port map( A1 => n24, A2 => n50, B1 => n25, B2 => n4, ZN => 
                           sel_34_port);
   U64 : OAI22_X1 port map( A1 => n26, A2 => n50, B1 => n27, B2 => n4, ZN => 
                           sel_33_port);
   U65 : OAI22_X1 port map( A1 => n28, A2 => n50, B1 => n29, B2 => n4, ZN => 
                           sel_32_port);
   U66 : OAI222_X1 port map( A1 => n30, A2 => n50, B1 => n31, B2 => n4, C1 => 
                           n10, C2 => n32, ZN => sel_31_port);
   U67 : OAI222_X1 port map( A1 => n34, A2 => n50, B1 => n35, B2 => n4, C1 => 
                           n10, C2 => n36, ZN => sel_30_port);
   U68 : OAI222_X1 port map( A1 => n37, A2 => n50, B1 => n38, B2 => n4, C1 => 
                           n10, C2 => n39, ZN => sel_29_port);
   U69 : OAI222_X1 port map( A1 => n40, A2 => n50, B1 => n41, B2 => n4, C1 => 
                           n10, C2 => n42, ZN => sel_28_port);
   U70 : OAI222_X1 port map( A1 => n43, A2 => n50, B1 => n44, B2 => n4, C1 => 
                           n10, C2 => n45, ZN => sel_27_port);
   U71 : OAI222_X1 port map( A1 => n46, A2 => n50, B1 => n47, B2 => n4, C1 => 
                           n10, C2 => n48, ZN => sel_26_port);
   U72 : OAI222_X1 port map( A1 => n6, A2 => n10, B1 => n8, B2 => n4, C1 => n9,
                           C2 => n50, ZN => sel_25_port);
   U73 : INV_X1 port map( A => dec(9), ZN => n9);
   U74 : INV_X1 port map( A => addr_pop(14), ZN => n8);
   U75 : INV_X1 port map( A => dec(25), ZN => n6);
   U76 : OAI222_X1 port map( A1 => n10, A2 => n11, B1 => n12, B2 => n4, C1 => 
                           n13, C2 => n50, ZN => sel_24_port);
   U77 : INV_X1 port map( A => win(1), ZN => n50);
   U78 : INV_X1 port map( A => dec(8), ZN => n13);
   U79 : INV_X1 port map( A => addr_pop(15), ZN => n12);
   U80 : INV_X1 port map( A => dec(24), ZN => n11);
   U81 : OAI22_X1 port map( A1 => n10, A2 => n14, B1 => n5, B2 => n15, ZN => 
                           sel_23_port);
   U82 : INV_X1 port map( A => addr_pop(0), ZN => n15);
   U83 : INV_X1 port map( A => dec(23), ZN => n14);
   U84 : OAI22_X1 port map( A1 => n10, A2 => n16, B1 => n5, B2 => n17, ZN => 
                           sel_22_port);
   U85 : INV_X1 port map( A => addr_pop(1), ZN => n17);
   U86 : INV_X1 port map( A => dec(22), ZN => n16);
   U87 : OAI22_X1 port map( A1 => n10, A2 => n18, B1 => n5, B2 => n19, ZN => 
                           sel_21_port);
   U88 : INV_X1 port map( A => addr_pop(2), ZN => n19);
   U89 : INV_X1 port map( A => dec(21), ZN => n18);
   U90 : OAI22_X1 port map( A1 => n10, A2 => n20, B1 => n5, B2 => n21, ZN => 
                           sel_20_port);
   U91 : INV_X1 port map( A => addr_pop(3), ZN => n21);
   U92 : INV_X1 port map( A => dec(20), ZN => n20);
   U93 : OAI22_X1 port map( A1 => n10, A2 => n22, B1 => n5, B2 => n23, ZN => 
                           sel_19_port);
   U94 : INV_X1 port map( A => addr_pop(4), ZN => n23);
   U95 : INV_X1 port map( A => dec(19), ZN => n22);
   U96 : OAI22_X1 port map( A1 => n10, A2 => n24, B1 => n5, B2 => n25, ZN => 
                           sel_18_port);
   U97 : INV_X1 port map( A => addr_pop(5), ZN => n25);
   U98 : INV_X1 port map( A => dec(18), ZN => n24);
   U99 : OAI22_X1 port map( A1 => n10, A2 => n26, B1 => n5, B2 => n27, ZN => 
                           sel_17_port);
   U100 : INV_X1 port map( A => addr_pop(6), ZN => n27);
   U101 : INV_X1 port map( A => dec(17), ZN => n26);
   U102 : OAI22_X1 port map( A1 => n10, A2 => n28, B1 => n5, B2 => n29, ZN => 
                           sel_16_port);
   U103 : INV_X1 port map( A => addr_pop(7), ZN => n29);
   U104 : INV_X1 port map( A => dec(16), ZN => n28);
   U105 : OAI222_X1 port map( A1 => n10, A2 => n30, B1 => n5, B2 => n31, C1 => 
                           n7, C2 => n32, ZN => sel_15_port);
   U106 : INV_X1 port map( A => dec(31), ZN => n32);
   U107 : INV_X1 port map( A => addr_pop(8), ZN => n31);
   U108 : INV_X1 port map( A => dec(15), ZN => n30);
   U109 : OAI222_X1 port map( A1 => n10, A2 => n34, B1 => n5, B2 => n35, C1 => 
                           n7, C2 => n36, ZN => sel_14_port);
   U110 : INV_X1 port map( A => dec(30), ZN => n36);
   U111 : INV_X1 port map( A => addr_pop(9), ZN => n35);
   U112 : INV_X1 port map( A => dec(14), ZN => n34);
   U113 : OAI222_X1 port map( A1 => n10, A2 => n37, B1 => n5, B2 => n38, C1 => 
                           n7, C2 => n39, ZN => sel_13_port);
   U114 : INV_X1 port map( A => dec(29), ZN => n39);
   U115 : INV_X1 port map( A => addr_pop(10), ZN => n38);
   U116 : INV_X1 port map( A => dec(13), ZN => n37);
   U117 : OAI222_X1 port map( A1 => n10, A2 => n40, B1 => n5, B2 => n41, C1 => 
                           n7, C2 => n42, ZN => sel_12_port);
   U118 : INV_X1 port map( A => dec(28), ZN => n42);
   U119 : INV_X1 port map( A => addr_pop(11), ZN => n41);
   U120 : INV_X1 port map( A => dec(12), ZN => n40);
   U121 : OAI222_X1 port map( A1 => n10, A2 => n43, B1 => n5, B2 => n44, C1 => 
                           n7, C2 => n45, ZN => sel_11_port);
   U122 : INV_X1 port map( A => dec(27), ZN => n45);
   U123 : INV_X1 port map( A => addr_pop(12), ZN => n44);
   U124 : INV_X1 port map( A => dec(11), ZN => n43);
   U125 : OAI222_X1 port map( A1 => n10, A2 => n46, B1 => n5, B2 => n47, C1 => 
                           n7, C2 => n48, ZN => sel_10_port);
   U126 : INV_X1 port map( A => dec(26), ZN => n48);
   U127 : INV_X1 port map( A => win(4), ZN => n7);
   U128 : INV_X1 port map( A => addr_pop(13), ZN => n47);
   U129 : INV_X1 port map( A => dec(10), ZN => n46);
   U130 : INV_X1 port map( A => win(0), ZN => n10);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity decoder_N5 is

   port( Q : in std_logic_vector (4 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end decoder_N5;

architecture SYN_Behavioural of decoder_N5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => Y(0));
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => Y(1));
   U3 : NOR2_X1 port map( A1 => n1, A2 => n4, ZN => Y(2));
   U4 : NOR2_X1 port map( A1 => n1, A2 => n5, ZN => Y(3));
   U5 : NOR2_X1 port map( A1 => n1, A2 => n6, ZN => Y(4));
   U6 : NOR2_X1 port map( A1 => n1, A2 => n7, ZN => Y(5));
   U7 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => Y(6));
   U8 : NOR2_X1 port map( A1 => n1, A2 => n9, ZN => Y(7));
   U9 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => n1);
   U10 : NOR2_X1 port map( A1 => n2, A2 => n12, ZN => Y(8));
   U11 : NOR2_X1 port map( A1 => n3, A2 => n12, ZN => Y(9));
   U12 : NOR2_X1 port map( A1 => n4, A2 => n12, ZN => Y(10));
   U13 : NOR2_X1 port map( A1 => n5, A2 => n12, ZN => Y(11));
   U14 : NOR2_X1 port map( A1 => n6, A2 => n12, ZN => Y(12));
   U15 : NOR2_X1 port map( A1 => n7, A2 => n12, ZN => Y(13));
   U16 : NOR2_X1 port map( A1 => n8, A2 => n12, ZN => Y(14));
   U17 : NOR2_X1 port map( A1 => n9, A2 => n12, ZN => Y(15));
   U18 : NAND2_X1 port map( A1 => Q(3), A2 => n10, ZN => n12);
   U19 : INV_X1 port map( A => Q(4), ZN => n10);
   U20 : NOR2_X1 port map( A1 => n2, A2 => n13, ZN => Y(16));
   U21 : NOR2_X1 port map( A1 => n3, A2 => n13, ZN => Y(17));
   U22 : NOR2_X1 port map( A1 => n4, A2 => n13, ZN => Y(18));
   U23 : NOR2_X1 port map( A1 => n5, A2 => n13, ZN => Y(19));
   U24 : NOR2_X1 port map( A1 => n6, A2 => n13, ZN => Y(20));
   U25 : NOR2_X1 port map( A1 => n7, A2 => n13, ZN => Y(21));
   U26 : NOR2_X1 port map( A1 => n8, A2 => n13, ZN => Y(22));
   U27 : NOR2_X1 port map( A1 => n9, A2 => n13, ZN => Y(23));
   U28 : NAND2_X1 port map( A1 => Q(4), A2 => n11, ZN => n13);
   U29 : INV_X1 port map( A => Q(3), ZN => n11);
   U30 : NOR2_X1 port map( A1 => n2, A2 => n14, ZN => Y(24));
   U31 : NAND3_X1 port map( A1 => n15, A2 => n16, A3 => n17, ZN => n2);
   U32 : NOR2_X1 port map( A1 => n3, A2 => n14, ZN => Y(25));
   U33 : NAND3_X1 port map( A1 => n15, A2 => n16, A3 => Q(0), ZN => n3);
   U34 : NOR2_X1 port map( A1 => n4, A2 => n14, ZN => Y(26));
   U35 : NAND3_X1 port map( A1 => n17, A2 => n16, A3 => Q(1), ZN => n4);
   U36 : NOR2_X1 port map( A1 => n5, A2 => n14, ZN => Y(27));
   U37 : NAND3_X1 port map( A1 => Q(0), A2 => n16, A3 => Q(1), ZN => n5);
   U38 : INV_X1 port map( A => Q(2), ZN => n16);
   U39 : NOR2_X1 port map( A1 => n6, A2 => n14, ZN => Y(28));
   U40 : NAND3_X1 port map( A1 => n17, A2 => n15, A3 => Q(2), ZN => n6);
   U41 : NOR2_X1 port map( A1 => n7, A2 => n14, ZN => Y(29));
   U42 : NAND3_X1 port map( A1 => Q(0), A2 => n15, A3 => Q(2), ZN => n7);
   U43 : INV_X1 port map( A => Q(1), ZN => n15);
   U44 : NOR2_X1 port map( A1 => n8, A2 => n14, ZN => Y(30));
   U45 : NAND3_X1 port map( A1 => Q(1), A2 => n17, A3 => Q(2), ZN => n8);
   U46 : INV_X1 port map( A => Q(0), ZN => n17);
   U47 : NOR2_X1 port map( A1 => n9, A2 => n14, ZN => Y(31));
   U48 : NAND2_X1 port map( A1 => Q(4), A2 => Q(3), ZN => n14);
   U49 : NAND3_X1 port map( A1 => Q(1), A2 => Q(0), A3 => Q(2), ZN => n9);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M1_0 is

   port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
         std_logic_vector (31 downto 0));

end mux_N32_M1_0;

architecture SYN_behav of mux_N32_M1_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => S, Z => n2);
   U3 : BUF_X1 port map( A => S, Z => n1);
   U4 : BUF_X1 port map( A => S, Z => n3);
   U5 : MUX2_X1 port map( A => Q(9), B => Q(41), S => n1, Z => Y(9));
   U6 : MUX2_X1 port map( A => Q(8), B => Q(40), S => n1, Z => Y(8));
   U7 : MUX2_X1 port map( A => Q(7), B => Q(39), S => n1, Z => Y(7));
   U8 : MUX2_X1 port map( A => Q(6), B => Q(38), S => n1, Z => Y(6));
   U9 : MUX2_X1 port map( A => Q(5), B => Q(37), S => n1, Z => Y(5));
   U10 : MUX2_X1 port map( A => Q(4), B => Q(36), S => n1, Z => Y(4));
   U11 : MUX2_X1 port map( A => Q(3), B => Q(35), S => n1, Z => Y(3));
   U12 : MUX2_X1 port map( A => Q(31), B => Q(63), S => n1, Z => Y(31));
   U13 : MUX2_X1 port map( A => Q(30), B => Q(62), S => n1, Z => Y(30));
   U14 : MUX2_X1 port map( A => Q(2), B => Q(34), S => n1, Z => Y(2));
   U15 : MUX2_X1 port map( A => Q(29), B => Q(61), S => n1, Z => Y(29));
   U16 : MUX2_X1 port map( A => Q(28), B => Q(60), S => n1, Z => Y(28));
   U17 : MUX2_X1 port map( A => Q(27), B => Q(59), S => n2, Z => Y(27));
   U18 : MUX2_X1 port map( A => Q(26), B => Q(58), S => n2, Z => Y(26));
   U19 : MUX2_X1 port map( A => Q(25), B => Q(57), S => n2, Z => Y(25));
   U20 : MUX2_X1 port map( A => Q(24), B => Q(56), S => n2, Z => Y(24));
   U21 : MUX2_X1 port map( A => Q(23), B => Q(55), S => n2, Z => Y(23));
   U22 : MUX2_X1 port map( A => Q(22), B => Q(54), S => n2, Z => Y(22));
   U23 : MUX2_X1 port map( A => Q(21), B => Q(53), S => n2, Z => Y(21));
   U24 : MUX2_X1 port map( A => Q(20), B => Q(52), S => n2, Z => Y(20));
   U25 : MUX2_X1 port map( A => Q(1), B => Q(33), S => n2, Z => Y(1));
   U26 : MUX2_X1 port map( A => Q(19), B => Q(51), S => n2, Z => Y(19));
   U27 : MUX2_X1 port map( A => Q(18), B => Q(50), S => n2, Z => Y(18));
   U28 : MUX2_X1 port map( A => Q(17), B => Q(49), S => n2, Z => Y(17));
   U29 : MUX2_X1 port map( A => Q(16), B => Q(48), S => n3, Z => Y(16));
   U30 : MUX2_X1 port map( A => Q(15), B => Q(47), S => n3, Z => Y(15));
   U31 : MUX2_X1 port map( A => Q(14), B => Q(46), S => n3, Z => Y(14));
   U32 : MUX2_X1 port map( A => Q(13), B => Q(45), S => n3, Z => Y(13));
   U33 : MUX2_X1 port map( A => Q(12), B => Q(44), S => n3, Z => Y(12));
   U34 : MUX2_X1 port map( A => Q(11), B => Q(43), S => n3, Z => Y(11));
   U35 : MUX2_X1 port map( A => Q(10), B => Q(42), S => n3, Z => Y(10));
   U36 : MUX2_X1 port map( A => Q(0), B => Q(32), S => n3, Z => Y(0));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N32_RSTVAL0_0 is

   port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector (31 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N32_RSTVAL0_0;

architecture SYN_Behavioural of reg_generic_N32_RSTVAL0_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   Q_reg_31_inst : DFF_X1 port map( D => n68, CK => Clk, Q => Q(31), QN => n67)
                           ;
   Q_reg_30_inst : DFF_X1 port map( D => n69, CK => Clk, Q => Q(30), QN => n66)
                           ;
   Q_reg_29_inst : DFF_X1 port map( D => n70, CK => Clk, Q => Q(29), QN => n65)
                           ;
   Q_reg_28_inst : DFF_X1 port map( D => n71, CK => Clk, Q => Q(28), QN => n64)
                           ;
   Q_reg_27_inst : DFF_X1 port map( D => n72, CK => Clk, Q => Q(27), QN => n63)
                           ;
   Q_reg_26_inst : DFF_X1 port map( D => n73, CK => Clk, Q => Q(26), QN => n62)
                           ;
   Q_reg_25_inst : DFF_X1 port map( D => n74, CK => Clk, Q => Q(25), QN => n61)
                           ;
   Q_reg_24_inst : DFF_X1 port map( D => n75, CK => Clk, Q => Q(24), QN => n60)
                           ;
   Q_reg_23_inst : DFF_X1 port map( D => n76, CK => Clk, Q => Q(23), QN => n59)
                           ;
   Q_reg_22_inst : DFF_X1 port map( D => n77, CK => Clk, Q => Q(22), QN => n58)
                           ;
   Q_reg_21_inst : DFF_X1 port map( D => n78, CK => Clk, Q => Q(21), QN => n57)
                           ;
   Q_reg_20_inst : DFF_X1 port map( D => n79, CK => Clk, Q => Q(20), QN => n56)
                           ;
   Q_reg_19_inst : DFF_X1 port map( D => n80, CK => Clk, Q => Q(19), QN => n55)
                           ;
   Q_reg_18_inst : DFF_X1 port map( D => n81, CK => Clk, Q => Q(18), QN => n54)
                           ;
   Q_reg_17_inst : DFF_X1 port map( D => n82, CK => Clk, Q => Q(17), QN => n53)
                           ;
   Q_reg_16_inst : DFF_X1 port map( D => n83, CK => Clk, Q => Q(16), QN => n52)
                           ;
   Q_reg_15_inst : DFF_X1 port map( D => n84, CK => Clk, Q => Q(15), QN => n51)
                           ;
   Q_reg_14_inst : DFF_X1 port map( D => n85, CK => Clk, Q => Q(14), QN => n50)
                           ;
   Q_reg_13_inst : DFF_X1 port map( D => n86, CK => Clk, Q => Q(13), QN => n49)
                           ;
   Q_reg_12_inst : DFF_X1 port map( D => n87, CK => Clk, Q => Q(12), QN => n48)
                           ;
   Q_reg_11_inst : DFF_X1 port map( D => n88, CK => Clk, Q => Q(11), QN => n47)
                           ;
   Q_reg_10_inst : DFF_X1 port map( D => n89, CK => Clk, Q => Q(10), QN => n46)
                           ;
   Q_reg_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => Q(9), QN => n45);
   Q_reg_8_inst : DFF_X1 port map( D => n91, CK => Clk, Q => Q(8), QN => n44);
   Q_reg_7_inst : DFF_X1 port map( D => n92, CK => Clk, Q => Q(7), QN => n43);
   Q_reg_6_inst : DFF_X1 port map( D => n93, CK => Clk, Q => Q(6), QN => n42);
   Q_reg_5_inst : DFF_X1 port map( D => n94, CK => Clk, Q => Q(5), QN => n41);
   Q_reg_4_inst : DFF_X1 port map( D => n95, CK => Clk, Q => Q(4), QN => n40);
   Q_reg_3_inst : DFF_X1 port map( D => n96, CK => Clk, Q => Q(3), QN => n39);
   Q_reg_2_inst : DFF_X1 port map( D => n97, CK => Clk, Q => Q(2), QN => n38);
   Q_reg_1_inst : DFF_X1 port map( D => n98, CK => Clk, Q => Q(1), QN => n37);
   Q_reg_0_inst : DFF_X1 port map( D => n99, CK => Clk, Q => Q(0), QN => n36);
   U3 : NAND2_X2 port map( A1 => n1, A2 => n35, ZN => n2);
   U4 : OR2_X2 port map( A1 => Rst, A2 => Enable, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n67, A2 => n1, B1 => n2, B2 => n3, ZN => n68);
   U6 : INV_X1 port map( A => D(31), ZN => n3);
   U7 : OAI22_X1 port map( A1 => n66, A2 => n1, B1 => n2, B2 => n4, ZN => n69);
   U8 : INV_X1 port map( A => D(30), ZN => n4);
   U9 : OAI22_X1 port map( A1 => n65, A2 => n1, B1 => n2, B2 => n5, ZN => n70);
   U10 : INV_X1 port map( A => D(29), ZN => n5);
   U11 : OAI22_X1 port map( A1 => n64, A2 => n1, B1 => n2, B2 => n6, ZN => n71)
                           ;
   U12 : INV_X1 port map( A => D(28), ZN => n6);
   U13 : OAI22_X1 port map( A1 => n63, A2 => n1, B1 => n2, B2 => n7, ZN => n72)
                           ;
   U14 : INV_X1 port map( A => D(27), ZN => n7);
   U15 : OAI22_X1 port map( A1 => n62, A2 => n1, B1 => n2, B2 => n8, ZN => n73)
                           ;
   U16 : INV_X1 port map( A => D(26), ZN => n8);
   U17 : OAI22_X1 port map( A1 => n61, A2 => n1, B1 => n2, B2 => n9, ZN => n74)
                           ;
   U18 : INV_X1 port map( A => D(25), ZN => n9);
   U19 : OAI22_X1 port map( A1 => n60, A2 => n1, B1 => n2, B2 => n10, ZN => n75
                           );
   U20 : INV_X1 port map( A => D(24), ZN => n10);
   U21 : OAI22_X1 port map( A1 => n59, A2 => n1, B1 => n2, B2 => n11, ZN => n76
                           );
   U22 : INV_X1 port map( A => D(23), ZN => n11);
   U23 : OAI22_X1 port map( A1 => n58, A2 => n1, B1 => n2, B2 => n12, ZN => n77
                           );
   U24 : INV_X1 port map( A => D(22), ZN => n12);
   U25 : OAI22_X1 port map( A1 => n57, A2 => n1, B1 => n2, B2 => n13, ZN => n78
                           );
   U26 : INV_X1 port map( A => D(21), ZN => n13);
   U27 : OAI22_X1 port map( A1 => n56, A2 => n1, B1 => n2, B2 => n14, ZN => n79
                           );
   U28 : INV_X1 port map( A => D(20), ZN => n14);
   U29 : OAI22_X1 port map( A1 => n55, A2 => n1, B1 => n2, B2 => n15, ZN => n80
                           );
   U30 : INV_X1 port map( A => D(19), ZN => n15);
   U31 : OAI22_X1 port map( A1 => n54, A2 => n1, B1 => n2, B2 => n16, ZN => n81
                           );
   U32 : INV_X1 port map( A => D(18), ZN => n16);
   U33 : OAI22_X1 port map( A1 => n53, A2 => n1, B1 => n2, B2 => n17, ZN => n82
                           );
   U34 : INV_X1 port map( A => D(17), ZN => n17);
   U35 : OAI22_X1 port map( A1 => n52, A2 => n1, B1 => n2, B2 => n18, ZN => n83
                           );
   U36 : INV_X1 port map( A => D(16), ZN => n18);
   U37 : OAI22_X1 port map( A1 => n51, A2 => n1, B1 => n2, B2 => n19, ZN => n84
                           );
   U38 : INV_X1 port map( A => D(15), ZN => n19);
   U39 : OAI22_X1 port map( A1 => n50, A2 => n1, B1 => n2, B2 => n20, ZN => n85
                           );
   U40 : INV_X1 port map( A => D(14), ZN => n20);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n1, B1 => n2, B2 => n21, ZN => n86
                           );
   U42 : INV_X1 port map( A => D(13), ZN => n21);
   U43 : OAI22_X1 port map( A1 => n48, A2 => n1, B1 => n2, B2 => n22, ZN => n87
                           );
   U44 : INV_X1 port map( A => D(12), ZN => n22);
   U45 : OAI22_X1 port map( A1 => n47, A2 => n1, B1 => n2, B2 => n23, ZN => n88
                           );
   U46 : INV_X1 port map( A => D(11), ZN => n23);
   U47 : OAI22_X1 port map( A1 => n46, A2 => n1, B1 => n2, B2 => n24, ZN => n89
                           );
   U48 : INV_X1 port map( A => D(10), ZN => n24);
   U49 : OAI22_X1 port map( A1 => n45, A2 => n1, B1 => n2, B2 => n25, ZN => n90
                           );
   U50 : INV_X1 port map( A => D(9), ZN => n25);
   U51 : OAI22_X1 port map( A1 => n44, A2 => n1, B1 => n2, B2 => n26, ZN => n91
                           );
   U52 : INV_X1 port map( A => D(8), ZN => n26);
   U53 : OAI22_X1 port map( A1 => n43, A2 => n1, B1 => n2, B2 => n27, ZN => n92
                           );
   U54 : INV_X1 port map( A => D(7), ZN => n27);
   U55 : OAI22_X1 port map( A1 => n42, A2 => n1, B1 => n2, B2 => n28, ZN => n93
                           );
   U56 : INV_X1 port map( A => D(6), ZN => n28);
   U57 : OAI22_X1 port map( A1 => n41, A2 => n1, B1 => n2, B2 => n29, ZN => n94
                           );
   U58 : INV_X1 port map( A => D(5), ZN => n29);
   U59 : OAI22_X1 port map( A1 => n40, A2 => n1, B1 => n2, B2 => n30, ZN => n95
                           );
   U60 : INV_X1 port map( A => D(4), ZN => n30);
   U61 : OAI22_X1 port map( A1 => n39, A2 => n1, B1 => n2, B2 => n31, ZN => n96
                           );
   U62 : INV_X1 port map( A => D(3), ZN => n31);
   U63 : OAI22_X1 port map( A1 => n38, A2 => n1, B1 => n2, B2 => n32, ZN => n97
                           );
   U64 : INV_X1 port map( A => D(2), ZN => n32);
   U65 : OAI22_X1 port map( A1 => n37, A2 => n1, B1 => n2, B2 => n33, ZN => n98
                           );
   U66 : INV_X1 port map( A => D(1), ZN => n33);
   U67 : OAI22_X1 port map( A1 => n36, A2 => n1, B1 => n2, B2 => n34, ZN => n99
                           );
   U68 : INV_X1 port map( A => D(0), ZN => n34);
   U69 : INV_X1 port map( A => Rst, ZN => n35);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity mux_N32_M5_0 is

   port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector (1023 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end mux_N32_M5_0;

architecture SYN_behav of mux_N32_M5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689 : 
      std_logic;

begin
   
   U2 : AND2_X2 port map( A1 => n661, A2 => n666, ZN => n16);
   U3 : AND2_X2 port map( A1 => n661, A2 => n664, ZN => n14);
   U4 : AND2_X2 port map( A1 => n663, A2 => n665, ZN => n12);
   U5 : AND2_X2 port map( A1 => n661, A2 => n662, ZN => n10);
   U6 : AND2_X2 port map( A1 => n666, A2 => n672, ZN => n22);
   U7 : AND2_X2 port map( A1 => n680, A2 => n665, ZN => n34);
   U8 : AND2_X2 port map( A1 => n662, A2 => n673, ZN => n28);
   U9 : AND2_X2 port map( A1 => n681, A2 => n664, ZN => n40);
   U10 : AND2_X2 port map( A1 => n665, A2 => n672, ZN => n26);
   U11 : AND2_X2 port map( A1 => n675, A2 => n664, ZN => n38);
   U12 : AND2_X2 port map( A1 => n681, A2 => n666, ZN => n52);
   U13 : AND2_X2 port map( A1 => n663, A2 => n662, ZN => n15);
   U14 : AND2_X2 port map( A1 => n662, A2 => n675, ZN => n46);
   U15 : AND2_X2 port map( A1 => n665, A2 => n673, ZN => n24);
   U16 : AND2_X2 port map( A1 => n680, A2 => n664, ZN => n36);
   U17 : AND2_X2 port map( A1 => n663, A2 => n666, ZN => n11);
   U18 : AND2_X2 port map( A1 => n682, A2 => n666, ZN => n50);
   U19 : AND2_X2 port map( A1 => n680, A2 => n662, ZN => n48);
   U20 : AND2_X2 port map( A1 => n661, A2 => n665, ZN => n13);
   U21 : AND2_X2 port map( A1 => n663, A2 => n664, ZN => n9);
   U22 : AND2_X2 port map( A1 => n664, A2 => n673, ZN => n21);
   U23 : AND2_X2 port map( A1 => n662, A2 => n672, ZN => n33);
   U24 : AND2_X2 port map( A1 => n675, A2 => n666, ZN => n27);
   U25 : AND2_X2 port map( A1 => n682, A2 => n665, ZN => n39);
   U26 : AND2_X2 port map( A1 => n682, A2 => n664, ZN => n45);
   U27 : AND2_X2 port map( A1 => n666, A2 => n673, ZN => n23);
   U28 : AND2_X2 port map( A1 => n675, A2 => n665, ZN => n35);
   U29 : AND2_X2 port map( A1 => n681, A2 => n662, ZN => n51);
   U30 : AND2_X2 port map( A1 => n672, A2 => n664, ZN => n25);
   U31 : AND2_X2 port map( A1 => n680, A2 => n666, ZN => n37);
   U32 : AND2_X2 port map( A1 => n682, A2 => n662, ZN => n49);
   U33 : AND2_X2 port map( A1 => n681, A2 => n665, ZN => n47);
   U34 : OR4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => Y(9));
   U35 : NAND4_X1 port map( A1 => n5, A2 => n6, A3 => n7, A4 => n8, ZN => n4);
   U36 : AOI22_X1 port map( A1 => Q(105), A2 => n9, B1 => Q(201), B2 => n10, ZN
                           => n8);
   U37 : AOI22_X1 port map( A1 => Q(169), A2 => n11, B1 => Q(41), B2 => n12, ZN
                           => n7);
   U38 : AOI22_X1 port map( A1 => Q(9), A2 => n13, B1 => Q(73), B2 => n14, ZN 
                           => n6);
   U39 : AOI22_X1 port map( A1 => Q(233), A2 => n15, B1 => Q(137), B2 => n16, 
                           ZN => n5);
   U40 : NAND4_X1 port map( A1 => n17, A2 => n18, A3 => n19, A4 => n20, ZN => 
                           n3);
   U41 : AOI22_X1 port map( A1 => Q(329), A2 => n21, B1 => Q(425), B2 => n22, 
                           ZN => n20);
   U42 : AOI22_X1 port map( A1 => Q(393), A2 => n23, B1 => Q(265), B2 => n24, 
                           ZN => n19);
   U43 : AOI22_X1 port map( A1 => Q(361), A2 => n25, B1 => Q(297), B2 => n26, 
                           ZN => n18);
   U44 : AOI22_X1 port map( A1 => Q(649), A2 => n27, B1 => Q(457), B2 => n28, 
                           ZN => n17);
   U45 : NAND4_X1 port map( A1 => n29, A2 => n30, A3 => n31, A4 => n32, ZN => 
                           n2);
   U46 : AOI22_X1 port map( A1 => Q(489), A2 => n33, B1 => Q(553), B2 => n34, 
                           ZN => n32);
   U47 : AOI22_X1 port map( A1 => Q(521), A2 => n35, B1 => Q(617), B2 => n36, 
                           ZN => n31);
   U48 : AOI22_X1 port map( A1 => Q(681), A2 => n37, B1 => Q(585), B2 => n38, 
                           ZN => n30);
   U49 : AOI22_X1 port map( A1 => Q(777), A2 => n39, B1 => Q(873), B2 => n40, 
                           ZN => n29);
   U50 : NAND4_X1 port map( A1 => n41, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           n1);
   U51 : AOI22_X1 port map( A1 => Q(841), A2 => n45, B1 => Q(713), B2 => n46, 
                           ZN => n44);
   U52 : AOI22_X1 port map( A1 => Q(809), A2 => n47, B1 => Q(745), B2 => n48, 
                           ZN => n43);
   U53 : AOI22_X1 port map( A1 => Q(969), A2 => n49, B1 => Q(905), B2 => n50, 
                           ZN => n42);
   U54 : AOI22_X1 port map( A1 => Q(1001), A2 => n51, B1 => Q(937), B2 => n52, 
                           ZN => n41);
   U55 : OR4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           Y(8));
   U56 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n56);
   U57 : AOI22_X1 port map( A1 => Q(104), A2 => n9, B1 => Q(200), B2 => n10, ZN
                           => n60);
   U58 : AOI22_X1 port map( A1 => Q(168), A2 => n11, B1 => Q(40), B2 => n12, ZN
                           => n59);
   U59 : AOI22_X1 port map( A1 => Q(8), A2 => n13, B1 => Q(72), B2 => n14, ZN 
                           => n58);
   U60 : AOI22_X1 port map( A1 => Q(232), A2 => n15, B1 => Q(136), B2 => n16, 
                           ZN => n57);
   U61 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           n55);
   U62 : AOI22_X1 port map( A1 => Q(328), A2 => n21, B1 => Q(424), B2 => n22, 
                           ZN => n64);
   U63 : AOI22_X1 port map( A1 => Q(392), A2 => n23, B1 => Q(264), B2 => n24, 
                           ZN => n63);
   U64 : AOI22_X1 port map( A1 => Q(360), A2 => n25, B1 => Q(296), B2 => n26, 
                           ZN => n62);
   U65 : AOI22_X1 port map( A1 => Q(648), A2 => n27, B1 => Q(456), B2 => n28, 
                           ZN => n61);
   U66 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           n54);
   U67 : AOI22_X1 port map( A1 => Q(488), A2 => n33, B1 => Q(552), B2 => n34, 
                           ZN => n68);
   U68 : AOI22_X1 port map( A1 => Q(520), A2 => n35, B1 => Q(616), B2 => n36, 
                           ZN => n67);
   U69 : AOI22_X1 port map( A1 => Q(680), A2 => n37, B1 => Q(584), B2 => n38, 
                           ZN => n66);
   U70 : AOI22_X1 port map( A1 => Q(776), A2 => n39, B1 => Q(872), B2 => n40, 
                           ZN => n65);
   U71 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n53);
   U72 : AOI22_X1 port map( A1 => Q(840), A2 => n45, B1 => Q(712), B2 => n46, 
                           ZN => n72);
   U73 : AOI22_X1 port map( A1 => Q(808), A2 => n47, B1 => Q(744), B2 => n48, 
                           ZN => n71);
   U74 : AOI22_X1 port map( A1 => Q(968), A2 => n49, B1 => Q(904), B2 => n50, 
                           ZN => n70);
   U75 : AOI22_X1 port map( A1 => Q(1000), A2 => n51, B1 => Q(936), B2 => n52, 
                           ZN => n69);
   U76 : OR4_X1 port map( A1 => n73, A2 => n74, A3 => n75, A4 => n76, ZN => 
                           Y(7));
   U77 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n79, A4 => n80, ZN => 
                           n76);
   U78 : AOI22_X1 port map( A1 => Q(103), A2 => n9, B1 => Q(199), B2 => n10, ZN
                           => n80);
   U79 : AOI22_X1 port map( A1 => Q(167), A2 => n11, B1 => Q(39), B2 => n12, ZN
                           => n79);
   U80 : AOI22_X1 port map( A1 => Q(7), A2 => n13, B1 => Q(71), B2 => n14, ZN 
                           => n78);
   U81 : AOI22_X1 port map( A1 => Q(231), A2 => n15, B1 => Q(135), B2 => n16, 
                           ZN => n77);
   U82 : NAND4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           n75);
   U83 : AOI22_X1 port map( A1 => Q(327), A2 => n21, B1 => Q(423), B2 => n22, 
                           ZN => n84);
   U84 : AOI22_X1 port map( A1 => Q(391), A2 => n23, B1 => Q(263), B2 => n24, 
                           ZN => n83);
   U85 : AOI22_X1 port map( A1 => Q(359), A2 => n25, B1 => Q(295), B2 => n26, 
                           ZN => n82);
   U86 : AOI22_X1 port map( A1 => Q(647), A2 => n27, B1 => Q(455), B2 => n28, 
                           ZN => n81);
   U87 : NAND4_X1 port map( A1 => n85, A2 => n86, A3 => n87, A4 => n88, ZN => 
                           n74);
   U88 : AOI22_X1 port map( A1 => Q(487), A2 => n33, B1 => Q(551), B2 => n34, 
                           ZN => n88);
   U89 : AOI22_X1 port map( A1 => Q(519), A2 => n35, B1 => Q(615), B2 => n36, 
                           ZN => n87);
   U90 : AOI22_X1 port map( A1 => Q(679), A2 => n37, B1 => Q(583), B2 => n38, 
                           ZN => n86);
   U91 : AOI22_X1 port map( A1 => Q(775), A2 => n39, B1 => Q(871), B2 => n40, 
                           ZN => n85);
   U92 : NAND4_X1 port map( A1 => n89, A2 => n90, A3 => n91, A4 => n92, ZN => 
                           n73);
   U93 : AOI22_X1 port map( A1 => Q(839), A2 => n45, B1 => Q(711), B2 => n46, 
                           ZN => n92);
   U94 : AOI22_X1 port map( A1 => Q(807), A2 => n47, B1 => Q(743), B2 => n48, 
                           ZN => n91);
   U95 : AOI22_X1 port map( A1 => Q(967), A2 => n49, B1 => Q(903), B2 => n50, 
                           ZN => n90);
   U96 : AOI22_X1 port map( A1 => Q(999), A2 => n51, B1 => Q(935), B2 => n52, 
                           ZN => n89);
   U97 : OR4_X1 port map( A1 => n93, A2 => n94, A3 => n95, A4 => n96, ZN => 
                           Y(6));
   U98 : NAND4_X1 port map( A1 => n97, A2 => n98, A3 => n99, A4 => n100, ZN => 
                           n96);
   U99 : AOI22_X1 port map( A1 => Q(102), A2 => n9, B1 => Q(198), B2 => n10, ZN
                           => n100);
   U100 : AOI22_X1 port map( A1 => Q(166), A2 => n11, B1 => Q(38), B2 => n12, 
                           ZN => n99);
   U101 : AOI22_X1 port map( A1 => Q(6), A2 => n13, B1 => Q(70), B2 => n14, ZN 
                           => n98);
   U102 : AOI22_X1 port map( A1 => Q(230), A2 => n15, B1 => Q(134), B2 => n16, 
                           ZN => n97);
   U103 : NAND4_X1 port map( A1 => n101, A2 => n102, A3 => n103, A4 => n104, ZN
                           => n95);
   U104 : AOI22_X1 port map( A1 => Q(326), A2 => n21, B1 => Q(422), B2 => n22, 
                           ZN => n104);
   U105 : AOI22_X1 port map( A1 => Q(390), A2 => n23, B1 => Q(262), B2 => n24, 
                           ZN => n103);
   U106 : AOI22_X1 port map( A1 => Q(358), A2 => n25, B1 => Q(294), B2 => n26, 
                           ZN => n102);
   U107 : AOI22_X1 port map( A1 => Q(646), A2 => n27, B1 => Q(454), B2 => n28, 
                           ZN => n101);
   U108 : NAND4_X1 port map( A1 => n105, A2 => n106, A3 => n107, A4 => n108, ZN
                           => n94);
   U109 : AOI22_X1 port map( A1 => Q(486), A2 => n33, B1 => Q(550), B2 => n34, 
                           ZN => n108);
   U110 : AOI22_X1 port map( A1 => Q(518), A2 => n35, B1 => Q(614), B2 => n36, 
                           ZN => n107);
   U111 : AOI22_X1 port map( A1 => Q(678), A2 => n37, B1 => Q(582), B2 => n38, 
                           ZN => n106);
   U112 : AOI22_X1 port map( A1 => Q(774), A2 => n39, B1 => Q(870), B2 => n40, 
                           ZN => n105);
   U113 : NAND4_X1 port map( A1 => n109, A2 => n110, A3 => n111, A4 => n112, ZN
                           => n93);
   U114 : AOI22_X1 port map( A1 => Q(838), A2 => n45, B1 => Q(710), B2 => n46, 
                           ZN => n112);
   U115 : AOI22_X1 port map( A1 => Q(806), A2 => n47, B1 => Q(742), B2 => n48, 
                           ZN => n111);
   U116 : AOI22_X1 port map( A1 => Q(966), A2 => n49, B1 => Q(902), B2 => n50, 
                           ZN => n110);
   U117 : AOI22_X1 port map( A1 => Q(998), A2 => n51, B1 => Q(934), B2 => n52, 
                           ZN => n109);
   U118 : OR4_X1 port map( A1 => n113, A2 => n114, A3 => n115, A4 => n116, ZN 
                           => Y(5));
   U119 : NAND4_X1 port map( A1 => n117, A2 => n118, A3 => n119, A4 => n120, ZN
                           => n116);
   U120 : AOI22_X1 port map( A1 => Q(101), A2 => n9, B1 => Q(197), B2 => n10, 
                           ZN => n120);
   U121 : AOI22_X1 port map( A1 => Q(165), A2 => n11, B1 => Q(37), B2 => n12, 
                           ZN => n119);
   U122 : AOI22_X1 port map( A1 => Q(5), A2 => n13, B1 => Q(69), B2 => n14, ZN 
                           => n118);
   U123 : AOI22_X1 port map( A1 => Q(229), A2 => n15, B1 => Q(133), B2 => n16, 
                           ZN => n117);
   U124 : NAND4_X1 port map( A1 => n121, A2 => n122, A3 => n123, A4 => n124, ZN
                           => n115);
   U125 : AOI22_X1 port map( A1 => Q(325), A2 => n21, B1 => Q(421), B2 => n22, 
                           ZN => n124);
   U126 : AOI22_X1 port map( A1 => Q(389), A2 => n23, B1 => Q(261), B2 => n24, 
                           ZN => n123);
   U127 : AOI22_X1 port map( A1 => Q(357), A2 => n25, B1 => Q(293), B2 => n26, 
                           ZN => n122);
   U128 : AOI22_X1 port map( A1 => Q(645), A2 => n27, B1 => Q(453), B2 => n28, 
                           ZN => n121);
   U129 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => n114);
   U130 : AOI22_X1 port map( A1 => Q(485), A2 => n33, B1 => Q(549), B2 => n34, 
                           ZN => n128);
   U131 : AOI22_X1 port map( A1 => Q(517), A2 => n35, B1 => Q(613), B2 => n36, 
                           ZN => n127);
   U132 : AOI22_X1 port map( A1 => Q(677), A2 => n37, B1 => Q(581), B2 => n38, 
                           ZN => n126);
   U133 : AOI22_X1 port map( A1 => Q(773), A2 => n39, B1 => Q(869), B2 => n40, 
                           ZN => n125);
   U134 : NAND4_X1 port map( A1 => n129, A2 => n130, A3 => n131, A4 => n132, ZN
                           => n113);
   U135 : AOI22_X1 port map( A1 => Q(837), A2 => n45, B1 => Q(709), B2 => n46, 
                           ZN => n132);
   U136 : AOI22_X1 port map( A1 => Q(805), A2 => n47, B1 => Q(741), B2 => n48, 
                           ZN => n131);
   U137 : AOI22_X1 port map( A1 => Q(965), A2 => n49, B1 => Q(901), B2 => n50, 
                           ZN => n130);
   U138 : AOI22_X1 port map( A1 => Q(997), A2 => n51, B1 => Q(933), B2 => n52, 
                           ZN => n129);
   U139 : OR4_X1 port map( A1 => n133, A2 => n134, A3 => n135, A4 => n136, ZN 
                           => Y(4));
   U140 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => n136);
   U141 : AOI22_X1 port map( A1 => Q(100), A2 => n9, B1 => Q(196), B2 => n10, 
                           ZN => n140);
   U142 : AOI22_X1 port map( A1 => Q(164), A2 => n11, B1 => Q(36), B2 => n12, 
                           ZN => n139);
   U143 : AOI22_X1 port map( A1 => Q(4), A2 => n13, B1 => Q(68), B2 => n14, ZN 
                           => n138);
   U144 : AOI22_X1 port map( A1 => Q(228), A2 => n15, B1 => Q(132), B2 => n16, 
                           ZN => n137);
   U145 : NAND4_X1 port map( A1 => n141, A2 => n142, A3 => n143, A4 => n144, ZN
                           => n135);
   U146 : AOI22_X1 port map( A1 => Q(324), A2 => n21, B1 => Q(420), B2 => n22, 
                           ZN => n144);
   U147 : AOI22_X1 port map( A1 => Q(388), A2 => n23, B1 => Q(260), B2 => n24, 
                           ZN => n143);
   U148 : AOI22_X1 port map( A1 => Q(356), A2 => n25, B1 => Q(292), B2 => n26, 
                           ZN => n142);
   U149 : AOI22_X1 port map( A1 => Q(644), A2 => n27, B1 => Q(452), B2 => n28, 
                           ZN => n141);
   U150 : NAND4_X1 port map( A1 => n145, A2 => n146, A3 => n147, A4 => n148, ZN
                           => n134);
   U151 : AOI22_X1 port map( A1 => Q(484), A2 => n33, B1 => Q(548), B2 => n34, 
                           ZN => n148);
   U152 : AOI22_X1 port map( A1 => Q(516), A2 => n35, B1 => Q(612), B2 => n36, 
                           ZN => n147);
   U153 : AOI22_X1 port map( A1 => Q(676), A2 => n37, B1 => Q(580), B2 => n38, 
                           ZN => n146);
   U154 : AOI22_X1 port map( A1 => Q(772), A2 => n39, B1 => Q(868), B2 => n40, 
                           ZN => n145);
   U155 : NAND4_X1 port map( A1 => n149, A2 => n150, A3 => n151, A4 => n152, ZN
                           => n133);
   U156 : AOI22_X1 port map( A1 => Q(836), A2 => n45, B1 => Q(708), B2 => n46, 
                           ZN => n152);
   U157 : AOI22_X1 port map( A1 => Q(804), A2 => n47, B1 => Q(740), B2 => n48, 
                           ZN => n151);
   U158 : AOI22_X1 port map( A1 => Q(964), A2 => n49, B1 => Q(900), B2 => n50, 
                           ZN => n150);
   U159 : AOI22_X1 port map( A1 => Q(996), A2 => n51, B1 => Q(932), B2 => n52, 
                           ZN => n149);
   U160 : OR4_X1 port map( A1 => n153, A2 => n154, A3 => n155, A4 => n156, ZN 
                           => Y(3));
   U161 : NAND4_X1 port map( A1 => n157, A2 => n158, A3 => n159, A4 => n160, ZN
                           => n156);
   U162 : AOI22_X1 port map( A1 => Q(99), A2 => n9, B1 => Q(195), B2 => n10, ZN
                           => n160);
   U163 : AOI22_X1 port map( A1 => Q(163), A2 => n11, B1 => Q(35), B2 => n12, 
                           ZN => n159);
   U164 : AOI22_X1 port map( A1 => Q(3), A2 => n13, B1 => Q(67), B2 => n14, ZN 
                           => n158);
   U165 : AOI22_X1 port map( A1 => Q(227), A2 => n15, B1 => Q(131), B2 => n16, 
                           ZN => n157);
   U166 : NAND4_X1 port map( A1 => n161, A2 => n162, A3 => n163, A4 => n164, ZN
                           => n155);
   U167 : AOI22_X1 port map( A1 => Q(323), A2 => n21, B1 => Q(419), B2 => n22, 
                           ZN => n164);
   U168 : AOI22_X1 port map( A1 => Q(387), A2 => n23, B1 => Q(259), B2 => n24, 
                           ZN => n163);
   U169 : AOI22_X1 port map( A1 => Q(355), A2 => n25, B1 => Q(291), B2 => n26, 
                           ZN => n162);
   U170 : AOI22_X1 port map( A1 => Q(643), A2 => n27, B1 => Q(451), B2 => n28, 
                           ZN => n161);
   U171 : NAND4_X1 port map( A1 => n165, A2 => n166, A3 => n167, A4 => n168, ZN
                           => n154);
   U172 : AOI22_X1 port map( A1 => Q(483), A2 => n33, B1 => Q(547), B2 => n34, 
                           ZN => n168);
   U173 : AOI22_X1 port map( A1 => Q(515), A2 => n35, B1 => Q(611), B2 => n36, 
                           ZN => n167);
   U174 : AOI22_X1 port map( A1 => Q(675), A2 => n37, B1 => Q(579), B2 => n38, 
                           ZN => n166);
   U175 : AOI22_X1 port map( A1 => Q(771), A2 => n39, B1 => Q(867), B2 => n40, 
                           ZN => n165);
   U176 : NAND4_X1 port map( A1 => n169, A2 => n170, A3 => n171, A4 => n172, ZN
                           => n153);
   U177 : AOI22_X1 port map( A1 => Q(835), A2 => n45, B1 => Q(707), B2 => n46, 
                           ZN => n172);
   U178 : AOI22_X1 port map( A1 => Q(803), A2 => n47, B1 => Q(739), B2 => n48, 
                           ZN => n171);
   U179 : AOI22_X1 port map( A1 => Q(963), A2 => n49, B1 => Q(899), B2 => n50, 
                           ZN => n170);
   U180 : AOI22_X1 port map( A1 => Q(995), A2 => n51, B1 => Q(931), B2 => n52, 
                           ZN => n169);
   U181 : OR4_X1 port map( A1 => n173, A2 => n174, A3 => n175, A4 => n176, ZN 
                           => Y(31));
   U182 : NAND4_X1 port map( A1 => n177, A2 => n178, A3 => n179, A4 => n180, ZN
                           => n176);
   U183 : AOI22_X1 port map( A1 => Q(127), A2 => n9, B1 => Q(223), B2 => n10, 
                           ZN => n180);
   U184 : AOI22_X1 port map( A1 => Q(191), A2 => n11, B1 => Q(63), B2 => n12, 
                           ZN => n179);
   U185 : AOI22_X1 port map( A1 => Q(31), A2 => n13, B1 => Q(95), B2 => n14, ZN
                           => n178);
   U186 : AOI22_X1 port map( A1 => Q(255), A2 => n15, B1 => Q(159), B2 => n16, 
                           ZN => n177);
   U187 : NAND4_X1 port map( A1 => n181, A2 => n182, A3 => n183, A4 => n184, ZN
                           => n175);
   U188 : AOI22_X1 port map( A1 => Q(351), A2 => n21, B1 => Q(447), B2 => n22, 
                           ZN => n184);
   U189 : AOI22_X1 port map( A1 => Q(415), A2 => n23, B1 => Q(287), B2 => n24, 
                           ZN => n183);
   U190 : AOI22_X1 port map( A1 => Q(383), A2 => n25, B1 => Q(319), B2 => n26, 
                           ZN => n182);
   U191 : AOI22_X1 port map( A1 => Q(671), A2 => n27, B1 => Q(479), B2 => n28, 
                           ZN => n181);
   U192 : NAND4_X1 port map( A1 => n185, A2 => n186, A3 => n187, A4 => n188, ZN
                           => n174);
   U193 : AOI22_X1 port map( A1 => Q(511), A2 => n33, B1 => Q(575), B2 => n34, 
                           ZN => n188);
   U194 : AOI22_X1 port map( A1 => Q(543), A2 => n35, B1 => Q(639), B2 => n36, 
                           ZN => n187);
   U195 : AOI22_X1 port map( A1 => Q(703), A2 => n37, B1 => Q(607), B2 => n38, 
                           ZN => n186);
   U196 : AOI22_X1 port map( A1 => Q(799), A2 => n39, B1 => Q(895), B2 => n40, 
                           ZN => n185);
   U197 : NAND4_X1 port map( A1 => n189, A2 => n190, A3 => n191, A4 => n192, ZN
                           => n173);
   U198 : AOI22_X1 port map( A1 => Q(863), A2 => n45, B1 => Q(735), B2 => n46, 
                           ZN => n192);
   U199 : AOI22_X1 port map( A1 => Q(831), A2 => n47, B1 => Q(767), B2 => n48, 
                           ZN => n191);
   U200 : AOI22_X1 port map( A1 => Q(991), A2 => n49, B1 => Q(927), B2 => n50, 
                           ZN => n190);
   U201 : AOI22_X1 port map( A1 => Q(1023), A2 => n51, B1 => Q(959), B2 => n52,
                           ZN => n189);
   U202 : OR4_X1 port map( A1 => n193, A2 => n194, A3 => n195, A4 => n196, ZN 
                           => Y(30));
   U203 : NAND4_X1 port map( A1 => n197, A2 => n198, A3 => n199, A4 => n200, ZN
                           => n196);
   U204 : AOI22_X1 port map( A1 => Q(126), A2 => n9, B1 => Q(222), B2 => n10, 
                           ZN => n200);
   U205 : AOI22_X1 port map( A1 => Q(190), A2 => n11, B1 => Q(62), B2 => n12, 
                           ZN => n199);
   U206 : AOI22_X1 port map( A1 => Q(30), A2 => n13, B1 => Q(94), B2 => n14, ZN
                           => n198);
   U207 : AOI22_X1 port map( A1 => Q(254), A2 => n15, B1 => Q(158), B2 => n16, 
                           ZN => n197);
   U208 : NAND4_X1 port map( A1 => n201, A2 => n202, A3 => n203, A4 => n204, ZN
                           => n195);
   U209 : AOI22_X1 port map( A1 => Q(350), A2 => n21, B1 => Q(446), B2 => n22, 
                           ZN => n204);
   U210 : AOI22_X1 port map( A1 => Q(414), A2 => n23, B1 => Q(286), B2 => n24, 
                           ZN => n203);
   U211 : AOI22_X1 port map( A1 => Q(382), A2 => n25, B1 => Q(318), B2 => n26, 
                           ZN => n202);
   U212 : AOI22_X1 port map( A1 => Q(670), A2 => n27, B1 => Q(478), B2 => n28, 
                           ZN => n201);
   U213 : NAND4_X1 port map( A1 => n205, A2 => n206, A3 => n207, A4 => n208, ZN
                           => n194);
   U214 : AOI22_X1 port map( A1 => Q(510), A2 => n33, B1 => Q(574), B2 => n34, 
                           ZN => n208);
   U215 : AOI22_X1 port map( A1 => Q(542), A2 => n35, B1 => Q(638), B2 => n36, 
                           ZN => n207);
   U216 : AOI22_X1 port map( A1 => Q(702), A2 => n37, B1 => Q(606), B2 => n38, 
                           ZN => n206);
   U217 : AOI22_X1 port map( A1 => Q(798), A2 => n39, B1 => Q(894), B2 => n40, 
                           ZN => n205);
   U218 : NAND4_X1 port map( A1 => n209, A2 => n210, A3 => n211, A4 => n212, ZN
                           => n193);
   U219 : AOI22_X1 port map( A1 => Q(862), A2 => n45, B1 => Q(734), B2 => n46, 
                           ZN => n212);
   U220 : AOI22_X1 port map( A1 => Q(830), A2 => n47, B1 => Q(766), B2 => n48, 
                           ZN => n211);
   U221 : AOI22_X1 port map( A1 => Q(990), A2 => n49, B1 => Q(926), B2 => n50, 
                           ZN => n210);
   U222 : AOI22_X1 port map( A1 => Q(1022), A2 => n51, B1 => Q(958), B2 => n52,
                           ZN => n209);
   U223 : OR4_X1 port map( A1 => n213, A2 => n214, A3 => n215, A4 => n216, ZN 
                           => Y(2));
   U224 : NAND4_X1 port map( A1 => n217, A2 => n218, A3 => n219, A4 => n220, ZN
                           => n216);
   U225 : AOI22_X1 port map( A1 => Q(98), A2 => n9, B1 => Q(194), B2 => n10, ZN
                           => n220);
   U226 : AOI22_X1 port map( A1 => Q(162), A2 => n11, B1 => Q(34), B2 => n12, 
                           ZN => n219);
   U227 : AOI22_X1 port map( A1 => Q(2), A2 => n13, B1 => Q(66), B2 => n14, ZN 
                           => n218);
   U228 : AOI22_X1 port map( A1 => Q(226), A2 => n15, B1 => Q(130), B2 => n16, 
                           ZN => n217);
   U229 : NAND4_X1 port map( A1 => n221, A2 => n222, A3 => n223, A4 => n224, ZN
                           => n215);
   U230 : AOI22_X1 port map( A1 => Q(322), A2 => n21, B1 => Q(418), B2 => n22, 
                           ZN => n224);
   U231 : AOI22_X1 port map( A1 => Q(386), A2 => n23, B1 => Q(258), B2 => n24, 
                           ZN => n223);
   U232 : AOI22_X1 port map( A1 => Q(354), A2 => n25, B1 => Q(290), B2 => n26, 
                           ZN => n222);
   U233 : AOI22_X1 port map( A1 => Q(642), A2 => n27, B1 => Q(450), B2 => n28, 
                           ZN => n221);
   U234 : NAND4_X1 port map( A1 => n225, A2 => n226, A3 => n227, A4 => n228, ZN
                           => n214);
   U235 : AOI22_X1 port map( A1 => Q(482), A2 => n33, B1 => Q(546), B2 => n34, 
                           ZN => n228);
   U236 : AOI22_X1 port map( A1 => Q(514), A2 => n35, B1 => Q(610), B2 => n36, 
                           ZN => n227);
   U237 : AOI22_X1 port map( A1 => Q(674), A2 => n37, B1 => Q(578), B2 => n38, 
                           ZN => n226);
   U238 : AOI22_X1 port map( A1 => Q(770), A2 => n39, B1 => Q(866), B2 => n40, 
                           ZN => n225);
   U239 : NAND4_X1 port map( A1 => n229, A2 => n230, A3 => n231, A4 => n232, ZN
                           => n213);
   U240 : AOI22_X1 port map( A1 => Q(834), A2 => n45, B1 => Q(706), B2 => n46, 
                           ZN => n232);
   U241 : AOI22_X1 port map( A1 => Q(802), A2 => n47, B1 => Q(738), B2 => n48, 
                           ZN => n231);
   U242 : AOI22_X1 port map( A1 => Q(962), A2 => n49, B1 => Q(898), B2 => n50, 
                           ZN => n230);
   U243 : AOI22_X1 port map( A1 => Q(994), A2 => n51, B1 => Q(930), B2 => n52, 
                           ZN => n229);
   U244 : OR4_X1 port map( A1 => n233, A2 => n234, A3 => n235, A4 => n236, ZN 
                           => Y(29));
   U245 : NAND4_X1 port map( A1 => n237, A2 => n238, A3 => n239, A4 => n240, ZN
                           => n236);
   U246 : AOI22_X1 port map( A1 => Q(125), A2 => n9, B1 => Q(221), B2 => n10, 
                           ZN => n240);
   U247 : AOI22_X1 port map( A1 => Q(189), A2 => n11, B1 => Q(61), B2 => n12, 
                           ZN => n239);
   U248 : AOI22_X1 port map( A1 => Q(29), A2 => n13, B1 => Q(93), B2 => n14, ZN
                           => n238);
   U249 : AOI22_X1 port map( A1 => Q(253), A2 => n15, B1 => Q(157), B2 => n16, 
                           ZN => n237);
   U250 : NAND4_X1 port map( A1 => n241, A2 => n242, A3 => n243, A4 => n244, ZN
                           => n235);
   U251 : AOI22_X1 port map( A1 => Q(349), A2 => n21, B1 => Q(445), B2 => n22, 
                           ZN => n244);
   U252 : AOI22_X1 port map( A1 => Q(413), A2 => n23, B1 => Q(285), B2 => n24, 
                           ZN => n243);
   U253 : AOI22_X1 port map( A1 => Q(381), A2 => n25, B1 => Q(317), B2 => n26, 
                           ZN => n242);
   U254 : AOI22_X1 port map( A1 => Q(669), A2 => n27, B1 => Q(477), B2 => n28, 
                           ZN => n241);
   U255 : NAND4_X1 port map( A1 => n245, A2 => n246, A3 => n247, A4 => n248, ZN
                           => n234);
   U256 : AOI22_X1 port map( A1 => Q(509), A2 => n33, B1 => Q(573), B2 => n34, 
                           ZN => n248);
   U257 : AOI22_X1 port map( A1 => Q(541), A2 => n35, B1 => Q(637), B2 => n36, 
                           ZN => n247);
   U258 : AOI22_X1 port map( A1 => Q(701), A2 => n37, B1 => Q(605), B2 => n38, 
                           ZN => n246);
   U259 : AOI22_X1 port map( A1 => Q(797), A2 => n39, B1 => Q(893), B2 => n40, 
                           ZN => n245);
   U260 : NAND4_X1 port map( A1 => n249, A2 => n250, A3 => n251, A4 => n252, ZN
                           => n233);
   U261 : AOI22_X1 port map( A1 => Q(861), A2 => n45, B1 => Q(733), B2 => n46, 
                           ZN => n252);
   U262 : AOI22_X1 port map( A1 => Q(829), A2 => n47, B1 => Q(765), B2 => n48, 
                           ZN => n251);
   U263 : AOI22_X1 port map( A1 => Q(989), A2 => n49, B1 => Q(925), B2 => n50, 
                           ZN => n250);
   U264 : AOI22_X1 port map( A1 => Q(1021), A2 => n51, B1 => Q(957), B2 => n52,
                           ZN => n249);
   U265 : OR4_X1 port map( A1 => n253, A2 => n254, A3 => n255, A4 => n256, ZN 
                           => Y(28));
   U266 : NAND4_X1 port map( A1 => n257, A2 => n258, A3 => n259, A4 => n260, ZN
                           => n256);
   U267 : AOI22_X1 port map( A1 => Q(124), A2 => n9, B1 => Q(220), B2 => n10, 
                           ZN => n260);
   U268 : AOI22_X1 port map( A1 => Q(188), A2 => n11, B1 => Q(60), B2 => n12, 
                           ZN => n259);
   U269 : AOI22_X1 port map( A1 => Q(28), A2 => n13, B1 => Q(92), B2 => n14, ZN
                           => n258);
   U270 : AOI22_X1 port map( A1 => Q(252), A2 => n15, B1 => Q(156), B2 => n16, 
                           ZN => n257);
   U271 : NAND4_X1 port map( A1 => n261, A2 => n262, A3 => n263, A4 => n264, ZN
                           => n255);
   U272 : AOI22_X1 port map( A1 => Q(348), A2 => n21, B1 => Q(444), B2 => n22, 
                           ZN => n264);
   U273 : AOI22_X1 port map( A1 => Q(412), A2 => n23, B1 => Q(284), B2 => n24, 
                           ZN => n263);
   U274 : AOI22_X1 port map( A1 => Q(380), A2 => n25, B1 => Q(316), B2 => n26, 
                           ZN => n262);
   U275 : AOI22_X1 port map( A1 => Q(668), A2 => n27, B1 => Q(476), B2 => n28, 
                           ZN => n261);
   U276 : NAND4_X1 port map( A1 => n265, A2 => n266, A3 => n267, A4 => n268, ZN
                           => n254);
   U277 : AOI22_X1 port map( A1 => Q(508), A2 => n33, B1 => Q(572), B2 => n34, 
                           ZN => n268);
   U278 : AOI22_X1 port map( A1 => Q(540), A2 => n35, B1 => Q(636), B2 => n36, 
                           ZN => n267);
   U279 : AOI22_X1 port map( A1 => Q(700), A2 => n37, B1 => Q(604), B2 => n38, 
                           ZN => n266);
   U280 : AOI22_X1 port map( A1 => Q(796), A2 => n39, B1 => Q(892), B2 => n40, 
                           ZN => n265);
   U281 : NAND4_X1 port map( A1 => n269, A2 => n270, A3 => n271, A4 => n272, ZN
                           => n253);
   U282 : AOI22_X1 port map( A1 => Q(860), A2 => n45, B1 => Q(732), B2 => n46, 
                           ZN => n272);
   U283 : AOI22_X1 port map( A1 => Q(828), A2 => n47, B1 => Q(764), B2 => n48, 
                           ZN => n271);
   U284 : AOI22_X1 port map( A1 => Q(988), A2 => n49, B1 => Q(924), B2 => n50, 
                           ZN => n270);
   U285 : AOI22_X1 port map( A1 => Q(1020), A2 => n51, B1 => Q(956), B2 => n52,
                           ZN => n269);
   U286 : OR4_X1 port map( A1 => n273, A2 => n274, A3 => n275, A4 => n276, ZN 
                           => Y(27));
   U287 : NAND4_X1 port map( A1 => n277, A2 => n278, A3 => n279, A4 => n280, ZN
                           => n276);
   U288 : AOI22_X1 port map( A1 => Q(123), A2 => n9, B1 => Q(219), B2 => n10, 
                           ZN => n280);
   U289 : AOI22_X1 port map( A1 => Q(187), A2 => n11, B1 => Q(59), B2 => n12, 
                           ZN => n279);
   U290 : AOI22_X1 port map( A1 => Q(27), A2 => n13, B1 => Q(91), B2 => n14, ZN
                           => n278);
   U291 : AOI22_X1 port map( A1 => Q(251), A2 => n15, B1 => Q(155), B2 => n16, 
                           ZN => n277);
   U292 : NAND4_X1 port map( A1 => n281, A2 => n282, A3 => n283, A4 => n284, ZN
                           => n275);
   U293 : AOI22_X1 port map( A1 => Q(347), A2 => n21, B1 => Q(443), B2 => n22, 
                           ZN => n284);
   U294 : AOI22_X1 port map( A1 => Q(411), A2 => n23, B1 => Q(283), B2 => n24, 
                           ZN => n283);
   U295 : AOI22_X1 port map( A1 => Q(379), A2 => n25, B1 => Q(315), B2 => n26, 
                           ZN => n282);
   U296 : AOI22_X1 port map( A1 => Q(667), A2 => n27, B1 => Q(475), B2 => n28, 
                           ZN => n281);
   U297 : NAND4_X1 port map( A1 => n285, A2 => n286, A3 => n287, A4 => n288, ZN
                           => n274);
   U298 : AOI22_X1 port map( A1 => Q(507), A2 => n33, B1 => Q(571), B2 => n34, 
                           ZN => n288);
   U299 : AOI22_X1 port map( A1 => Q(539), A2 => n35, B1 => Q(635), B2 => n36, 
                           ZN => n287);
   U300 : AOI22_X1 port map( A1 => Q(699), A2 => n37, B1 => Q(603), B2 => n38, 
                           ZN => n286);
   U301 : AOI22_X1 port map( A1 => Q(795), A2 => n39, B1 => Q(891), B2 => n40, 
                           ZN => n285);
   U302 : NAND4_X1 port map( A1 => n289, A2 => n290, A3 => n291, A4 => n292, ZN
                           => n273);
   U303 : AOI22_X1 port map( A1 => Q(859), A2 => n45, B1 => Q(731), B2 => n46, 
                           ZN => n292);
   U304 : AOI22_X1 port map( A1 => Q(827), A2 => n47, B1 => Q(763), B2 => n48, 
                           ZN => n291);
   U305 : AOI22_X1 port map( A1 => Q(987), A2 => n49, B1 => Q(923), B2 => n50, 
                           ZN => n290);
   U306 : AOI22_X1 port map( A1 => Q(1019), A2 => n51, B1 => Q(955), B2 => n52,
                           ZN => n289);
   U307 : OR4_X1 port map( A1 => n293, A2 => n294, A3 => n295, A4 => n296, ZN 
                           => Y(26));
   U308 : NAND4_X1 port map( A1 => n297, A2 => n298, A3 => n299, A4 => n300, ZN
                           => n296);
   U309 : AOI22_X1 port map( A1 => Q(122), A2 => n9, B1 => Q(218), B2 => n10, 
                           ZN => n300);
   U310 : AOI22_X1 port map( A1 => Q(186), A2 => n11, B1 => Q(58), B2 => n12, 
                           ZN => n299);
   U311 : AOI22_X1 port map( A1 => Q(26), A2 => n13, B1 => Q(90), B2 => n14, ZN
                           => n298);
   U312 : AOI22_X1 port map( A1 => Q(250), A2 => n15, B1 => Q(154), B2 => n16, 
                           ZN => n297);
   U313 : NAND4_X1 port map( A1 => n301, A2 => n302, A3 => n303, A4 => n304, ZN
                           => n295);
   U314 : AOI22_X1 port map( A1 => Q(346), A2 => n21, B1 => Q(442), B2 => n22, 
                           ZN => n304);
   U315 : AOI22_X1 port map( A1 => Q(410), A2 => n23, B1 => Q(282), B2 => n24, 
                           ZN => n303);
   U316 : AOI22_X1 port map( A1 => Q(378), A2 => n25, B1 => Q(314), B2 => n26, 
                           ZN => n302);
   U317 : AOI22_X1 port map( A1 => Q(666), A2 => n27, B1 => Q(474), B2 => n28, 
                           ZN => n301);
   U318 : NAND4_X1 port map( A1 => n305, A2 => n306, A3 => n307, A4 => n308, ZN
                           => n294);
   U319 : AOI22_X1 port map( A1 => Q(506), A2 => n33, B1 => Q(570), B2 => n34, 
                           ZN => n308);
   U320 : AOI22_X1 port map( A1 => Q(538), A2 => n35, B1 => Q(634), B2 => n36, 
                           ZN => n307);
   U321 : AOI22_X1 port map( A1 => Q(698), A2 => n37, B1 => Q(602), B2 => n38, 
                           ZN => n306);
   U322 : AOI22_X1 port map( A1 => Q(794), A2 => n39, B1 => Q(890), B2 => n40, 
                           ZN => n305);
   U323 : NAND4_X1 port map( A1 => n309, A2 => n310, A3 => n311, A4 => n312, ZN
                           => n293);
   U324 : AOI22_X1 port map( A1 => Q(858), A2 => n45, B1 => Q(730), B2 => n46, 
                           ZN => n312);
   U325 : AOI22_X1 port map( A1 => Q(826), A2 => n47, B1 => Q(762), B2 => n48, 
                           ZN => n311);
   U326 : AOI22_X1 port map( A1 => Q(986), A2 => n49, B1 => Q(922), B2 => n50, 
                           ZN => n310);
   U327 : AOI22_X1 port map( A1 => Q(1018), A2 => n51, B1 => Q(954), B2 => n52,
                           ZN => n309);
   U328 : OR4_X1 port map( A1 => n313, A2 => n314, A3 => n315, A4 => n316, ZN 
                           => Y(25));
   U329 : NAND4_X1 port map( A1 => n317, A2 => n318, A3 => n319, A4 => n320, ZN
                           => n316);
   U330 : AOI22_X1 port map( A1 => Q(121), A2 => n9, B1 => Q(217), B2 => n10, 
                           ZN => n320);
   U331 : AOI22_X1 port map( A1 => Q(185), A2 => n11, B1 => Q(57), B2 => n12, 
                           ZN => n319);
   U332 : AOI22_X1 port map( A1 => Q(25), A2 => n13, B1 => Q(89), B2 => n14, ZN
                           => n318);
   U333 : AOI22_X1 port map( A1 => Q(249), A2 => n15, B1 => Q(153), B2 => n16, 
                           ZN => n317);
   U334 : NAND4_X1 port map( A1 => n321, A2 => n322, A3 => n323, A4 => n324, ZN
                           => n315);
   U335 : AOI22_X1 port map( A1 => Q(345), A2 => n21, B1 => Q(441), B2 => n22, 
                           ZN => n324);
   U336 : AOI22_X1 port map( A1 => Q(409), A2 => n23, B1 => Q(281), B2 => n24, 
                           ZN => n323);
   U337 : AOI22_X1 port map( A1 => Q(377), A2 => n25, B1 => Q(313), B2 => n26, 
                           ZN => n322);
   U338 : AOI22_X1 port map( A1 => Q(665), A2 => n27, B1 => Q(473), B2 => n28, 
                           ZN => n321);
   U339 : NAND4_X1 port map( A1 => n325, A2 => n326, A3 => n327, A4 => n328, ZN
                           => n314);
   U340 : AOI22_X1 port map( A1 => Q(505), A2 => n33, B1 => Q(569), B2 => n34, 
                           ZN => n328);
   U341 : AOI22_X1 port map( A1 => Q(537), A2 => n35, B1 => Q(633), B2 => n36, 
                           ZN => n327);
   U342 : AOI22_X1 port map( A1 => Q(697), A2 => n37, B1 => Q(601), B2 => n38, 
                           ZN => n326);
   U343 : AOI22_X1 port map( A1 => Q(793), A2 => n39, B1 => Q(889), B2 => n40, 
                           ZN => n325);
   U344 : NAND4_X1 port map( A1 => n329, A2 => n330, A3 => n331, A4 => n332, ZN
                           => n313);
   U345 : AOI22_X1 port map( A1 => Q(857), A2 => n45, B1 => Q(729), B2 => n46, 
                           ZN => n332);
   U346 : AOI22_X1 port map( A1 => Q(825), A2 => n47, B1 => Q(761), B2 => n48, 
                           ZN => n331);
   U347 : AOI22_X1 port map( A1 => Q(985), A2 => n49, B1 => Q(921), B2 => n50, 
                           ZN => n330);
   U348 : AOI22_X1 port map( A1 => Q(1017), A2 => n51, B1 => Q(953), B2 => n52,
                           ZN => n329);
   U349 : OR4_X1 port map( A1 => n333, A2 => n334, A3 => n335, A4 => n336, ZN 
                           => Y(24));
   U350 : NAND4_X1 port map( A1 => n337, A2 => n338, A3 => n339, A4 => n340, ZN
                           => n336);
   U351 : AOI22_X1 port map( A1 => Q(120), A2 => n9, B1 => Q(216), B2 => n10, 
                           ZN => n340);
   U352 : AOI22_X1 port map( A1 => Q(184), A2 => n11, B1 => Q(56), B2 => n12, 
                           ZN => n339);
   U353 : AOI22_X1 port map( A1 => Q(24), A2 => n13, B1 => Q(88), B2 => n14, ZN
                           => n338);
   U354 : AOI22_X1 port map( A1 => Q(248), A2 => n15, B1 => Q(152), B2 => n16, 
                           ZN => n337);
   U355 : NAND4_X1 port map( A1 => n341, A2 => n342, A3 => n343, A4 => n344, ZN
                           => n335);
   U356 : AOI22_X1 port map( A1 => Q(344), A2 => n21, B1 => Q(440), B2 => n22, 
                           ZN => n344);
   U357 : AOI22_X1 port map( A1 => Q(408), A2 => n23, B1 => Q(280), B2 => n24, 
                           ZN => n343);
   U358 : AOI22_X1 port map( A1 => Q(376), A2 => n25, B1 => Q(312), B2 => n26, 
                           ZN => n342);
   U359 : AOI22_X1 port map( A1 => Q(664), A2 => n27, B1 => Q(472), B2 => n28, 
                           ZN => n341);
   U360 : NAND4_X1 port map( A1 => n345, A2 => n346, A3 => n347, A4 => n348, ZN
                           => n334);
   U361 : AOI22_X1 port map( A1 => Q(504), A2 => n33, B1 => Q(568), B2 => n34, 
                           ZN => n348);
   U362 : AOI22_X1 port map( A1 => Q(536), A2 => n35, B1 => Q(632), B2 => n36, 
                           ZN => n347);
   U363 : AOI22_X1 port map( A1 => Q(696), A2 => n37, B1 => Q(600), B2 => n38, 
                           ZN => n346);
   U364 : AOI22_X1 port map( A1 => Q(792), A2 => n39, B1 => Q(888), B2 => n40, 
                           ZN => n345);
   U365 : NAND4_X1 port map( A1 => n349, A2 => n350, A3 => n351, A4 => n352, ZN
                           => n333);
   U366 : AOI22_X1 port map( A1 => Q(856), A2 => n45, B1 => Q(728), B2 => n46, 
                           ZN => n352);
   U367 : AOI22_X1 port map( A1 => Q(824), A2 => n47, B1 => Q(760), B2 => n48, 
                           ZN => n351);
   U368 : AOI22_X1 port map( A1 => Q(984), A2 => n49, B1 => Q(920), B2 => n50, 
                           ZN => n350);
   U369 : AOI22_X1 port map( A1 => Q(1016), A2 => n51, B1 => Q(952), B2 => n52,
                           ZN => n349);
   U370 : OR4_X1 port map( A1 => n353, A2 => n354, A3 => n355, A4 => n356, ZN 
                           => Y(23));
   U371 : NAND4_X1 port map( A1 => n357, A2 => n358, A3 => n359, A4 => n360, ZN
                           => n356);
   U372 : AOI22_X1 port map( A1 => Q(119), A2 => n9, B1 => Q(215), B2 => n10, 
                           ZN => n360);
   U373 : AOI22_X1 port map( A1 => Q(183), A2 => n11, B1 => Q(55), B2 => n12, 
                           ZN => n359);
   U374 : AOI22_X1 port map( A1 => Q(23), A2 => n13, B1 => Q(87), B2 => n14, ZN
                           => n358);
   U375 : AOI22_X1 port map( A1 => Q(247), A2 => n15, B1 => Q(151), B2 => n16, 
                           ZN => n357);
   U376 : NAND4_X1 port map( A1 => n361, A2 => n362, A3 => n363, A4 => n364, ZN
                           => n355);
   U377 : AOI22_X1 port map( A1 => Q(343), A2 => n21, B1 => Q(439), B2 => n22, 
                           ZN => n364);
   U378 : AOI22_X1 port map( A1 => Q(407), A2 => n23, B1 => Q(279), B2 => n24, 
                           ZN => n363);
   U379 : AOI22_X1 port map( A1 => Q(375), A2 => n25, B1 => Q(311), B2 => n26, 
                           ZN => n362);
   U380 : AOI22_X1 port map( A1 => Q(663), A2 => n27, B1 => Q(471), B2 => n28, 
                           ZN => n361);
   U381 : NAND4_X1 port map( A1 => n365, A2 => n366, A3 => n367, A4 => n368, ZN
                           => n354);
   U382 : AOI22_X1 port map( A1 => Q(503), A2 => n33, B1 => Q(567), B2 => n34, 
                           ZN => n368);
   U383 : AOI22_X1 port map( A1 => Q(535), A2 => n35, B1 => Q(631), B2 => n36, 
                           ZN => n367);
   U384 : AOI22_X1 port map( A1 => Q(695), A2 => n37, B1 => Q(599), B2 => n38, 
                           ZN => n366);
   U385 : AOI22_X1 port map( A1 => Q(791), A2 => n39, B1 => Q(887), B2 => n40, 
                           ZN => n365);
   U386 : NAND4_X1 port map( A1 => n369, A2 => n370, A3 => n371, A4 => n372, ZN
                           => n353);
   U387 : AOI22_X1 port map( A1 => Q(855), A2 => n45, B1 => Q(727), B2 => n46, 
                           ZN => n372);
   U388 : AOI22_X1 port map( A1 => Q(823), A2 => n47, B1 => Q(759), B2 => n48, 
                           ZN => n371);
   U389 : AOI22_X1 port map( A1 => Q(983), A2 => n49, B1 => Q(919), B2 => n50, 
                           ZN => n370);
   U390 : AOI22_X1 port map( A1 => Q(1015), A2 => n51, B1 => Q(951), B2 => n52,
                           ZN => n369);
   U391 : OR4_X1 port map( A1 => n373, A2 => n374, A3 => n375, A4 => n376, ZN 
                           => Y(22));
   U392 : NAND4_X1 port map( A1 => n377, A2 => n378, A3 => n379, A4 => n380, ZN
                           => n376);
   U393 : AOI22_X1 port map( A1 => Q(118), A2 => n9, B1 => Q(214), B2 => n10, 
                           ZN => n380);
   U394 : AOI22_X1 port map( A1 => Q(182), A2 => n11, B1 => Q(54), B2 => n12, 
                           ZN => n379);
   U395 : AOI22_X1 port map( A1 => Q(22), A2 => n13, B1 => Q(86), B2 => n14, ZN
                           => n378);
   U396 : AOI22_X1 port map( A1 => Q(246), A2 => n15, B1 => Q(150), B2 => n16, 
                           ZN => n377);
   U397 : NAND4_X1 port map( A1 => n381, A2 => n382, A3 => n383, A4 => n384, ZN
                           => n375);
   U398 : AOI22_X1 port map( A1 => Q(342), A2 => n21, B1 => Q(438), B2 => n22, 
                           ZN => n384);
   U399 : AOI22_X1 port map( A1 => Q(406), A2 => n23, B1 => Q(278), B2 => n24, 
                           ZN => n383);
   U400 : AOI22_X1 port map( A1 => Q(374), A2 => n25, B1 => Q(310), B2 => n26, 
                           ZN => n382);
   U401 : AOI22_X1 port map( A1 => Q(662), A2 => n27, B1 => Q(470), B2 => n28, 
                           ZN => n381);
   U402 : NAND4_X1 port map( A1 => n385, A2 => n386, A3 => n387, A4 => n388, ZN
                           => n374);
   U403 : AOI22_X1 port map( A1 => Q(502), A2 => n33, B1 => Q(566), B2 => n34, 
                           ZN => n388);
   U404 : AOI22_X1 port map( A1 => Q(534), A2 => n35, B1 => Q(630), B2 => n36, 
                           ZN => n387);
   U405 : AOI22_X1 port map( A1 => Q(694), A2 => n37, B1 => Q(598), B2 => n38, 
                           ZN => n386);
   U406 : AOI22_X1 port map( A1 => Q(790), A2 => n39, B1 => Q(886), B2 => n40, 
                           ZN => n385);
   U407 : NAND4_X1 port map( A1 => n389, A2 => n390, A3 => n391, A4 => n392, ZN
                           => n373);
   U408 : AOI22_X1 port map( A1 => Q(854), A2 => n45, B1 => Q(726), B2 => n46, 
                           ZN => n392);
   U409 : AOI22_X1 port map( A1 => Q(822), A2 => n47, B1 => Q(758), B2 => n48, 
                           ZN => n391);
   U410 : AOI22_X1 port map( A1 => Q(982), A2 => n49, B1 => Q(918), B2 => n50, 
                           ZN => n390);
   U411 : AOI22_X1 port map( A1 => Q(1014), A2 => n51, B1 => Q(950), B2 => n52,
                           ZN => n389);
   U412 : OR4_X1 port map( A1 => n393, A2 => n394, A3 => n395, A4 => n396, ZN 
                           => Y(21));
   U413 : NAND4_X1 port map( A1 => n397, A2 => n398, A3 => n399, A4 => n400, ZN
                           => n396);
   U414 : AOI22_X1 port map( A1 => Q(117), A2 => n9, B1 => Q(213), B2 => n10, 
                           ZN => n400);
   U415 : AOI22_X1 port map( A1 => Q(181), A2 => n11, B1 => Q(53), B2 => n12, 
                           ZN => n399);
   U416 : AOI22_X1 port map( A1 => Q(21), A2 => n13, B1 => Q(85), B2 => n14, ZN
                           => n398);
   U417 : AOI22_X1 port map( A1 => Q(245), A2 => n15, B1 => Q(149), B2 => n16, 
                           ZN => n397);
   U418 : NAND4_X1 port map( A1 => n401, A2 => n402, A3 => n403, A4 => n404, ZN
                           => n395);
   U419 : AOI22_X1 port map( A1 => Q(341), A2 => n21, B1 => Q(437), B2 => n22, 
                           ZN => n404);
   U420 : AOI22_X1 port map( A1 => Q(405), A2 => n23, B1 => Q(277), B2 => n24, 
                           ZN => n403);
   U421 : AOI22_X1 port map( A1 => Q(373), A2 => n25, B1 => Q(309), B2 => n26, 
                           ZN => n402);
   U422 : AOI22_X1 port map( A1 => Q(661), A2 => n27, B1 => Q(469), B2 => n28, 
                           ZN => n401);
   U423 : NAND4_X1 port map( A1 => n405, A2 => n406, A3 => n407, A4 => n408, ZN
                           => n394);
   U424 : AOI22_X1 port map( A1 => Q(501), A2 => n33, B1 => Q(565), B2 => n34, 
                           ZN => n408);
   U425 : AOI22_X1 port map( A1 => Q(533), A2 => n35, B1 => Q(629), B2 => n36, 
                           ZN => n407);
   U426 : AOI22_X1 port map( A1 => Q(693), A2 => n37, B1 => Q(597), B2 => n38, 
                           ZN => n406);
   U427 : AOI22_X1 port map( A1 => Q(789), A2 => n39, B1 => Q(885), B2 => n40, 
                           ZN => n405);
   U428 : NAND4_X1 port map( A1 => n409, A2 => n410, A3 => n411, A4 => n412, ZN
                           => n393);
   U429 : AOI22_X1 port map( A1 => Q(853), A2 => n45, B1 => Q(725), B2 => n46, 
                           ZN => n412);
   U430 : AOI22_X1 port map( A1 => Q(821), A2 => n47, B1 => Q(757), B2 => n48, 
                           ZN => n411);
   U431 : AOI22_X1 port map( A1 => Q(981), A2 => n49, B1 => Q(917), B2 => n50, 
                           ZN => n410);
   U432 : AOI22_X1 port map( A1 => Q(1013), A2 => n51, B1 => Q(949), B2 => n52,
                           ZN => n409);
   U433 : OR4_X1 port map( A1 => n413, A2 => n414, A3 => n415, A4 => n416, ZN 
                           => Y(20));
   U434 : NAND4_X1 port map( A1 => n417, A2 => n418, A3 => n419, A4 => n420, ZN
                           => n416);
   U435 : AOI22_X1 port map( A1 => Q(116), A2 => n9, B1 => Q(212), B2 => n10, 
                           ZN => n420);
   U436 : AOI22_X1 port map( A1 => Q(180), A2 => n11, B1 => Q(52), B2 => n12, 
                           ZN => n419);
   U437 : AOI22_X1 port map( A1 => Q(20), A2 => n13, B1 => Q(84), B2 => n14, ZN
                           => n418);
   U438 : AOI22_X1 port map( A1 => Q(244), A2 => n15, B1 => Q(148), B2 => n16, 
                           ZN => n417);
   U439 : NAND4_X1 port map( A1 => n421, A2 => n422, A3 => n423, A4 => n424, ZN
                           => n415);
   U440 : AOI22_X1 port map( A1 => Q(340), A2 => n21, B1 => Q(436), B2 => n22, 
                           ZN => n424);
   U441 : AOI22_X1 port map( A1 => Q(404), A2 => n23, B1 => Q(276), B2 => n24, 
                           ZN => n423);
   U442 : AOI22_X1 port map( A1 => Q(372), A2 => n25, B1 => Q(308), B2 => n26, 
                           ZN => n422);
   U443 : AOI22_X1 port map( A1 => Q(660), A2 => n27, B1 => Q(468), B2 => n28, 
                           ZN => n421);
   U444 : NAND4_X1 port map( A1 => n425, A2 => n426, A3 => n427, A4 => n428, ZN
                           => n414);
   U445 : AOI22_X1 port map( A1 => Q(500), A2 => n33, B1 => Q(564), B2 => n34, 
                           ZN => n428);
   U446 : AOI22_X1 port map( A1 => Q(532), A2 => n35, B1 => Q(628), B2 => n36, 
                           ZN => n427);
   U447 : AOI22_X1 port map( A1 => Q(692), A2 => n37, B1 => Q(596), B2 => n38, 
                           ZN => n426);
   U448 : AOI22_X1 port map( A1 => Q(788), A2 => n39, B1 => Q(884), B2 => n40, 
                           ZN => n425);
   U449 : NAND4_X1 port map( A1 => n429, A2 => n430, A3 => n431, A4 => n432, ZN
                           => n413);
   U450 : AOI22_X1 port map( A1 => Q(852), A2 => n45, B1 => Q(724), B2 => n46, 
                           ZN => n432);
   U451 : AOI22_X1 port map( A1 => Q(820), A2 => n47, B1 => Q(756), B2 => n48, 
                           ZN => n431);
   U452 : AOI22_X1 port map( A1 => Q(980), A2 => n49, B1 => Q(916), B2 => n50, 
                           ZN => n430);
   U453 : AOI22_X1 port map( A1 => Q(1012), A2 => n51, B1 => Q(948), B2 => n52,
                           ZN => n429);
   U454 : OR4_X1 port map( A1 => n433, A2 => n434, A3 => n435, A4 => n436, ZN 
                           => Y(1));
   U455 : NAND4_X1 port map( A1 => n437, A2 => n438, A3 => n439, A4 => n440, ZN
                           => n436);
   U456 : AOI22_X1 port map( A1 => Q(97), A2 => n9, B1 => Q(193), B2 => n10, ZN
                           => n440);
   U457 : AOI22_X1 port map( A1 => Q(161), A2 => n11, B1 => Q(33), B2 => n12, 
                           ZN => n439);
   U458 : AOI22_X1 port map( A1 => Q(1), A2 => n13, B1 => Q(65), B2 => n14, ZN 
                           => n438);
   U459 : AOI22_X1 port map( A1 => Q(225), A2 => n15, B1 => Q(129), B2 => n16, 
                           ZN => n437);
   U460 : NAND4_X1 port map( A1 => n441, A2 => n442, A3 => n443, A4 => n444, ZN
                           => n435);
   U461 : AOI22_X1 port map( A1 => Q(321), A2 => n21, B1 => Q(417), B2 => n22, 
                           ZN => n444);
   U462 : AOI22_X1 port map( A1 => Q(385), A2 => n23, B1 => Q(257), B2 => n24, 
                           ZN => n443);
   U463 : AOI22_X1 port map( A1 => Q(353), A2 => n25, B1 => Q(289), B2 => n26, 
                           ZN => n442);
   U464 : AOI22_X1 port map( A1 => Q(641), A2 => n27, B1 => Q(449), B2 => n28, 
                           ZN => n441);
   U465 : NAND4_X1 port map( A1 => n445, A2 => n446, A3 => n447, A4 => n448, ZN
                           => n434);
   U466 : AOI22_X1 port map( A1 => Q(481), A2 => n33, B1 => Q(545), B2 => n34, 
                           ZN => n448);
   U467 : AOI22_X1 port map( A1 => Q(513), A2 => n35, B1 => Q(609), B2 => n36, 
                           ZN => n447);
   U468 : AOI22_X1 port map( A1 => Q(673), A2 => n37, B1 => Q(577), B2 => n38, 
                           ZN => n446);
   U469 : AOI22_X1 port map( A1 => Q(769), A2 => n39, B1 => Q(865), B2 => n40, 
                           ZN => n445);
   U470 : NAND4_X1 port map( A1 => n449, A2 => n450, A3 => n451, A4 => n452, ZN
                           => n433);
   U471 : AOI22_X1 port map( A1 => Q(833), A2 => n45, B1 => Q(705), B2 => n46, 
                           ZN => n452);
   U472 : AOI22_X1 port map( A1 => Q(801), A2 => n47, B1 => Q(737), B2 => n48, 
                           ZN => n451);
   U473 : AOI22_X1 port map( A1 => Q(961), A2 => n49, B1 => Q(897), B2 => n50, 
                           ZN => n450);
   U474 : AOI22_X1 port map( A1 => Q(993), A2 => n51, B1 => Q(929), B2 => n52, 
                           ZN => n449);
   U475 : OR4_X1 port map( A1 => n453, A2 => n454, A3 => n455, A4 => n456, ZN 
                           => Y(19));
   U476 : NAND4_X1 port map( A1 => n457, A2 => n458, A3 => n459, A4 => n460, ZN
                           => n456);
   U477 : AOI22_X1 port map( A1 => Q(115), A2 => n9, B1 => Q(211), B2 => n10, 
                           ZN => n460);
   U478 : AOI22_X1 port map( A1 => Q(179), A2 => n11, B1 => Q(51), B2 => n12, 
                           ZN => n459);
   U479 : AOI22_X1 port map( A1 => Q(19), A2 => n13, B1 => Q(83), B2 => n14, ZN
                           => n458);
   U480 : AOI22_X1 port map( A1 => Q(243), A2 => n15, B1 => Q(147), B2 => n16, 
                           ZN => n457);
   U481 : NAND4_X1 port map( A1 => n461, A2 => n462, A3 => n463, A4 => n464, ZN
                           => n455);
   U482 : AOI22_X1 port map( A1 => Q(339), A2 => n21, B1 => Q(435), B2 => n22, 
                           ZN => n464);
   U483 : AOI22_X1 port map( A1 => Q(403), A2 => n23, B1 => Q(275), B2 => n24, 
                           ZN => n463);
   U484 : AOI22_X1 port map( A1 => Q(371), A2 => n25, B1 => Q(307), B2 => n26, 
                           ZN => n462);
   U485 : AOI22_X1 port map( A1 => Q(659), A2 => n27, B1 => Q(467), B2 => n28, 
                           ZN => n461);
   U486 : NAND4_X1 port map( A1 => n465, A2 => n466, A3 => n467, A4 => n468, ZN
                           => n454);
   U487 : AOI22_X1 port map( A1 => Q(499), A2 => n33, B1 => Q(563), B2 => n34, 
                           ZN => n468);
   U488 : AOI22_X1 port map( A1 => Q(531), A2 => n35, B1 => Q(627), B2 => n36, 
                           ZN => n467);
   U489 : AOI22_X1 port map( A1 => Q(691), A2 => n37, B1 => Q(595), B2 => n38, 
                           ZN => n466);
   U490 : AOI22_X1 port map( A1 => Q(787), A2 => n39, B1 => Q(883), B2 => n40, 
                           ZN => n465);
   U491 : NAND4_X1 port map( A1 => n469, A2 => n470, A3 => n471, A4 => n472, ZN
                           => n453);
   U492 : AOI22_X1 port map( A1 => Q(851), A2 => n45, B1 => Q(723), B2 => n46, 
                           ZN => n472);
   U493 : AOI22_X1 port map( A1 => Q(819), A2 => n47, B1 => Q(755), B2 => n48, 
                           ZN => n471);
   U494 : AOI22_X1 port map( A1 => Q(979), A2 => n49, B1 => Q(915), B2 => n50, 
                           ZN => n470);
   U495 : AOI22_X1 port map( A1 => Q(1011), A2 => n51, B1 => Q(947), B2 => n52,
                           ZN => n469);
   U496 : OR4_X1 port map( A1 => n473, A2 => n474, A3 => n475, A4 => n476, ZN 
                           => Y(18));
   U497 : NAND4_X1 port map( A1 => n477, A2 => n478, A3 => n479, A4 => n480, ZN
                           => n476);
   U498 : AOI22_X1 port map( A1 => Q(114), A2 => n9, B1 => Q(210), B2 => n10, 
                           ZN => n480);
   U499 : AOI22_X1 port map( A1 => Q(178), A2 => n11, B1 => Q(50), B2 => n12, 
                           ZN => n479);
   U500 : AOI22_X1 port map( A1 => Q(18), A2 => n13, B1 => Q(82), B2 => n14, ZN
                           => n478);
   U501 : AOI22_X1 port map( A1 => Q(242), A2 => n15, B1 => Q(146), B2 => n16, 
                           ZN => n477);
   U502 : NAND4_X1 port map( A1 => n481, A2 => n482, A3 => n483, A4 => n484, ZN
                           => n475);
   U503 : AOI22_X1 port map( A1 => Q(338), A2 => n21, B1 => Q(434), B2 => n22, 
                           ZN => n484);
   U504 : AOI22_X1 port map( A1 => Q(402), A2 => n23, B1 => Q(274), B2 => n24, 
                           ZN => n483);
   U505 : AOI22_X1 port map( A1 => Q(370), A2 => n25, B1 => Q(306), B2 => n26, 
                           ZN => n482);
   U506 : AOI22_X1 port map( A1 => Q(658), A2 => n27, B1 => Q(466), B2 => n28, 
                           ZN => n481);
   U507 : NAND4_X1 port map( A1 => n485, A2 => n486, A3 => n487, A4 => n488, ZN
                           => n474);
   U508 : AOI22_X1 port map( A1 => Q(498), A2 => n33, B1 => Q(562), B2 => n34, 
                           ZN => n488);
   U509 : AOI22_X1 port map( A1 => Q(530), A2 => n35, B1 => Q(626), B2 => n36, 
                           ZN => n487);
   U510 : AOI22_X1 port map( A1 => Q(690), A2 => n37, B1 => Q(594), B2 => n38, 
                           ZN => n486);
   U511 : AOI22_X1 port map( A1 => Q(786), A2 => n39, B1 => Q(882), B2 => n40, 
                           ZN => n485);
   U512 : NAND4_X1 port map( A1 => n489, A2 => n490, A3 => n491, A4 => n492, ZN
                           => n473);
   U513 : AOI22_X1 port map( A1 => Q(850), A2 => n45, B1 => Q(722), B2 => n46, 
                           ZN => n492);
   U514 : AOI22_X1 port map( A1 => Q(818), A2 => n47, B1 => Q(754), B2 => n48, 
                           ZN => n491);
   U515 : AOI22_X1 port map( A1 => Q(978), A2 => n49, B1 => Q(914), B2 => n50, 
                           ZN => n490);
   U516 : AOI22_X1 port map( A1 => Q(1010), A2 => n51, B1 => Q(946), B2 => n52,
                           ZN => n489);
   U517 : OR4_X1 port map( A1 => n493, A2 => n494, A3 => n495, A4 => n496, ZN 
                           => Y(17));
   U518 : NAND4_X1 port map( A1 => n497, A2 => n498, A3 => n499, A4 => n500, ZN
                           => n496);
   U519 : AOI22_X1 port map( A1 => Q(113), A2 => n9, B1 => Q(209), B2 => n10, 
                           ZN => n500);
   U520 : AOI22_X1 port map( A1 => Q(177), A2 => n11, B1 => Q(49), B2 => n12, 
                           ZN => n499);
   U521 : AOI22_X1 port map( A1 => Q(17), A2 => n13, B1 => Q(81), B2 => n14, ZN
                           => n498);
   U522 : AOI22_X1 port map( A1 => Q(241), A2 => n15, B1 => Q(145), B2 => n16, 
                           ZN => n497);
   U523 : NAND4_X1 port map( A1 => n501, A2 => n502, A3 => n503, A4 => n504, ZN
                           => n495);
   U524 : AOI22_X1 port map( A1 => Q(337), A2 => n21, B1 => Q(433), B2 => n22, 
                           ZN => n504);
   U525 : AOI22_X1 port map( A1 => Q(401), A2 => n23, B1 => Q(273), B2 => n24, 
                           ZN => n503);
   U526 : AOI22_X1 port map( A1 => Q(369), A2 => n25, B1 => Q(305), B2 => n26, 
                           ZN => n502);
   U527 : AOI22_X1 port map( A1 => Q(657), A2 => n27, B1 => Q(465), B2 => n28, 
                           ZN => n501);
   U528 : NAND4_X1 port map( A1 => n505, A2 => n506, A3 => n507, A4 => n508, ZN
                           => n494);
   U529 : AOI22_X1 port map( A1 => Q(497), A2 => n33, B1 => Q(561), B2 => n34, 
                           ZN => n508);
   U530 : AOI22_X1 port map( A1 => Q(529), A2 => n35, B1 => Q(625), B2 => n36, 
                           ZN => n507);
   U531 : AOI22_X1 port map( A1 => Q(689), A2 => n37, B1 => Q(593), B2 => n38, 
                           ZN => n506);
   U532 : AOI22_X1 port map( A1 => Q(785), A2 => n39, B1 => Q(881), B2 => n40, 
                           ZN => n505);
   U533 : NAND4_X1 port map( A1 => n509, A2 => n510, A3 => n511, A4 => n512, ZN
                           => n493);
   U534 : AOI22_X1 port map( A1 => Q(849), A2 => n45, B1 => Q(721), B2 => n46, 
                           ZN => n512);
   U535 : AOI22_X1 port map( A1 => Q(817), A2 => n47, B1 => Q(753), B2 => n48, 
                           ZN => n511);
   U536 : AOI22_X1 port map( A1 => Q(977), A2 => n49, B1 => Q(913), B2 => n50, 
                           ZN => n510);
   U537 : AOI22_X1 port map( A1 => Q(1009), A2 => n51, B1 => Q(945), B2 => n52,
                           ZN => n509);
   U538 : OR4_X1 port map( A1 => n513, A2 => n514, A3 => n515, A4 => n516, ZN 
                           => Y(16));
   U539 : NAND4_X1 port map( A1 => n517, A2 => n518, A3 => n519, A4 => n520, ZN
                           => n516);
   U540 : AOI22_X1 port map( A1 => Q(112), A2 => n9, B1 => Q(208), B2 => n10, 
                           ZN => n520);
   U541 : AOI22_X1 port map( A1 => Q(176), A2 => n11, B1 => Q(48), B2 => n12, 
                           ZN => n519);
   U542 : AOI22_X1 port map( A1 => Q(16), A2 => n13, B1 => Q(80), B2 => n14, ZN
                           => n518);
   U543 : AOI22_X1 port map( A1 => Q(240), A2 => n15, B1 => Q(144), B2 => n16, 
                           ZN => n517);
   U544 : NAND4_X1 port map( A1 => n521, A2 => n522, A3 => n523, A4 => n524, ZN
                           => n515);
   U545 : AOI22_X1 port map( A1 => Q(336), A2 => n21, B1 => Q(432), B2 => n22, 
                           ZN => n524);
   U546 : AOI22_X1 port map( A1 => Q(400), A2 => n23, B1 => Q(272), B2 => n24, 
                           ZN => n523);
   U547 : AOI22_X1 port map( A1 => Q(368), A2 => n25, B1 => Q(304), B2 => n26, 
                           ZN => n522);
   U548 : AOI22_X1 port map( A1 => Q(656), A2 => n27, B1 => Q(464), B2 => n28, 
                           ZN => n521);
   U549 : NAND4_X1 port map( A1 => n525, A2 => n526, A3 => n527, A4 => n528, ZN
                           => n514);
   U550 : AOI22_X1 port map( A1 => Q(496), A2 => n33, B1 => Q(560), B2 => n34, 
                           ZN => n528);
   U551 : AOI22_X1 port map( A1 => Q(528), A2 => n35, B1 => Q(624), B2 => n36, 
                           ZN => n527);
   U552 : AOI22_X1 port map( A1 => Q(688), A2 => n37, B1 => Q(592), B2 => n38, 
                           ZN => n526);
   U553 : AOI22_X1 port map( A1 => Q(784), A2 => n39, B1 => Q(880), B2 => n40, 
                           ZN => n525);
   U554 : NAND4_X1 port map( A1 => n529, A2 => n530, A3 => n531, A4 => n532, ZN
                           => n513);
   U555 : AOI22_X1 port map( A1 => Q(848), A2 => n45, B1 => Q(720), B2 => n46, 
                           ZN => n532);
   U556 : AOI22_X1 port map( A1 => Q(816), A2 => n47, B1 => Q(752), B2 => n48, 
                           ZN => n531);
   U557 : AOI22_X1 port map( A1 => Q(976), A2 => n49, B1 => Q(912), B2 => n50, 
                           ZN => n530);
   U558 : AOI22_X1 port map( A1 => Q(1008), A2 => n51, B1 => Q(944), B2 => n52,
                           ZN => n529);
   U559 : OR4_X1 port map( A1 => n533, A2 => n534, A3 => n535, A4 => n536, ZN 
                           => Y(15));
   U560 : NAND4_X1 port map( A1 => n537, A2 => n538, A3 => n539, A4 => n540, ZN
                           => n536);
   U561 : AOI22_X1 port map( A1 => Q(111), A2 => n9, B1 => Q(207), B2 => n10, 
                           ZN => n540);
   U562 : AOI22_X1 port map( A1 => Q(175), A2 => n11, B1 => Q(47), B2 => n12, 
                           ZN => n539);
   U563 : AOI22_X1 port map( A1 => Q(15), A2 => n13, B1 => Q(79), B2 => n14, ZN
                           => n538);
   U564 : AOI22_X1 port map( A1 => Q(239), A2 => n15, B1 => Q(143), B2 => n16, 
                           ZN => n537);
   U565 : NAND4_X1 port map( A1 => n541, A2 => n542, A3 => n543, A4 => n544, ZN
                           => n535);
   U566 : AOI22_X1 port map( A1 => Q(335), A2 => n21, B1 => Q(431), B2 => n22, 
                           ZN => n544);
   U567 : AOI22_X1 port map( A1 => Q(399), A2 => n23, B1 => Q(271), B2 => n24, 
                           ZN => n543);
   U568 : AOI22_X1 port map( A1 => Q(367), A2 => n25, B1 => Q(303), B2 => n26, 
                           ZN => n542);
   U569 : AOI22_X1 port map( A1 => Q(655), A2 => n27, B1 => Q(463), B2 => n28, 
                           ZN => n541);
   U570 : NAND4_X1 port map( A1 => n545, A2 => n546, A3 => n547, A4 => n548, ZN
                           => n534);
   U571 : AOI22_X1 port map( A1 => Q(495), A2 => n33, B1 => Q(559), B2 => n34, 
                           ZN => n548);
   U572 : AOI22_X1 port map( A1 => Q(527), A2 => n35, B1 => Q(623), B2 => n36, 
                           ZN => n547);
   U573 : AOI22_X1 port map( A1 => Q(687), A2 => n37, B1 => Q(591), B2 => n38, 
                           ZN => n546);
   U574 : AOI22_X1 port map( A1 => Q(783), A2 => n39, B1 => Q(879), B2 => n40, 
                           ZN => n545);
   U575 : NAND4_X1 port map( A1 => n549, A2 => n550, A3 => n551, A4 => n552, ZN
                           => n533);
   U576 : AOI22_X1 port map( A1 => Q(847), A2 => n45, B1 => Q(719), B2 => n46, 
                           ZN => n552);
   U577 : AOI22_X1 port map( A1 => Q(815), A2 => n47, B1 => Q(751), B2 => n48, 
                           ZN => n551);
   U578 : AOI22_X1 port map( A1 => Q(975), A2 => n49, B1 => Q(911), B2 => n50, 
                           ZN => n550);
   U579 : AOI22_X1 port map( A1 => Q(1007), A2 => n51, B1 => Q(943), B2 => n52,
                           ZN => n549);
   U580 : OR4_X1 port map( A1 => n553, A2 => n554, A3 => n555, A4 => n556, ZN 
                           => Y(14));
   U581 : NAND4_X1 port map( A1 => n557, A2 => n558, A3 => n559, A4 => n560, ZN
                           => n556);
   U582 : AOI22_X1 port map( A1 => Q(110), A2 => n9, B1 => Q(206), B2 => n10, 
                           ZN => n560);
   U583 : AOI22_X1 port map( A1 => Q(174), A2 => n11, B1 => Q(46), B2 => n12, 
                           ZN => n559);
   U584 : AOI22_X1 port map( A1 => Q(14), A2 => n13, B1 => Q(78), B2 => n14, ZN
                           => n558);
   U585 : AOI22_X1 port map( A1 => Q(238), A2 => n15, B1 => Q(142), B2 => n16, 
                           ZN => n557);
   U586 : NAND4_X1 port map( A1 => n561, A2 => n562, A3 => n563, A4 => n564, ZN
                           => n555);
   U587 : AOI22_X1 port map( A1 => Q(334), A2 => n21, B1 => Q(430), B2 => n22, 
                           ZN => n564);
   U588 : AOI22_X1 port map( A1 => Q(398), A2 => n23, B1 => Q(270), B2 => n24, 
                           ZN => n563);
   U589 : AOI22_X1 port map( A1 => Q(366), A2 => n25, B1 => Q(302), B2 => n26, 
                           ZN => n562);
   U590 : AOI22_X1 port map( A1 => Q(654), A2 => n27, B1 => Q(462), B2 => n28, 
                           ZN => n561);
   U591 : NAND4_X1 port map( A1 => n565, A2 => n566, A3 => n567, A4 => n568, ZN
                           => n554);
   U592 : AOI22_X1 port map( A1 => Q(494), A2 => n33, B1 => Q(558), B2 => n34, 
                           ZN => n568);
   U593 : AOI22_X1 port map( A1 => Q(526), A2 => n35, B1 => Q(622), B2 => n36, 
                           ZN => n567);
   U594 : AOI22_X1 port map( A1 => Q(686), A2 => n37, B1 => Q(590), B2 => n38, 
                           ZN => n566);
   U595 : AOI22_X1 port map( A1 => Q(782), A2 => n39, B1 => Q(878), B2 => n40, 
                           ZN => n565);
   U596 : NAND4_X1 port map( A1 => n569, A2 => n570, A3 => n571, A4 => n572, ZN
                           => n553);
   U597 : AOI22_X1 port map( A1 => Q(846), A2 => n45, B1 => Q(718), B2 => n46, 
                           ZN => n572);
   U598 : AOI22_X1 port map( A1 => Q(814), A2 => n47, B1 => Q(750), B2 => n48, 
                           ZN => n571);
   U599 : AOI22_X1 port map( A1 => Q(974), A2 => n49, B1 => Q(910), B2 => n50, 
                           ZN => n570);
   U600 : AOI22_X1 port map( A1 => Q(1006), A2 => n51, B1 => Q(942), B2 => n52,
                           ZN => n569);
   U601 : OR4_X1 port map( A1 => n573, A2 => n574, A3 => n575, A4 => n576, ZN 
                           => Y(13));
   U602 : NAND4_X1 port map( A1 => n577, A2 => n578, A3 => n579, A4 => n580, ZN
                           => n576);
   U603 : AOI22_X1 port map( A1 => Q(109), A2 => n9, B1 => Q(205), B2 => n10, 
                           ZN => n580);
   U604 : AOI22_X1 port map( A1 => Q(173), A2 => n11, B1 => Q(45), B2 => n12, 
                           ZN => n579);
   U605 : AOI22_X1 port map( A1 => Q(13), A2 => n13, B1 => Q(77), B2 => n14, ZN
                           => n578);
   U606 : AOI22_X1 port map( A1 => Q(237), A2 => n15, B1 => Q(141), B2 => n16, 
                           ZN => n577);
   U607 : NAND4_X1 port map( A1 => n581, A2 => n582, A3 => n583, A4 => n584, ZN
                           => n575);
   U608 : AOI22_X1 port map( A1 => Q(333), A2 => n21, B1 => Q(429), B2 => n22, 
                           ZN => n584);
   U609 : AOI22_X1 port map( A1 => Q(397), A2 => n23, B1 => Q(269), B2 => n24, 
                           ZN => n583);
   U610 : AOI22_X1 port map( A1 => Q(365), A2 => n25, B1 => Q(301), B2 => n26, 
                           ZN => n582);
   U611 : AOI22_X1 port map( A1 => Q(653), A2 => n27, B1 => Q(461), B2 => n28, 
                           ZN => n581);
   U612 : NAND4_X1 port map( A1 => n585, A2 => n586, A3 => n587, A4 => n588, ZN
                           => n574);
   U613 : AOI22_X1 port map( A1 => Q(493), A2 => n33, B1 => Q(557), B2 => n34, 
                           ZN => n588);
   U614 : AOI22_X1 port map( A1 => Q(525), A2 => n35, B1 => Q(621), B2 => n36, 
                           ZN => n587);
   U615 : AOI22_X1 port map( A1 => Q(685), A2 => n37, B1 => Q(589), B2 => n38, 
                           ZN => n586);
   U616 : AOI22_X1 port map( A1 => Q(781), A2 => n39, B1 => Q(877), B2 => n40, 
                           ZN => n585);
   U617 : NAND4_X1 port map( A1 => n589, A2 => n590, A3 => n591, A4 => n592, ZN
                           => n573);
   U618 : AOI22_X1 port map( A1 => Q(845), A2 => n45, B1 => Q(717), B2 => n46, 
                           ZN => n592);
   U619 : AOI22_X1 port map( A1 => Q(813), A2 => n47, B1 => Q(749), B2 => n48, 
                           ZN => n591);
   U620 : AOI22_X1 port map( A1 => Q(973), A2 => n49, B1 => Q(909), B2 => n50, 
                           ZN => n590);
   U621 : AOI22_X1 port map( A1 => Q(1005), A2 => n51, B1 => Q(941), B2 => n52,
                           ZN => n589);
   U622 : OR4_X1 port map( A1 => n593, A2 => n594, A3 => n595, A4 => n596, ZN 
                           => Y(12));
   U623 : NAND4_X1 port map( A1 => n597, A2 => n598, A3 => n599, A4 => n600, ZN
                           => n596);
   U624 : AOI22_X1 port map( A1 => Q(108), A2 => n9, B1 => Q(204), B2 => n10, 
                           ZN => n600);
   U625 : AOI22_X1 port map( A1 => Q(172), A2 => n11, B1 => Q(44), B2 => n12, 
                           ZN => n599);
   U626 : AOI22_X1 port map( A1 => Q(12), A2 => n13, B1 => Q(76), B2 => n14, ZN
                           => n598);
   U627 : AOI22_X1 port map( A1 => Q(236), A2 => n15, B1 => Q(140), B2 => n16, 
                           ZN => n597);
   U628 : NAND4_X1 port map( A1 => n601, A2 => n602, A3 => n603, A4 => n604, ZN
                           => n595);
   U629 : AOI22_X1 port map( A1 => Q(332), A2 => n21, B1 => Q(428), B2 => n22, 
                           ZN => n604);
   U630 : AOI22_X1 port map( A1 => Q(396), A2 => n23, B1 => Q(268), B2 => n24, 
                           ZN => n603);
   U631 : AOI22_X1 port map( A1 => Q(364), A2 => n25, B1 => Q(300), B2 => n26, 
                           ZN => n602);
   U632 : AOI22_X1 port map( A1 => Q(652), A2 => n27, B1 => Q(460), B2 => n28, 
                           ZN => n601);
   U633 : NAND4_X1 port map( A1 => n605, A2 => n606, A3 => n607, A4 => n608, ZN
                           => n594);
   U634 : AOI22_X1 port map( A1 => Q(492), A2 => n33, B1 => Q(556), B2 => n34, 
                           ZN => n608);
   U635 : AOI22_X1 port map( A1 => Q(524), A2 => n35, B1 => Q(620), B2 => n36, 
                           ZN => n607);
   U636 : AOI22_X1 port map( A1 => Q(684), A2 => n37, B1 => Q(588), B2 => n38, 
                           ZN => n606);
   U637 : AOI22_X1 port map( A1 => Q(780), A2 => n39, B1 => Q(876), B2 => n40, 
                           ZN => n605);
   U638 : NAND4_X1 port map( A1 => n609, A2 => n610, A3 => n611, A4 => n612, ZN
                           => n593);
   U639 : AOI22_X1 port map( A1 => Q(844), A2 => n45, B1 => Q(716), B2 => n46, 
                           ZN => n612);
   U640 : AOI22_X1 port map( A1 => Q(812), A2 => n47, B1 => Q(748), B2 => n48, 
                           ZN => n611);
   U641 : AOI22_X1 port map( A1 => Q(972), A2 => n49, B1 => Q(908), B2 => n50, 
                           ZN => n610);
   U642 : AOI22_X1 port map( A1 => Q(1004), A2 => n51, B1 => Q(940), B2 => n52,
                           ZN => n609);
   U643 : OR4_X1 port map( A1 => n613, A2 => n614, A3 => n615, A4 => n616, ZN 
                           => Y(11));
   U644 : NAND4_X1 port map( A1 => n617, A2 => n618, A3 => n619, A4 => n620, ZN
                           => n616);
   U645 : AOI22_X1 port map( A1 => Q(107), A2 => n9, B1 => Q(203), B2 => n10, 
                           ZN => n620);
   U646 : AOI22_X1 port map( A1 => Q(171), A2 => n11, B1 => Q(43), B2 => n12, 
                           ZN => n619);
   U647 : AOI22_X1 port map( A1 => Q(11), A2 => n13, B1 => Q(75), B2 => n14, ZN
                           => n618);
   U648 : AOI22_X1 port map( A1 => Q(235), A2 => n15, B1 => Q(139), B2 => n16, 
                           ZN => n617);
   U649 : NAND4_X1 port map( A1 => n621, A2 => n622, A3 => n623, A4 => n624, ZN
                           => n615);
   U650 : AOI22_X1 port map( A1 => Q(331), A2 => n21, B1 => Q(427), B2 => n22, 
                           ZN => n624);
   U651 : AOI22_X1 port map( A1 => Q(395), A2 => n23, B1 => Q(267), B2 => n24, 
                           ZN => n623);
   U652 : AOI22_X1 port map( A1 => Q(363), A2 => n25, B1 => Q(299), B2 => n26, 
                           ZN => n622);
   U653 : AOI22_X1 port map( A1 => Q(651), A2 => n27, B1 => Q(459), B2 => n28, 
                           ZN => n621);
   U654 : NAND4_X1 port map( A1 => n625, A2 => n626, A3 => n627, A4 => n628, ZN
                           => n614);
   U655 : AOI22_X1 port map( A1 => Q(491), A2 => n33, B1 => Q(555), B2 => n34, 
                           ZN => n628);
   U656 : AOI22_X1 port map( A1 => Q(523), A2 => n35, B1 => Q(619), B2 => n36, 
                           ZN => n627);
   U657 : AOI22_X1 port map( A1 => Q(683), A2 => n37, B1 => Q(587), B2 => n38, 
                           ZN => n626);
   U658 : AOI22_X1 port map( A1 => Q(779), A2 => n39, B1 => Q(875), B2 => n40, 
                           ZN => n625);
   U659 : NAND4_X1 port map( A1 => n629, A2 => n630, A3 => n631, A4 => n632, ZN
                           => n613);
   U660 : AOI22_X1 port map( A1 => Q(843), A2 => n45, B1 => Q(715), B2 => n46, 
                           ZN => n632);
   U661 : AOI22_X1 port map( A1 => Q(811), A2 => n47, B1 => Q(747), B2 => n48, 
                           ZN => n631);
   U662 : AOI22_X1 port map( A1 => Q(971), A2 => n49, B1 => Q(907), B2 => n50, 
                           ZN => n630);
   U663 : AOI22_X1 port map( A1 => Q(1003), A2 => n51, B1 => Q(939), B2 => n52,
                           ZN => n629);
   U664 : OR4_X1 port map( A1 => n633, A2 => n634, A3 => n635, A4 => n636, ZN 
                           => Y(10));
   U665 : NAND4_X1 port map( A1 => n637, A2 => n638, A3 => n639, A4 => n640, ZN
                           => n636);
   U666 : AOI22_X1 port map( A1 => Q(106), A2 => n9, B1 => Q(202), B2 => n10, 
                           ZN => n640);
   U667 : AOI22_X1 port map( A1 => Q(170), A2 => n11, B1 => Q(42), B2 => n12, 
                           ZN => n639);
   U668 : AOI22_X1 port map( A1 => Q(10), A2 => n13, B1 => Q(74), B2 => n14, ZN
                           => n638);
   U669 : AOI22_X1 port map( A1 => Q(234), A2 => n15, B1 => Q(138), B2 => n16, 
                           ZN => n637);
   U670 : NAND4_X1 port map( A1 => n641, A2 => n642, A3 => n643, A4 => n644, ZN
                           => n635);
   U671 : AOI22_X1 port map( A1 => Q(330), A2 => n21, B1 => Q(426), B2 => n22, 
                           ZN => n644);
   U672 : AOI22_X1 port map( A1 => Q(394), A2 => n23, B1 => Q(266), B2 => n24, 
                           ZN => n643);
   U673 : AOI22_X1 port map( A1 => Q(362), A2 => n25, B1 => Q(298), B2 => n26, 
                           ZN => n642);
   U674 : AOI22_X1 port map( A1 => Q(650), A2 => n27, B1 => Q(458), B2 => n28, 
                           ZN => n641);
   U675 : NAND4_X1 port map( A1 => n645, A2 => n646, A3 => n647, A4 => n648, ZN
                           => n634);
   U676 : AOI22_X1 port map( A1 => Q(490), A2 => n33, B1 => Q(554), B2 => n34, 
                           ZN => n648);
   U677 : AOI22_X1 port map( A1 => Q(522), A2 => n35, B1 => Q(618), B2 => n36, 
                           ZN => n647);
   U678 : AOI22_X1 port map( A1 => Q(682), A2 => n37, B1 => Q(586), B2 => n38, 
                           ZN => n646);
   U679 : AOI22_X1 port map( A1 => Q(778), A2 => n39, B1 => Q(874), B2 => n40, 
                           ZN => n645);
   U680 : NAND4_X1 port map( A1 => n649, A2 => n650, A3 => n651, A4 => n652, ZN
                           => n633);
   U681 : AOI22_X1 port map( A1 => Q(842), A2 => n45, B1 => Q(714), B2 => n46, 
                           ZN => n652);
   U682 : AOI22_X1 port map( A1 => Q(810), A2 => n47, B1 => Q(746), B2 => n48, 
                           ZN => n651);
   U683 : AOI22_X1 port map( A1 => Q(970), A2 => n49, B1 => Q(906), B2 => n50, 
                           ZN => n650);
   U684 : AOI22_X1 port map( A1 => Q(1002), A2 => n51, B1 => Q(938), B2 => n52,
                           ZN => n649);
   U685 : OR4_X1 port map( A1 => n653, A2 => n654, A3 => n655, A4 => n656, ZN 
                           => Y(0));
   U686 : NAND4_X1 port map( A1 => n657, A2 => n658, A3 => n659, A4 => n660, ZN
                           => n656);
   U687 : AOI22_X1 port map( A1 => Q(96), A2 => n9, B1 => Q(192), B2 => n10, ZN
                           => n660);
   U688 : AOI22_X1 port map( A1 => Q(160), A2 => n11, B1 => Q(32), B2 => n12, 
                           ZN => n659);
   U689 : AOI22_X1 port map( A1 => Q(0), A2 => n13, B1 => Q(64), B2 => n14, ZN 
                           => n658);
   U690 : AOI22_X1 port map( A1 => Q(224), A2 => n15, B1 => Q(128), B2 => n16, 
                           ZN => n657);
   U691 : NOR3_X1 port map( A1 => S(3), A2 => S(4), A3 => S(0), ZN => n661);
   U692 : NOR3_X1 port map( A1 => S(3), A2 => S(4), A3 => n667, ZN => n663);
   U693 : NAND4_X1 port map( A1 => n668, A2 => n669, A3 => n670, A4 => n671, ZN
                           => n655);
   U694 : AOI22_X1 port map( A1 => Q(320), A2 => n21, B1 => Q(416), B2 => n22, 
                           ZN => n671);
   U695 : AOI22_X1 port map( A1 => Q(384), A2 => n23, B1 => Q(256), B2 => n24, 
                           ZN => n670);
   U696 : AOI22_X1 port map( A1 => Q(352), A2 => n25, B1 => Q(288), B2 => n26, 
                           ZN => n669);
   U697 : AOI22_X1 port map( A1 => Q(640), A2 => n27, B1 => Q(448), B2 => n28, 
                           ZN => n668);
   U698 : NOR3_X1 port map( A1 => S(0), A2 => S(4), A3 => n674, ZN => n673);
   U699 : NAND4_X1 port map( A1 => n676, A2 => n677, A3 => n678, A4 => n679, ZN
                           => n654);
   U700 : AOI22_X1 port map( A1 => Q(480), A2 => n33, B1 => Q(544), B2 => n34, 
                           ZN => n679);
   U701 : NOR3_X1 port map( A1 => n674, A2 => S(4), A3 => n667, ZN => n672);
   U702 : AOI22_X1 port map( A1 => Q(512), A2 => n35, B1 => Q(608), B2 => n36, 
                           ZN => n678);
   U703 : AOI22_X1 port map( A1 => Q(672), A2 => n37, B1 => Q(576), B2 => n38, 
                           ZN => n677);
   U704 : AOI22_X1 port map( A1 => Q(768), A2 => n39, B1 => Q(864), B2 => n40, 
                           ZN => n676);
   U705 : NAND4_X1 port map( A1 => n683, A2 => n684, A3 => n685, A4 => n686, ZN
                           => n653);
   U706 : AOI22_X1 port map( A1 => Q(832), A2 => n45, B1 => Q(704), B2 => n46, 
                           ZN => n686);
   U707 : NOR3_X1 port map( A1 => S(0), A2 => S(3), A3 => n687, ZN => n675);
   U708 : NOR2_X1 port map( A1 => n688, A2 => S(2), ZN => n664);
   U709 : AOI22_X1 port map( A1 => Q(800), A2 => n47, B1 => Q(736), B2 => n48, 
                           ZN => n685);
   U710 : NOR3_X1 port map( A1 => n667, A2 => S(3), A3 => n687, ZN => n680);
   U711 : NOR2_X1 port map( A1 => S(1), A2 => S(2), ZN => n665);
   U712 : AOI22_X1 port map( A1 => Q(960), A2 => n49, B1 => Q(896), B2 => n50, 
                           ZN => n684);
   U713 : NOR3_X1 port map( A1 => n674, A2 => S(0), A3 => n687, ZN => n682);
   U714 : AOI22_X1 port map( A1 => Q(992), A2 => n51, B1 => Q(928), B2 => n52, 
                           ZN => n683);
   U715 : NOR2_X1 port map( A1 => n689, A2 => S(1), ZN => n666);
   U716 : NOR2_X1 port map( A1 => n689, A2 => n688, ZN => n662);
   U717 : INV_X1 port map( A => S(1), ZN => n688);
   U718 : INV_X1 port map( A => S(2), ZN => n689);
   U719 : NOR3_X1 port map( A1 => n667, A2 => n674, A3 => n687, ZN => n681);
   U720 : INV_X1 port map( A => S(4), ZN => n687);
   U721 : INV_X1 port map( A => S(3), ZN => n674);
   U722 : INV_X1 port map( A => S(0), ZN => n667);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity select_block_NBIT_DATA32_N8_F5 is

   port( regs : in std_logic_vector (2559 downto 0);  win : in std_logic_vector
         (4 downto 0);  curr_proc_regs : out std_logic_vector (767 downto 0));

end select_block_NBIT_DATA32_N8_F5;

architecture SYN_behav of select_block_NBIT_DATA32_N8_F5 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
      n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
      n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
      n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
      n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
      n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
      n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
      n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
      n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
      n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
      n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
      n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
      n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
      n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
      n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
      n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
      n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
      n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432 : 
      std_logic;

begin
   
   U2 : BUF_X1 port map( A => n382, Z => n221);
   U3 : BUF_X1 port map( A => n382, Z => n216);
   U4 : BUF_X1 port map( A => n382, Z => n219);
   U5 : BUF_X1 port map( A => n382, Z => n218);
   U6 : BUF_X1 port map( A => n382, Z => n217);
   U7 : BUF_X1 port map( A => n382, Z => n215);
   U8 : BUF_X1 port map( A => n382, Z => n220);
   U9 : BUF_X1 port map( A => n382, Z => n222);
   U10 : BUF_X1 port map( A => n382, Z => n224);
   U11 : BUF_X1 port map( A => n382, Z => n223);
   U12 : BUF_X1 port map( A => n382, Z => n225);
   U13 : BUF_X1 port map( A => n381, Z => n146);
   U14 : BUF_X1 port map( A => n381, Z => n148);
   U15 : BUF_X1 port map( A => n381, Z => n149);
   U16 : BUF_X1 port map( A => n381, Z => n145);
   U17 : BUF_X1 port map( A => n381, Z => n147);
   U18 : BUF_X1 port map( A => n381, Z => n141);
   U19 : BUF_X1 port map( A => n381, Z => n142);
   U20 : BUF_X1 port map( A => n381, Z => n140);
   U21 : BUF_X1 port map( A => n381, Z => n143);
   U22 : BUF_X1 port map( A => n381, Z => n144);
   U23 : BUF_X1 port map( A => n383, Z => n296);
   U24 : BUF_X1 port map( A => n383, Z => n291);
   U25 : BUF_X1 port map( A => n383, Z => n294);
   U26 : BUF_X1 port map( A => n383, Z => n293);
   U27 : BUF_X1 port map( A => n383, Z => n292);
   U28 : BUF_X1 port map( A => n383, Z => n290);
   U29 : BUF_X1 port map( A => n383, Z => n295);
   U30 : BUF_X1 port map( A => n383, Z => n297);
   U31 : BUF_X1 port map( A => n383, Z => n299);
   U32 : BUF_X1 port map( A => n383, Z => n298);
   U33 : BUF_X1 port map( A => n378, Z => n70);
   U34 : BUF_X1 port map( A => n378, Z => n66);
   U35 : BUF_X1 port map( A => n378, Z => n67);
   U36 : BUF_X1 port map( A => n378, Z => n73);
   U37 : BUF_X1 port map( A => n378, Z => n74);
   U38 : BUF_X1 port map( A => n378, Z => n72);
   U39 : BUF_X1 port map( A => n378, Z => n65);
   U40 : BUF_X1 port map( A => n378, Z => n71);
   U41 : BUF_X1 port map( A => n378, Z => n69);
   U42 : BUF_X1 port map( A => n378, Z => n68);
   U43 : BUF_X1 port map( A => n381, Z => n150);
   U44 : BUF_X1 port map( A => n383, Z => n300);
   U45 : BUF_X1 port map( A => n378, Z => n75);
   U46 : BUF_X1 port map( A => win(4), Z => n374);
   U47 : BUF_X1 port map( A => win(4), Z => n368);
   U48 : BUF_X1 port map( A => win(4), Z => n367);
   U49 : BUF_X1 port map( A => win(4), Z => n369);
   U50 : BUF_X1 port map( A => win(4), Z => n373);
   U51 : BUF_X1 port map( A => win(4), Z => n371);
   U52 : BUF_X1 port map( A => win(4), Z => n370);
   U53 : BUF_X1 port map( A => win(4), Z => n372);
   U54 : BUF_X1 port map( A => win(4), Z => n366);
   U55 : BUF_X1 port map( A => win(4), Z => n375);
   U56 : BUF_X1 port map( A => win(4), Z => n376);
   U57 : CLKBUF_X1 port map( A => n75, Z => n1);
   U58 : CLKBUF_X1 port map( A => n75, Z => n2);
   U59 : CLKBUF_X1 port map( A => n75, Z => n3);
   U60 : CLKBUF_X1 port map( A => n75, Z => n4);
   U61 : CLKBUF_X1 port map( A => n74, Z => n5);
   U62 : CLKBUF_X1 port map( A => n74, Z => n6);
   U63 : CLKBUF_X1 port map( A => n74, Z => n7);
   U64 : CLKBUF_X1 port map( A => n74, Z => n8);
   U65 : CLKBUF_X1 port map( A => n74, Z => n9);
   U66 : CLKBUF_X1 port map( A => n74, Z => n10);
   U67 : CLKBUF_X1 port map( A => n73, Z => n11);
   U68 : CLKBUF_X1 port map( A => n73, Z => n12);
   U69 : CLKBUF_X1 port map( A => n73, Z => n13);
   U70 : CLKBUF_X1 port map( A => n73, Z => n14);
   U71 : CLKBUF_X1 port map( A => n73, Z => n15);
   U72 : CLKBUF_X1 port map( A => n73, Z => n16);
   U73 : CLKBUF_X1 port map( A => n72, Z => n17);
   U74 : CLKBUF_X1 port map( A => n72, Z => n18);
   U75 : CLKBUF_X1 port map( A => n72, Z => n19);
   U76 : CLKBUF_X1 port map( A => n72, Z => n20);
   U77 : CLKBUF_X1 port map( A => n72, Z => n21);
   U78 : CLKBUF_X1 port map( A => n72, Z => n22);
   U79 : CLKBUF_X1 port map( A => n71, Z => n23);
   U80 : CLKBUF_X1 port map( A => n71, Z => n24);
   U81 : CLKBUF_X1 port map( A => n71, Z => n25);
   U82 : CLKBUF_X1 port map( A => n71, Z => n26);
   U83 : CLKBUF_X1 port map( A => n71, Z => n27);
   U84 : CLKBUF_X1 port map( A => n71, Z => n28);
   U85 : CLKBUF_X1 port map( A => n70, Z => n29);
   U86 : CLKBUF_X1 port map( A => n70, Z => n30);
   U87 : CLKBUF_X1 port map( A => n70, Z => n31);
   U88 : CLKBUF_X1 port map( A => n70, Z => n32);
   U89 : CLKBUF_X1 port map( A => n70, Z => n33);
   U90 : CLKBUF_X1 port map( A => n70, Z => n34);
   U91 : CLKBUF_X1 port map( A => n69, Z => n35);
   U92 : CLKBUF_X1 port map( A => n69, Z => n36);
   U93 : CLKBUF_X1 port map( A => n69, Z => n37);
   U94 : CLKBUF_X1 port map( A => n69, Z => n38);
   U95 : CLKBUF_X1 port map( A => n69, Z => n39);
   U96 : CLKBUF_X1 port map( A => n69, Z => n40);
   U97 : CLKBUF_X1 port map( A => n68, Z => n41);
   U98 : CLKBUF_X1 port map( A => n68, Z => n42);
   U99 : CLKBUF_X1 port map( A => n68, Z => n43);
   U100 : CLKBUF_X1 port map( A => n68, Z => n44);
   U101 : CLKBUF_X1 port map( A => n68, Z => n45);
   U102 : CLKBUF_X1 port map( A => n68, Z => n46);
   U103 : CLKBUF_X1 port map( A => n67, Z => n47);
   U104 : CLKBUF_X1 port map( A => n67, Z => n48);
   U105 : CLKBUF_X1 port map( A => n67, Z => n49);
   U106 : CLKBUF_X1 port map( A => n67, Z => n50);
   U107 : CLKBUF_X1 port map( A => n67, Z => n51);
   U108 : CLKBUF_X1 port map( A => n67, Z => n52);
   U109 : CLKBUF_X1 port map( A => n66, Z => n53);
   U110 : CLKBUF_X1 port map( A => n66, Z => n54);
   U111 : CLKBUF_X1 port map( A => n66, Z => n55);
   U112 : CLKBUF_X1 port map( A => n66, Z => n56);
   U113 : CLKBUF_X1 port map( A => n66, Z => n57);
   U114 : CLKBUF_X1 port map( A => n66, Z => n58);
   U115 : CLKBUF_X1 port map( A => n65, Z => n59);
   U116 : CLKBUF_X1 port map( A => n65, Z => n60);
   U117 : CLKBUF_X1 port map( A => n65, Z => n61);
   U118 : CLKBUF_X1 port map( A => n65, Z => n62);
   U119 : CLKBUF_X1 port map( A => n65, Z => n63);
   U120 : CLKBUF_X1 port map( A => n65, Z => n64);
   U121 : CLKBUF_X1 port map( A => n150, Z => n76);
   U122 : CLKBUF_X1 port map( A => n150, Z => n77);
   U123 : CLKBUF_X1 port map( A => n150, Z => n78);
   U124 : CLKBUF_X1 port map( A => n150, Z => n79);
   U125 : CLKBUF_X1 port map( A => n149, Z => n80);
   U126 : CLKBUF_X1 port map( A => n149, Z => n81);
   U127 : CLKBUF_X1 port map( A => n149, Z => n82);
   U128 : CLKBUF_X1 port map( A => n149, Z => n83);
   U129 : CLKBUF_X1 port map( A => n149, Z => n84);
   U130 : CLKBUF_X1 port map( A => n149, Z => n85);
   U131 : CLKBUF_X1 port map( A => n148, Z => n86);
   U132 : CLKBUF_X1 port map( A => n148, Z => n87);
   U133 : CLKBUF_X1 port map( A => n148, Z => n88);
   U134 : CLKBUF_X1 port map( A => n148, Z => n89);
   U135 : CLKBUF_X1 port map( A => n148, Z => n90);
   U136 : CLKBUF_X1 port map( A => n148, Z => n91);
   U137 : CLKBUF_X1 port map( A => n147, Z => n92);
   U138 : CLKBUF_X1 port map( A => n147, Z => n93);
   U139 : CLKBUF_X1 port map( A => n147, Z => n94);
   U140 : CLKBUF_X1 port map( A => n147, Z => n95);
   U141 : CLKBUF_X1 port map( A => n147, Z => n96);
   U142 : CLKBUF_X1 port map( A => n147, Z => n97);
   U143 : CLKBUF_X1 port map( A => n146, Z => n98);
   U144 : CLKBUF_X1 port map( A => n146, Z => n99);
   U145 : CLKBUF_X1 port map( A => n146, Z => n100);
   U146 : CLKBUF_X1 port map( A => n146, Z => n101);
   U147 : CLKBUF_X1 port map( A => n146, Z => n102);
   U148 : CLKBUF_X1 port map( A => n146, Z => n103);
   U149 : CLKBUF_X1 port map( A => n145, Z => n104);
   U150 : CLKBUF_X1 port map( A => n145, Z => n105);
   U151 : CLKBUF_X1 port map( A => n145, Z => n106);
   U152 : CLKBUF_X1 port map( A => n145, Z => n107);
   U153 : CLKBUF_X1 port map( A => n145, Z => n108);
   U154 : CLKBUF_X1 port map( A => n145, Z => n109);
   U155 : CLKBUF_X1 port map( A => n144, Z => n110);
   U156 : CLKBUF_X1 port map( A => n144, Z => n111);
   U157 : CLKBUF_X1 port map( A => n144, Z => n112);
   U158 : CLKBUF_X1 port map( A => n144, Z => n113);
   U159 : CLKBUF_X1 port map( A => n144, Z => n114);
   U160 : CLKBUF_X1 port map( A => n144, Z => n115);
   U161 : CLKBUF_X1 port map( A => n143, Z => n116);
   U162 : CLKBUF_X1 port map( A => n143, Z => n117);
   U163 : CLKBUF_X1 port map( A => n143, Z => n118);
   U164 : CLKBUF_X1 port map( A => n143, Z => n119);
   U165 : CLKBUF_X1 port map( A => n143, Z => n120);
   U166 : CLKBUF_X1 port map( A => n143, Z => n121);
   U167 : CLKBUF_X1 port map( A => n142, Z => n122);
   U168 : CLKBUF_X1 port map( A => n142, Z => n123);
   U169 : CLKBUF_X1 port map( A => n142, Z => n124);
   U170 : CLKBUF_X1 port map( A => n142, Z => n125);
   U171 : CLKBUF_X1 port map( A => n142, Z => n126);
   U172 : CLKBUF_X1 port map( A => n142, Z => n127);
   U173 : CLKBUF_X1 port map( A => n141, Z => n128);
   U174 : CLKBUF_X1 port map( A => n141, Z => n129);
   U175 : CLKBUF_X1 port map( A => n141, Z => n130);
   U176 : CLKBUF_X1 port map( A => n141, Z => n131);
   U177 : CLKBUF_X1 port map( A => n141, Z => n132);
   U178 : CLKBUF_X1 port map( A => n141, Z => n133);
   U179 : CLKBUF_X1 port map( A => n140, Z => n134);
   U180 : CLKBUF_X1 port map( A => n140, Z => n135);
   U181 : CLKBUF_X1 port map( A => n140, Z => n136);
   U182 : CLKBUF_X1 port map( A => n140, Z => n137);
   U183 : CLKBUF_X1 port map( A => n140, Z => n138);
   U184 : CLKBUF_X1 port map( A => n140, Z => n139);
   U185 : CLKBUF_X1 port map( A => n225, Z => n151);
   U186 : CLKBUF_X1 port map( A => n225, Z => n152);
   U187 : CLKBUF_X1 port map( A => n225, Z => n153);
   U188 : CLKBUF_X1 port map( A => n225, Z => n154);
   U189 : CLKBUF_X1 port map( A => n224, Z => n155);
   U190 : CLKBUF_X1 port map( A => n224, Z => n156);
   U191 : CLKBUF_X1 port map( A => n224, Z => n157);
   U192 : CLKBUF_X1 port map( A => n224, Z => n158);
   U193 : CLKBUF_X1 port map( A => n224, Z => n159);
   U194 : CLKBUF_X1 port map( A => n224, Z => n160);
   U195 : CLKBUF_X1 port map( A => n223, Z => n161);
   U196 : CLKBUF_X1 port map( A => n223, Z => n162);
   U197 : CLKBUF_X1 port map( A => n223, Z => n163);
   U198 : CLKBUF_X1 port map( A => n223, Z => n164);
   U199 : CLKBUF_X1 port map( A => n223, Z => n165);
   U200 : CLKBUF_X1 port map( A => n223, Z => n166);
   U201 : CLKBUF_X1 port map( A => n222, Z => n167);
   U202 : CLKBUF_X1 port map( A => n222, Z => n168);
   U203 : CLKBUF_X1 port map( A => n222, Z => n169);
   U204 : CLKBUF_X1 port map( A => n222, Z => n170);
   U205 : CLKBUF_X1 port map( A => n222, Z => n171);
   U206 : CLKBUF_X1 port map( A => n222, Z => n172);
   U207 : CLKBUF_X1 port map( A => n221, Z => n173);
   U208 : CLKBUF_X1 port map( A => n221, Z => n174);
   U209 : CLKBUF_X1 port map( A => n221, Z => n175);
   U210 : CLKBUF_X1 port map( A => n221, Z => n176);
   U211 : CLKBUF_X1 port map( A => n221, Z => n177);
   U212 : CLKBUF_X1 port map( A => n221, Z => n178);
   U213 : CLKBUF_X1 port map( A => n220, Z => n179);
   U214 : CLKBUF_X1 port map( A => n220, Z => n180);
   U215 : CLKBUF_X1 port map( A => n220, Z => n181);
   U216 : CLKBUF_X1 port map( A => n220, Z => n182);
   U217 : CLKBUF_X1 port map( A => n220, Z => n183);
   U218 : CLKBUF_X1 port map( A => n220, Z => n184);
   U219 : CLKBUF_X1 port map( A => n219, Z => n185);
   U220 : CLKBUF_X1 port map( A => n219, Z => n186);
   U221 : CLKBUF_X1 port map( A => n219, Z => n187);
   U222 : CLKBUF_X1 port map( A => n219, Z => n188);
   U223 : CLKBUF_X1 port map( A => n219, Z => n189);
   U224 : CLKBUF_X1 port map( A => n219, Z => n190);
   U225 : CLKBUF_X1 port map( A => n218, Z => n191);
   U226 : CLKBUF_X1 port map( A => n218, Z => n192);
   U227 : CLKBUF_X1 port map( A => n218, Z => n193);
   U228 : CLKBUF_X1 port map( A => n218, Z => n194);
   U229 : CLKBUF_X1 port map( A => n218, Z => n195);
   U230 : CLKBUF_X1 port map( A => n218, Z => n196);
   U231 : CLKBUF_X1 port map( A => n217, Z => n197);
   U232 : CLKBUF_X1 port map( A => n217, Z => n198);
   U233 : CLKBUF_X1 port map( A => n217, Z => n199);
   U234 : CLKBUF_X1 port map( A => n217, Z => n200);
   U235 : CLKBUF_X1 port map( A => n217, Z => n201);
   U236 : CLKBUF_X1 port map( A => n217, Z => n202);
   U237 : CLKBUF_X1 port map( A => n216, Z => n203);
   U238 : CLKBUF_X1 port map( A => n216, Z => n204);
   U239 : CLKBUF_X1 port map( A => n216, Z => n205);
   U240 : CLKBUF_X1 port map( A => n216, Z => n206);
   U241 : CLKBUF_X1 port map( A => n216, Z => n207);
   U242 : CLKBUF_X1 port map( A => n216, Z => n208);
   U243 : CLKBUF_X1 port map( A => n215, Z => n209);
   U244 : CLKBUF_X1 port map( A => n215, Z => n210);
   U245 : CLKBUF_X1 port map( A => n215, Z => n211);
   U246 : CLKBUF_X1 port map( A => n215, Z => n212);
   U247 : CLKBUF_X1 port map( A => n215, Z => n213);
   U248 : CLKBUF_X1 port map( A => n215, Z => n214);
   U249 : CLKBUF_X1 port map( A => n300, Z => n226);
   U250 : CLKBUF_X1 port map( A => n300, Z => n227);
   U251 : CLKBUF_X1 port map( A => n300, Z => n228);
   U252 : CLKBUF_X1 port map( A => n300, Z => n229);
   U253 : CLKBUF_X1 port map( A => n299, Z => n230);
   U254 : CLKBUF_X1 port map( A => n299, Z => n231);
   U255 : CLKBUF_X1 port map( A => n299, Z => n232);
   U256 : CLKBUF_X1 port map( A => n299, Z => n233);
   U257 : CLKBUF_X1 port map( A => n299, Z => n234);
   U258 : CLKBUF_X1 port map( A => n299, Z => n235);
   U259 : CLKBUF_X1 port map( A => n298, Z => n236);
   U260 : CLKBUF_X1 port map( A => n298, Z => n237);
   U261 : CLKBUF_X1 port map( A => n298, Z => n238);
   U262 : CLKBUF_X1 port map( A => n298, Z => n239);
   U263 : CLKBUF_X1 port map( A => n298, Z => n240);
   U264 : CLKBUF_X1 port map( A => n298, Z => n241);
   U265 : CLKBUF_X1 port map( A => n297, Z => n242);
   U266 : CLKBUF_X1 port map( A => n297, Z => n243);
   U267 : CLKBUF_X1 port map( A => n297, Z => n244);
   U268 : CLKBUF_X1 port map( A => n297, Z => n245);
   U269 : CLKBUF_X1 port map( A => n297, Z => n246);
   U270 : CLKBUF_X1 port map( A => n297, Z => n247);
   U271 : CLKBUF_X1 port map( A => n296, Z => n248);
   U272 : CLKBUF_X1 port map( A => n296, Z => n249);
   U273 : CLKBUF_X1 port map( A => n296, Z => n250);
   U274 : CLKBUF_X1 port map( A => n296, Z => n251);
   U275 : CLKBUF_X1 port map( A => n296, Z => n252);
   U276 : CLKBUF_X1 port map( A => n296, Z => n253);
   U277 : CLKBUF_X1 port map( A => n295, Z => n254);
   U278 : CLKBUF_X1 port map( A => n295, Z => n255);
   U279 : CLKBUF_X1 port map( A => n295, Z => n256);
   U280 : CLKBUF_X1 port map( A => n295, Z => n257);
   U281 : CLKBUF_X1 port map( A => n295, Z => n258);
   U282 : CLKBUF_X1 port map( A => n295, Z => n259);
   U283 : CLKBUF_X1 port map( A => n294, Z => n260);
   U284 : CLKBUF_X1 port map( A => n294, Z => n261);
   U285 : CLKBUF_X1 port map( A => n294, Z => n262);
   U286 : CLKBUF_X1 port map( A => n294, Z => n263);
   U287 : CLKBUF_X1 port map( A => n294, Z => n264);
   U288 : CLKBUF_X1 port map( A => n294, Z => n265);
   U289 : CLKBUF_X1 port map( A => n293, Z => n266);
   U290 : CLKBUF_X1 port map( A => n293, Z => n267);
   U291 : CLKBUF_X1 port map( A => n293, Z => n268);
   U292 : CLKBUF_X1 port map( A => n293, Z => n269);
   U293 : CLKBUF_X1 port map( A => n293, Z => n270);
   U294 : CLKBUF_X1 port map( A => n293, Z => n271);
   U295 : CLKBUF_X1 port map( A => n292, Z => n272);
   U296 : CLKBUF_X1 port map( A => n292, Z => n273);
   U297 : CLKBUF_X1 port map( A => n292, Z => n274);
   U298 : CLKBUF_X1 port map( A => n292, Z => n275);
   U299 : CLKBUF_X1 port map( A => n292, Z => n276);
   U300 : CLKBUF_X1 port map( A => n292, Z => n277);
   U301 : CLKBUF_X1 port map( A => n291, Z => n278);
   U302 : CLKBUF_X1 port map( A => n291, Z => n279);
   U303 : CLKBUF_X1 port map( A => n291, Z => n280);
   U304 : CLKBUF_X1 port map( A => n291, Z => n281);
   U305 : CLKBUF_X1 port map( A => n291, Z => n282);
   U306 : CLKBUF_X1 port map( A => n291, Z => n283);
   U307 : CLKBUF_X1 port map( A => n290, Z => n284);
   U308 : CLKBUF_X1 port map( A => n290, Z => n285);
   U309 : CLKBUF_X1 port map( A => n290, Z => n286);
   U310 : CLKBUF_X1 port map( A => n290, Z => n287);
   U311 : CLKBUF_X1 port map( A => n290, Z => n288);
   U312 : CLKBUF_X1 port map( A => n290, Z => n289);
   U313 : CLKBUF_X1 port map( A => n376, Z => n301);
   U314 : CLKBUF_X1 port map( A => n376, Z => n302);
   U315 : CLKBUF_X1 port map( A => n376, Z => n303);
   U316 : CLKBUF_X1 port map( A => n376, Z => n304);
   U317 : CLKBUF_X1 port map( A => n376, Z => n305);
   U318 : CLKBUF_X1 port map( A => n375, Z => n306);
   U319 : CLKBUF_X1 port map( A => n375, Z => n307);
   U320 : CLKBUF_X1 port map( A => n375, Z => n308);
   U321 : CLKBUF_X1 port map( A => n375, Z => n309);
   U322 : CLKBUF_X1 port map( A => n375, Z => n310);
   U323 : CLKBUF_X1 port map( A => n375, Z => n311);
   U324 : CLKBUF_X1 port map( A => n374, Z => n312);
   U325 : CLKBUF_X1 port map( A => n374, Z => n313);
   U326 : CLKBUF_X1 port map( A => n374, Z => n314);
   U327 : CLKBUF_X1 port map( A => n374, Z => n315);
   U328 : CLKBUF_X1 port map( A => n374, Z => n316);
   U329 : CLKBUF_X1 port map( A => n374, Z => n317);
   U330 : CLKBUF_X1 port map( A => n373, Z => n318);
   U331 : CLKBUF_X1 port map( A => n373, Z => n319);
   U332 : CLKBUF_X1 port map( A => n373, Z => n320);
   U333 : CLKBUF_X1 port map( A => n373, Z => n321);
   U334 : CLKBUF_X1 port map( A => n373, Z => n322);
   U335 : CLKBUF_X1 port map( A => n373, Z => n323);
   U336 : CLKBUF_X1 port map( A => n372, Z => n324);
   U337 : CLKBUF_X1 port map( A => n372, Z => n325);
   U338 : CLKBUF_X1 port map( A => n372, Z => n326);
   U339 : CLKBUF_X1 port map( A => n372, Z => n327);
   U340 : CLKBUF_X1 port map( A => n372, Z => n328);
   U341 : CLKBUF_X1 port map( A => n372, Z => n329);
   U342 : CLKBUF_X1 port map( A => n371, Z => n330);
   U343 : CLKBUF_X1 port map( A => n371, Z => n331);
   U344 : CLKBUF_X1 port map( A => n371, Z => n332);
   U345 : CLKBUF_X1 port map( A => n371, Z => n333);
   U346 : CLKBUF_X1 port map( A => n371, Z => n334);
   U347 : CLKBUF_X1 port map( A => n371, Z => n335);
   U348 : CLKBUF_X1 port map( A => n370, Z => n336);
   U349 : CLKBUF_X1 port map( A => n370, Z => n337);
   U350 : CLKBUF_X1 port map( A => n370, Z => n338);
   U351 : CLKBUF_X1 port map( A => n370, Z => n339);
   U352 : CLKBUF_X1 port map( A => n370, Z => n340);
   U353 : CLKBUF_X1 port map( A => n370, Z => n341);
   U354 : CLKBUF_X1 port map( A => n369, Z => n342);
   U355 : CLKBUF_X1 port map( A => n369, Z => n343);
   U356 : CLKBUF_X1 port map( A => n369, Z => n344);
   U357 : CLKBUF_X1 port map( A => n369, Z => n345);
   U358 : CLKBUF_X1 port map( A => n369, Z => n346);
   U359 : CLKBUF_X1 port map( A => n369, Z => n347);
   U360 : CLKBUF_X1 port map( A => n368, Z => n348);
   U361 : CLKBUF_X1 port map( A => n368, Z => n349);
   U362 : CLKBUF_X1 port map( A => n368, Z => n350);
   U363 : CLKBUF_X1 port map( A => n368, Z => n351);
   U364 : CLKBUF_X1 port map( A => n368, Z => n352);
   U365 : CLKBUF_X1 port map( A => n368, Z => n353);
   U366 : CLKBUF_X1 port map( A => n367, Z => n354);
   U367 : CLKBUF_X1 port map( A => n367, Z => n355);
   U368 : CLKBUF_X1 port map( A => n367, Z => n356);
   U369 : CLKBUF_X1 port map( A => n367, Z => n357);
   U370 : CLKBUF_X1 port map( A => n367, Z => n358);
   U371 : CLKBUF_X1 port map( A => n367, Z => n359);
   U372 : CLKBUF_X1 port map( A => n366, Z => n360);
   U373 : CLKBUF_X1 port map( A => n366, Z => n361);
   U374 : CLKBUF_X1 port map( A => n366, Z => n362);
   U375 : CLKBUF_X1 port map( A => n366, Z => n363);
   U376 : CLKBUF_X1 port map( A => n366, Z => n364);
   U377 : CLKBUF_X1 port map( A => n366, Z => n365);
   U378 : INV_X1 port map( A => n377, ZN => curr_proc_regs(31));
   U379 : AOI221_X1 port map( B1 => n43, B2 => regs(1055), C1 => regs(2079), C2
                           => n301, A => n379, ZN => n377);
   U380 : INV_X1 port map( A => n380, ZN => n379);
   U381 : AOI222_X1 port map( A1 => regs(31), A2 => n107, B1 => regs(1567), B2 
                           => n214, C1 => regs(543), C2 => n289, ZN => n380);
   U382 : INV_X1 port map( A => n384, ZN => curr_proc_regs(543));
   U383 : AOI221_X1 port map( B1 => regs(1567), B2 => n22, C1 => regs(31), C2 
                           => n301, A => n385, ZN => n384);
   U384 : INV_X1 port map( A => n386, ZN => n385);
   U385 : AOI222_X1 port map( A1 => n139, A2 => regs(543), B1 => regs(2079), B2
                           => n214, C1 => regs(1055), C2 => n289, ZN => n386);
   U386 : INV_X1 port map( A => n387, ZN => curr_proc_regs(30));
   U387 : AOI221_X1 port map( B1 => n38, B2 => regs(1054), C1 => n301, C2 => 
                           regs(2078), A => n388, ZN => n387);
   U388 : INV_X1 port map( A => n389, ZN => n388);
   U389 : AOI222_X1 port map( A1 => regs(30), A2 => n99, B1 => regs(1566), B2 
                           => n214, C1 => regs(542), C2 => n289, ZN => n389);
   U390 : INV_X1 port map( A => n390, ZN => curr_proc_regs(542));
   U391 : AOI221_X1 port map( B1 => n33, B2 => regs(1566), C1 => n322, C2 => 
                           regs(30), A => n391, ZN => n390);
   U392 : INV_X1 port map( A => n392, ZN => n391);
   U393 : AOI222_X1 port map( A1 => regs(542), A2 => n92, B1 => regs(2078), B2 
                           => n214, C1 => regs(1054), C2 => n289, ZN => n392);
   U394 : INV_X1 port map( A => n393, ZN => curr_proc_regs(29));
   U395 : AOI221_X1 port map( B1 => n33, B2 => regs(1053), C1 => n333, C2 => 
                           regs(2077), A => n394, ZN => n393);
   U396 : INV_X1 port map( A => n395, ZN => n394);
   U397 : AOI222_X1 port map( A1 => regs(29), A2 => n92, B1 => regs(1565), B2 
                           => n214, C1 => regs(541), C2 => n289, ZN => n395);
   U398 : INV_X1 port map( A => n396, ZN => curr_proc_regs(541));
   U399 : AOI221_X1 port map( B1 => n33, B2 => regs(1565), C1 => n333, C2 => 
                           regs(29), A => n397, ZN => n396);
   U400 : INV_X1 port map( A => n398, ZN => n397);
   U401 : AOI222_X1 port map( A1 => regs(541), A2 => n92, B1 => regs(2077), B2 
                           => n214, C1 => regs(1053), C2 => n289, ZN => n398);
   U402 : INV_X1 port map( A => n399, ZN => curr_proc_regs(28));
   U403 : AOI221_X1 port map( B1 => n33, B2 => regs(1052), C1 => n332, C2 => 
                           regs(2076), A => n400, ZN => n399);
   U404 : INV_X1 port map( A => n401, ZN => n400);
   U405 : AOI222_X1 port map( A1 => regs(28), A2 => n92, B1 => regs(1564), B2 
                           => n214, C1 => regs(540), C2 => n289, ZN => n401);
   U406 : INV_X1 port map( A => n402, ZN => curr_proc_regs(540));
   U407 : AOI221_X1 port map( B1 => n33, B2 => regs(1564), C1 => n332, C2 => 
                           regs(28), A => n403, ZN => n402);
   U408 : INV_X1 port map( A => n404, ZN => n403);
   U409 : AOI222_X1 port map( A1 => regs(540), A2 => n92, B1 => regs(2076), B2 
                           => n214, C1 => regs(1052), C2 => n289, ZN => n404);
   U410 : INV_X1 port map( A => n405, ZN => curr_proc_regs(27));
   U411 : AOI221_X1 port map( B1 => n33, B2 => regs(1051), C1 => n332, C2 => 
                           regs(2075), A => n406, ZN => n405);
   U412 : INV_X1 port map( A => n407, ZN => n406);
   U413 : AOI222_X1 port map( A1 => regs(27), A2 => n92, B1 => regs(1563), B2 
                           => n214, C1 => regs(539), C2 => n289, ZN => n407);
   U414 : INV_X1 port map( A => n408, ZN => curr_proc_regs(539));
   U415 : AOI221_X1 port map( B1 => n33, B2 => regs(1563), C1 => n332, C2 => 
                           regs(27), A => n409, ZN => n408);
   U416 : INV_X1 port map( A => n410, ZN => n409);
   U417 : AOI222_X1 port map( A1 => regs(539), A2 => n92, B1 => regs(2075), B2 
                           => n214, C1 => regs(1051), C2 => n289, ZN => n410);
   U418 : INV_X1 port map( A => n411, ZN => curr_proc_regs(26));
   U419 : AOI221_X1 port map( B1 => n33, B2 => regs(1050), C1 => n332, C2 => 
                           regs(2074), A => n412, ZN => n411);
   U420 : INV_X1 port map( A => n413, ZN => n412);
   U421 : AOI222_X1 port map( A1 => regs(26), A2 => n92, B1 => regs(1562), B2 
                           => n214, C1 => regs(538), C2 => n289, ZN => n413);
   U422 : INV_X1 port map( A => n414, ZN => curr_proc_regs(538));
   U423 : AOI221_X1 port map( B1 => n33, B2 => regs(1562), C1 => n332, C2 => 
                           regs(26), A => n415, ZN => n414);
   U424 : INV_X1 port map( A => n416, ZN => n415);
   U425 : AOI222_X1 port map( A1 => regs(538), A2 => n92, B1 => regs(2074), B2 
                           => n214, C1 => regs(1050), C2 => n289, ZN => n416);
   U426 : INV_X1 port map( A => n417, ZN => curr_proc_regs(25));
   U427 : AOI221_X1 port map( B1 => n33, B2 => regs(1049), C1 => n332, C2 => 
                           regs(2073), A => n418, ZN => n417);
   U428 : INV_X1 port map( A => n419, ZN => n418);
   U429 : AOI222_X1 port map( A1 => regs(25), A2 => n92, B1 => regs(1561), B2 
                           => n213, C1 => regs(537), C2 => n288, ZN => n419);
   U430 : INV_X1 port map( A => n420, ZN => curr_proc_regs(537));
   U431 : AOI221_X1 port map( B1 => n33, B2 => regs(1561), C1 => n332, C2 => 
                           regs(25), A => n421, ZN => n420);
   U432 : INV_X1 port map( A => n422, ZN => n421);
   U433 : AOI222_X1 port map( A1 => regs(537), A2 => n92, B1 => regs(2073), B2 
                           => n213, C1 => regs(1049), C2 => n288, ZN => n422);
   U434 : INV_X1 port map( A => n423, ZN => curr_proc_regs(24));
   U435 : AOI221_X1 port map( B1 => n34, B2 => regs(1048), C1 => n332, C2 => 
                           regs(2072), A => n424, ZN => n423);
   U436 : INV_X1 port map( A => n425, ZN => n424);
   U437 : AOI222_X1 port map( A1 => regs(24), A2 => n92, B1 => regs(1560), B2 
                           => n213, C1 => regs(536), C2 => n288, ZN => n425);
   U438 : INV_X1 port map( A => n426, ZN => curr_proc_regs(536));
   U439 : AOI221_X1 port map( B1 => n34, B2 => regs(1560), C1 => n332, C2 => 
                           regs(24), A => n427, ZN => n426);
   U440 : INV_X1 port map( A => n428, ZN => n427);
   U441 : AOI222_X1 port map( A1 => regs(536), A2 => n93, B1 => regs(2072), B2 
                           => n213, C1 => regs(1048), C2 => n288, ZN => n428);
   U442 : INV_X1 port map( A => n429, ZN => curr_proc_regs(23));
   U443 : AOI221_X1 port map( B1 => n34, B2 => regs(1047), C1 => n332, C2 => 
                           regs(2071), A => n430, ZN => n429);
   U444 : INV_X1 port map( A => n431, ZN => n430);
   U445 : AOI222_X1 port map( A1 => regs(23), A2 => n93, B1 => regs(1559), B2 
                           => n213, C1 => regs(535), C2 => n288, ZN => n431);
   U446 : INV_X1 port map( A => n432, ZN => curr_proc_regs(535));
   U447 : AOI221_X1 port map( B1 => n34, B2 => regs(1559), C1 => n332, C2 => 
                           regs(23), A => n433, ZN => n432);
   U448 : INV_X1 port map( A => n434, ZN => n433);
   U449 : AOI222_X1 port map( A1 => regs(535), A2 => n93, B1 => regs(2071), B2 
                           => n213, C1 => regs(1047), C2 => n288, ZN => n434);
   U450 : INV_X1 port map( A => n435, ZN => curr_proc_regs(22));
   U451 : AOI221_X1 port map( B1 => n34, B2 => regs(1046), C1 => n331, C2 => 
                           regs(2070), A => n436, ZN => n435);
   U452 : INV_X1 port map( A => n437, ZN => n436);
   U453 : AOI222_X1 port map( A1 => regs(22), A2 => n93, B1 => regs(1558), B2 
                           => n213, C1 => regs(534), C2 => n288, ZN => n437);
   U454 : INV_X1 port map( A => n438, ZN => curr_proc_regs(534));
   U455 : AOI221_X1 port map( B1 => n34, B2 => regs(1558), C1 => n331, C2 => 
                           regs(22), A => n439, ZN => n438);
   U456 : INV_X1 port map( A => n440, ZN => n439);
   U457 : AOI222_X1 port map( A1 => regs(534), A2 => n93, B1 => regs(2070), B2 
                           => n213, C1 => regs(1046), C2 => n288, ZN => n440);
   U458 : INV_X1 port map( A => n441, ZN => curr_proc_regs(21));
   U459 : AOI221_X1 port map( B1 => n34, B2 => regs(1045), C1 => n331, C2 => 
                           regs(2069), A => n442, ZN => n441);
   U460 : INV_X1 port map( A => n443, ZN => n442);
   U461 : AOI222_X1 port map( A1 => regs(21), A2 => n93, B1 => regs(1557), B2 
                           => n213, C1 => regs(533), C2 => n288, ZN => n443);
   U462 : INV_X1 port map( A => n444, ZN => curr_proc_regs(533));
   U463 : AOI221_X1 port map( B1 => n34, B2 => regs(1557), C1 => n331, C2 => 
                           regs(21), A => n445, ZN => n444);
   U464 : INV_X1 port map( A => n446, ZN => n445);
   U465 : AOI222_X1 port map( A1 => regs(533), A2 => n93, B1 => regs(2069), B2 
                           => n213, C1 => regs(1045), C2 => n288, ZN => n446);
   U466 : INV_X1 port map( A => n447, ZN => curr_proc_regs(20));
   U467 : AOI221_X1 port map( B1 => n34, B2 => regs(1044), C1 => n331, C2 => 
                           regs(2068), A => n448, ZN => n447);
   U468 : INV_X1 port map( A => n449, ZN => n448);
   U469 : AOI222_X1 port map( A1 => regs(20), A2 => n93, B1 => regs(1556), B2 
                           => n213, C1 => regs(532), C2 => n288, ZN => n449);
   U470 : INV_X1 port map( A => n450, ZN => curr_proc_regs(532));
   U471 : AOI221_X1 port map( B1 => n34, B2 => regs(1556), C1 => n331, C2 => 
                           regs(20), A => n451, ZN => n450);
   U472 : INV_X1 port map( A => n452, ZN => n451);
   U473 : AOI222_X1 port map( A1 => regs(532), A2 => n93, B1 => regs(2068), B2 
                           => n213, C1 => regs(1044), C2 => n288, ZN => n452);
   U474 : INV_X1 port map( A => n453, ZN => curr_proc_regs(19));
   U475 : AOI221_X1 port map( B1 => n34, B2 => regs(1043), C1 => n331, C2 => 
                           regs(2067), A => n454, ZN => n453);
   U476 : INV_X1 port map( A => n455, ZN => n454);
   U477 : AOI222_X1 port map( A1 => regs(19), A2 => n93, B1 => regs(1555), B2 
                           => n212, C1 => regs(531), C2 => n287, ZN => n455);
   U478 : INV_X1 port map( A => n456, ZN => curr_proc_regs(531));
   U479 : AOI221_X1 port map( B1 => n34, B2 => regs(1555), C1 => n331, C2 => 
                           regs(19), A => n457, ZN => n456);
   U480 : INV_X1 port map( A => n458, ZN => n457);
   U481 : AOI222_X1 port map( A1 => regs(531), A2 => n93, B1 => regs(2067), B2 
                           => n212, C1 => regs(1043), C2 => n287, ZN => n458);
   U482 : INV_X1 port map( A => n459, ZN => curr_proc_regs(18));
   U483 : AOI221_X1 port map( B1 => n35, B2 => regs(1042), C1 => n331, C2 => 
                           regs(2066), A => n460, ZN => n459);
   U484 : INV_X1 port map( A => n461, ZN => n460);
   U485 : AOI222_X1 port map( A1 => regs(18), A2 => n93, B1 => regs(1554), B2 
                           => n212, C1 => regs(530), C2 => n287, ZN => n461);
   U486 : INV_X1 port map( A => n462, ZN => curr_proc_regs(530));
   U487 : AOI221_X1 port map( B1 => n35, B2 => regs(1554), C1 => n331, C2 => 
                           regs(18), A => n463, ZN => n462);
   U488 : INV_X1 port map( A => n464, ZN => n463);
   U489 : AOI222_X1 port map( A1 => regs(530), A2 => n94, B1 => regs(2066), B2 
                           => n212, C1 => regs(1042), C2 => n287, ZN => n464);
   U490 : INV_X1 port map( A => n465, ZN => curr_proc_regs(17));
   U491 : AOI221_X1 port map( B1 => n35, B2 => regs(1041), C1 => n331, C2 => 
                           regs(2065), A => n466, ZN => n465);
   U492 : INV_X1 port map( A => n467, ZN => n466);
   U493 : AOI222_X1 port map( A1 => regs(17), A2 => n94, B1 => regs(1553), B2 
                           => n212, C1 => regs(529), C2 => n287, ZN => n467);
   U494 : INV_X1 port map( A => n468, ZN => curr_proc_regs(529));
   U495 : AOI221_X1 port map( B1 => n35, B2 => regs(1553), C1 => n331, C2 => 
                           regs(17), A => n469, ZN => n468);
   U496 : INV_X1 port map( A => n470, ZN => n469);
   U497 : AOI222_X1 port map( A1 => regs(529), A2 => n94, B1 => regs(2065), B2 
                           => n212, C1 => regs(1041), C2 => n287, ZN => n470);
   U498 : INV_X1 port map( A => n471, ZN => curr_proc_regs(16));
   U499 : AOI221_X1 port map( B1 => n35, B2 => regs(1040), C1 => n330, C2 => 
                           regs(2064), A => n472, ZN => n471);
   U500 : INV_X1 port map( A => n473, ZN => n472);
   U501 : AOI222_X1 port map( A1 => regs(16), A2 => n94, B1 => regs(1552), B2 
                           => n212, C1 => regs(528), C2 => n287, ZN => n473);
   U502 : INV_X1 port map( A => n474, ZN => curr_proc_regs(528));
   U503 : AOI221_X1 port map( B1 => n35, B2 => regs(1552), C1 => n330, C2 => 
                           regs(16), A => n475, ZN => n474);
   U504 : INV_X1 port map( A => n476, ZN => n475);
   U505 : AOI222_X1 port map( A1 => regs(528), A2 => n94, B1 => regs(2064), B2 
                           => n212, C1 => regs(1040), C2 => n287, ZN => n476);
   U506 : INV_X1 port map( A => n477, ZN => curr_proc_regs(15));
   U507 : AOI221_X1 port map( B1 => n35, B2 => regs(1039), C1 => n330, C2 => 
                           regs(2063), A => n478, ZN => n477);
   U508 : INV_X1 port map( A => n479, ZN => n478);
   U509 : AOI222_X1 port map( A1 => regs(15), A2 => n94, B1 => regs(1551), B2 
                           => n212, C1 => regs(527), C2 => n287, ZN => n479);
   U510 : INV_X1 port map( A => n480, ZN => curr_proc_regs(527));
   U511 : AOI221_X1 port map( B1 => n35, B2 => regs(1551), C1 => n330, C2 => 
                           regs(15), A => n481, ZN => n480);
   U512 : INV_X1 port map( A => n482, ZN => n481);
   U513 : AOI222_X1 port map( A1 => regs(527), A2 => n94, B1 => regs(2063), B2 
                           => n212, C1 => regs(1039), C2 => n287, ZN => n482);
   U514 : INV_X1 port map( A => n483, ZN => curr_proc_regs(14));
   U515 : AOI221_X1 port map( B1 => n35, B2 => regs(1038), C1 => n330, C2 => 
                           regs(2062), A => n484, ZN => n483);
   U516 : INV_X1 port map( A => n485, ZN => n484);
   U517 : AOI222_X1 port map( A1 => regs(14), A2 => n94, B1 => regs(1550), B2 
                           => n212, C1 => regs(526), C2 => n287, ZN => n485);
   U518 : INV_X1 port map( A => n486, ZN => curr_proc_regs(526));
   U519 : AOI221_X1 port map( B1 => n35, B2 => regs(1550), C1 => n330, C2 => 
                           regs(14), A => n487, ZN => n486);
   U520 : INV_X1 port map( A => n488, ZN => n487);
   U521 : AOI222_X1 port map( A1 => regs(526), A2 => n94, B1 => regs(2062), B2 
                           => n212, C1 => regs(1038), C2 => n287, ZN => n488);
   U522 : INV_X1 port map( A => n489, ZN => curr_proc_regs(13));
   U523 : AOI221_X1 port map( B1 => n35, B2 => regs(1037), C1 => n330, C2 => 
                           regs(2061), A => n490, ZN => n489);
   U524 : INV_X1 port map( A => n491, ZN => n490);
   U525 : AOI222_X1 port map( A1 => regs(13), A2 => n94, B1 => regs(1549), B2 
                           => n211, C1 => regs(525), C2 => n286, ZN => n491);
   U526 : INV_X1 port map( A => n492, ZN => curr_proc_regs(525));
   U527 : AOI221_X1 port map( B1 => n35, B2 => regs(1549), C1 => n330, C2 => 
                           regs(13), A => n493, ZN => n492);
   U528 : INV_X1 port map( A => n494, ZN => n493);
   U529 : AOI222_X1 port map( A1 => regs(525), A2 => n94, B1 => regs(2061), B2 
                           => n211, C1 => regs(1037), C2 => n286, ZN => n494);
   U530 : INV_X1 port map( A => n495, ZN => curr_proc_regs(12));
   U531 : AOI221_X1 port map( B1 => n36, B2 => regs(1036), C1 => n330, C2 => 
                           regs(2060), A => n496, ZN => n495);
   U532 : INV_X1 port map( A => n497, ZN => n496);
   U533 : AOI222_X1 port map( A1 => regs(12), A2 => n94, B1 => regs(1548), B2 
                           => n211, C1 => regs(524), C2 => n286, ZN => n497);
   U534 : INV_X1 port map( A => n498, ZN => curr_proc_regs(524));
   U535 : AOI221_X1 port map( B1 => n36, B2 => regs(1548), C1 => n330, C2 => 
                           regs(12), A => n499, ZN => n498);
   U536 : INV_X1 port map( A => n500, ZN => n499);
   U537 : AOI222_X1 port map( A1 => regs(524), A2 => n95, B1 => regs(2060), B2 
                           => n211, C1 => regs(1036), C2 => n286, ZN => n500);
   U538 : INV_X1 port map( A => n501, ZN => curr_proc_regs(11));
   U539 : AOI221_X1 port map( B1 => n36, B2 => regs(1035), C1 => n330, C2 => 
                           regs(2059), A => n502, ZN => n501);
   U540 : INV_X1 port map( A => n503, ZN => n502);
   U541 : AOI222_X1 port map( A1 => regs(11), A2 => n95, B1 => regs(1547), B2 
                           => n211, C1 => regs(523), C2 => n286, ZN => n503);
   U542 : INV_X1 port map( A => n504, ZN => curr_proc_regs(523));
   U543 : AOI221_X1 port map( B1 => n36, B2 => regs(1547), C1 => n330, C2 => 
                           regs(11), A => n505, ZN => n504);
   U544 : INV_X1 port map( A => n506, ZN => n505);
   U545 : AOI222_X1 port map( A1 => regs(523), A2 => n95, B1 => regs(2059), B2 
                           => n211, C1 => regs(1035), C2 => n286, ZN => n506);
   U546 : INV_X1 port map( A => n507, ZN => curr_proc_regs(10));
   U547 : AOI221_X1 port map( B1 => n36, B2 => regs(1034), C1 => n329, C2 => 
                           regs(2058), A => n508, ZN => n507);
   U548 : INV_X1 port map( A => n509, ZN => n508);
   U549 : AOI222_X1 port map( A1 => regs(10), A2 => n95, B1 => regs(1546), B2 
                           => n211, C1 => regs(522), C2 => n286, ZN => n509);
   U550 : INV_X1 port map( A => n510, ZN => curr_proc_regs(522));
   U551 : AOI221_X1 port map( B1 => n36, B2 => regs(1546), C1 => n329, C2 => 
                           regs(10), A => n511, ZN => n510);
   U552 : INV_X1 port map( A => n512, ZN => n511);
   U553 : AOI222_X1 port map( A1 => regs(522), A2 => n95, B1 => regs(2058), B2 
                           => n211, C1 => regs(1034), C2 => n286, ZN => n512);
   U554 : INV_X1 port map( A => n513, ZN => curr_proc_regs(521));
   U555 : AOI221_X1 port map( B1 => n36, B2 => regs(1545), C1 => n329, C2 => 
                           regs(9), A => n514, ZN => n513);
   U556 : INV_X1 port map( A => n515, ZN => n514);
   U557 : AOI222_X1 port map( A1 => regs(521), A2 => n95, B1 => regs(2057), B2 
                           => n211, C1 => regs(1033), C2 => n286, ZN => n515);
   U558 : INV_X1 port map( A => n516, ZN => curr_proc_regs(9));
   U559 : AOI221_X1 port map( B1 => n36, B2 => regs(1033), C1 => n329, C2 => 
                           regs(2057), A => n517, ZN => n516);
   U560 : INV_X1 port map( A => n518, ZN => n517);
   U561 : AOI222_X1 port map( A1 => regs(9), A2 => n95, B1 => regs(1545), B2 =>
                           n211, C1 => regs(521), C2 => n286, ZN => n518);
   U562 : INV_X1 port map( A => n519, ZN => curr_proc_regs(520));
   U563 : AOI221_X1 port map( B1 => n36, B2 => regs(1544), C1 => n329, C2 => 
                           regs(8), A => n520, ZN => n519);
   U564 : INV_X1 port map( A => n521, ZN => n520);
   U565 : AOI222_X1 port map( A1 => regs(520), A2 => n95, B1 => regs(2056), B2 
                           => n211, C1 => regs(1032), C2 => n286, ZN => n521);
   U566 : INV_X1 port map( A => n522, ZN => curr_proc_regs(8));
   U567 : AOI221_X1 port map( B1 => n36, B2 => regs(1032), C1 => n329, C2 => 
                           regs(2056), A => n523, ZN => n522);
   U568 : INV_X1 port map( A => n524, ZN => n523);
   U569 : AOI222_X1 port map( A1 => regs(8), A2 => n95, B1 => regs(1544), B2 =>
                           n211, C1 => regs(520), C2 => n286, ZN => n524);
   U570 : INV_X1 port map( A => n525, ZN => curr_proc_regs(519));
   U571 : AOI221_X1 port map( B1 => n36, B2 => regs(1543), C1 => n329, C2 => 
                           regs(7), A => n526, ZN => n525);
   U572 : INV_X1 port map( A => n527, ZN => n526);
   U573 : AOI222_X1 port map( A1 => regs(519), A2 => n95, B1 => regs(2055), B2 
                           => n210, C1 => regs(1031), C2 => n285, ZN => n527);
   U574 : INV_X1 port map( A => n528, ZN => curr_proc_regs(7));
   U575 : AOI221_X1 port map( B1 => n36, B2 => regs(1031), C1 => n329, C2 => 
                           regs(2055), A => n529, ZN => n528);
   U576 : INV_X1 port map( A => n530, ZN => n529);
   U577 : AOI222_X1 port map( A1 => regs(7), A2 => n95, B1 => regs(1543), B2 =>
                           n210, C1 => regs(519), C2 => n285, ZN => n530);
   U578 : INV_X1 port map( A => n531, ZN => curr_proc_regs(518));
   U579 : AOI221_X1 port map( B1 => n37, B2 => regs(1542), C1 => n329, C2 => 
                           regs(6), A => n532, ZN => n531);
   U580 : INV_X1 port map( A => n533, ZN => n532);
   U581 : AOI222_X1 port map( A1 => regs(518), A2 => n95, B1 => regs(2054), B2 
                           => n210, C1 => regs(1030), C2 => n285, ZN => n533);
   U582 : INV_X1 port map( A => n534, ZN => curr_proc_regs(6));
   U583 : AOI221_X1 port map( B1 => n37, B2 => regs(1030), C1 => n329, C2 => 
                           regs(2054), A => n535, ZN => n534);
   U584 : INV_X1 port map( A => n536, ZN => n535);
   U585 : AOI222_X1 port map( A1 => regs(6), A2 => n96, B1 => regs(1542), B2 =>
                           n210, C1 => regs(518), C2 => n285, ZN => n536);
   U586 : INV_X1 port map( A => n537, ZN => curr_proc_regs(517));
   U587 : AOI221_X1 port map( B1 => n37, B2 => regs(1541), C1 => n329, C2 => 
                           regs(5), A => n538, ZN => n537);
   U588 : INV_X1 port map( A => n539, ZN => n538);
   U589 : AOI222_X1 port map( A1 => regs(517), A2 => n96, B1 => regs(2053), B2 
                           => n210, C1 => regs(1029), C2 => n285, ZN => n539);
   U590 : INV_X1 port map( A => n540, ZN => curr_proc_regs(5));
   U591 : AOI221_X1 port map( B1 => n37, B2 => regs(1029), C1 => n329, C2 => 
                           regs(2053), A => n541, ZN => n540);
   U592 : INV_X1 port map( A => n542, ZN => n541);
   U593 : AOI222_X1 port map( A1 => regs(5), A2 => n96, B1 => regs(1541), B2 =>
                           n210, C1 => regs(517), C2 => n285, ZN => n542);
   U594 : INV_X1 port map( A => n543, ZN => curr_proc_regs(4));
   U595 : AOI221_X1 port map( B1 => n37, B2 => regs(1028), C1 => n328, C2 => 
                           regs(2052), A => n544, ZN => n543);
   U596 : INV_X1 port map( A => n545, ZN => n544);
   U597 : AOI222_X1 port map( A1 => regs(4), A2 => n96, B1 => regs(1540), B2 =>
                           n210, C1 => regs(516), C2 => n285, ZN => n545);
   U598 : INV_X1 port map( A => n546, ZN => curr_proc_regs(516));
   U599 : AOI221_X1 port map( B1 => n37, B2 => regs(1540), C1 => n328, C2 => 
                           regs(4), A => n547, ZN => n546);
   U600 : INV_X1 port map( A => n548, ZN => n547);
   U601 : AOI222_X1 port map( A1 => regs(516), A2 => n96, B1 => regs(2052), B2 
                           => n210, C1 => regs(1028), C2 => n285, ZN => n548);
   U602 : INV_X1 port map( A => n549, ZN => curr_proc_regs(3));
   U603 : AOI221_X1 port map( B1 => n37, B2 => regs(1027), C1 => n328, C2 => 
                           regs(2051), A => n550, ZN => n549);
   U604 : INV_X1 port map( A => n551, ZN => n550);
   U605 : AOI222_X1 port map( A1 => regs(3), A2 => n96, B1 => regs(1539), B2 =>
                           n210, C1 => regs(515), C2 => n285, ZN => n551);
   U606 : INV_X1 port map( A => n552, ZN => curr_proc_regs(515));
   U607 : AOI221_X1 port map( B1 => n37, B2 => regs(1539), C1 => n328, C2 => 
                           regs(3), A => n553, ZN => n552);
   U608 : INV_X1 port map( A => n554, ZN => n553);
   U609 : AOI222_X1 port map( A1 => regs(515), A2 => n96, B1 => regs(2051), B2 
                           => n210, C1 => regs(1027), C2 => n285, ZN => n554);
   U610 : INV_X1 port map( A => n555, ZN => curr_proc_regs(2));
   U611 : AOI221_X1 port map( B1 => n37, B2 => regs(1026), C1 => n328, C2 => 
                           regs(2050), A => n556, ZN => n555);
   U612 : INV_X1 port map( A => n557, ZN => n556);
   U613 : AOI222_X1 port map( A1 => regs(2), A2 => n96, B1 => regs(1538), B2 =>
                           n210, C1 => regs(514), C2 => n285, ZN => n557);
   U614 : INV_X1 port map( A => n558, ZN => curr_proc_regs(514));
   U615 : AOI221_X1 port map( B1 => n37, B2 => regs(1538), C1 => n328, C2 => 
                           regs(2), A => n559, ZN => n558);
   U616 : INV_X1 port map( A => n560, ZN => n559);
   U617 : AOI222_X1 port map( A1 => regs(514), A2 => n96, B1 => regs(2050), B2 
                           => n210, C1 => regs(1026), C2 => n285, ZN => n560);
   U618 : INV_X1 port map( A => n561, ZN => curr_proc_regs(1));
   U619 : AOI221_X1 port map( B1 => n37, B2 => regs(1025), C1 => n328, C2 => 
                           regs(2049), A => n562, ZN => n561);
   U620 : INV_X1 port map( A => n563, ZN => n562);
   U621 : AOI222_X1 port map( A1 => regs(1), A2 => n96, B1 => regs(1537), B2 =>
                           n209, C1 => regs(513), C2 => n284, ZN => n563);
   U622 : INV_X1 port map( A => n564, ZN => curr_proc_regs(513));
   U623 : AOI221_X1 port map( B1 => n37, B2 => regs(1537), C1 => n328, C2 => 
                           regs(1), A => n565, ZN => n564);
   U624 : INV_X1 port map( A => n566, ZN => n565);
   U625 : AOI222_X1 port map( A1 => regs(513), A2 => n96, B1 => regs(2049), B2 
                           => n209, C1 => regs(1025), C2 => n284, ZN => n566);
   U626 : INV_X1 port map( A => n567, ZN => curr_proc_regs(0));
   U627 : AOI221_X1 port map( B1 => n38, B2 => regs(1024), C1 => n328, C2 => 
                           regs(2048), A => n568, ZN => n567);
   U628 : INV_X1 port map( A => n569, ZN => n568);
   U629 : AOI222_X1 port map( A1 => regs(0), A2 => n96, B1 => regs(1536), B2 =>
                           n209, C1 => regs(512), C2 => n284, ZN => n569);
   U630 : INV_X1 port map( A => n570, ZN => curr_proc_regs(512));
   U631 : AOI221_X1 port map( B1 => n38, B2 => regs(1536), C1 => n328, C2 => 
                           regs(0), A => n571, ZN => n570);
   U632 : INV_X1 port map( A => n572, ZN => n571);
   U633 : AOI222_X1 port map( A1 => regs(512), A2 => n97, B1 => regs(2048), B2 
                           => n209, C1 => regs(1024), C2 => n284, ZN => n572);
   U634 : INV_X1 port map( A => n573, ZN => curr_proc_regs(575));
   U635 : AOI221_X1 port map( B1 => n38, B2 => regs(1599), C1 => n328, C2 => 
                           regs(63), A => n574, ZN => n573);
   U636 : INV_X1 port map( A => n575, ZN => n574);
   U637 : AOI222_X1 port map( A1 => regs(575), A2 => n97, B1 => regs(2111), B2 
                           => n209, C1 => regs(1087), C2 => n284, ZN => n575);
   U638 : INV_X1 port map( A => n576, ZN => curr_proc_regs(63));
   U639 : AOI221_X1 port map( B1 => n38, B2 => regs(1087), C1 => n328, C2 => 
                           regs(2111), A => n577, ZN => n576);
   U640 : INV_X1 port map( A => n578, ZN => n577);
   U641 : AOI222_X1 port map( A1 => regs(63), A2 => n97, B1 => regs(1599), B2 
                           => n209, C1 => regs(575), C2 => n284, ZN => n578);
   U642 : INV_X1 port map( A => n579, ZN => curr_proc_regs(574));
   U643 : AOI221_X1 port map( B1 => n38, B2 => regs(1598), C1 => n327, C2 => 
                           regs(62), A => n580, ZN => n579);
   U644 : INV_X1 port map( A => n581, ZN => n580);
   U645 : AOI222_X1 port map( A1 => regs(574), A2 => n97, B1 => regs(2110), B2 
                           => n209, C1 => regs(1086), C2 => n284, ZN => n581);
   U646 : INV_X1 port map( A => n582, ZN => curr_proc_regs(62));
   U647 : AOI221_X1 port map( B1 => n38, B2 => regs(1086), C1 => n327, C2 => 
                           regs(2110), A => n583, ZN => n582);
   U648 : INV_X1 port map( A => n584, ZN => n583);
   U649 : AOI222_X1 port map( A1 => regs(62), A2 => n97, B1 => regs(1598), B2 
                           => n209, C1 => regs(574), C2 => n284, ZN => n584);
   U650 : INV_X1 port map( A => n585, ZN => curr_proc_regs(573));
   U651 : AOI221_X1 port map( B1 => n38, B2 => regs(1597), C1 => n327, C2 => 
                           regs(61), A => n586, ZN => n585);
   U652 : INV_X1 port map( A => n587, ZN => n586);
   U653 : AOI222_X1 port map( A1 => regs(573), A2 => n97, B1 => regs(2109), B2 
                           => n209, C1 => regs(1085), C2 => n284, ZN => n587);
   U654 : INV_X1 port map( A => n588, ZN => curr_proc_regs(61));
   U655 : AOI221_X1 port map( B1 => n38, B2 => regs(1085), C1 => n327, C2 => 
                           regs(2109), A => n589, ZN => n588);
   U656 : INV_X1 port map( A => n590, ZN => n589);
   U657 : AOI222_X1 port map( A1 => regs(61), A2 => n97, B1 => regs(1597), B2 
                           => n209, C1 => regs(573), C2 => n284, ZN => n590);
   U658 : INV_X1 port map( A => n591, ZN => curr_proc_regs(572));
   U659 : AOI221_X1 port map( B1 => n38, B2 => regs(1596), C1 => n327, C2 => 
                           regs(60), A => n592, ZN => n591);
   U660 : INV_X1 port map( A => n593, ZN => n592);
   U661 : AOI222_X1 port map( A1 => regs(572), A2 => n97, B1 => regs(2108), B2 
                           => n209, C1 => regs(1084), C2 => n284, ZN => n593);
   U662 : INV_X1 port map( A => n594, ZN => curr_proc_regs(60));
   U663 : AOI221_X1 port map( B1 => n38, B2 => regs(1084), C1 => n327, C2 => 
                           regs(2108), A => n595, ZN => n594);
   U664 : INV_X1 port map( A => n596, ZN => n595);
   U665 : AOI222_X1 port map( A1 => regs(60), A2 => n97, B1 => regs(1596), B2 
                           => n209, C1 => regs(572), C2 => n284, ZN => n596);
   U666 : INV_X1 port map( A => n597, ZN => curr_proc_regs(571));
   U667 : AOI221_X1 port map( B1 => n38, B2 => regs(1595), C1 => n327, C2 => 
                           regs(59), A => n598, ZN => n597);
   U668 : INV_X1 port map( A => n599, ZN => n598);
   U669 : AOI222_X1 port map( A1 => regs(571), A2 => n97, B1 => regs(2107), B2 
                           => n208, C1 => regs(1083), C2 => n283, ZN => n599);
   U670 : INV_X1 port map( A => n600, ZN => curr_proc_regs(59));
   U671 : AOI221_X1 port map( B1 => n39, B2 => regs(1083), C1 => n327, C2 => 
                           regs(2107), A => n601, ZN => n600);
   U672 : INV_X1 port map( A => n602, ZN => n601);
   U673 : AOI222_X1 port map( A1 => regs(59), A2 => n97, B1 => regs(1595), B2 
                           => n208, C1 => regs(571), C2 => n283, ZN => n602);
   U674 : INV_X1 port map( A => n603, ZN => curr_proc_regs(570));
   U675 : AOI221_X1 port map( B1 => n39, B2 => regs(1594), C1 => n327, C2 => 
                           regs(58), A => n604, ZN => n603);
   U676 : INV_X1 port map( A => n605, ZN => n604);
   U677 : AOI222_X1 port map( A1 => regs(570), A2 => n97, B1 => regs(2106), B2 
                           => n208, C1 => regs(1082), C2 => n283, ZN => n605);
   U678 : INV_X1 port map( A => n606, ZN => curr_proc_regs(58));
   U679 : AOI221_X1 port map( B1 => n39, B2 => regs(1082), C1 => n327, C2 => 
                           regs(2106), A => n607, ZN => n606);
   U680 : INV_X1 port map( A => n608, ZN => n607);
   U681 : AOI222_X1 port map( A1 => regs(58), A2 => n98, B1 => regs(1594), B2 
                           => n208, C1 => regs(570), C2 => n283, ZN => n608);
   U682 : INV_X1 port map( A => n609, ZN => curr_proc_regs(569));
   U683 : AOI221_X1 port map( B1 => n39, B2 => regs(1593), C1 => n327, C2 => 
                           regs(57), A => n610, ZN => n609);
   U684 : INV_X1 port map( A => n611, ZN => n610);
   U685 : AOI222_X1 port map( A1 => regs(569), A2 => n98, B1 => regs(2105), B2 
                           => n208, C1 => regs(1081), C2 => n283, ZN => n611);
   U686 : INV_X1 port map( A => n612, ZN => curr_proc_regs(57));
   U687 : AOI221_X1 port map( B1 => n39, B2 => regs(1081), C1 => n326, C2 => 
                           regs(2105), A => n613, ZN => n612);
   U688 : INV_X1 port map( A => n614, ZN => n613);
   U689 : AOI222_X1 port map( A1 => regs(57), A2 => n98, B1 => regs(1593), B2 
                           => n208, C1 => regs(569), C2 => n283, ZN => n614);
   U690 : INV_X1 port map( A => n615, ZN => curr_proc_regs(568));
   U691 : AOI221_X1 port map( B1 => n39, B2 => regs(1592), C1 => n326, C2 => 
                           regs(56), A => n616, ZN => n615);
   U692 : INV_X1 port map( A => n617, ZN => n616);
   U693 : AOI222_X1 port map( A1 => regs(568), A2 => n98, B1 => regs(2104), B2 
                           => n208, C1 => regs(1080), C2 => n283, ZN => n617);
   U694 : INV_X1 port map( A => n618, ZN => curr_proc_regs(56));
   U695 : AOI221_X1 port map( B1 => n39, B2 => regs(1080), C1 => n326, C2 => 
                           regs(2104), A => n619, ZN => n618);
   U696 : INV_X1 port map( A => n620, ZN => n619);
   U697 : AOI222_X1 port map( A1 => regs(56), A2 => n98, B1 => regs(1592), B2 
                           => n208, C1 => regs(568), C2 => n283, ZN => n620);
   U698 : INV_X1 port map( A => n621, ZN => curr_proc_regs(55));
   U699 : AOI221_X1 port map( B1 => n39, B2 => regs(1079), C1 => n326, C2 => 
                           regs(2103), A => n622, ZN => n621);
   U700 : INV_X1 port map( A => n623, ZN => n622);
   U701 : AOI222_X1 port map( A1 => regs(55), A2 => n98, B1 => regs(1591), B2 
                           => n208, C1 => regs(567), C2 => n283, ZN => n623);
   U702 : INV_X1 port map( A => n624, ZN => curr_proc_regs(567));
   U703 : AOI221_X1 port map( B1 => n39, B2 => regs(1591), C1 => n326, C2 => 
                           regs(55), A => n625, ZN => n624);
   U704 : INV_X1 port map( A => n626, ZN => n625);
   U705 : AOI222_X1 port map( A1 => regs(567), A2 => n98, B1 => regs(2103), B2 
                           => n208, C1 => regs(1079), C2 => n283, ZN => n626);
   U706 : INV_X1 port map( A => n627, ZN => curr_proc_regs(54));
   U707 : AOI221_X1 port map( B1 => n39, B2 => regs(1078), C1 => n326, C2 => 
                           regs(2102), A => n628, ZN => n627);
   U708 : INV_X1 port map( A => n629, ZN => n628);
   U709 : AOI222_X1 port map( A1 => regs(54), A2 => n98, B1 => regs(1590), B2 
                           => n208, C1 => regs(566), C2 => n283, ZN => n629);
   U710 : INV_X1 port map( A => n630, ZN => curr_proc_regs(566));
   U711 : AOI221_X1 port map( B1 => n39, B2 => regs(1590), C1 => n326, C2 => 
                           regs(54), A => n631, ZN => n630);
   U712 : INV_X1 port map( A => n632, ZN => n631);
   U713 : AOI222_X1 port map( A1 => regs(566), A2 => n98, B1 => regs(2102), B2 
                           => n208, C1 => regs(1078), C2 => n283, ZN => n632);
   U714 : INV_X1 port map( A => n633, ZN => curr_proc_regs(53));
   U715 : AOI221_X1 port map( B1 => n39, B2 => regs(1077), C1 => n326, C2 => 
                           regs(2101), A => n634, ZN => n633);
   U716 : INV_X1 port map( A => n635, ZN => n634);
   U717 : AOI222_X1 port map( A1 => regs(53), A2 => n98, B1 => regs(1589), B2 
                           => n207, C1 => regs(565), C2 => n282, ZN => n635);
   U718 : INV_X1 port map( A => n636, ZN => curr_proc_regs(565));
   U719 : AOI221_X1 port map( B1 => n40, B2 => regs(1589), C1 => n326, C2 => 
                           regs(53), A => n637, ZN => n636);
   U720 : INV_X1 port map( A => n638, ZN => n637);
   U721 : AOI222_X1 port map( A1 => regs(565), A2 => n98, B1 => regs(2101), B2 
                           => n207, C1 => regs(1077), C2 => n282, ZN => n638);
   U722 : INV_X1 port map( A => n639, ZN => curr_proc_regs(52));
   U723 : AOI221_X1 port map( B1 => n40, B2 => regs(1076), C1 => n326, C2 => 
                           regs(2100), A => n640, ZN => n639);
   U724 : INV_X1 port map( A => n641, ZN => n640);
   U725 : AOI222_X1 port map( A1 => regs(52), A2 => n98, B1 => regs(1588), B2 
                           => n207, C1 => regs(564), C2 => n282, ZN => n641);
   U726 : INV_X1 port map( A => n642, ZN => curr_proc_regs(564));
   U727 : AOI221_X1 port map( B1 => n40, B2 => regs(1588), C1 => n326, C2 => 
                           regs(52), A => n643, ZN => n642);
   U728 : INV_X1 port map( A => n644, ZN => n643);
   U729 : AOI222_X1 port map( A1 => regs(564), A2 => n99, B1 => regs(2100), B2 
                           => n207, C1 => regs(1076), C2 => n282, ZN => n644);
   U730 : INV_X1 port map( A => n645, ZN => curr_proc_regs(51));
   U731 : AOI221_X1 port map( B1 => n40, B2 => regs(1075), C1 => n326, C2 => 
                           regs(2099), A => n646, ZN => n645);
   U732 : INV_X1 port map( A => n647, ZN => n646);
   U733 : AOI222_X1 port map( A1 => regs(51), A2 => n99, B1 => regs(1587), B2 
                           => n207, C1 => regs(563), C2 => n282, ZN => n647);
   U734 : INV_X1 port map( A => n648, ZN => curr_proc_regs(563));
   U735 : AOI221_X1 port map( B1 => n40, B2 => regs(1587), C1 => n325, C2 => 
                           regs(51), A => n649, ZN => n648);
   U736 : INV_X1 port map( A => n650, ZN => n649);
   U737 : AOI222_X1 port map( A1 => regs(563), A2 => n99, B1 => regs(2099), B2 
                           => n207, C1 => regs(1075), C2 => n282, ZN => n650);
   U738 : INV_X1 port map( A => n651, ZN => curr_proc_regs(50));
   U739 : AOI221_X1 port map( B1 => n40, B2 => regs(1074), C1 => n325, C2 => 
                           regs(2098), A => n652, ZN => n651);
   U740 : INV_X1 port map( A => n653, ZN => n652);
   U741 : AOI222_X1 port map( A1 => regs(50), A2 => n99, B1 => regs(1586), B2 
                           => n207, C1 => regs(562), C2 => n282, ZN => n653);
   U742 : INV_X1 port map( A => n654, ZN => curr_proc_regs(562));
   U743 : AOI221_X1 port map( B1 => n40, B2 => regs(1586), C1 => n325, C2 => 
                           regs(50), A => n655, ZN => n654);
   U744 : INV_X1 port map( A => n656, ZN => n655);
   U745 : AOI222_X1 port map( A1 => regs(562), A2 => n99, B1 => regs(2098), B2 
                           => n207, C1 => regs(1074), C2 => n282, ZN => n656);
   U746 : INV_X1 port map( A => n657, ZN => curr_proc_regs(49));
   U747 : AOI221_X1 port map( B1 => n40, B2 => regs(1073), C1 => n325, C2 => 
                           regs(2097), A => n658, ZN => n657);
   U748 : INV_X1 port map( A => n659, ZN => n658);
   U749 : AOI222_X1 port map( A1 => regs(49), A2 => n99, B1 => regs(1585), B2 
                           => n207, C1 => regs(561), C2 => n282, ZN => n659);
   U750 : INV_X1 port map( A => n660, ZN => curr_proc_regs(561));
   U751 : AOI221_X1 port map( B1 => n40, B2 => regs(1585), C1 => n325, C2 => 
                           regs(49), A => n661, ZN => n660);
   U752 : INV_X1 port map( A => n662, ZN => n661);
   U753 : AOI222_X1 port map( A1 => regs(561), A2 => n99, B1 => regs(2097), B2 
                           => n207, C1 => regs(1073), C2 => n282, ZN => n662);
   U754 : INV_X1 port map( A => n663, ZN => curr_proc_regs(48));
   U755 : AOI221_X1 port map( B1 => n40, B2 => regs(1072), C1 => n325, C2 => 
                           regs(2096), A => n664, ZN => n663);
   U756 : INV_X1 port map( A => n665, ZN => n664);
   U757 : AOI222_X1 port map( A1 => regs(48), A2 => n99, B1 => regs(1584), B2 
                           => n207, C1 => regs(560), C2 => n282, ZN => n665);
   U758 : INV_X1 port map( A => n666, ZN => curr_proc_regs(560));
   U759 : AOI221_X1 port map( B1 => n40, B2 => regs(1584), C1 => n325, C2 => 
                           regs(48), A => n667, ZN => n666);
   U760 : INV_X1 port map( A => n668, ZN => n667);
   U761 : AOI222_X1 port map( A1 => regs(560), A2 => n99, B1 => regs(2096), B2 
                           => n207, C1 => regs(1072), C2 => n282, ZN => n668);
   U762 : INV_X1 port map( A => n669, ZN => curr_proc_regs(47));
   U763 : AOI221_X1 port map( B1 => n40, B2 => regs(1071), C1 => n325, C2 => 
                           regs(2095), A => n670, ZN => n669);
   U764 : INV_X1 port map( A => n671, ZN => n670);
   U765 : AOI222_X1 port map( A1 => regs(47), A2 => n99, B1 => regs(1583), B2 
                           => n206, C1 => regs(559), C2 => n281, ZN => n671);
   U766 : INV_X1 port map( A => n672, ZN => curr_proc_regs(559));
   U767 : AOI221_X1 port map( B1 => n41, B2 => regs(1583), C1 => n325, C2 => 
                           regs(47), A => n673, ZN => n672);
   U768 : INV_X1 port map( A => n674, ZN => n673);
   U769 : AOI222_X1 port map( A1 => regs(559), A2 => n99, B1 => regs(2095), B2 
                           => n206, C1 => regs(1071), C2 => n281, ZN => n674);
   U770 : INV_X1 port map( A => n675, ZN => curr_proc_regs(46));
   U771 : AOI221_X1 port map( B1 => n41, B2 => regs(1070), C1 => n325, C2 => 
                           regs(2094), A => n676, ZN => n675);
   U772 : INV_X1 port map( A => n677, ZN => n676);
   U773 : AOI222_X1 port map( A1 => regs(46), A2 => n100, B1 => regs(1582), B2 
                           => n206, C1 => regs(558), C2 => n281, ZN => n677);
   U774 : INV_X1 port map( A => n678, ZN => curr_proc_regs(558));
   U775 : AOI221_X1 port map( B1 => n41, B2 => regs(1582), C1 => n325, C2 => 
                           regs(46), A => n679, ZN => n678);
   U776 : INV_X1 port map( A => n680, ZN => n679);
   U777 : AOI222_X1 port map( A1 => regs(558), A2 => n100, B1 => regs(2094), B2
                           => n206, C1 => regs(1070), C2 => n281, ZN => n680);
   U778 : INV_X1 port map( A => n681, ZN => curr_proc_regs(45));
   U779 : AOI221_X1 port map( B1 => n41, B2 => regs(1069), C1 => n325, C2 => 
                           regs(2093), A => n682, ZN => n681);
   U780 : INV_X1 port map( A => n683, ZN => n682);
   U781 : AOI222_X1 port map( A1 => regs(45), A2 => n100, B1 => regs(1581), B2 
                           => n206, C1 => regs(557), C2 => n281, ZN => n683);
   U782 : INV_X1 port map( A => n684, ZN => curr_proc_regs(557));
   U783 : AOI221_X1 port map( B1 => n41, B2 => regs(1581), C1 => n324, C2 => 
                           regs(45), A => n685, ZN => n684);
   U784 : INV_X1 port map( A => n686, ZN => n685);
   U785 : AOI222_X1 port map( A1 => regs(557), A2 => n100, B1 => regs(2093), B2
                           => n206, C1 => regs(1069), C2 => n281, ZN => n686);
   U786 : INV_X1 port map( A => n687, ZN => curr_proc_regs(44));
   U787 : AOI221_X1 port map( B1 => n41, B2 => regs(1068), C1 => n324, C2 => 
                           regs(2092), A => n688, ZN => n687);
   U788 : INV_X1 port map( A => n689, ZN => n688);
   U789 : AOI222_X1 port map( A1 => regs(44), A2 => n100, B1 => regs(1580), B2 
                           => n206, C1 => regs(556), C2 => n281, ZN => n689);
   U790 : INV_X1 port map( A => n690, ZN => curr_proc_regs(556));
   U791 : AOI221_X1 port map( B1 => n41, B2 => regs(1580), C1 => n324, C2 => 
                           regs(44), A => n691, ZN => n690);
   U792 : INV_X1 port map( A => n692, ZN => n691);
   U793 : AOI222_X1 port map( A1 => regs(556), A2 => n100, B1 => regs(2092), B2
                           => n206, C1 => regs(1068), C2 => n281, ZN => n692);
   U794 : INV_X1 port map( A => n693, ZN => curr_proc_regs(43));
   U795 : AOI221_X1 port map( B1 => n41, B2 => regs(1067), C1 => n324, C2 => 
                           regs(2091), A => n694, ZN => n693);
   U796 : INV_X1 port map( A => n695, ZN => n694);
   U797 : AOI222_X1 port map( A1 => regs(43), A2 => n100, B1 => regs(1579), B2 
                           => n206, C1 => regs(555), C2 => n281, ZN => n695);
   U798 : INV_X1 port map( A => n696, ZN => curr_proc_regs(555));
   U799 : AOI221_X1 port map( B1 => n41, B2 => regs(1579), C1 => n324, C2 => 
                           regs(43), A => n697, ZN => n696);
   U800 : INV_X1 port map( A => n698, ZN => n697);
   U801 : AOI222_X1 port map( A1 => regs(555), A2 => n100, B1 => regs(2091), B2
                           => n206, C1 => regs(1067), C2 => n281, ZN => n698);
   U802 : INV_X1 port map( A => n699, ZN => curr_proc_regs(42));
   U803 : AOI221_X1 port map( B1 => n41, B2 => regs(1066), C1 => n324, C2 => 
                           regs(2090), A => n700, ZN => n699);
   U804 : INV_X1 port map( A => n701, ZN => n700);
   U805 : AOI222_X1 port map( A1 => regs(42), A2 => n100, B1 => regs(1578), B2 
                           => n206, C1 => regs(554), C2 => n281, ZN => n701);
   U806 : INV_X1 port map( A => n702, ZN => curr_proc_regs(554));
   U807 : AOI221_X1 port map( B1 => n41, B2 => regs(1578), C1 => n324, C2 => 
                           regs(42), A => n703, ZN => n702);
   U808 : INV_X1 port map( A => n704, ZN => n703);
   U809 : AOI222_X1 port map( A1 => regs(554), A2 => n100, B1 => regs(2090), B2
                           => n206, C1 => regs(1066), C2 => n281, ZN => n704);
   U810 : INV_X1 port map( A => n705, ZN => curr_proc_regs(41));
   U811 : AOI221_X1 port map( B1 => n41, B2 => regs(1065), C1 => n324, C2 => 
                           regs(2089), A => n706, ZN => n705);
   U812 : INV_X1 port map( A => n707, ZN => n706);
   U813 : AOI222_X1 port map( A1 => regs(41), A2 => n100, B1 => regs(1577), B2 
                           => n205, C1 => regs(553), C2 => n280, ZN => n707);
   U814 : INV_X1 port map( A => n708, ZN => curr_proc_regs(553));
   U815 : AOI221_X1 port map( B1 => n42, B2 => regs(1577), C1 => n324, C2 => 
                           regs(41), A => n709, ZN => n708);
   U816 : INV_X1 port map( A => n710, ZN => n709);
   U817 : AOI222_X1 port map( A1 => regs(553), A2 => n100, B1 => regs(2089), B2
                           => n205, C1 => regs(1065), C2 => n280, ZN => n710);
   U818 : INV_X1 port map( A => n711, ZN => curr_proc_regs(40));
   U819 : AOI221_X1 port map( B1 => n42, B2 => regs(1064), C1 => n324, C2 => 
                           regs(2088), A => n712, ZN => n711);
   U820 : INV_X1 port map( A => n713, ZN => n712);
   U821 : AOI222_X1 port map( A1 => regs(40), A2 => n101, B1 => regs(1576), B2 
                           => n205, C1 => regs(552), C2 => n280, ZN => n713);
   U822 : INV_X1 port map( A => n714, ZN => curr_proc_regs(552));
   U823 : AOI221_X1 port map( B1 => n42, B2 => regs(1576), C1 => n324, C2 => 
                           regs(40), A => n715, ZN => n714);
   U824 : INV_X1 port map( A => n716, ZN => n715);
   U825 : AOI222_X1 port map( A1 => regs(552), A2 => n101, B1 => regs(2088), B2
                           => n205, C1 => regs(1064), C2 => n280, ZN => n716);
   U826 : INV_X1 port map( A => n717, ZN => curr_proc_regs(39));
   U827 : AOI221_X1 port map( B1 => n42, B2 => regs(1063), C1 => n324, C2 => 
                           regs(2087), A => n718, ZN => n717);
   U828 : INV_X1 port map( A => n719, ZN => n718);
   U829 : AOI222_X1 port map( A1 => regs(39), A2 => n101, B1 => regs(1575), B2 
                           => n205, C1 => regs(551), C2 => n280, ZN => n719);
   U830 : INV_X1 port map( A => n720, ZN => curr_proc_regs(551));
   U831 : AOI221_X1 port map( B1 => n42, B2 => regs(1575), C1 => n323, C2 => 
                           regs(39), A => n721, ZN => n720);
   U832 : INV_X1 port map( A => n722, ZN => n721);
   U833 : AOI222_X1 port map( A1 => regs(551), A2 => n101, B1 => regs(2087), B2
                           => n205, C1 => regs(1063), C2 => n280, ZN => n722);
   U834 : INV_X1 port map( A => n723, ZN => curr_proc_regs(38));
   U835 : AOI221_X1 port map( B1 => n42, B2 => regs(1062), C1 => n323, C2 => 
                           regs(2086), A => n724, ZN => n723);
   U836 : INV_X1 port map( A => n725, ZN => n724);
   U837 : AOI222_X1 port map( A1 => regs(38), A2 => n101, B1 => regs(1574), B2 
                           => n205, C1 => regs(550), C2 => n280, ZN => n725);
   U838 : INV_X1 port map( A => n726, ZN => curr_proc_regs(550));
   U839 : AOI221_X1 port map( B1 => n42, B2 => regs(1574), C1 => n323, C2 => 
                           regs(38), A => n727, ZN => n726);
   U840 : INV_X1 port map( A => n728, ZN => n727);
   U841 : AOI222_X1 port map( A1 => regs(550), A2 => n101, B1 => regs(2086), B2
                           => n205, C1 => regs(1062), C2 => n280, ZN => n728);
   U842 : INV_X1 port map( A => n729, ZN => curr_proc_regs(37));
   U843 : AOI221_X1 port map( B1 => n42, B2 => regs(1061), C1 => n323, C2 => 
                           regs(2085), A => n730, ZN => n729);
   U844 : INV_X1 port map( A => n731, ZN => n730);
   U845 : AOI222_X1 port map( A1 => regs(37), A2 => n101, B1 => regs(1573), B2 
                           => n205, C1 => regs(549), C2 => n280, ZN => n731);
   U846 : INV_X1 port map( A => n732, ZN => curr_proc_regs(549));
   U847 : AOI221_X1 port map( B1 => n42, B2 => regs(1573), C1 => n323, C2 => 
                           regs(37), A => n733, ZN => n732);
   U848 : INV_X1 port map( A => n734, ZN => n733);
   U849 : AOI222_X1 port map( A1 => regs(549), A2 => n101, B1 => regs(2085), B2
                           => n205, C1 => regs(1061), C2 => n280, ZN => n734);
   U850 : INV_X1 port map( A => n735, ZN => curr_proc_regs(36));
   U851 : AOI221_X1 port map( B1 => n42, B2 => regs(1060), C1 => n323, C2 => 
                           regs(2084), A => n736, ZN => n735);
   U852 : INV_X1 port map( A => n737, ZN => n736);
   U853 : AOI222_X1 port map( A1 => regs(36), A2 => n101, B1 => regs(1572), B2 
                           => n205, C1 => regs(548), C2 => n280, ZN => n737);
   U854 : INV_X1 port map( A => n738, ZN => curr_proc_regs(548));
   U855 : AOI221_X1 port map( B1 => n42, B2 => regs(1572), C1 => n323, C2 => 
                           regs(36), A => n739, ZN => n738);
   U856 : INV_X1 port map( A => n740, ZN => n739);
   U857 : AOI222_X1 port map( A1 => regs(548), A2 => n101, B1 => regs(2084), B2
                           => n205, C1 => regs(1060), C2 => n280, ZN => n740);
   U858 : INV_X1 port map( A => n741, ZN => curr_proc_regs(35));
   U859 : AOI221_X1 port map( B1 => n42, B2 => regs(1059), C1 => n323, C2 => 
                           regs(2083), A => n742, ZN => n741);
   U860 : INV_X1 port map( A => n743, ZN => n742);
   U861 : AOI222_X1 port map( A1 => regs(35), A2 => n101, B1 => regs(1571), B2 
                           => n204, C1 => regs(547), C2 => n279, ZN => n743);
   U862 : INV_X1 port map( A => n744, ZN => curr_proc_regs(547));
   U863 : AOI221_X1 port map( B1 => n43, B2 => regs(1571), C1 => n323, C2 => 
                           regs(35), A => n745, ZN => n744);
   U864 : INV_X1 port map( A => n746, ZN => n745);
   U865 : AOI222_X1 port map( A1 => regs(547), A2 => n101, B1 => regs(2083), B2
                           => n204, C1 => regs(1059), C2 => n279, ZN => n746);
   U866 : INV_X1 port map( A => n747, ZN => curr_proc_regs(34));
   U867 : AOI221_X1 port map( B1 => n43, B2 => regs(1058), C1 => n323, C2 => 
                           regs(2082), A => n748, ZN => n747);
   U868 : INV_X1 port map( A => n749, ZN => n748);
   U869 : AOI222_X1 port map( A1 => regs(34), A2 => n102, B1 => regs(1570), B2 
                           => n204, C1 => regs(546), C2 => n279, ZN => n749);
   U870 : INV_X1 port map( A => n750, ZN => curr_proc_regs(546));
   U871 : AOI221_X1 port map( B1 => n43, B2 => regs(1570), C1 => n323, C2 => 
                           regs(34), A => n751, ZN => n750);
   U872 : INV_X1 port map( A => n752, ZN => n751);
   U873 : AOI222_X1 port map( A1 => regs(546), A2 => n102, B1 => regs(2082), B2
                           => n204, C1 => regs(1058), C2 => n279, ZN => n752);
   U874 : INV_X1 port map( A => n753, ZN => curr_proc_regs(33));
   U875 : AOI221_X1 port map( B1 => n43, B2 => regs(1057), C1 => n323, C2 => 
                           regs(2081), A => n754, ZN => n753);
   U876 : INV_X1 port map( A => n755, ZN => n754);
   U877 : AOI222_X1 port map( A1 => regs(33), A2 => n102, B1 => regs(1569), B2 
                           => n204, C1 => regs(545), C2 => n279, ZN => n755);
   U878 : INV_X1 port map( A => n756, ZN => curr_proc_regs(545));
   U879 : AOI221_X1 port map( B1 => n43, B2 => regs(1569), C1 => n322, C2 => 
                           regs(33), A => n757, ZN => n756);
   U880 : INV_X1 port map( A => n758, ZN => n757);
   U881 : AOI222_X1 port map( A1 => regs(545), A2 => n102, B1 => regs(2081), B2
                           => n204, C1 => regs(1057), C2 => n279, ZN => n758);
   U882 : INV_X1 port map( A => n759, ZN => curr_proc_regs(32));
   U883 : AOI221_X1 port map( B1 => n43, B2 => regs(1056), C1 => n322, C2 => 
                           regs(2080), A => n760, ZN => n759);
   U884 : INV_X1 port map( A => n761, ZN => n760);
   U885 : AOI222_X1 port map( A1 => regs(32), A2 => n102, B1 => regs(1568), B2 
                           => n204, C1 => regs(544), C2 => n279, ZN => n761);
   U886 : INV_X1 port map( A => n762, ZN => curr_proc_regs(544));
   U887 : AOI221_X1 port map( B1 => n43, B2 => regs(1568), C1 => n322, C2 => 
                           regs(32), A => n763, ZN => n762);
   U888 : INV_X1 port map( A => n764, ZN => n763);
   U889 : AOI222_X1 port map( A1 => regs(544), A2 => n102, B1 => regs(2080), B2
                           => n204, C1 => regs(1056), C2 => n279, ZN => n764);
   U890 : INV_X1 port map( A => n765, ZN => curr_proc_regs(607));
   U891 : AOI221_X1 port map( B1 => n43, B2 => regs(1631), C1 => n322, C2 => 
                           regs(95), A => n766, ZN => n765);
   U892 : INV_X1 port map( A => n767, ZN => n766);
   U893 : AOI222_X1 port map( A1 => regs(607), A2 => n102, B1 => regs(2143), B2
                           => n204, C1 => regs(1119), C2 => n279, ZN => n767);
   U894 : INV_X1 port map( A => n768, ZN => curr_proc_regs(95));
   U895 : AOI221_X1 port map( B1 => n27, B2 => regs(1119), C1 => n322, C2 => 
                           regs(2143), A => n769, ZN => n768);
   U896 : INV_X1 port map( A => n770, ZN => n769);
   U897 : AOI222_X1 port map( A1 => regs(95), A2 => n102, B1 => regs(1631), B2 
                           => n204, C1 => regs(607), C2 => n279, ZN => n770);
   U898 : INV_X1 port map( A => n771, ZN => curr_proc_regs(606));
   U899 : AOI221_X1 port map( B1 => n22, B2 => regs(1630), C1 => n327, C2 => 
                           regs(94), A => n772, ZN => n771);
   U900 : INV_X1 port map( A => n773, ZN => n772);
   U901 : AOI222_X1 port map( A1 => regs(606), A2 => n102, B1 => regs(2142), B2
                           => n204, C1 => regs(1118), C2 => n279, ZN => n773);
   U902 : INV_X1 port map( A => n774, ZN => curr_proc_regs(94));
   U903 : AOI221_X1 port map( B1 => n22, B2 => regs(1118), C1 => n343, C2 => 
                           regs(2142), A => n775, ZN => n774);
   U904 : INV_X1 port map( A => n776, ZN => n775);
   U905 : AOI222_X1 port map( A1 => regs(94), A2 => n102, B1 => regs(1630), B2 
                           => n204, C1 => regs(606), C2 => n279, ZN => n776);
   U906 : INV_X1 port map( A => n777, ZN => curr_proc_regs(605));
   U907 : AOI221_X1 port map( B1 => n22, B2 => regs(1629), C1 => n343, C2 => 
                           regs(93), A => n778, ZN => n777);
   U908 : INV_X1 port map( A => n779, ZN => n778);
   U909 : AOI222_X1 port map( A1 => regs(605), A2 => n102, B1 => regs(2141), B2
                           => n203, C1 => regs(1117), C2 => n278, ZN => n779);
   U910 : INV_X1 port map( A => n780, ZN => curr_proc_regs(93));
   U911 : AOI221_X1 port map( B1 => n22, B2 => regs(1117), C1 => n343, C2 => 
                           regs(2141), A => n781, ZN => n780);
   U912 : INV_X1 port map( A => n782, ZN => n781);
   U913 : AOI222_X1 port map( A1 => regs(93), A2 => n102, B1 => regs(1629), B2 
                           => n203, C1 => regs(605), C2 => n278, ZN => n782);
   U914 : INV_X1 port map( A => n783, ZN => curr_proc_regs(604));
   U915 : AOI221_X1 port map( B1 => n22, B2 => regs(1628), C1 => n343, C2 => 
                           regs(92), A => n784, ZN => n783);
   U916 : INV_X1 port map( A => n785, ZN => n784);
   U917 : AOI222_X1 port map( A1 => regs(604), A2 => n103, B1 => regs(2140), B2
                           => n203, C1 => regs(1116), C2 => n278, ZN => n785);
   U918 : INV_X1 port map( A => n786, ZN => curr_proc_regs(92));
   U919 : AOI221_X1 port map( B1 => n22, B2 => regs(1116), C1 => n343, C2 => 
                           regs(2140), A => n787, ZN => n786);
   U920 : INV_X1 port map( A => n788, ZN => n787);
   U921 : AOI222_X1 port map( A1 => regs(92), A2 => n103, B1 => regs(1628), B2 
                           => n203, C1 => regs(604), C2 => n278, ZN => n788);
   U922 : INV_X1 port map( A => n789, ZN => curr_proc_regs(603));
   U923 : AOI221_X1 port map( B1 => n23, B2 => regs(1627), C1 => n343, C2 => 
                           regs(91), A => n790, ZN => n789);
   U924 : INV_X1 port map( A => n791, ZN => n790);
   U925 : AOI222_X1 port map( A1 => regs(603), A2 => n103, B1 => regs(2139), B2
                           => n203, C1 => regs(1115), C2 => n278, ZN => n791);
   U926 : INV_X1 port map( A => n792, ZN => curr_proc_regs(91));
   U927 : AOI221_X1 port map( B1 => n23, B2 => regs(1115), C1 => n343, C2 => 
                           regs(2139), A => n793, ZN => n792);
   U928 : INV_X1 port map( A => n794, ZN => n793);
   U929 : AOI222_X1 port map( A1 => regs(91), A2 => n103, B1 => regs(1627), B2 
                           => n203, C1 => regs(603), C2 => n278, ZN => n794);
   U930 : INV_X1 port map( A => n795, ZN => curr_proc_regs(602));
   U931 : AOI221_X1 port map( B1 => n23, B2 => regs(1626), C1 => n343, C2 => 
                           regs(90), A => n796, ZN => n795);
   U932 : INV_X1 port map( A => n797, ZN => n796);
   U933 : AOI222_X1 port map( A1 => regs(602), A2 => n103, B1 => regs(2138), B2
                           => n203, C1 => regs(1114), C2 => n278, ZN => n797);
   U934 : INV_X1 port map( A => n798, ZN => curr_proc_regs(90));
   U935 : AOI221_X1 port map( B1 => n23, B2 => regs(1114), C1 => n343, C2 => 
                           regs(2138), A => n799, ZN => n798);
   U936 : INV_X1 port map( A => n800, ZN => n799);
   U937 : AOI222_X1 port map( A1 => regs(90), A2 => n103, B1 => regs(1626), B2 
                           => n203, C1 => regs(602), C2 => n278, ZN => n800);
   U938 : INV_X1 port map( A => n801, ZN => curr_proc_regs(601));
   U939 : AOI221_X1 port map( B1 => n23, B2 => regs(1625), C1 => n343, C2 => 
                           regs(89), A => n802, ZN => n801);
   U940 : INV_X1 port map( A => n803, ZN => n802);
   U941 : AOI222_X1 port map( A1 => regs(601), A2 => n103, B1 => regs(2137), B2
                           => n203, C1 => regs(1113), C2 => n278, ZN => n803);
   U942 : INV_X1 port map( A => n804, ZN => curr_proc_regs(89));
   U943 : AOI221_X1 port map( B1 => n23, B2 => regs(1113), C1 => n342, C2 => 
                           regs(2137), A => n805, ZN => n804);
   U944 : INV_X1 port map( A => n806, ZN => n805);
   U945 : AOI222_X1 port map( A1 => regs(89), A2 => n103, B1 => regs(1625), B2 
                           => n203, C1 => regs(601), C2 => n278, ZN => n806);
   U946 : INV_X1 port map( A => n807, ZN => curr_proc_regs(600));
   U947 : AOI221_X1 port map( B1 => n23, B2 => regs(1624), C1 => n342, C2 => 
                           regs(88), A => n808, ZN => n807);
   U948 : INV_X1 port map( A => n809, ZN => n808);
   U949 : AOI222_X1 port map( A1 => regs(600), A2 => n103, B1 => regs(2136), B2
                           => n203, C1 => regs(1112), C2 => n278, ZN => n809);
   U950 : INV_X1 port map( A => n810, ZN => curr_proc_regs(88));
   U951 : AOI221_X1 port map( B1 => n23, B2 => regs(1112), C1 => n342, C2 => 
                           regs(2136), A => n811, ZN => n810);
   U952 : INV_X1 port map( A => n812, ZN => n811);
   U953 : AOI222_X1 port map( A1 => regs(88), A2 => n103, B1 => regs(1624), B2 
                           => n203, C1 => regs(600), C2 => n278, ZN => n812);
   U954 : INV_X1 port map( A => n813, ZN => curr_proc_regs(599));
   U955 : AOI221_X1 port map( B1 => n23, B2 => regs(1623), C1 => n342, C2 => 
                           regs(87), A => n814, ZN => n813);
   U956 : INV_X1 port map( A => n815, ZN => n814);
   U957 : AOI222_X1 port map( A1 => regs(599), A2 => n103, B1 => regs(2135), B2
                           => n202, C1 => regs(1111), C2 => n277, ZN => n815);
   U958 : INV_X1 port map( A => n816, ZN => curr_proc_regs(87));
   U959 : AOI221_X1 port map( B1 => n23, B2 => regs(1111), C1 => n342, C2 => 
                           regs(2135), A => n817, ZN => n816);
   U960 : INV_X1 port map( A => n818, ZN => n817);
   U961 : AOI222_X1 port map( A1 => regs(87), A2 => n103, B1 => regs(1623), B2 
                           => n202, C1 => regs(599), C2 => n277, ZN => n818);
   U962 : INV_X1 port map( A => n819, ZN => curr_proc_regs(598));
   U963 : AOI221_X1 port map( B1 => n23, B2 => regs(1622), C1 => n342, C2 => 
                           regs(86), A => n820, ZN => n819);
   U964 : INV_X1 port map( A => n821, ZN => n820);
   U965 : AOI222_X1 port map( A1 => regs(598), A2 => n104, B1 => regs(2134), B2
                           => n202, C1 => regs(1110), C2 => n277, ZN => n821);
   U966 : INV_X1 port map( A => n822, ZN => curr_proc_regs(86));
   U967 : AOI221_X1 port map( B1 => n23, B2 => regs(1110), C1 => n342, C2 => 
                           regs(2134), A => n823, ZN => n822);
   U968 : INV_X1 port map( A => n824, ZN => n823);
   U969 : AOI222_X1 port map( A1 => regs(86), A2 => n104, B1 => regs(1622), B2 
                           => n202, C1 => regs(598), C2 => n277, ZN => n824);
   U970 : INV_X1 port map( A => n825, ZN => curr_proc_regs(597));
   U971 : AOI221_X1 port map( B1 => n24, B2 => regs(1621), C1 => n342, C2 => 
                           regs(85), A => n826, ZN => n825);
   U972 : INV_X1 port map( A => n827, ZN => n826);
   U973 : AOI222_X1 port map( A1 => regs(597), A2 => n104, B1 => regs(2133), B2
                           => n202, C1 => regs(1109), C2 => n277, ZN => n827);
   U974 : INV_X1 port map( A => n828, ZN => curr_proc_regs(85));
   U975 : AOI221_X1 port map( B1 => n24, B2 => regs(1109), C1 => n342, C2 => 
                           regs(2133), A => n829, ZN => n828);
   U976 : INV_X1 port map( A => n830, ZN => n829);
   U977 : AOI222_X1 port map( A1 => regs(85), A2 => n104, B1 => regs(1621), B2 
                           => n202, C1 => regs(597), C2 => n277, ZN => n830);
   U978 : INV_X1 port map( A => n831, ZN => curr_proc_regs(596));
   U979 : AOI221_X1 port map( B1 => n24, B2 => regs(1620), C1 => n342, C2 => 
                           regs(84), A => n832, ZN => n831);
   U980 : INV_X1 port map( A => n833, ZN => n832);
   U981 : AOI222_X1 port map( A1 => regs(596), A2 => n104, B1 => regs(2132), B2
                           => n202, C1 => regs(1108), C2 => n277, ZN => n833);
   U982 : INV_X1 port map( A => n834, ZN => curr_proc_regs(84));
   U983 : AOI221_X1 port map( B1 => n24, B2 => regs(1108), C1 => n342, C2 => 
                           regs(2132), A => n835, ZN => n834);
   U984 : INV_X1 port map( A => n836, ZN => n835);
   U985 : AOI222_X1 port map( A1 => regs(84), A2 => n104, B1 => regs(1620), B2 
                           => n202, C1 => regs(596), C2 => n277, ZN => n836);
   U986 : INV_X1 port map( A => n837, ZN => curr_proc_regs(595));
   U987 : AOI221_X1 port map( B1 => n24, B2 => regs(1619), C1 => n342, C2 => 
                           regs(83), A => n838, ZN => n837);
   U988 : INV_X1 port map( A => n839, ZN => n838);
   U989 : AOI222_X1 port map( A1 => regs(595), A2 => n104, B1 => regs(2131), B2
                           => n202, C1 => regs(1107), C2 => n277, ZN => n839);
   U990 : INV_X1 port map( A => n840, ZN => curr_proc_regs(83));
   U991 : AOI221_X1 port map( B1 => n24, B2 => regs(1107), C1 => n341, C2 => 
                           regs(2131), A => n841, ZN => n840);
   U992 : INV_X1 port map( A => n842, ZN => n841);
   U993 : AOI222_X1 port map( A1 => regs(83), A2 => n104, B1 => regs(1619), B2 
                           => n202, C1 => regs(595), C2 => n277, ZN => n842);
   U994 : INV_X1 port map( A => n843, ZN => curr_proc_regs(594));
   U995 : AOI221_X1 port map( B1 => n24, B2 => regs(1618), C1 => n341, C2 => 
                           regs(82), A => n844, ZN => n843);
   U996 : INV_X1 port map( A => n845, ZN => n844);
   U997 : AOI222_X1 port map( A1 => regs(594), A2 => n104, B1 => regs(2130), B2
                           => n202, C1 => regs(1106), C2 => n277, ZN => n845);
   U998 : INV_X1 port map( A => n846, ZN => curr_proc_regs(82));
   U999 : AOI221_X1 port map( B1 => n24, B2 => regs(1106), C1 => n341, C2 => 
                           regs(2130), A => n847, ZN => n846);
   U1000 : INV_X1 port map( A => n848, ZN => n847);
   U1001 : AOI222_X1 port map( A1 => regs(82), A2 => n104, B1 => regs(1618), B2
                           => n202, C1 => regs(594), C2 => n277, ZN => n848);
   U1002 : INV_X1 port map( A => n849, ZN => curr_proc_regs(593));
   U1003 : AOI221_X1 port map( B1 => n24, B2 => regs(1617), C1 => n341, C2 => 
                           regs(81), A => n850, ZN => n849);
   U1004 : INV_X1 port map( A => n851, ZN => n850);
   U1005 : AOI222_X1 port map( A1 => regs(593), A2 => n104, B1 => regs(2129), 
                           B2 => n201, C1 => regs(1105), C2 => n276, ZN => n851
                           );
   U1006 : INV_X1 port map( A => n852, ZN => curr_proc_regs(81));
   U1007 : AOI221_X1 port map( B1 => n24, B2 => regs(1105), C1 => n341, C2 => 
                           regs(2129), A => n853, ZN => n852);
   U1008 : INV_X1 port map( A => n854, ZN => n853);
   U1009 : AOI222_X1 port map( A1 => regs(81), A2 => n104, B1 => regs(1617), B2
                           => n201, C1 => regs(593), C2 => n276, ZN => n854);
   U1010 : INV_X1 port map( A => n855, ZN => curr_proc_regs(592));
   U1011 : AOI221_X1 port map( B1 => n24, B2 => regs(1616), C1 => n341, C2 => 
                           regs(80), A => n856, ZN => n855);
   U1012 : INV_X1 port map( A => n857, ZN => n856);
   U1013 : AOI222_X1 port map( A1 => regs(592), A2 => n105, B1 => regs(2128), 
                           B2 => n201, C1 => regs(1104), C2 => n276, ZN => n857
                           );
   U1014 : INV_X1 port map( A => n858, ZN => curr_proc_regs(80));
   U1015 : AOI221_X1 port map( B1 => n24, B2 => regs(1104), C1 => n341, C2 => 
                           regs(2128), A => n859, ZN => n858);
   U1016 : INV_X1 port map( A => n860, ZN => n859);
   U1017 : AOI222_X1 port map( A1 => regs(80), A2 => n105, B1 => regs(1616), B2
                           => n201, C1 => regs(592), C2 => n276, ZN => n860);
   U1018 : INV_X1 port map( A => n861, ZN => curr_proc_regs(591));
   U1019 : AOI221_X1 port map( B1 => n25, B2 => regs(1615), C1 => n341, C2 => 
                           regs(79), A => n862, ZN => n861);
   U1020 : INV_X1 port map( A => n863, ZN => n862);
   U1021 : AOI222_X1 port map( A1 => regs(591), A2 => n105, B1 => regs(2127), 
                           B2 => n201, C1 => regs(1103), C2 => n276, ZN => n863
                           );
   U1022 : INV_X1 port map( A => n864, ZN => curr_proc_regs(79));
   U1023 : AOI221_X1 port map( B1 => n25, B2 => regs(1103), C1 => n341, C2 => 
                           regs(2127), A => n865, ZN => n864);
   U1024 : INV_X1 port map( A => n866, ZN => n865);
   U1025 : AOI222_X1 port map( A1 => regs(79), A2 => n105, B1 => regs(1615), B2
                           => n201, C1 => regs(591), C2 => n276, ZN => n866);
   U1026 : INV_X1 port map( A => n867, ZN => curr_proc_regs(590));
   U1027 : AOI221_X1 port map( B1 => n25, B2 => regs(1614), C1 => n341, C2 => 
                           regs(78), A => n868, ZN => n867);
   U1028 : INV_X1 port map( A => n869, ZN => n868);
   U1029 : AOI222_X1 port map( A1 => regs(590), A2 => n105, B1 => regs(2126), 
                           B2 => n201, C1 => regs(1102), C2 => n276, ZN => n869
                           );
   U1030 : INV_X1 port map( A => n870, ZN => curr_proc_regs(78));
   U1031 : AOI221_X1 port map( B1 => n25, B2 => regs(1102), C1 => n341, C2 => 
                           regs(2126), A => n871, ZN => n870);
   U1032 : INV_X1 port map( A => n872, ZN => n871);
   U1033 : AOI222_X1 port map( A1 => regs(78), A2 => n105, B1 => regs(1614), B2
                           => n201, C1 => regs(590), C2 => n276, ZN => n872);
   U1034 : INV_X1 port map( A => n873, ZN => curr_proc_regs(589));
   U1035 : AOI221_X1 port map( B1 => n25, B2 => regs(1613), C1 => n341, C2 => 
                           regs(77), A => n874, ZN => n873);
   U1036 : INV_X1 port map( A => n875, ZN => n874);
   U1037 : AOI222_X1 port map( A1 => regs(589), A2 => n105, B1 => regs(2125), 
                           B2 => n201, C1 => regs(1101), C2 => n276, ZN => n875
                           );
   U1038 : INV_X1 port map( A => n876, ZN => curr_proc_regs(77));
   U1039 : AOI221_X1 port map( B1 => n25, B2 => regs(1101), C1 => n340, C2 => 
                           regs(2125), A => n877, ZN => n876);
   U1040 : INV_X1 port map( A => n878, ZN => n877);
   U1041 : AOI222_X1 port map( A1 => regs(77), A2 => n105, B1 => regs(1613), B2
                           => n201, C1 => regs(589), C2 => n276, ZN => n878);
   U1042 : INV_X1 port map( A => n879, ZN => curr_proc_regs(588));
   U1043 : AOI221_X1 port map( B1 => n25, B2 => regs(1612), C1 => n340, C2 => 
                           regs(76), A => n880, ZN => n879);
   U1044 : INV_X1 port map( A => n881, ZN => n880);
   U1045 : AOI222_X1 port map( A1 => regs(588), A2 => n105, B1 => regs(2124), 
                           B2 => n201, C1 => regs(1100), C2 => n276, ZN => n881
                           );
   U1046 : INV_X1 port map( A => n882, ZN => curr_proc_regs(76));
   U1047 : AOI221_X1 port map( B1 => n25, B2 => regs(1100), C1 => n340, C2 => 
                           regs(2124), A => n883, ZN => n882);
   U1048 : INV_X1 port map( A => n884, ZN => n883);
   U1049 : AOI222_X1 port map( A1 => regs(76), A2 => n105, B1 => regs(1612), B2
                           => n201, C1 => regs(588), C2 => n276, ZN => n884);
   U1050 : INV_X1 port map( A => n885, ZN => curr_proc_regs(587));
   U1051 : AOI221_X1 port map( B1 => n25, B2 => regs(1611), C1 => n340, C2 => 
                           regs(75), A => n886, ZN => n885);
   U1052 : INV_X1 port map( A => n887, ZN => n886);
   U1053 : AOI222_X1 port map( A1 => regs(587), A2 => n105, B1 => regs(2123), 
                           B2 => n200, C1 => regs(1099), C2 => n275, ZN => n887
                           );
   U1054 : INV_X1 port map( A => n888, ZN => curr_proc_regs(75));
   U1055 : AOI221_X1 port map( B1 => n25, B2 => regs(1099), C1 => n340, C2 => 
                           regs(2123), A => n889, ZN => n888);
   U1056 : INV_X1 port map( A => n890, ZN => n889);
   U1057 : AOI222_X1 port map( A1 => regs(75), A2 => n105, B1 => regs(1611), B2
                           => n200, C1 => regs(587), C2 => n275, ZN => n890);
   U1058 : INV_X1 port map( A => n891, ZN => curr_proc_regs(586));
   U1059 : AOI221_X1 port map( B1 => n25, B2 => regs(1610), C1 => n340, C2 => 
                           regs(74), A => n892, ZN => n891);
   U1060 : INV_X1 port map( A => n893, ZN => n892);
   U1061 : AOI222_X1 port map( A1 => regs(586), A2 => n106, B1 => regs(2122), 
                           B2 => n200, C1 => regs(1098), C2 => n275, ZN => n893
                           );
   U1062 : INV_X1 port map( A => n894, ZN => curr_proc_regs(74));
   U1063 : AOI221_X1 port map( B1 => n25, B2 => regs(1098), C1 => n340, C2 => 
                           regs(2122), A => n895, ZN => n894);
   U1064 : INV_X1 port map( A => n896, ZN => n895);
   U1065 : AOI222_X1 port map( A1 => regs(74), A2 => n106, B1 => regs(1610), B2
                           => n200, C1 => regs(586), C2 => n275, ZN => n896);
   U1066 : INV_X1 port map( A => n897, ZN => curr_proc_regs(585));
   U1067 : AOI221_X1 port map( B1 => n26, B2 => regs(1609), C1 => n340, C2 => 
                           regs(73), A => n898, ZN => n897);
   U1068 : INV_X1 port map( A => n899, ZN => n898);
   U1069 : AOI222_X1 port map( A1 => regs(585), A2 => n106, B1 => regs(2121), 
                           B2 => n200, C1 => regs(1097), C2 => n275, ZN => n899
                           );
   U1070 : INV_X1 port map( A => n900, ZN => curr_proc_regs(73));
   U1071 : AOI221_X1 port map( B1 => n26, B2 => regs(1097), C1 => n340, C2 => 
                           regs(2121), A => n901, ZN => n900);
   U1072 : INV_X1 port map( A => n902, ZN => n901);
   U1073 : AOI222_X1 port map( A1 => regs(73), A2 => n106, B1 => regs(1609), B2
                           => n200, C1 => regs(585), C2 => n275, ZN => n902);
   U1074 : INV_X1 port map( A => n903, ZN => curr_proc_regs(584));
   U1075 : AOI221_X1 port map( B1 => n26, B2 => regs(1608), C1 => n340, C2 => 
                           regs(72), A => n904, ZN => n903);
   U1076 : INV_X1 port map( A => n905, ZN => n904);
   U1077 : AOI222_X1 port map( A1 => regs(584), A2 => n106, B1 => regs(2120), 
                           B2 => n200, C1 => regs(1096), C2 => n275, ZN => n905
                           );
   U1078 : INV_X1 port map( A => n906, ZN => curr_proc_regs(72));
   U1079 : AOI221_X1 port map( B1 => n26, B2 => regs(1096), C1 => n340, C2 => 
                           regs(2120), A => n907, ZN => n906);
   U1080 : INV_X1 port map( A => n908, ZN => n907);
   U1081 : AOI222_X1 port map( A1 => regs(72), A2 => n106, B1 => regs(1608), B2
                           => n200, C1 => regs(584), C2 => n275, ZN => n908);
   U1082 : INV_X1 port map( A => n909, ZN => curr_proc_regs(583));
   U1083 : AOI221_X1 port map( B1 => n26, B2 => regs(1607), C1 => n340, C2 => 
                           regs(71), A => n910, ZN => n909);
   U1084 : INV_X1 port map( A => n911, ZN => n910);
   U1085 : AOI222_X1 port map( A1 => regs(583), A2 => n106, B1 => regs(2119), 
                           B2 => n200, C1 => regs(1095), C2 => n275, ZN => n911
                           );
   U1086 : INV_X1 port map( A => n912, ZN => curr_proc_regs(71));
   U1087 : AOI221_X1 port map( B1 => n26, B2 => regs(1095), C1 => n339, C2 => 
                           regs(2119), A => n913, ZN => n912);
   U1088 : INV_X1 port map( A => n914, ZN => n913);
   U1089 : AOI222_X1 port map( A1 => regs(71), A2 => n106, B1 => regs(1607), B2
                           => n200, C1 => regs(583), C2 => n275, ZN => n914);
   U1090 : INV_X1 port map( A => n915, ZN => curr_proc_regs(582));
   U1091 : AOI221_X1 port map( B1 => n26, B2 => regs(1606), C1 => n339, C2 => 
                           regs(70), A => n916, ZN => n915);
   U1092 : INV_X1 port map( A => n917, ZN => n916);
   U1093 : AOI222_X1 port map( A1 => regs(582), A2 => n106, B1 => regs(2118), 
                           B2 => n200, C1 => regs(1094), C2 => n275, ZN => n917
                           );
   U1094 : INV_X1 port map( A => n918, ZN => curr_proc_regs(70));
   U1095 : AOI221_X1 port map( B1 => n26, B2 => regs(1094), C1 => n339, C2 => 
                           regs(2118), A => n919, ZN => n918);
   U1096 : INV_X1 port map( A => n920, ZN => n919);
   U1097 : AOI222_X1 port map( A1 => regs(70), A2 => n106, B1 => regs(1606), B2
                           => n200, C1 => regs(582), C2 => n275, ZN => n920);
   U1098 : INV_X1 port map( A => n921, ZN => curr_proc_regs(581));
   U1099 : AOI221_X1 port map( B1 => n26, B2 => regs(1605), C1 => n339, C2 => 
                           regs(69), A => n922, ZN => n921);
   U1100 : INV_X1 port map( A => n923, ZN => n922);
   U1101 : AOI222_X1 port map( A1 => regs(581), A2 => n106, B1 => regs(2117), 
                           B2 => n199, C1 => regs(1093), C2 => n274, ZN => n923
                           );
   U1102 : INV_X1 port map( A => n924, ZN => curr_proc_regs(69));
   U1103 : AOI221_X1 port map( B1 => n26, B2 => regs(1093), C1 => n339, C2 => 
                           regs(2117), A => n925, ZN => n924);
   U1104 : INV_X1 port map( A => n926, ZN => n925);
   U1105 : AOI222_X1 port map( A1 => regs(69), A2 => n106, B1 => regs(1605), B2
                           => n199, C1 => regs(581), C2 => n274, ZN => n926);
   U1106 : INV_X1 port map( A => n927, ZN => curr_proc_regs(580));
   U1107 : AOI221_X1 port map( B1 => n26, B2 => regs(1604), C1 => n339, C2 => 
                           regs(68), A => n928, ZN => n927);
   U1108 : INV_X1 port map( A => n929, ZN => n928);
   U1109 : AOI222_X1 port map( A1 => regs(580), A2 => n107, B1 => regs(2116), 
                           B2 => n199, C1 => regs(1092), C2 => n274, ZN => n929
                           );
   U1110 : INV_X1 port map( A => n930, ZN => curr_proc_regs(68));
   U1111 : AOI221_X1 port map( B1 => n26, B2 => regs(1092), C1 => n339, C2 => 
                           regs(2116), A => n931, ZN => n930);
   U1112 : INV_X1 port map( A => n932, ZN => n931);
   U1113 : AOI222_X1 port map( A1 => regs(68), A2 => n107, B1 => regs(1604), B2
                           => n199, C1 => regs(580), C2 => n274, ZN => n932);
   U1114 : INV_X1 port map( A => n933, ZN => curr_proc_regs(579));
   U1115 : AOI221_X1 port map( B1 => n27, B2 => regs(1603), C1 => n339, C2 => 
                           regs(67), A => n934, ZN => n933);
   U1116 : INV_X1 port map( A => n935, ZN => n934);
   U1117 : AOI222_X1 port map( A1 => regs(579), A2 => n107, B1 => regs(2115), 
                           B2 => n199, C1 => regs(1091), C2 => n274, ZN => n935
                           );
   U1118 : INV_X1 port map( A => n936, ZN => curr_proc_regs(67));
   U1119 : AOI221_X1 port map( B1 => n27, B2 => regs(1091), C1 => n339, C2 => 
                           regs(2115), A => n937, ZN => n936);
   U1120 : INV_X1 port map( A => n938, ZN => n937);
   U1121 : AOI222_X1 port map( A1 => regs(67), A2 => n107, B1 => regs(1603), B2
                           => n199, C1 => regs(579), C2 => n274, ZN => n938);
   U1122 : INV_X1 port map( A => n939, ZN => curr_proc_regs(578));
   U1123 : AOI221_X1 port map( B1 => n27, B2 => regs(1602), C1 => n339, C2 => 
                           regs(66), A => n940, ZN => n939);
   U1124 : INV_X1 port map( A => n941, ZN => n940);
   U1125 : AOI222_X1 port map( A1 => regs(578), A2 => n107, B1 => regs(2114), 
                           B2 => n199, C1 => regs(1090), C2 => n274, ZN => n941
                           );
   U1126 : INV_X1 port map( A => n942, ZN => curr_proc_regs(66));
   U1127 : AOI221_X1 port map( B1 => n27, B2 => regs(1090), C1 => n339, C2 => 
                           regs(2114), A => n943, ZN => n942);
   U1128 : INV_X1 port map( A => n944, ZN => n943);
   U1129 : AOI222_X1 port map( A1 => regs(66), A2 => n107, B1 => regs(1602), B2
                           => n199, C1 => regs(578), C2 => n274, ZN => n944);
   U1130 : INV_X1 port map( A => n945, ZN => curr_proc_regs(577));
   U1131 : AOI221_X1 port map( B1 => n27, B2 => regs(1601), C1 => n339, C2 => 
                           regs(65), A => n946, ZN => n945);
   U1132 : INV_X1 port map( A => n947, ZN => n946);
   U1133 : AOI222_X1 port map( A1 => regs(577), A2 => n107, B1 => regs(2113), 
                           B2 => n199, C1 => regs(1089), C2 => n274, ZN => n947
                           );
   U1134 : INV_X1 port map( A => n948, ZN => curr_proc_regs(65));
   U1135 : AOI221_X1 port map( B1 => n27, B2 => regs(1089), C1 => n338, C2 => 
                           regs(2113), A => n949, ZN => n948);
   U1136 : INV_X1 port map( A => n950, ZN => n949);
   U1137 : AOI222_X1 port map( A1 => regs(65), A2 => n107, B1 => regs(1601), B2
                           => n199, C1 => regs(577), C2 => n274, ZN => n950);
   U1138 : INV_X1 port map( A => n951, ZN => curr_proc_regs(576));
   U1139 : AOI221_X1 port map( B1 => n27, B2 => regs(1600), C1 => n338, C2 => 
                           regs(64), A => n952, ZN => n951);
   U1140 : INV_X1 port map( A => n953, ZN => n952);
   U1141 : AOI222_X1 port map( A1 => regs(576), A2 => n107, B1 => regs(2112), 
                           B2 => n199, C1 => regs(1088), C2 => n274, ZN => n953
                           );
   U1142 : INV_X1 port map( A => n954, ZN => curr_proc_regs(64));
   U1143 : AOI221_X1 port map( B1 => n27, B2 => regs(1088), C1 => n338, C2 => 
                           regs(2112), A => n955, ZN => n954);
   U1144 : INV_X1 port map( A => n956, ZN => n955);
   U1145 : AOI222_X1 port map( A1 => regs(64), A2 => n107, B1 => regs(1600), B2
                           => n199, C1 => regs(576), C2 => n274, ZN => n956);
   U1146 : INV_X1 port map( A => n957, ZN => curr_proc_regs(127));
   U1147 : AOI221_X1 port map( B1 => n27, B2 => regs(1151), C1 => n338, C2 => 
                           regs(2175), A => n958, ZN => n957);
   U1148 : INV_X1 port map( A => n959, ZN => n958);
   U1149 : AOI222_X1 port map( A1 => regs(127), A2 => n107, B1 => regs(1663), 
                           B2 => n198, C1 => regs(639), C2 => n273, ZN => n959)
                           ;
   U1150 : INV_X1 port map( A => n960, ZN => curr_proc_regs(639));
   U1151 : AOI221_X1 port map( B1 => n27, B2 => regs(1663), C1 => n338, C2 => 
                           regs(127), A => n961, ZN => n960);
   U1152 : INV_X1 port map( A => n962, ZN => n961);
   U1153 : AOI222_X1 port map( A1 => regs(639), A2 => n83, B1 => regs(2175), B2
                           => n198, C1 => regs(1151), C2 => n273, ZN => n962);
   U1154 : INV_X1 port map( A => n963, ZN => curr_proc_regs(126));
   U1155 : AOI221_X1 port map( B1 => n27, B2 => regs(1150), C1 => n338, C2 => 
                           regs(2174), A => n964, ZN => n963);
   U1156 : INV_X1 port map( A => n965, ZN => n964);
   U1157 : AOI222_X1 port map( A1 => regs(126), A2 => n76, B1 => regs(1662), B2
                           => n198, C1 => regs(638), C2 => n273, ZN => n965);
   U1158 : INV_X1 port map( A => n966, ZN => curr_proc_regs(638));
   U1159 : AOI221_X1 port map( B1 => n28, B2 => regs(1662), C1 => n338, C2 => 
                           regs(126), A => n967, ZN => n966);
   U1160 : INV_X1 port map( A => n968, ZN => n967);
   U1161 : AOI222_X1 port map( A1 => regs(638), A2 => n76, B1 => regs(2174), B2
                           => n198, C1 => regs(1150), C2 => n273, ZN => n968);
   U1162 : INV_X1 port map( A => n969, ZN => curr_proc_regs(125));
   U1163 : AOI221_X1 port map( B1 => n28, B2 => regs(1149), C1 => n338, C2 => 
                           regs(2173), A => n970, ZN => n969);
   U1164 : INV_X1 port map( A => n971, ZN => n970);
   U1165 : AOI222_X1 port map( A1 => regs(125), A2 => n76, B1 => regs(1661), B2
                           => n198, C1 => regs(637), C2 => n273, ZN => n971);
   U1166 : INV_X1 port map( A => n972, ZN => curr_proc_regs(637));
   U1167 : AOI221_X1 port map( B1 => n28, B2 => regs(1661), C1 => n338, C2 => 
                           regs(125), A => n973, ZN => n972);
   U1168 : INV_X1 port map( A => n974, ZN => n973);
   U1169 : AOI222_X1 port map( A1 => regs(637), A2 => n76, B1 => regs(2173), B2
                           => n198, C1 => regs(1149), C2 => n273, ZN => n974);
   U1170 : INV_X1 port map( A => n975, ZN => curr_proc_regs(124));
   U1171 : AOI221_X1 port map( B1 => n28, B2 => regs(1148), C1 => n338, C2 => 
                           regs(2172), A => n976, ZN => n975);
   U1172 : INV_X1 port map( A => n977, ZN => n976);
   U1173 : AOI222_X1 port map( A1 => regs(124), A2 => n76, B1 => regs(1660), B2
                           => n198, C1 => regs(636), C2 => n273, ZN => n977);
   U1174 : INV_X1 port map( A => n978, ZN => curr_proc_regs(636));
   U1175 : AOI221_X1 port map( B1 => n28, B2 => regs(1660), C1 => n338, C2 => 
                           regs(124), A => n979, ZN => n978);
   U1176 : INV_X1 port map( A => n980, ZN => n979);
   U1177 : AOI222_X1 port map( A1 => regs(636), A2 => n76, B1 => regs(2172), B2
                           => n198, C1 => regs(1148), C2 => n273, ZN => n980);
   U1178 : INV_X1 port map( A => n981, ZN => curr_proc_regs(123));
   U1179 : AOI221_X1 port map( B1 => n28, B2 => regs(1147), C1 => n338, C2 => 
                           regs(2171), A => n982, ZN => n981);
   U1180 : INV_X1 port map( A => n983, ZN => n982);
   U1181 : AOI222_X1 port map( A1 => regs(123), A2 => n76, B1 => regs(1659), B2
                           => n198, C1 => regs(635), C2 => n273, ZN => n983);
   U1182 : INV_X1 port map( A => n984, ZN => curr_proc_regs(635));
   U1183 : AOI221_X1 port map( B1 => n28, B2 => regs(1659), C1 => n337, C2 => 
                           regs(123), A => n985, ZN => n984);
   U1184 : INV_X1 port map( A => n986, ZN => n985);
   U1185 : AOI222_X1 port map( A1 => regs(635), A2 => n76, B1 => regs(2171), B2
                           => n198, C1 => regs(1147), C2 => n273, ZN => n986);
   U1186 : INV_X1 port map( A => n987, ZN => curr_proc_regs(122));
   U1187 : AOI221_X1 port map( B1 => n28, B2 => regs(1146), C1 => n337, C2 => 
                           regs(2170), A => n988, ZN => n987);
   U1188 : INV_X1 port map( A => n989, ZN => n988);
   U1189 : AOI222_X1 port map( A1 => regs(122), A2 => n76, B1 => regs(1658), B2
                           => n198, C1 => regs(634), C2 => n273, ZN => n989);
   U1190 : INV_X1 port map( A => n990, ZN => curr_proc_regs(634));
   U1191 : AOI221_X1 port map( B1 => n28, B2 => regs(1658), C1 => n337, C2 => 
                           regs(122), A => n991, ZN => n990);
   U1192 : INV_X1 port map( A => n992, ZN => n991);
   U1193 : AOI222_X1 port map( A1 => regs(634), A2 => n76, B1 => regs(2170), B2
                           => n198, C1 => regs(1146), C2 => n273, ZN => n992);
   U1194 : INV_X1 port map( A => n993, ZN => curr_proc_regs(121));
   U1195 : AOI221_X1 port map( B1 => n28, B2 => regs(1145), C1 => n337, C2 => 
                           regs(2169), A => n994, ZN => n993);
   U1196 : INV_X1 port map( A => n995, ZN => n994);
   U1197 : AOI222_X1 port map( A1 => regs(121), A2 => n76, B1 => regs(1657), B2
                           => n197, C1 => regs(633), C2 => n272, ZN => n995);
   U1198 : INV_X1 port map( A => n996, ZN => curr_proc_regs(633));
   U1199 : AOI221_X1 port map( B1 => n28, B2 => regs(1657), C1 => n337, C2 => 
                           regs(121), A => n997, ZN => n996);
   U1200 : INV_X1 port map( A => n998, ZN => n997);
   U1201 : AOI222_X1 port map( A1 => regs(633), A2 => n77, B1 => regs(2169), B2
                           => n197, C1 => regs(1145), C2 => n272, ZN => n998);
   U1202 : INV_X1 port map( A => n999, ZN => curr_proc_regs(120));
   U1203 : AOI221_X1 port map( B1 => n28, B2 => regs(1144), C1 => n337, C2 => 
                           regs(2168), A => n1000, ZN => n999);
   U1204 : INV_X1 port map( A => n1001, ZN => n1000);
   U1205 : AOI222_X1 port map( A1 => regs(120), A2 => n77, B1 => regs(1656), B2
                           => n197, C1 => regs(632), C2 => n272, ZN => n1001);
   U1206 : INV_X1 port map( A => n1002, ZN => curr_proc_regs(632));
   U1207 : AOI221_X1 port map( B1 => n29, B2 => regs(1656), C1 => n337, C2 => 
                           regs(120), A => n1003, ZN => n1002);
   U1208 : INV_X1 port map( A => n1004, ZN => n1003);
   U1209 : AOI222_X1 port map( A1 => regs(632), A2 => n77, B1 => regs(2168), B2
                           => n197, C1 => regs(1144), C2 => n272, ZN => n1004);
   U1210 : INV_X1 port map( A => n1005, ZN => curr_proc_regs(119));
   U1211 : AOI221_X1 port map( B1 => n29, B2 => regs(1143), C1 => n337, C2 => 
                           regs(2167), A => n1006, ZN => n1005);
   U1212 : INV_X1 port map( A => n1007, ZN => n1006);
   U1213 : AOI222_X1 port map( A1 => regs(119), A2 => n77, B1 => regs(1655), B2
                           => n197, C1 => regs(631), C2 => n272, ZN => n1007);
   U1214 : INV_X1 port map( A => n1008, ZN => curr_proc_regs(631));
   U1215 : AOI221_X1 port map( B1 => n29, B2 => regs(1655), C1 => n337, C2 => 
                           regs(119), A => n1009, ZN => n1008);
   U1216 : INV_X1 port map( A => n1010, ZN => n1009);
   U1217 : AOI222_X1 port map( A1 => regs(631), A2 => n77, B1 => regs(2167), B2
                           => n197, C1 => regs(1143), C2 => n272, ZN => n1010);
   U1218 : INV_X1 port map( A => n1011, ZN => curr_proc_regs(118));
   U1219 : AOI221_X1 port map( B1 => n29, B2 => regs(1142), C1 => n337, C2 => 
                           regs(2166), A => n1012, ZN => n1011);
   U1220 : INV_X1 port map( A => n1013, ZN => n1012);
   U1221 : AOI222_X1 port map( A1 => regs(118), A2 => n77, B1 => regs(1654), B2
                           => n197, C1 => regs(630), C2 => n272, ZN => n1013);
   U1222 : INV_X1 port map( A => n1014, ZN => curr_proc_regs(630));
   U1223 : AOI221_X1 port map( B1 => n29, B2 => regs(1654), C1 => n337, C2 => 
                           regs(118), A => n1015, ZN => n1014);
   U1224 : INV_X1 port map( A => n1016, ZN => n1015);
   U1225 : AOI222_X1 port map( A1 => regs(630), A2 => n77, B1 => regs(2166), B2
                           => n197, C1 => regs(1142), C2 => n272, ZN => n1016);
   U1226 : INV_X1 port map( A => n1017, ZN => curr_proc_regs(117));
   U1227 : AOI221_X1 port map( B1 => n29, B2 => regs(1141), C1 => n337, C2 => 
                           regs(2165), A => n1018, ZN => n1017);
   U1228 : INV_X1 port map( A => n1019, ZN => n1018);
   U1229 : AOI222_X1 port map( A1 => regs(117), A2 => n77, B1 => regs(1653), B2
                           => n197, C1 => regs(629), C2 => n272, ZN => n1019);
   U1230 : INV_X1 port map( A => n1020, ZN => curr_proc_regs(629));
   U1231 : AOI221_X1 port map( B1 => n29, B2 => regs(1653), C1 => n336, C2 => 
                           regs(117), A => n1021, ZN => n1020);
   U1232 : INV_X1 port map( A => n1022, ZN => n1021);
   U1233 : AOI222_X1 port map( A1 => regs(629), A2 => n77, B1 => regs(2165), B2
                           => n197, C1 => regs(1141), C2 => n272, ZN => n1022);
   U1234 : INV_X1 port map( A => n1023, ZN => curr_proc_regs(116));
   U1235 : AOI221_X1 port map( B1 => n29, B2 => regs(1140), C1 => n336, C2 => 
                           regs(2164), A => n1024, ZN => n1023);
   U1236 : INV_X1 port map( A => n1025, ZN => n1024);
   U1237 : AOI222_X1 port map( A1 => regs(116), A2 => n77, B1 => regs(1652), B2
                           => n197, C1 => regs(628), C2 => n272, ZN => n1025);
   U1238 : INV_X1 port map( A => n1026, ZN => curr_proc_regs(628));
   U1239 : AOI221_X1 port map( B1 => n29, B2 => regs(1652), C1 => n336, C2 => 
                           regs(116), A => n1027, ZN => n1026);
   U1240 : INV_X1 port map( A => n1028, ZN => n1027);
   U1241 : AOI222_X1 port map( A1 => regs(628), A2 => n77, B1 => regs(2164), B2
                           => n197, C1 => regs(1140), C2 => n272, ZN => n1028);
   U1242 : INV_X1 port map( A => n1029, ZN => curr_proc_regs(115));
   U1243 : AOI221_X1 port map( B1 => n29, B2 => regs(1139), C1 => n336, C2 => 
                           regs(2163), A => n1030, ZN => n1029);
   U1244 : INV_X1 port map( A => n1031, ZN => n1030);
   U1245 : AOI222_X1 port map( A1 => regs(115), A2 => n77, B1 => regs(1651), B2
                           => n196, C1 => regs(627), C2 => n271, ZN => n1031);
   U1246 : INV_X1 port map( A => n1032, ZN => curr_proc_regs(627));
   U1247 : AOI221_X1 port map( B1 => n29, B2 => regs(1651), C1 => n336, C2 => 
                           regs(115), A => n1033, ZN => n1032);
   U1248 : INV_X1 port map( A => n1034, ZN => n1033);
   U1249 : AOI222_X1 port map( A1 => regs(627), A2 => n78, B1 => regs(2163), B2
                           => n196, C1 => regs(1139), C2 => n271, ZN => n1034);
   U1250 : INV_X1 port map( A => n1035, ZN => curr_proc_regs(114));
   U1251 : AOI221_X1 port map( B1 => n29, B2 => regs(1138), C1 => n336, C2 => 
                           regs(2162), A => n1036, ZN => n1035);
   U1252 : INV_X1 port map( A => n1037, ZN => n1036);
   U1253 : AOI222_X1 port map( A1 => regs(114), A2 => n78, B1 => regs(1650), B2
                           => n196, C1 => regs(626), C2 => n271, ZN => n1037);
   U1254 : INV_X1 port map( A => n1038, ZN => curr_proc_regs(626));
   U1255 : AOI221_X1 port map( B1 => n30, B2 => regs(1650), C1 => n336, C2 => 
                           regs(114), A => n1039, ZN => n1038);
   U1256 : INV_X1 port map( A => n1040, ZN => n1039);
   U1257 : AOI222_X1 port map( A1 => regs(626), A2 => n78, B1 => regs(2162), B2
                           => n196, C1 => regs(1138), C2 => n271, ZN => n1040);
   U1258 : INV_X1 port map( A => n1041, ZN => curr_proc_regs(113));
   U1259 : AOI221_X1 port map( B1 => n30, B2 => regs(1137), C1 => n336, C2 => 
                           regs(2161), A => n1042, ZN => n1041);
   U1260 : INV_X1 port map( A => n1043, ZN => n1042);
   U1261 : AOI222_X1 port map( A1 => regs(113), A2 => n78, B1 => regs(1649), B2
                           => n196, C1 => regs(625), C2 => n271, ZN => n1043);
   U1262 : INV_X1 port map( A => n1044, ZN => curr_proc_regs(625));
   U1263 : AOI221_X1 port map( B1 => n30, B2 => regs(1649), C1 => n336, C2 => 
                           regs(113), A => n1045, ZN => n1044);
   U1264 : INV_X1 port map( A => n1046, ZN => n1045);
   U1265 : AOI222_X1 port map( A1 => regs(625), A2 => n78, B1 => regs(2161), B2
                           => n196, C1 => regs(1137), C2 => n271, ZN => n1046);
   U1266 : INV_X1 port map( A => n1047, ZN => curr_proc_regs(112));
   U1267 : AOI221_X1 port map( B1 => n30, B2 => regs(1136), C1 => n336, C2 => 
                           regs(2160), A => n1048, ZN => n1047);
   U1268 : INV_X1 port map( A => n1049, ZN => n1048);
   U1269 : AOI222_X1 port map( A1 => regs(112), A2 => n78, B1 => regs(1648), B2
                           => n196, C1 => regs(624), C2 => n271, ZN => n1049);
   U1270 : INV_X1 port map( A => n1050, ZN => curr_proc_regs(624));
   U1271 : AOI221_X1 port map( B1 => n30, B2 => regs(1648), C1 => n336, C2 => 
                           regs(112), A => n1051, ZN => n1050);
   U1272 : INV_X1 port map( A => n1052, ZN => n1051);
   U1273 : AOI222_X1 port map( A1 => regs(624), A2 => n78, B1 => regs(2160), B2
                           => n196, C1 => regs(1136), C2 => n271, ZN => n1052);
   U1274 : INV_X1 port map( A => n1053, ZN => curr_proc_regs(111));
   U1275 : AOI221_X1 port map( B1 => n30, B2 => regs(1135), C1 => n336, C2 => 
                           regs(2159), A => n1054, ZN => n1053);
   U1276 : INV_X1 port map( A => n1055, ZN => n1054);
   U1277 : AOI222_X1 port map( A1 => regs(111), A2 => n78, B1 => regs(1647), B2
                           => n196, C1 => regs(623), C2 => n271, ZN => n1055);
   U1278 : INV_X1 port map( A => n1056, ZN => curr_proc_regs(623));
   U1279 : AOI221_X1 port map( B1 => n30, B2 => regs(1647), C1 => n335, C2 => 
                           regs(111), A => n1057, ZN => n1056);
   U1280 : INV_X1 port map( A => n1058, ZN => n1057);
   U1281 : AOI222_X1 port map( A1 => regs(623), A2 => n78, B1 => regs(2159), B2
                           => n196, C1 => regs(1135), C2 => n271, ZN => n1058);
   U1282 : INV_X1 port map( A => n1059, ZN => curr_proc_regs(110));
   U1283 : AOI221_X1 port map( B1 => n30, B2 => regs(1134), C1 => n335, C2 => 
                           regs(2158), A => n1060, ZN => n1059);
   U1284 : INV_X1 port map( A => n1061, ZN => n1060);
   U1285 : AOI222_X1 port map( A1 => regs(110), A2 => n78, B1 => regs(1646), B2
                           => n196, C1 => regs(622), C2 => n271, ZN => n1061);
   U1286 : INV_X1 port map( A => n1062, ZN => curr_proc_regs(622));
   U1287 : AOI221_X1 port map( B1 => n30, B2 => regs(1646), C1 => n335, C2 => 
                           regs(110), A => n1063, ZN => n1062);
   U1288 : INV_X1 port map( A => n1064, ZN => n1063);
   U1289 : AOI222_X1 port map( A1 => regs(622), A2 => n78, B1 => regs(2158), B2
                           => n196, C1 => regs(1134), C2 => n271, ZN => n1064);
   U1290 : INV_X1 port map( A => n1065, ZN => curr_proc_regs(109));
   U1291 : AOI221_X1 port map( B1 => n30, B2 => regs(1133), C1 => n335, C2 => 
                           regs(2157), A => n1066, ZN => n1065);
   U1292 : INV_X1 port map( A => n1067, ZN => n1066);
   U1293 : AOI222_X1 port map( A1 => regs(109), A2 => n78, B1 => regs(1645), B2
                           => n195, C1 => regs(621), C2 => n270, ZN => n1067);
   U1294 : INV_X1 port map( A => n1068, ZN => curr_proc_regs(621));
   U1295 : AOI221_X1 port map( B1 => n30, B2 => regs(1645), C1 => n335, C2 => 
                           regs(109), A => n1069, ZN => n1068);
   U1296 : INV_X1 port map( A => n1070, ZN => n1069);
   U1297 : AOI222_X1 port map( A1 => regs(621), A2 => n79, B1 => regs(2157), B2
                           => n195, C1 => regs(1133), C2 => n270, ZN => n1070);
   U1298 : INV_X1 port map( A => n1071, ZN => curr_proc_regs(108));
   U1299 : AOI221_X1 port map( B1 => n30, B2 => regs(1132), C1 => n335, C2 => 
                           regs(2156), A => n1072, ZN => n1071);
   U1300 : INV_X1 port map( A => n1073, ZN => n1072);
   U1301 : AOI222_X1 port map( A1 => regs(108), A2 => n79, B1 => regs(1644), B2
                           => n195, C1 => regs(620), C2 => n270, ZN => n1073);
   U1302 : INV_X1 port map( A => n1074, ZN => curr_proc_regs(620));
   U1303 : AOI221_X1 port map( B1 => n31, B2 => regs(1644), C1 => n335, C2 => 
                           regs(108), A => n1075, ZN => n1074);
   U1304 : INV_X1 port map( A => n1076, ZN => n1075);
   U1305 : AOI222_X1 port map( A1 => regs(620), A2 => n79, B1 => regs(2156), B2
                           => n195, C1 => regs(1132), C2 => n270, ZN => n1076);
   U1306 : INV_X1 port map( A => n1077, ZN => curr_proc_regs(107));
   U1307 : AOI221_X1 port map( B1 => n31, B2 => regs(1131), C1 => n335, C2 => 
                           regs(2155), A => n1078, ZN => n1077);
   U1308 : INV_X1 port map( A => n1079, ZN => n1078);
   U1309 : AOI222_X1 port map( A1 => regs(107), A2 => n79, B1 => regs(1643), B2
                           => n195, C1 => regs(619), C2 => n270, ZN => n1079);
   U1310 : INV_X1 port map( A => n1080, ZN => curr_proc_regs(619));
   U1311 : AOI221_X1 port map( B1 => n31, B2 => regs(1643), C1 => n335, C2 => 
                           regs(107), A => n1081, ZN => n1080);
   U1312 : INV_X1 port map( A => n1082, ZN => n1081);
   U1313 : AOI222_X1 port map( A1 => regs(619), A2 => n79, B1 => regs(2155), B2
                           => n195, C1 => regs(1131), C2 => n270, ZN => n1082);
   U1314 : INV_X1 port map( A => n1083, ZN => curr_proc_regs(106));
   U1315 : AOI221_X1 port map( B1 => n31, B2 => regs(1130), C1 => n335, C2 => 
                           regs(2154), A => n1084, ZN => n1083);
   U1316 : INV_X1 port map( A => n1085, ZN => n1084);
   U1317 : AOI222_X1 port map( A1 => regs(106), A2 => n79, B1 => regs(1642), B2
                           => n195, C1 => regs(618), C2 => n270, ZN => n1085);
   U1318 : INV_X1 port map( A => n1086, ZN => curr_proc_regs(618));
   U1319 : AOI221_X1 port map( B1 => n31, B2 => regs(1642), C1 => n335, C2 => 
                           regs(106), A => n1087, ZN => n1086);
   U1320 : INV_X1 port map( A => n1088, ZN => n1087);
   U1321 : AOI222_X1 port map( A1 => regs(618), A2 => n79, B1 => regs(2154), B2
                           => n195, C1 => regs(1130), C2 => n270, ZN => n1088);
   U1322 : INV_X1 port map( A => n1089, ZN => curr_proc_regs(105));
   U1323 : AOI221_X1 port map( B1 => n31, B2 => regs(1129), C1 => n335, C2 => 
                           regs(2153), A => n1090, ZN => n1089);
   U1324 : INV_X1 port map( A => n1091, ZN => n1090);
   U1325 : AOI222_X1 port map( A1 => regs(105), A2 => n79, B1 => regs(1641), B2
                           => n195, C1 => regs(617), C2 => n270, ZN => n1091);
   U1326 : INV_X1 port map( A => n1092, ZN => curr_proc_regs(617));
   U1327 : AOI221_X1 port map( B1 => n31, B2 => regs(1641), C1 => n334, C2 => 
                           regs(105), A => n1093, ZN => n1092);
   U1328 : INV_X1 port map( A => n1094, ZN => n1093);
   U1329 : AOI222_X1 port map( A1 => regs(617), A2 => n79, B1 => regs(2153), B2
                           => n195, C1 => regs(1129), C2 => n270, ZN => n1094);
   U1330 : INV_X1 port map( A => n1095, ZN => curr_proc_regs(104));
   U1331 : AOI221_X1 port map( B1 => n31, B2 => regs(1128), C1 => n334, C2 => 
                           regs(2152), A => n1096, ZN => n1095);
   U1332 : INV_X1 port map( A => n1097, ZN => n1096);
   U1333 : AOI222_X1 port map( A1 => regs(104), A2 => n79, B1 => regs(1640), B2
                           => n195, C1 => regs(616), C2 => n270, ZN => n1097);
   U1334 : INV_X1 port map( A => n1098, ZN => curr_proc_regs(616));
   U1335 : AOI221_X1 port map( B1 => n31, B2 => regs(1640), C1 => n334, C2 => 
                           regs(104), A => n1099, ZN => n1098);
   U1336 : INV_X1 port map( A => n1100, ZN => n1099);
   U1337 : AOI222_X1 port map( A1 => regs(616), A2 => n79, B1 => regs(2152), B2
                           => n195, C1 => regs(1128), C2 => n270, ZN => n1100);
   U1338 : INV_X1 port map( A => n1101, ZN => curr_proc_regs(103));
   U1339 : AOI221_X1 port map( B1 => n31, B2 => regs(1127), C1 => n334, C2 => 
                           regs(2151), A => n1102, ZN => n1101);
   U1340 : INV_X1 port map( A => n1103, ZN => n1102);
   U1341 : AOI222_X1 port map( A1 => regs(103), A2 => n79, B1 => regs(1639), B2
                           => n194, C1 => regs(615), C2 => n269, ZN => n1103);
   U1342 : INV_X1 port map( A => n1104, ZN => curr_proc_regs(615));
   U1343 : AOI221_X1 port map( B1 => n31, B2 => regs(1639), C1 => n334, C2 => 
                           regs(103), A => n1105, ZN => n1104);
   U1344 : INV_X1 port map( A => n1106, ZN => n1105);
   U1345 : AOI222_X1 port map( A1 => regs(615), A2 => n80, B1 => regs(2151), B2
                           => n194, C1 => regs(1127), C2 => n269, ZN => n1106);
   U1346 : INV_X1 port map( A => n1107, ZN => curr_proc_regs(102));
   U1347 : AOI221_X1 port map( B1 => n31, B2 => regs(1126), C1 => n334, C2 => 
                           regs(2150), A => n1108, ZN => n1107);
   U1348 : INV_X1 port map( A => n1109, ZN => n1108);
   U1349 : AOI222_X1 port map( A1 => regs(102), A2 => n80, B1 => regs(1638), B2
                           => n194, C1 => regs(614), C2 => n269, ZN => n1109);
   U1350 : INV_X1 port map( A => n1110, ZN => curr_proc_regs(614));
   U1351 : AOI221_X1 port map( B1 => n32, B2 => regs(1638), C1 => n334, C2 => 
                           regs(102), A => n1111, ZN => n1110);
   U1352 : INV_X1 port map( A => n1112, ZN => n1111);
   U1353 : AOI222_X1 port map( A1 => regs(614), A2 => n80, B1 => regs(2150), B2
                           => n194, C1 => regs(1126), C2 => n269, ZN => n1112);
   U1354 : INV_X1 port map( A => n1113, ZN => curr_proc_regs(101));
   U1355 : AOI221_X1 port map( B1 => n32, B2 => regs(1125), C1 => n334, C2 => 
                           regs(2149), A => n1114, ZN => n1113);
   U1356 : INV_X1 port map( A => n1115, ZN => n1114);
   U1357 : AOI222_X1 port map( A1 => regs(101), A2 => n80, B1 => regs(1637), B2
                           => n194, C1 => regs(613), C2 => n269, ZN => n1115);
   U1358 : INV_X1 port map( A => n1116, ZN => curr_proc_regs(613));
   U1359 : AOI221_X1 port map( B1 => n32, B2 => regs(1637), C1 => n334, C2 => 
                           regs(101), A => n1117, ZN => n1116);
   U1360 : INV_X1 port map( A => n1118, ZN => n1117);
   U1361 : AOI222_X1 port map( A1 => regs(613), A2 => n80, B1 => regs(2149), B2
                           => n194, C1 => regs(1125), C2 => n269, ZN => n1118);
   U1362 : INV_X1 port map( A => n1119, ZN => curr_proc_regs(100));
   U1363 : AOI221_X1 port map( B1 => n32, B2 => regs(1124), C1 => n334, C2 => 
                           regs(2148), A => n1120, ZN => n1119);
   U1364 : INV_X1 port map( A => n1121, ZN => n1120);
   U1365 : AOI222_X1 port map( A1 => regs(100), A2 => n80, B1 => regs(1636), B2
                           => n194, C1 => regs(612), C2 => n269, ZN => n1121);
   U1366 : INV_X1 port map( A => n1122, ZN => curr_proc_regs(612));
   U1367 : AOI221_X1 port map( B1 => n32, B2 => regs(1636), C1 => n334, C2 => 
                           regs(100), A => n1123, ZN => n1122);
   U1368 : INV_X1 port map( A => n1124, ZN => n1123);
   U1369 : AOI222_X1 port map( A1 => regs(612), A2 => n80, B1 => regs(2148), B2
                           => n194, C1 => regs(1124), C2 => n269, ZN => n1124);
   U1370 : INV_X1 port map( A => n1125, ZN => curr_proc_regs(611));
   U1371 : AOI221_X1 port map( B1 => n32, B2 => regs(1635), C1 => n334, C2 => 
                           regs(99), A => n1126, ZN => n1125);
   U1372 : INV_X1 port map( A => n1127, ZN => n1126);
   U1373 : AOI222_X1 port map( A1 => regs(611), A2 => n80, B1 => regs(2147), B2
                           => n194, C1 => regs(1123), C2 => n269, ZN => n1127);
   U1374 : INV_X1 port map( A => n1128, ZN => curr_proc_regs(99));
   U1375 : AOI221_X1 port map( B1 => n32, B2 => regs(1123), C1 => n333, C2 => 
                           regs(2147), A => n1129, ZN => n1128);
   U1376 : INV_X1 port map( A => n1130, ZN => n1129);
   U1377 : AOI222_X1 port map( A1 => regs(99), A2 => n80, B1 => regs(1635), B2 
                           => n194, C1 => regs(611), C2 => n269, ZN => n1130);
   U1378 : INV_X1 port map( A => n1131, ZN => curr_proc_regs(610));
   U1379 : AOI221_X1 port map( B1 => n32, B2 => regs(1634), C1 => n333, C2 => 
                           regs(98), A => n1132, ZN => n1131);
   U1380 : INV_X1 port map( A => n1133, ZN => n1132);
   U1381 : AOI222_X1 port map( A1 => regs(610), A2 => n80, B1 => regs(2146), B2
                           => n194, C1 => regs(1122), C2 => n269, ZN => n1133);
   U1382 : INV_X1 port map( A => n1134, ZN => curr_proc_regs(98));
   U1383 : AOI221_X1 port map( B1 => n32, B2 => regs(1122), C1 => n333, C2 => 
                           regs(2146), A => n1135, ZN => n1134);
   U1384 : INV_X1 port map( A => n1136, ZN => n1135);
   U1385 : AOI222_X1 port map( A1 => regs(98), A2 => n80, B1 => regs(1634), B2 
                           => n194, C1 => regs(610), C2 => n269, ZN => n1136);
   U1386 : INV_X1 port map( A => n1137, ZN => curr_proc_regs(609));
   U1387 : AOI221_X1 port map( B1 => n32, B2 => regs(1633), C1 => n333, C2 => 
                           regs(97), A => n1138, ZN => n1137);
   U1388 : INV_X1 port map( A => n1139, ZN => n1138);
   U1389 : AOI222_X1 port map( A1 => regs(609), A2 => n80, B1 => regs(2145), B2
                           => n193, C1 => regs(1121), C2 => n268, ZN => n1139);
   U1390 : INV_X1 port map( A => n1140, ZN => curr_proc_regs(97));
   U1391 : AOI221_X1 port map( B1 => n32, B2 => regs(1121), C1 => n333, C2 => 
                           regs(2145), A => n1141, ZN => n1140);
   U1392 : INV_X1 port map( A => n1142, ZN => n1141);
   U1393 : AOI222_X1 port map( A1 => regs(97), A2 => n81, B1 => regs(1633), B2 
                           => n193, C1 => regs(609), C2 => n268, ZN => n1142);
   U1394 : INV_X1 port map( A => n1143, ZN => curr_proc_regs(608));
   U1395 : AOI221_X1 port map( B1 => n32, B2 => regs(1632), C1 => n333, C2 => 
                           regs(96), A => n1144, ZN => n1143);
   U1396 : INV_X1 port map( A => n1145, ZN => n1144);
   U1397 : AOI222_X1 port map( A1 => regs(608), A2 => n81, B1 => regs(2144), B2
                           => n193, C1 => regs(1120), C2 => n268, ZN => n1145);
   U1398 : INV_X1 port map( A => n1146, ZN => curr_proc_regs(96));
   U1399 : AOI221_X1 port map( B1 => n33, B2 => regs(1120), C1 => n333, C2 => 
                           regs(2144), A => n1147, ZN => n1146);
   U1400 : INV_X1 port map( A => n1148, ZN => n1147);
   U1401 : AOI222_X1 port map( A1 => regs(96), A2 => n81, B1 => regs(1632), B2 
                           => n193, C1 => regs(608), C2 => n268, ZN => n1148);
   U1402 : INV_X1 port map( A => n1149, ZN => curr_proc_regs(159));
   U1403 : AOI221_X1 port map( B1 => n59, B2 => regs(1183), C1 => n333, C2 => 
                           regs(2207), A => n1150, ZN => n1149);
   U1404 : INV_X1 port map( A => n1151, ZN => n1150);
   U1405 : AOI222_X1 port map( A1 => regs(159), A2 => n81, B1 => regs(1695), B2
                           => n193, C1 => regs(671), C2 => n268, ZN => n1151);
   U1406 : INV_X1 port map( A => n1152, ZN => curr_proc_regs(671));
   U1407 : AOI221_X1 port map( B1 => n54, B2 => regs(1695), C1 => n333, C2 => 
                           regs(159), A => n1153, ZN => n1152);
   U1408 : INV_X1 port map( A => n1154, ZN => n1153);
   U1409 : AOI222_X1 port map( A1 => regs(671), A2 => n81, B1 => regs(2207), B2
                           => n193, C1 => regs(1183), C2 => n268, ZN => n1154);
   U1410 : INV_X1 port map( A => n1155, ZN => curr_proc_regs(158));
   U1411 : AOI221_X1 port map( B1 => n54, B2 => regs(1182), C1 => n333, C2 => 
                           regs(2206), A => n1156, ZN => n1155);
   U1412 : INV_X1 port map( A => n1157, ZN => n1156);
   U1413 : AOI222_X1 port map( A1 => regs(158), A2 => n81, B1 => regs(1694), B2
                           => n193, C1 => regs(670), C2 => n268, ZN => n1157);
   U1414 : INV_X1 port map( A => n1158, ZN => curr_proc_regs(670));
   U1415 : AOI221_X1 port map( B1 => n54, B2 => regs(1694), C1 => n311, C2 => 
                           regs(158), A => n1159, ZN => n1158);
   U1416 : INV_X1 port map( A => n1160, ZN => n1159);
   U1417 : AOI222_X1 port map( A1 => regs(670), A2 => n81, B1 => regs(2206), B2
                           => n193, C1 => regs(1182), C2 => n268, ZN => n1160);
   U1418 : INV_X1 port map( A => n1161, ZN => curr_proc_regs(157));
   U1419 : AOI221_X1 port map( B1 => n54, B2 => regs(1181), C1 => n311, C2 => 
                           regs(2205), A => n1162, ZN => n1161);
   U1420 : INV_X1 port map( A => n1163, ZN => n1162);
   U1421 : AOI222_X1 port map( A1 => regs(157), A2 => n81, B1 => regs(1693), B2
                           => n193, C1 => regs(669), C2 => n268, ZN => n1163);
   U1422 : INV_X1 port map( A => n1164, ZN => curr_proc_regs(669));
   U1423 : AOI221_X1 port map( B1 => n54, B2 => regs(1693), C1 => n311, C2 => 
                           regs(157), A => n1165, ZN => n1164);
   U1424 : INV_X1 port map( A => n1166, ZN => n1165);
   U1425 : AOI222_X1 port map( A1 => regs(669), A2 => n81, B1 => regs(2205), B2
                           => n193, C1 => regs(1181), C2 => n268, ZN => n1166);
   U1426 : INV_X1 port map( A => n1167, ZN => curr_proc_regs(156));
   U1427 : AOI221_X1 port map( B1 => n54, B2 => regs(1180), C1 => n311, C2 => 
                           regs(2204), A => n1168, ZN => n1167);
   U1428 : INV_X1 port map( A => n1169, ZN => n1168);
   U1429 : AOI222_X1 port map( A1 => regs(156), A2 => n81, B1 => regs(1692), B2
                           => n193, C1 => regs(668), C2 => n268, ZN => n1169);
   U1430 : INV_X1 port map( A => n1170, ZN => curr_proc_regs(668));
   U1431 : AOI221_X1 port map( B1 => n54, B2 => regs(1692), C1 => n311, C2 => 
                           regs(156), A => n1171, ZN => n1170);
   U1432 : INV_X1 port map( A => n1172, ZN => n1171);
   U1433 : AOI222_X1 port map( A1 => regs(668), A2 => n81, B1 => regs(2204), B2
                           => n193, C1 => regs(1180), C2 => n268, ZN => n1172);
   U1434 : INV_X1 port map( A => n1173, ZN => curr_proc_regs(155));
   U1435 : AOI221_X1 port map( B1 => n55, B2 => regs(1179), C1 => n311, C2 => 
                           regs(2203), A => n1174, ZN => n1173);
   U1436 : INV_X1 port map( A => n1175, ZN => n1174);
   U1437 : AOI222_X1 port map( A1 => regs(155), A2 => n81, B1 => regs(1691), B2
                           => n192, C1 => regs(667), C2 => n267, ZN => n1175);
   U1438 : INV_X1 port map( A => n1176, ZN => curr_proc_regs(667));
   U1439 : AOI221_X1 port map( B1 => n55, B2 => regs(1691), C1 => n311, C2 => 
                           regs(155), A => n1177, ZN => n1176);
   U1440 : INV_X1 port map( A => n1178, ZN => n1177);
   U1441 : AOI222_X1 port map( A1 => regs(667), A2 => n82, B1 => regs(2203), B2
                           => n192, C1 => regs(1179), C2 => n267, ZN => n1178);
   U1442 : INV_X1 port map( A => n1179, ZN => curr_proc_regs(154));
   U1443 : AOI221_X1 port map( B1 => n55, B2 => regs(1178), C1 => n311, C2 => 
                           regs(2202), A => n1180, ZN => n1179);
   U1444 : INV_X1 port map( A => n1181, ZN => n1180);
   U1445 : AOI222_X1 port map( A1 => regs(154), A2 => n82, B1 => regs(1690), B2
                           => n192, C1 => regs(666), C2 => n267, ZN => n1181);
   U1446 : INV_X1 port map( A => n1182, ZN => curr_proc_regs(666));
   U1447 : AOI221_X1 port map( B1 => n55, B2 => regs(1690), C1 => n311, C2 => 
                           regs(154), A => n1183, ZN => n1182);
   U1448 : INV_X1 port map( A => n1184, ZN => n1183);
   U1449 : AOI222_X1 port map( A1 => regs(666), A2 => n82, B1 => regs(2202), B2
                           => n192, C1 => regs(1178), C2 => n267, ZN => n1184);
   U1450 : INV_X1 port map( A => n1185, ZN => curr_proc_regs(153));
   U1451 : AOI221_X1 port map( B1 => n55, B2 => regs(1177), C1 => n311, C2 => 
                           regs(2201), A => n1186, ZN => n1185);
   U1452 : INV_X1 port map( A => n1187, ZN => n1186);
   U1453 : AOI222_X1 port map( A1 => regs(153), A2 => n82, B1 => regs(1689), B2
                           => n192, C1 => regs(665), C2 => n267, ZN => n1187);
   U1454 : INV_X1 port map( A => n1188, ZN => curr_proc_regs(665));
   U1455 : AOI221_X1 port map( B1 => n55, B2 => regs(1689), C1 => n311, C2 => 
                           regs(153), A => n1189, ZN => n1188);
   U1456 : INV_X1 port map( A => n1190, ZN => n1189);
   U1457 : AOI222_X1 port map( A1 => regs(665), A2 => n82, B1 => regs(2201), B2
                           => n192, C1 => regs(1177), C2 => n267, ZN => n1190);
   U1458 : INV_X1 port map( A => n1191, ZN => curr_proc_regs(152));
   U1459 : AOI221_X1 port map( B1 => n55, B2 => regs(1176), C1 => n310, C2 => 
                           regs(2200), A => n1192, ZN => n1191);
   U1460 : INV_X1 port map( A => n1193, ZN => n1192);
   U1461 : AOI222_X1 port map( A1 => regs(152), A2 => n82, B1 => regs(1688), B2
                           => n192, C1 => regs(664), C2 => n267, ZN => n1193);
   U1462 : INV_X1 port map( A => n1194, ZN => curr_proc_regs(664));
   U1463 : AOI221_X1 port map( B1 => n55, B2 => regs(1688), C1 => n310, C2 => 
                           regs(152), A => n1195, ZN => n1194);
   U1464 : INV_X1 port map( A => n1196, ZN => n1195);
   U1465 : AOI222_X1 port map( A1 => regs(664), A2 => n82, B1 => regs(2200), B2
                           => n192, C1 => regs(1176), C2 => n267, ZN => n1196);
   U1466 : INV_X1 port map( A => n1197, ZN => curr_proc_regs(151));
   U1467 : AOI221_X1 port map( B1 => n55, B2 => regs(1175), C1 => n310, C2 => 
                           regs(2199), A => n1198, ZN => n1197);
   U1468 : INV_X1 port map( A => n1199, ZN => n1198);
   U1469 : AOI222_X1 port map( A1 => regs(151), A2 => n82, B1 => regs(1687), B2
                           => n192, C1 => regs(663), C2 => n267, ZN => n1199);
   U1470 : INV_X1 port map( A => n1200, ZN => curr_proc_regs(663));
   U1471 : AOI221_X1 port map( B1 => n55, B2 => regs(1687), C1 => n310, C2 => 
                           regs(151), A => n1201, ZN => n1200);
   U1472 : INV_X1 port map( A => n1202, ZN => n1201);
   U1473 : AOI222_X1 port map( A1 => regs(663), A2 => n82, B1 => regs(2199), B2
                           => n192, C1 => regs(1175), C2 => n267, ZN => n1202);
   U1474 : INV_X1 port map( A => n1203, ZN => curr_proc_regs(150));
   U1475 : AOI221_X1 port map( B1 => n55, B2 => regs(1174), C1 => n310, C2 => 
                           regs(2198), A => n1204, ZN => n1203);
   U1476 : INV_X1 port map( A => n1205, ZN => n1204);
   U1477 : AOI222_X1 port map( A1 => regs(150), A2 => n82, B1 => regs(1686), B2
                           => n192, C1 => regs(662), C2 => n267, ZN => n1205);
   U1478 : INV_X1 port map( A => n1206, ZN => curr_proc_regs(662));
   U1479 : AOI221_X1 port map( B1 => n55, B2 => regs(1686), C1 => n310, C2 => 
                           regs(150), A => n1207, ZN => n1206);
   U1480 : INV_X1 port map( A => n1208, ZN => n1207);
   U1481 : AOI222_X1 port map( A1 => regs(662), A2 => n82, B1 => regs(2198), B2
                           => n192, C1 => regs(1174), C2 => n267, ZN => n1208);
   U1482 : INV_X1 port map( A => n1209, ZN => curr_proc_regs(149));
   U1483 : AOI221_X1 port map( B1 => n56, B2 => regs(1173), C1 => n310, C2 => 
                           regs(2197), A => n1210, ZN => n1209);
   U1484 : INV_X1 port map( A => n1211, ZN => n1210);
   U1485 : AOI222_X1 port map( A1 => regs(149), A2 => n82, B1 => regs(1685), B2
                           => n191, C1 => regs(661), C2 => n266, ZN => n1211);
   U1486 : INV_X1 port map( A => n1212, ZN => curr_proc_regs(661));
   U1487 : AOI221_X1 port map( B1 => n56, B2 => regs(1685), C1 => n310, C2 => 
                           regs(149), A => n1213, ZN => n1212);
   U1488 : INV_X1 port map( A => n1214, ZN => n1213);
   U1489 : AOI222_X1 port map( A1 => regs(661), A2 => n83, B1 => regs(2197), B2
                           => n191, C1 => regs(1173), C2 => n266, ZN => n1214);
   U1490 : INV_X1 port map( A => n1215, ZN => curr_proc_regs(148));
   U1491 : AOI221_X1 port map( B1 => n56, B2 => regs(1172), C1 => n310, C2 => 
                           regs(2196), A => n1216, ZN => n1215);
   U1492 : INV_X1 port map( A => n1217, ZN => n1216);
   U1493 : AOI222_X1 port map( A1 => regs(148), A2 => n83, B1 => regs(1684), B2
                           => n191, C1 => regs(660), C2 => n266, ZN => n1217);
   U1494 : INV_X1 port map( A => n1218, ZN => curr_proc_regs(660));
   U1495 : AOI221_X1 port map( B1 => n56, B2 => regs(1684), C1 => n310, C2 => 
                           regs(148), A => n1219, ZN => n1218);
   U1496 : INV_X1 port map( A => n1220, ZN => n1219);
   U1497 : AOI222_X1 port map( A1 => regs(660), A2 => n83, B1 => regs(2196), B2
                           => n191, C1 => regs(1172), C2 => n266, ZN => n1220);
   U1498 : INV_X1 port map( A => n1221, ZN => curr_proc_regs(147));
   U1499 : AOI221_X1 port map( B1 => n56, B2 => regs(1171), C1 => n310, C2 => 
                           regs(2195), A => n1222, ZN => n1221);
   U1500 : INV_X1 port map( A => n1223, ZN => n1222);
   U1501 : AOI222_X1 port map( A1 => regs(147), A2 => n83, B1 => regs(1683), B2
                           => n191, C1 => regs(659), C2 => n266, ZN => n1223);
   U1502 : INV_X1 port map( A => n1224, ZN => curr_proc_regs(659));
   U1503 : AOI221_X1 port map( B1 => n56, B2 => regs(1683), C1 => n310, C2 => 
                           regs(147), A => n1225, ZN => n1224);
   U1504 : INV_X1 port map( A => n1226, ZN => n1225);
   U1505 : AOI222_X1 port map( A1 => regs(659), A2 => n83, B1 => regs(2195), B2
                           => n191, C1 => regs(1171), C2 => n266, ZN => n1226);
   U1506 : INV_X1 port map( A => n1227, ZN => curr_proc_regs(146));
   U1507 : AOI221_X1 port map( B1 => n56, B2 => regs(1170), C1 => n309, C2 => 
                           regs(2194), A => n1228, ZN => n1227);
   U1508 : INV_X1 port map( A => n1229, ZN => n1228);
   U1509 : AOI222_X1 port map( A1 => regs(146), A2 => n83, B1 => regs(1682), B2
                           => n191, C1 => regs(658), C2 => n266, ZN => n1229);
   U1510 : INV_X1 port map( A => n1230, ZN => curr_proc_regs(658));
   U1511 : AOI221_X1 port map( B1 => n56, B2 => regs(1682), C1 => n309, C2 => 
                           regs(146), A => n1231, ZN => n1230);
   U1512 : INV_X1 port map( A => n1232, ZN => n1231);
   U1513 : AOI222_X1 port map( A1 => regs(658), A2 => n83, B1 => regs(2194), B2
                           => n191, C1 => regs(1170), C2 => n266, ZN => n1232);
   U1514 : INV_X1 port map( A => n1233, ZN => curr_proc_regs(145));
   U1515 : AOI221_X1 port map( B1 => n56, B2 => regs(1169), C1 => n309, C2 => 
                           regs(2193), A => n1234, ZN => n1233);
   U1516 : INV_X1 port map( A => n1235, ZN => n1234);
   U1517 : AOI222_X1 port map( A1 => regs(145), A2 => n83, B1 => regs(1681), B2
                           => n191, C1 => regs(657), C2 => n266, ZN => n1235);
   U1518 : INV_X1 port map( A => n1236, ZN => curr_proc_regs(657));
   U1519 : AOI221_X1 port map( B1 => n56, B2 => regs(1681), C1 => n309, C2 => 
                           regs(145), A => n1237, ZN => n1236);
   U1520 : INV_X1 port map( A => n1238, ZN => n1237);
   U1521 : AOI222_X1 port map( A1 => regs(657), A2 => n83, B1 => regs(2193), B2
                           => n191, C1 => regs(1169), C2 => n266, ZN => n1238);
   U1522 : INV_X1 port map( A => n1239, ZN => curr_proc_regs(144));
   U1523 : AOI221_X1 port map( B1 => n56, B2 => regs(1168), C1 => n309, C2 => 
                           regs(2192), A => n1240, ZN => n1239);
   U1524 : INV_X1 port map( A => n1241, ZN => n1240);
   U1525 : AOI222_X1 port map( A1 => regs(144), A2 => n83, B1 => regs(1680), B2
                           => n191, C1 => regs(656), C2 => n266, ZN => n1241);
   U1526 : INV_X1 port map( A => n1242, ZN => curr_proc_regs(656));
   U1527 : AOI221_X1 port map( B1 => n56, B2 => regs(1680), C1 => n309, C2 => 
                           regs(144), A => n1243, ZN => n1242);
   U1528 : INV_X1 port map( A => n1244, ZN => n1243);
   U1529 : AOI222_X1 port map( A1 => regs(656), A2 => n83, B1 => regs(2192), B2
                           => n191, C1 => regs(1168), C2 => n266, ZN => n1244);
   U1530 : INV_X1 port map( A => n1245, ZN => curr_proc_regs(143));
   U1531 : AOI221_X1 port map( B1 => n57, B2 => regs(1167), C1 => n309, C2 => 
                           regs(2191), A => n1246, ZN => n1245);
   U1532 : INV_X1 port map( A => n1247, ZN => n1246);
   U1533 : AOI222_X1 port map( A1 => regs(143), A2 => n84, B1 => regs(1679), B2
                           => n190, C1 => regs(655), C2 => n265, ZN => n1247);
   U1534 : INV_X1 port map( A => n1248, ZN => curr_proc_regs(655));
   U1535 : AOI221_X1 port map( B1 => n57, B2 => regs(1679), C1 => n309, C2 => 
                           regs(143), A => n1249, ZN => n1248);
   U1536 : INV_X1 port map( A => n1250, ZN => n1249);
   U1537 : AOI222_X1 port map( A1 => regs(655), A2 => n84, B1 => regs(2191), B2
                           => n190, C1 => regs(1167), C2 => n265, ZN => n1250);
   U1538 : INV_X1 port map( A => n1251, ZN => curr_proc_regs(142));
   U1539 : AOI221_X1 port map( B1 => n57, B2 => regs(1166), C1 => n309, C2 => 
                           regs(2190), A => n1252, ZN => n1251);
   U1540 : INV_X1 port map( A => n1253, ZN => n1252);
   U1541 : AOI222_X1 port map( A1 => regs(142), A2 => n84, B1 => regs(1678), B2
                           => n190, C1 => regs(654), C2 => n265, ZN => n1253);
   U1542 : INV_X1 port map( A => n1254, ZN => curr_proc_regs(654));
   U1543 : AOI221_X1 port map( B1 => n57, B2 => regs(1678), C1 => n309, C2 => 
                           regs(142), A => n1255, ZN => n1254);
   U1544 : INV_X1 port map( A => n1256, ZN => n1255);
   U1545 : AOI222_X1 port map( A1 => regs(654), A2 => n84, B1 => regs(2190), B2
                           => n190, C1 => regs(1166), C2 => n265, ZN => n1256);
   U1546 : INV_X1 port map( A => n1257, ZN => curr_proc_regs(141));
   U1547 : AOI221_X1 port map( B1 => n57, B2 => regs(1165), C1 => n309, C2 => 
                           regs(2189), A => n1258, ZN => n1257);
   U1548 : INV_X1 port map( A => n1259, ZN => n1258);
   U1549 : AOI222_X1 port map( A1 => regs(141), A2 => n84, B1 => regs(1677), B2
                           => n190, C1 => regs(653), C2 => n265, ZN => n1259);
   U1550 : INV_X1 port map( A => n1260, ZN => curr_proc_regs(653));
   U1551 : AOI221_X1 port map( B1 => n57, B2 => regs(1677), C1 => n309, C2 => 
                           regs(141), A => n1261, ZN => n1260);
   U1552 : INV_X1 port map( A => n1262, ZN => n1261);
   U1553 : AOI222_X1 port map( A1 => regs(653), A2 => n84, B1 => regs(2189), B2
                           => n190, C1 => regs(1165), C2 => n265, ZN => n1262);
   U1554 : INV_X1 port map( A => n1263, ZN => curr_proc_regs(140));
   U1555 : AOI221_X1 port map( B1 => n57, B2 => regs(1164), C1 => n308, C2 => 
                           regs(2188), A => n1264, ZN => n1263);
   U1556 : INV_X1 port map( A => n1265, ZN => n1264);
   U1557 : AOI222_X1 port map( A1 => regs(140), A2 => n84, B1 => regs(1676), B2
                           => n190, C1 => regs(652), C2 => n265, ZN => n1265);
   U1558 : INV_X1 port map( A => n1266, ZN => curr_proc_regs(652));
   U1559 : AOI221_X1 port map( B1 => n57, B2 => regs(1676), C1 => n308, C2 => 
                           regs(140), A => n1267, ZN => n1266);
   U1560 : INV_X1 port map( A => n1268, ZN => n1267);
   U1561 : AOI222_X1 port map( A1 => regs(652), A2 => n84, B1 => regs(2188), B2
                           => n190, C1 => regs(1164), C2 => n265, ZN => n1268);
   U1562 : INV_X1 port map( A => n1269, ZN => curr_proc_regs(139));
   U1563 : AOI221_X1 port map( B1 => n57, B2 => regs(1163), C1 => n308, C2 => 
                           regs(2187), A => n1270, ZN => n1269);
   U1564 : INV_X1 port map( A => n1271, ZN => n1270);
   U1565 : AOI222_X1 port map( A1 => regs(139), A2 => n84, B1 => regs(1675), B2
                           => n190, C1 => regs(651), C2 => n265, ZN => n1271);
   U1566 : INV_X1 port map( A => n1272, ZN => curr_proc_regs(651));
   U1567 : AOI221_X1 port map( B1 => n57, B2 => regs(1675), C1 => n308, C2 => 
                           regs(139), A => n1273, ZN => n1272);
   U1568 : INV_X1 port map( A => n1274, ZN => n1273);
   U1569 : AOI222_X1 port map( A1 => regs(651), A2 => n84, B1 => regs(2187), B2
                           => n190, C1 => regs(1163), C2 => n265, ZN => n1274);
   U1570 : INV_X1 port map( A => n1275, ZN => curr_proc_regs(138));
   U1571 : AOI221_X1 port map( B1 => n57, B2 => regs(1162), C1 => n308, C2 => 
                           regs(2186), A => n1276, ZN => n1275);
   U1572 : INV_X1 port map( A => n1277, ZN => n1276);
   U1573 : AOI222_X1 port map( A1 => regs(138), A2 => n84, B1 => regs(1674), B2
                           => n190, C1 => regs(650), C2 => n265, ZN => n1277);
   U1574 : INV_X1 port map( A => n1278, ZN => curr_proc_regs(650));
   U1575 : AOI221_X1 port map( B1 => n57, B2 => regs(1674), C1 => n308, C2 => 
                           regs(138), A => n1279, ZN => n1278);
   U1576 : INV_X1 port map( A => n1280, ZN => n1279);
   U1577 : AOI222_X1 port map( A1 => regs(650), A2 => n84, B1 => regs(2186), B2
                           => n190, C1 => regs(1162), C2 => n265, ZN => n1280);
   U1578 : INV_X1 port map( A => n1281, ZN => curr_proc_regs(137));
   U1579 : AOI221_X1 port map( B1 => n58, B2 => regs(1161), C1 => n308, C2 => 
                           regs(2185), A => n1282, ZN => n1281);
   U1580 : INV_X1 port map( A => n1283, ZN => n1282);
   U1581 : AOI222_X1 port map( A1 => regs(137), A2 => n85, B1 => regs(1673), B2
                           => n189, C1 => regs(649), C2 => n264, ZN => n1283);
   U1582 : INV_X1 port map( A => n1284, ZN => curr_proc_regs(649));
   U1583 : AOI221_X1 port map( B1 => n58, B2 => regs(1673), C1 => n308, C2 => 
                           regs(137), A => n1285, ZN => n1284);
   U1584 : INV_X1 port map( A => n1286, ZN => n1285);
   U1585 : AOI222_X1 port map( A1 => regs(649), A2 => n85, B1 => regs(2185), B2
                           => n189, C1 => regs(1161), C2 => n264, ZN => n1286);
   U1586 : INV_X1 port map( A => n1287, ZN => curr_proc_regs(136));
   U1587 : AOI221_X1 port map( B1 => n58, B2 => regs(1160), C1 => n308, C2 => 
                           regs(2184), A => n1288, ZN => n1287);
   U1588 : INV_X1 port map( A => n1289, ZN => n1288);
   U1589 : AOI222_X1 port map( A1 => regs(136), A2 => n85, B1 => regs(1672), B2
                           => n189, C1 => regs(648), C2 => n264, ZN => n1289);
   U1590 : INV_X1 port map( A => n1290, ZN => curr_proc_regs(648));
   U1591 : AOI221_X1 port map( B1 => n58, B2 => regs(1672), C1 => n308, C2 => 
                           regs(136), A => n1291, ZN => n1290);
   U1592 : INV_X1 port map( A => n1292, ZN => n1291);
   U1593 : AOI222_X1 port map( A1 => regs(648), A2 => n85, B1 => regs(2184), B2
                           => n189, C1 => regs(1160), C2 => n264, ZN => n1292);
   U1594 : INV_X1 port map( A => n1293, ZN => curr_proc_regs(135));
   U1595 : AOI221_X1 port map( B1 => n58, B2 => regs(1159), C1 => n308, C2 => 
                           regs(2183), A => n1294, ZN => n1293);
   U1596 : INV_X1 port map( A => n1295, ZN => n1294);
   U1597 : AOI222_X1 port map( A1 => regs(135), A2 => n85, B1 => regs(1671), B2
                           => n189, C1 => regs(647), C2 => n264, ZN => n1295);
   U1598 : INV_X1 port map( A => n1296, ZN => curr_proc_regs(647));
   U1599 : AOI221_X1 port map( B1 => n58, B2 => regs(1671), C1 => n308, C2 => 
                           regs(135), A => n1297, ZN => n1296);
   U1600 : INV_X1 port map( A => n1298, ZN => n1297);
   U1601 : AOI222_X1 port map( A1 => regs(647), A2 => n85, B1 => regs(2183), B2
                           => n189, C1 => regs(1159), C2 => n264, ZN => n1298);
   U1602 : INV_X1 port map( A => n1299, ZN => curr_proc_regs(134));
   U1603 : AOI221_X1 port map( B1 => n58, B2 => regs(1158), C1 => n307, C2 => 
                           regs(2182), A => n1300, ZN => n1299);
   U1604 : INV_X1 port map( A => n1301, ZN => n1300);
   U1605 : AOI222_X1 port map( A1 => regs(134), A2 => n85, B1 => regs(1670), B2
                           => n189, C1 => regs(646), C2 => n264, ZN => n1301);
   U1606 : INV_X1 port map( A => n1302, ZN => curr_proc_regs(646));
   U1607 : AOI221_X1 port map( B1 => n58, B2 => regs(1670), C1 => n307, C2 => 
                           regs(134), A => n1303, ZN => n1302);
   U1608 : INV_X1 port map( A => n1304, ZN => n1303);
   U1609 : AOI222_X1 port map( A1 => regs(646), A2 => n85, B1 => regs(2182), B2
                           => n189, C1 => regs(1158), C2 => n264, ZN => n1304);
   U1610 : INV_X1 port map( A => n1305, ZN => curr_proc_regs(133));
   U1611 : AOI221_X1 port map( B1 => n58, B2 => regs(1157), C1 => n307, C2 => 
                           regs(2181), A => n1306, ZN => n1305);
   U1612 : INV_X1 port map( A => n1307, ZN => n1306);
   U1613 : AOI222_X1 port map( A1 => regs(133), A2 => n85, B1 => regs(1669), B2
                           => n189, C1 => regs(645), C2 => n264, ZN => n1307);
   U1614 : INV_X1 port map( A => n1308, ZN => curr_proc_regs(645));
   U1615 : AOI221_X1 port map( B1 => n58, B2 => regs(1669), C1 => n307, C2 => 
                           regs(133), A => n1309, ZN => n1308);
   U1616 : INV_X1 port map( A => n1310, ZN => n1309);
   U1617 : AOI222_X1 port map( A1 => regs(645), A2 => n85, B1 => regs(2181), B2
                           => n189, C1 => regs(1157), C2 => n264, ZN => n1310);
   U1618 : INV_X1 port map( A => n1311, ZN => curr_proc_regs(132));
   U1619 : AOI221_X1 port map( B1 => n58, B2 => regs(1156), C1 => n307, C2 => 
                           regs(2180), A => n1312, ZN => n1311);
   U1620 : INV_X1 port map( A => n1313, ZN => n1312);
   U1621 : AOI222_X1 port map( A1 => regs(132), A2 => n85, B1 => regs(1668), B2
                           => n189, C1 => regs(644), C2 => n264, ZN => n1313);
   U1622 : INV_X1 port map( A => n1314, ZN => curr_proc_regs(644));
   U1623 : AOI221_X1 port map( B1 => n58, B2 => regs(1668), C1 => n307, C2 => 
                           regs(132), A => n1315, ZN => n1314);
   U1624 : INV_X1 port map( A => n1316, ZN => n1315);
   U1625 : AOI222_X1 port map( A1 => regs(644), A2 => n85, B1 => regs(2180), B2
                           => n189, C1 => regs(1156), C2 => n264, ZN => n1316);
   U1626 : INV_X1 port map( A => n1317, ZN => curr_proc_regs(131));
   U1627 : AOI221_X1 port map( B1 => n59, B2 => regs(1155), C1 => n307, C2 => 
                           regs(2179), A => n1318, ZN => n1317);
   U1628 : INV_X1 port map( A => n1319, ZN => n1318);
   U1629 : AOI222_X1 port map( A1 => regs(131), A2 => n86, B1 => regs(1667), B2
                           => n188, C1 => regs(643), C2 => n263, ZN => n1319);
   U1630 : INV_X1 port map( A => n1320, ZN => curr_proc_regs(643));
   U1631 : AOI221_X1 port map( B1 => n59, B2 => regs(1667), C1 => n307, C2 => 
                           regs(131), A => n1321, ZN => n1320);
   U1632 : INV_X1 port map( A => n1322, ZN => n1321);
   U1633 : AOI222_X1 port map( A1 => regs(643), A2 => n86, B1 => regs(2179), B2
                           => n188, C1 => regs(1155), C2 => n263, ZN => n1322);
   U1634 : INV_X1 port map( A => n1323, ZN => curr_proc_regs(130));
   U1635 : AOI221_X1 port map( B1 => n59, B2 => regs(1154), C1 => n307, C2 => 
                           regs(2178), A => n1324, ZN => n1323);
   U1636 : INV_X1 port map( A => n1325, ZN => n1324);
   U1637 : AOI222_X1 port map( A1 => regs(130), A2 => n86, B1 => regs(1666), B2
                           => n188, C1 => regs(642), C2 => n263, ZN => n1325);
   U1638 : INV_X1 port map( A => n1326, ZN => curr_proc_regs(642));
   U1639 : AOI221_X1 port map( B1 => n59, B2 => regs(1666), C1 => n307, C2 => 
                           regs(130), A => n1327, ZN => n1326);
   U1640 : INV_X1 port map( A => n1328, ZN => n1327);
   U1641 : AOI222_X1 port map( A1 => regs(642), A2 => n86, B1 => regs(2178), B2
                           => n188, C1 => regs(1154), C2 => n263, ZN => n1328);
   U1642 : INV_X1 port map( A => n1329, ZN => curr_proc_regs(129));
   U1643 : AOI221_X1 port map( B1 => n59, B2 => regs(1153), C1 => n307, C2 => 
                           regs(2177), A => n1330, ZN => n1329);
   U1644 : INV_X1 port map( A => n1331, ZN => n1330);
   U1645 : AOI222_X1 port map( A1 => regs(129), A2 => n86, B1 => regs(1665), B2
                           => n188, C1 => regs(641), C2 => n263, ZN => n1331);
   U1646 : INV_X1 port map( A => n1332, ZN => curr_proc_regs(641));
   U1647 : AOI221_X1 port map( B1 => n59, B2 => regs(1665), C1 => n307, C2 => 
                           regs(129), A => n1333, ZN => n1332);
   U1648 : INV_X1 port map( A => n1334, ZN => n1333);
   U1649 : AOI222_X1 port map( A1 => regs(641), A2 => n86, B1 => regs(2177), B2
                           => n188, C1 => regs(1153), C2 => n263, ZN => n1334);
   U1650 : INV_X1 port map( A => n1335, ZN => curr_proc_regs(128));
   U1651 : AOI221_X1 port map( B1 => n59, B2 => regs(1152), C1 => n306, C2 => 
                           regs(2176), A => n1336, ZN => n1335);
   U1652 : INV_X1 port map( A => n1337, ZN => n1336);
   U1653 : AOI222_X1 port map( A1 => regs(128), A2 => n86, B1 => regs(1664), B2
                           => n188, C1 => regs(640), C2 => n263, ZN => n1337);
   U1654 : INV_X1 port map( A => n1338, ZN => curr_proc_regs(640));
   U1655 : AOI221_X1 port map( B1 => n59, B2 => regs(1664), C1 => n306, C2 => 
                           regs(128), A => n1339, ZN => n1338);
   U1656 : INV_X1 port map( A => n1340, ZN => n1339);
   U1657 : AOI222_X1 port map( A1 => regs(640), A2 => n86, B1 => regs(2176), B2
                           => n188, C1 => regs(1152), C2 => n263, ZN => n1340);
   U1658 : INV_X1 port map( A => n1341, ZN => curr_proc_regs(191));
   U1659 : AOI221_X1 port map( B1 => n59, B2 => regs(1215), C1 => n306, C2 => 
                           regs(2239), A => n1342, ZN => n1341);
   U1660 : INV_X1 port map( A => n1343, ZN => n1342);
   U1661 : AOI222_X1 port map( A1 => regs(191), A2 => n86, B1 => regs(1727), B2
                           => n188, C1 => regs(703), C2 => n263, ZN => n1343);
   U1662 : INV_X1 port map( A => n1344, ZN => curr_proc_regs(703));
   U1663 : AOI221_X1 port map( B1 => n59, B2 => regs(1727), C1 => n306, C2 => 
                           regs(191), A => n1345, ZN => n1344);
   U1664 : INV_X1 port map( A => n1346, ZN => n1345);
   U1665 : AOI222_X1 port map( A1 => regs(703), A2 => n86, B1 => regs(2239), B2
                           => n188, C1 => regs(1215), C2 => n263, ZN => n1346);
   U1666 : INV_X1 port map( A => n1347, ZN => curr_proc_regs(190));
   U1667 : AOI221_X1 port map( B1 => n59, B2 => regs(1214), C1 => n306, C2 => 
                           regs(2238), A => n1348, ZN => n1347);
   U1668 : INV_X1 port map( A => n1349, ZN => n1348);
   U1669 : AOI222_X1 port map( A1 => regs(190), A2 => n86, B1 => regs(1726), B2
                           => n188, C1 => regs(702), C2 => n263, ZN => n1349);
   U1670 : INV_X1 port map( A => n1350, ZN => curr_proc_regs(702));
   U1671 : AOI221_X1 port map( B1 => n60, B2 => regs(1726), C1 => n306, C2 => 
                           regs(190), A => n1351, ZN => n1350);
   U1672 : INV_X1 port map( A => n1352, ZN => n1351);
   U1673 : AOI222_X1 port map( A1 => regs(702), A2 => n86, B1 => regs(2238), B2
                           => n188, C1 => regs(1214), C2 => n263, ZN => n1352);
   U1674 : INV_X1 port map( A => n1353, ZN => curr_proc_regs(189));
   U1675 : AOI221_X1 port map( B1 => n60, B2 => regs(1213), C1 => n306, C2 => 
                           regs(2237), A => n1354, ZN => n1353);
   U1676 : INV_X1 port map( A => n1355, ZN => n1354);
   U1677 : AOI222_X1 port map( A1 => regs(189), A2 => n87, B1 => regs(1725), B2
                           => n187, C1 => regs(701), C2 => n262, ZN => n1355);
   U1678 : INV_X1 port map( A => n1356, ZN => curr_proc_regs(701));
   U1679 : AOI221_X1 port map( B1 => n60, B2 => regs(1725), C1 => n306, C2 => 
                           regs(189), A => n1357, ZN => n1356);
   U1680 : INV_X1 port map( A => n1358, ZN => n1357);
   U1681 : AOI222_X1 port map( A1 => regs(701), A2 => n87, B1 => regs(2237), B2
                           => n187, C1 => regs(1213), C2 => n262, ZN => n1358);
   U1682 : INV_X1 port map( A => n1359, ZN => curr_proc_regs(188));
   U1683 : AOI221_X1 port map( B1 => n60, B2 => regs(1212), C1 => n306, C2 => 
                           regs(2236), A => n1360, ZN => n1359);
   U1684 : INV_X1 port map( A => n1361, ZN => n1360);
   U1685 : AOI222_X1 port map( A1 => regs(188), A2 => n87, B1 => regs(1724), B2
                           => n187, C1 => regs(700), C2 => n262, ZN => n1361);
   U1686 : INV_X1 port map( A => n1362, ZN => curr_proc_regs(700));
   U1687 : AOI221_X1 port map( B1 => n60, B2 => regs(1724), C1 => n306, C2 => 
                           regs(188), A => n1363, ZN => n1362);
   U1688 : INV_X1 port map( A => n1364, ZN => n1363);
   U1689 : AOI222_X1 port map( A1 => regs(700), A2 => n87, B1 => regs(2236), B2
                           => n187, C1 => regs(1212), C2 => n262, ZN => n1364);
   U1690 : INV_X1 port map( A => n1365, ZN => curr_proc_regs(187));
   U1691 : AOI221_X1 port map( B1 => n60, B2 => regs(1211), C1 => n306, C2 => 
                           regs(2235), A => n1366, ZN => n1365);
   U1692 : INV_X1 port map( A => n1367, ZN => n1366);
   U1693 : AOI222_X1 port map( A1 => regs(187), A2 => n87, B1 => regs(1723), B2
                           => n187, C1 => regs(699), C2 => n262, ZN => n1367);
   U1694 : INV_X1 port map( A => n1368, ZN => curr_proc_regs(699));
   U1695 : AOI221_X1 port map( B1 => n60, B2 => regs(1723), C1 => n305, C2 => 
                           regs(187), A => n1369, ZN => n1368);
   U1696 : INV_X1 port map( A => n1370, ZN => n1369);
   U1697 : AOI222_X1 port map( A1 => regs(699), A2 => n87, B1 => regs(2235), B2
                           => n187, C1 => regs(1211), C2 => n262, ZN => n1370);
   U1698 : INV_X1 port map( A => n1371, ZN => curr_proc_regs(186));
   U1699 : AOI221_X1 port map( B1 => n60, B2 => regs(1210), C1 => n305, C2 => 
                           regs(2234), A => n1372, ZN => n1371);
   U1700 : INV_X1 port map( A => n1373, ZN => n1372);
   U1701 : AOI222_X1 port map( A1 => regs(186), A2 => n87, B1 => regs(1722), B2
                           => n187, C1 => regs(698), C2 => n262, ZN => n1373);
   U1702 : INV_X1 port map( A => n1374, ZN => curr_proc_regs(698));
   U1703 : AOI221_X1 port map( B1 => n60, B2 => regs(1722), C1 => n305, C2 => 
                           regs(186), A => n1375, ZN => n1374);
   U1704 : INV_X1 port map( A => n1376, ZN => n1375);
   U1705 : AOI222_X1 port map( A1 => regs(698), A2 => n87, B1 => regs(2234), B2
                           => n187, C1 => regs(1210), C2 => n262, ZN => n1376);
   U1706 : INV_X1 port map( A => n1377, ZN => curr_proc_regs(185));
   U1707 : AOI221_X1 port map( B1 => n60, B2 => regs(1209), C1 => n305, C2 => 
                           regs(2233), A => n1378, ZN => n1377);
   U1708 : INV_X1 port map( A => n1379, ZN => n1378);
   U1709 : AOI222_X1 port map( A1 => regs(185), A2 => n87, B1 => regs(1721), B2
                           => n187, C1 => regs(697), C2 => n262, ZN => n1379);
   U1710 : INV_X1 port map( A => n1380, ZN => curr_proc_regs(697));
   U1711 : AOI221_X1 port map( B1 => n60, B2 => regs(1721), C1 => n305, C2 => 
                           regs(185), A => n1381, ZN => n1380);
   U1712 : INV_X1 port map( A => n1382, ZN => n1381);
   U1713 : AOI222_X1 port map( A1 => regs(697), A2 => n87, B1 => regs(2233), B2
                           => n187, C1 => regs(1209), C2 => n262, ZN => n1382);
   U1714 : INV_X1 port map( A => n1383, ZN => curr_proc_regs(184));
   U1715 : AOI221_X1 port map( B1 => n60, B2 => regs(1208), C1 => n305, C2 => 
                           regs(2232), A => n1384, ZN => n1383);
   U1716 : INV_X1 port map( A => n1385, ZN => n1384);
   U1717 : AOI222_X1 port map( A1 => regs(184), A2 => n87, B1 => regs(1720), B2
                           => n187, C1 => regs(696), C2 => n262, ZN => n1385);
   U1718 : INV_X1 port map( A => n1386, ZN => curr_proc_regs(696));
   U1719 : AOI221_X1 port map( B1 => n61, B2 => regs(1720), C1 => n305, C2 => 
                           regs(184), A => n1387, ZN => n1386);
   U1720 : INV_X1 port map( A => n1388, ZN => n1387);
   U1721 : AOI222_X1 port map( A1 => regs(696), A2 => n87, B1 => regs(2232), B2
                           => n187, C1 => regs(1208), C2 => n262, ZN => n1388);
   U1722 : INV_X1 port map( A => n1389, ZN => curr_proc_regs(183));
   U1723 : AOI221_X1 port map( B1 => n61, B2 => regs(1207), C1 => n305, C2 => 
                           regs(2231), A => n1390, ZN => n1389);
   U1724 : INV_X1 port map( A => n1391, ZN => n1390);
   U1725 : AOI222_X1 port map( A1 => regs(183), A2 => n88, B1 => regs(1719), B2
                           => n186, C1 => regs(695), C2 => n261, ZN => n1391);
   U1726 : INV_X1 port map( A => n1392, ZN => curr_proc_regs(695));
   U1727 : AOI221_X1 port map( B1 => n61, B2 => regs(1719), C1 => n305, C2 => 
                           regs(183), A => n1393, ZN => n1392);
   U1728 : INV_X1 port map( A => n1394, ZN => n1393);
   U1729 : AOI222_X1 port map( A1 => regs(695), A2 => n88, B1 => regs(2231), B2
                           => n186, C1 => regs(1207), C2 => n261, ZN => n1394);
   U1730 : INV_X1 port map( A => n1395, ZN => curr_proc_regs(182));
   U1731 : AOI221_X1 port map( B1 => n61, B2 => regs(1206), C1 => n305, C2 => 
                           regs(2230), A => n1396, ZN => n1395);
   U1732 : INV_X1 port map( A => n1397, ZN => n1396);
   U1733 : AOI222_X1 port map( A1 => regs(182), A2 => n88, B1 => regs(1718), B2
                           => n186, C1 => regs(694), C2 => n261, ZN => n1397);
   U1734 : INV_X1 port map( A => n1398, ZN => curr_proc_regs(694));
   U1735 : AOI221_X1 port map( B1 => n61, B2 => regs(1718), C1 => n305, C2 => 
                           regs(182), A => n1399, ZN => n1398);
   U1736 : INV_X1 port map( A => n1400, ZN => n1399);
   U1737 : AOI222_X1 port map( A1 => regs(694), A2 => n88, B1 => regs(2230), B2
                           => n186, C1 => regs(1206), C2 => n261, ZN => n1400);
   U1738 : INV_X1 port map( A => n1401, ZN => curr_proc_regs(181));
   U1739 : AOI221_X1 port map( B1 => n61, B2 => regs(1205), C1 => n305, C2 => 
                           regs(2229), A => n1402, ZN => n1401);
   U1740 : INV_X1 port map( A => n1403, ZN => n1402);
   U1741 : AOI222_X1 port map( A1 => regs(181), A2 => n88, B1 => regs(1717), B2
                           => n186, C1 => regs(693), C2 => n261, ZN => n1403);
   U1742 : INV_X1 port map( A => n1404, ZN => curr_proc_regs(693));
   U1743 : AOI221_X1 port map( B1 => n61, B2 => regs(1717), C1 => n304, C2 => 
                           regs(181), A => n1405, ZN => n1404);
   U1744 : INV_X1 port map( A => n1406, ZN => n1405);
   U1745 : AOI222_X1 port map( A1 => regs(693), A2 => n88, B1 => regs(2229), B2
                           => n186, C1 => regs(1205), C2 => n261, ZN => n1406);
   U1746 : INV_X1 port map( A => n1407, ZN => curr_proc_regs(180));
   U1747 : AOI221_X1 port map( B1 => n61, B2 => regs(1204), C1 => n304, C2 => 
                           regs(2228), A => n1408, ZN => n1407);
   U1748 : INV_X1 port map( A => n1409, ZN => n1408);
   U1749 : AOI222_X1 port map( A1 => regs(180), A2 => n88, B1 => regs(1716), B2
                           => n186, C1 => regs(692), C2 => n261, ZN => n1409);
   U1750 : INV_X1 port map( A => n1410, ZN => curr_proc_regs(692));
   U1751 : AOI221_X1 port map( B1 => n61, B2 => regs(1716), C1 => n304, C2 => 
                           regs(180), A => n1411, ZN => n1410);
   U1752 : INV_X1 port map( A => n1412, ZN => n1411);
   U1753 : AOI222_X1 port map( A1 => regs(692), A2 => n88, B1 => regs(2228), B2
                           => n186, C1 => regs(1204), C2 => n261, ZN => n1412);
   U1754 : INV_X1 port map( A => n1413, ZN => curr_proc_regs(179));
   U1755 : AOI221_X1 port map( B1 => n61, B2 => regs(1203), C1 => n304, C2 => 
                           regs(2227), A => n1414, ZN => n1413);
   U1756 : INV_X1 port map( A => n1415, ZN => n1414);
   U1757 : AOI222_X1 port map( A1 => regs(179), A2 => n88, B1 => regs(1715), B2
                           => n186, C1 => regs(691), C2 => n261, ZN => n1415);
   U1758 : INV_X1 port map( A => n1416, ZN => curr_proc_regs(691));
   U1759 : AOI221_X1 port map( B1 => n61, B2 => regs(1715), C1 => n304, C2 => 
                           regs(179), A => n1417, ZN => n1416);
   U1760 : INV_X1 port map( A => n1418, ZN => n1417);
   U1761 : AOI222_X1 port map( A1 => regs(691), A2 => n88, B1 => regs(2227), B2
                           => n186, C1 => regs(1203), C2 => n261, ZN => n1418);
   U1762 : INV_X1 port map( A => n1419, ZN => curr_proc_regs(178));
   U1763 : AOI221_X1 port map( B1 => n61, B2 => regs(1202), C1 => n304, C2 => 
                           regs(2226), A => n1420, ZN => n1419);
   U1764 : INV_X1 port map( A => n1421, ZN => n1420);
   U1765 : AOI222_X1 port map( A1 => regs(178), A2 => n88, B1 => regs(1714), B2
                           => n186, C1 => regs(690), C2 => n261, ZN => n1421);
   U1766 : INV_X1 port map( A => n1422, ZN => curr_proc_regs(690));
   U1767 : AOI221_X1 port map( B1 => n62, B2 => regs(1714), C1 => n304, C2 => 
                           regs(178), A => n1423, ZN => n1422);
   U1768 : INV_X1 port map( A => n1424, ZN => n1423);
   U1769 : AOI222_X1 port map( A1 => regs(690), A2 => n88, B1 => regs(2226), B2
                           => n186, C1 => regs(1202), C2 => n261, ZN => n1424);
   U1770 : INV_X1 port map( A => n1425, ZN => curr_proc_regs(177));
   U1771 : AOI221_X1 port map( B1 => n62, B2 => regs(1201), C1 => n304, C2 => 
                           regs(2225), A => n1426, ZN => n1425);
   U1772 : INV_X1 port map( A => n1427, ZN => n1426);
   U1773 : AOI222_X1 port map( A1 => regs(177), A2 => n89, B1 => regs(1713), B2
                           => n185, C1 => regs(689), C2 => n260, ZN => n1427);
   U1774 : INV_X1 port map( A => n1428, ZN => curr_proc_regs(689));
   U1775 : AOI221_X1 port map( B1 => n62, B2 => regs(1713), C1 => n304, C2 => 
                           regs(177), A => n1429, ZN => n1428);
   U1776 : INV_X1 port map( A => n1430, ZN => n1429);
   U1777 : AOI222_X1 port map( A1 => regs(689), A2 => n89, B1 => regs(2225), B2
                           => n185, C1 => regs(1201), C2 => n260, ZN => n1430);
   U1778 : INV_X1 port map( A => n1431, ZN => curr_proc_regs(176));
   U1779 : AOI221_X1 port map( B1 => n62, B2 => regs(1200), C1 => n304, C2 => 
                           regs(2224), A => n1432, ZN => n1431);
   U1780 : INV_X1 port map( A => n1433, ZN => n1432);
   U1781 : AOI222_X1 port map( A1 => regs(176), A2 => n89, B1 => regs(1712), B2
                           => n185, C1 => regs(688), C2 => n260, ZN => n1433);
   U1782 : INV_X1 port map( A => n1434, ZN => curr_proc_regs(688));
   U1783 : AOI221_X1 port map( B1 => n62, B2 => regs(1712), C1 => n304, C2 => 
                           regs(176), A => n1435, ZN => n1434);
   U1784 : INV_X1 port map( A => n1436, ZN => n1435);
   U1785 : AOI222_X1 port map( A1 => regs(688), A2 => n89, B1 => regs(2224), B2
                           => n185, C1 => regs(1200), C2 => n260, ZN => n1436);
   U1786 : INV_X1 port map( A => n1437, ZN => curr_proc_regs(175));
   U1787 : AOI221_X1 port map( B1 => n62, B2 => regs(1199), C1 => n304, C2 => 
                           regs(2223), A => n1438, ZN => n1437);
   U1788 : INV_X1 port map( A => n1439, ZN => n1438);
   U1789 : AOI222_X1 port map( A1 => regs(175), A2 => n89, B1 => regs(1711), B2
                           => n185, C1 => regs(687), C2 => n260, ZN => n1439);
   U1790 : INV_X1 port map( A => n1440, ZN => curr_proc_regs(687));
   U1791 : AOI221_X1 port map( B1 => n62, B2 => regs(1711), C1 => n303, C2 => 
                           regs(175), A => n1441, ZN => n1440);
   U1792 : INV_X1 port map( A => n1442, ZN => n1441);
   U1793 : AOI222_X1 port map( A1 => regs(687), A2 => n89, B1 => regs(2223), B2
                           => n185, C1 => regs(1199), C2 => n260, ZN => n1442);
   U1794 : INV_X1 port map( A => n1443, ZN => curr_proc_regs(174));
   U1795 : AOI221_X1 port map( B1 => n62, B2 => regs(1198), C1 => n303, C2 => 
                           regs(2222), A => n1444, ZN => n1443);
   U1796 : INV_X1 port map( A => n1445, ZN => n1444);
   U1797 : AOI222_X1 port map( A1 => regs(174), A2 => n89, B1 => regs(1710), B2
                           => n185, C1 => regs(686), C2 => n260, ZN => n1445);
   U1798 : INV_X1 port map( A => n1446, ZN => curr_proc_regs(686));
   U1799 : AOI221_X1 port map( B1 => n62, B2 => regs(1710), C1 => n303, C2 => 
                           regs(174), A => n1447, ZN => n1446);
   U1800 : INV_X1 port map( A => n1448, ZN => n1447);
   U1801 : AOI222_X1 port map( A1 => regs(686), A2 => n89, B1 => regs(2222), B2
                           => n185, C1 => regs(1198), C2 => n260, ZN => n1448);
   U1802 : INV_X1 port map( A => n1449, ZN => curr_proc_regs(173));
   U1803 : AOI221_X1 port map( B1 => n62, B2 => regs(1197), C1 => n303, C2 => 
                           regs(2221), A => n1450, ZN => n1449);
   U1804 : INV_X1 port map( A => n1451, ZN => n1450);
   U1805 : AOI222_X1 port map( A1 => regs(173), A2 => n89, B1 => regs(1709), B2
                           => n185, C1 => regs(685), C2 => n260, ZN => n1451);
   U1806 : INV_X1 port map( A => n1452, ZN => curr_proc_regs(685));
   U1807 : AOI221_X1 port map( B1 => n62, B2 => regs(1709), C1 => n303, C2 => 
                           regs(173), A => n1453, ZN => n1452);
   U1808 : INV_X1 port map( A => n1454, ZN => n1453);
   U1809 : AOI222_X1 port map( A1 => regs(685), A2 => n89, B1 => regs(2221), B2
                           => n185, C1 => regs(1197), C2 => n260, ZN => n1454);
   U1810 : INV_X1 port map( A => n1455, ZN => curr_proc_regs(172));
   U1811 : AOI221_X1 port map( B1 => n62, B2 => regs(1196), C1 => n303, C2 => 
                           regs(2220), A => n1456, ZN => n1455);
   U1812 : INV_X1 port map( A => n1457, ZN => n1456);
   U1813 : AOI222_X1 port map( A1 => regs(172), A2 => n89, B1 => regs(1708), B2
                           => n185, C1 => regs(684), C2 => n260, ZN => n1457);
   U1814 : INV_X1 port map( A => n1458, ZN => curr_proc_regs(684));
   U1815 : AOI221_X1 port map( B1 => n63, B2 => regs(1708), C1 => n303, C2 => 
                           regs(172), A => n1459, ZN => n1458);
   U1816 : INV_X1 port map( A => n1460, ZN => n1459);
   U1817 : AOI222_X1 port map( A1 => regs(684), A2 => n89, B1 => regs(2220), B2
                           => n185, C1 => regs(1196), C2 => n260, ZN => n1460);
   U1818 : INV_X1 port map( A => n1461, ZN => curr_proc_regs(171));
   U1819 : AOI221_X1 port map( B1 => n63, B2 => regs(1195), C1 => n303, C2 => 
                           regs(2219), A => n1462, ZN => n1461);
   U1820 : INV_X1 port map( A => n1463, ZN => n1462);
   U1821 : AOI222_X1 port map( A1 => regs(171), A2 => n90, B1 => regs(1707), B2
                           => n184, C1 => regs(683), C2 => n259, ZN => n1463);
   U1822 : INV_X1 port map( A => n1464, ZN => curr_proc_regs(683));
   U1823 : AOI221_X1 port map( B1 => n63, B2 => regs(1707), C1 => n303, C2 => 
                           regs(171), A => n1465, ZN => n1464);
   U1824 : INV_X1 port map( A => n1466, ZN => n1465);
   U1825 : AOI222_X1 port map( A1 => regs(683), A2 => n90, B1 => regs(2219), B2
                           => n184, C1 => regs(1195), C2 => n259, ZN => n1466);
   U1826 : INV_X1 port map( A => n1467, ZN => curr_proc_regs(170));
   U1827 : AOI221_X1 port map( B1 => n63, B2 => regs(1194), C1 => n303, C2 => 
                           regs(2218), A => n1468, ZN => n1467);
   U1828 : INV_X1 port map( A => n1469, ZN => n1468);
   U1829 : AOI222_X1 port map( A1 => regs(170), A2 => n90, B1 => regs(1706), B2
                           => n184, C1 => regs(682), C2 => n259, ZN => n1469);
   U1830 : INV_X1 port map( A => n1470, ZN => curr_proc_regs(682));
   U1831 : AOI221_X1 port map( B1 => n63, B2 => regs(1706), C1 => n303, C2 => 
                           regs(170), A => n1471, ZN => n1470);
   U1832 : INV_X1 port map( A => n1472, ZN => n1471);
   U1833 : AOI222_X1 port map( A1 => regs(682), A2 => n90, B1 => regs(2218), B2
                           => n184, C1 => regs(1194), C2 => n259, ZN => n1472);
   U1834 : INV_X1 port map( A => n1473, ZN => curr_proc_regs(169));
   U1835 : AOI221_X1 port map( B1 => n63, B2 => regs(1193), C1 => n303, C2 => 
                           regs(2217), A => n1474, ZN => n1473);
   U1836 : INV_X1 port map( A => n1475, ZN => n1474);
   U1837 : AOI222_X1 port map( A1 => regs(169), A2 => n90, B1 => regs(1705), B2
                           => n184, C1 => regs(681), C2 => n259, ZN => n1475);
   U1838 : INV_X1 port map( A => n1476, ZN => curr_proc_regs(681));
   U1839 : AOI221_X1 port map( B1 => n63, B2 => regs(1705), C1 => n302, C2 => 
                           regs(169), A => n1477, ZN => n1476);
   U1840 : INV_X1 port map( A => n1478, ZN => n1477);
   U1841 : AOI222_X1 port map( A1 => regs(681), A2 => n90, B1 => regs(2217), B2
                           => n184, C1 => regs(1193), C2 => n259, ZN => n1478);
   U1842 : INV_X1 port map( A => n1479, ZN => curr_proc_regs(168));
   U1843 : AOI221_X1 port map( B1 => n63, B2 => regs(1192), C1 => n302, C2 => 
                           regs(2216), A => n1480, ZN => n1479);
   U1844 : INV_X1 port map( A => n1481, ZN => n1480);
   U1845 : AOI222_X1 port map( A1 => regs(168), A2 => n90, B1 => regs(1704), B2
                           => n184, C1 => regs(680), C2 => n259, ZN => n1481);
   U1846 : INV_X1 port map( A => n1482, ZN => curr_proc_regs(680));
   U1847 : AOI221_X1 port map( B1 => n63, B2 => regs(1704), C1 => n302, C2 => 
                           regs(168), A => n1483, ZN => n1482);
   U1848 : INV_X1 port map( A => n1484, ZN => n1483);
   U1849 : AOI222_X1 port map( A1 => regs(680), A2 => n90, B1 => regs(2216), B2
                           => n184, C1 => regs(1192), C2 => n259, ZN => n1484);
   U1850 : INV_X1 port map( A => n1485, ZN => curr_proc_regs(167));
   U1851 : AOI221_X1 port map( B1 => n63, B2 => regs(1191), C1 => n302, C2 => 
                           regs(2215), A => n1486, ZN => n1485);
   U1852 : INV_X1 port map( A => n1487, ZN => n1486);
   U1853 : AOI222_X1 port map( A1 => regs(167), A2 => n90, B1 => regs(1703), B2
                           => n184, C1 => regs(679), C2 => n259, ZN => n1487);
   U1854 : INV_X1 port map( A => n1488, ZN => curr_proc_regs(679));
   U1855 : AOI221_X1 port map( B1 => n63, B2 => regs(1703), C1 => n302, C2 => 
                           regs(167), A => n1489, ZN => n1488);
   U1856 : INV_X1 port map( A => n1490, ZN => n1489);
   U1857 : AOI222_X1 port map( A1 => regs(679), A2 => n90, B1 => regs(2215), B2
                           => n184, C1 => regs(1191), C2 => n259, ZN => n1490);
   U1858 : INV_X1 port map( A => n1491, ZN => curr_proc_regs(166));
   U1859 : AOI221_X1 port map( B1 => n63, B2 => regs(1190), C1 => n302, C2 => 
                           regs(2214), A => n1492, ZN => n1491);
   U1860 : INV_X1 port map( A => n1493, ZN => n1492);
   U1861 : AOI222_X1 port map( A1 => regs(166), A2 => n90, B1 => regs(1702), B2
                           => n184, C1 => regs(678), C2 => n259, ZN => n1493);
   U1862 : INV_X1 port map( A => n1494, ZN => curr_proc_regs(678));
   U1863 : AOI221_X1 port map( B1 => n64, B2 => regs(1702), C1 => n302, C2 => 
                           regs(166), A => n1495, ZN => n1494);
   U1864 : INV_X1 port map( A => n1496, ZN => n1495);
   U1865 : AOI222_X1 port map( A1 => regs(678), A2 => n90, B1 => regs(2214), B2
                           => n184, C1 => regs(1190), C2 => n259, ZN => n1496);
   U1866 : INV_X1 port map( A => n1497, ZN => curr_proc_regs(165));
   U1867 : AOI221_X1 port map( B1 => n64, B2 => regs(1189), C1 => n302, C2 => 
                           regs(2213), A => n1498, ZN => n1497);
   U1868 : INV_X1 port map( A => n1499, ZN => n1498);
   U1869 : AOI222_X1 port map( A1 => regs(165), A2 => n91, B1 => regs(1701), B2
                           => n183, C1 => regs(677), C2 => n258, ZN => n1499);
   U1870 : INV_X1 port map( A => n1500, ZN => curr_proc_regs(677));
   U1871 : AOI221_X1 port map( B1 => n64, B2 => regs(1701), C1 => n302, C2 => 
                           regs(165), A => n1501, ZN => n1500);
   U1872 : INV_X1 port map( A => n1502, ZN => n1501);
   U1873 : AOI222_X1 port map( A1 => regs(677), A2 => n91, B1 => regs(2213), B2
                           => n183, C1 => regs(1189), C2 => n258, ZN => n1502);
   U1874 : INV_X1 port map( A => n1503, ZN => curr_proc_regs(164));
   U1875 : AOI221_X1 port map( B1 => n64, B2 => regs(1188), C1 => n302, C2 => 
                           regs(2212), A => n1504, ZN => n1503);
   U1876 : INV_X1 port map( A => n1505, ZN => n1504);
   U1877 : AOI222_X1 port map( A1 => regs(164), A2 => n91, B1 => regs(1700), B2
                           => n183, C1 => regs(676), C2 => n258, ZN => n1505);
   U1878 : INV_X1 port map( A => n1506, ZN => curr_proc_regs(676));
   U1879 : AOI221_X1 port map( B1 => n64, B2 => regs(1700), C1 => n302, C2 => 
                           regs(164), A => n1507, ZN => n1506);
   U1880 : INV_X1 port map( A => n1508, ZN => n1507);
   U1881 : AOI222_X1 port map( A1 => regs(676), A2 => n91, B1 => regs(2212), B2
                           => n183, C1 => regs(1188), C2 => n258, ZN => n1508);
   U1882 : INV_X1 port map( A => n1509, ZN => curr_proc_regs(163));
   U1883 : AOI221_X1 port map( B1 => n64, B2 => regs(1187), C1 => n302, C2 => 
                           regs(2211), A => n1510, ZN => n1509);
   U1884 : INV_X1 port map( A => n1511, ZN => n1510);
   U1885 : AOI222_X1 port map( A1 => regs(163), A2 => n91, B1 => regs(1699), B2
                           => n183, C1 => regs(675), C2 => n258, ZN => n1511);
   U1886 : INV_X1 port map( A => n1512, ZN => curr_proc_regs(675));
   U1887 : AOI221_X1 port map( B1 => n64, B2 => regs(1699), C1 => n301, C2 => 
                           regs(163), A => n1513, ZN => n1512);
   U1888 : INV_X1 port map( A => n1514, ZN => n1513);
   U1889 : AOI222_X1 port map( A1 => regs(675), A2 => n91, B1 => regs(2211), B2
                           => n183, C1 => regs(1187), C2 => n258, ZN => n1514);
   U1890 : INV_X1 port map( A => n1515, ZN => curr_proc_regs(162));
   U1891 : AOI221_X1 port map( B1 => n64, B2 => regs(1186), C1 => n301, C2 => 
                           regs(2210), A => n1516, ZN => n1515);
   U1892 : INV_X1 port map( A => n1517, ZN => n1516);
   U1893 : AOI222_X1 port map( A1 => regs(162), A2 => n91, B1 => regs(1698), B2
                           => n183, C1 => regs(674), C2 => n258, ZN => n1517);
   U1894 : INV_X1 port map( A => n1518, ZN => curr_proc_regs(674));
   U1895 : AOI221_X1 port map( B1 => n64, B2 => regs(1698), C1 => n301, C2 => 
                           regs(162), A => n1519, ZN => n1518);
   U1896 : INV_X1 port map( A => n1520, ZN => n1519);
   U1897 : AOI222_X1 port map( A1 => regs(674), A2 => n91, B1 => regs(2210), B2
                           => n183, C1 => regs(1186), C2 => n258, ZN => n1520);
   U1898 : INV_X1 port map( A => n1521, ZN => curr_proc_regs(161));
   U1899 : AOI221_X1 port map( B1 => n64, B2 => regs(1185), C1 => n301, C2 => 
                           regs(2209), A => n1522, ZN => n1521);
   U1900 : INV_X1 port map( A => n1523, ZN => n1522);
   U1901 : AOI222_X1 port map( A1 => regs(161), A2 => n91, B1 => regs(1697), B2
                           => n183, C1 => regs(673), C2 => n258, ZN => n1523);
   U1902 : INV_X1 port map( A => n1524, ZN => curr_proc_regs(673));
   U1903 : AOI221_X1 port map( B1 => n64, B2 => regs(1697), C1 => n301, C2 => 
                           regs(161), A => n1525, ZN => n1524);
   U1904 : INV_X1 port map( A => n1526, ZN => n1525);
   U1905 : AOI222_X1 port map( A1 => regs(673), A2 => n91, B1 => regs(2209), B2
                           => n183, C1 => regs(1185), C2 => n258, ZN => n1526);
   U1906 : INV_X1 port map( A => n1527, ZN => curr_proc_regs(160));
   U1907 : AOI221_X1 port map( B1 => n64, B2 => regs(1184), C1 => n301, C2 => 
                           regs(2208), A => n1528, ZN => n1527);
   U1908 : INV_X1 port map( A => n1529, ZN => n1528);
   U1909 : AOI222_X1 port map( A1 => regs(160), A2 => n91, B1 => regs(1696), B2
                           => n183, C1 => regs(672), C2 => n258, ZN => n1529);
   U1910 : INV_X1 port map( A => n1530, ZN => curr_proc_regs(672));
   U1911 : AOI221_X1 port map( B1 => n49, B2 => regs(1696), C1 => n301, C2 => 
                           regs(160), A => n1531, ZN => n1530);
   U1912 : INV_X1 port map( A => n1532, ZN => n1531);
   U1913 : AOI222_X1 port map( A1 => regs(672), A2 => n91, B1 => regs(2208), B2
                           => n183, C1 => regs(1184), C2 => n258, ZN => n1532);
   U1914 : INV_X1 port map( A => n1533, ZN => curr_proc_regs(223));
   U1915 : AOI221_X1 port map( B1 => n43, B2 => regs(1247), C1 => n306, C2 => 
                           regs(2271), A => n1534, ZN => n1533);
   U1916 : INV_X1 port map( A => n1535, ZN => n1534);
   U1917 : AOI222_X1 port map( A1 => regs(223), A2 => n131, B1 => regs(1759), 
                           B2 => n182, C1 => regs(735), C2 => n257, ZN => n1535
                           );
   U1918 : INV_X1 port map( A => n1536, ZN => curr_proc_regs(735));
   U1919 : AOI221_X1 port map( B1 => n43, B2 => regs(1759), C1 => n322, C2 => 
                           regs(223), A => n1537, ZN => n1536);
   U1920 : INV_X1 port map( A => n1538, ZN => n1537);
   U1921 : AOI222_X1 port map( A1 => regs(735), A2 => n124, B1 => regs(2271), 
                           B2 => n182, C1 => regs(1247), C2 => n257, ZN => 
                           n1538);
   U1922 : INV_X1 port map( A => n1539, ZN => curr_proc_regs(222));
   U1923 : AOI221_X1 port map( B1 => n43, B2 => regs(1246), C1 => n322, C2 => 
                           regs(2270), A => n1540, ZN => n1539);
   U1924 : INV_X1 port map( A => n1541, ZN => n1540);
   U1925 : AOI222_X1 port map( A1 => regs(222), A2 => n124, B1 => regs(1758), 
                           B2 => n182, C1 => regs(734), C2 => n257, ZN => n1541
                           );
   U1926 : INV_X1 port map( A => n1542, ZN => curr_proc_regs(734));
   U1927 : AOI221_X1 port map( B1 => n44, B2 => regs(1758), C1 => n322, C2 => 
                           regs(222), A => n1543, ZN => n1542);
   U1928 : INV_X1 port map( A => n1544, ZN => n1543);
   U1929 : AOI222_X1 port map( A1 => regs(734), A2 => n124, B1 => regs(2270), 
                           B2 => n182, C1 => regs(1246), C2 => n257, ZN => 
                           n1544);
   U1930 : INV_X1 port map( A => n1545, ZN => curr_proc_regs(221));
   U1931 : AOI221_X1 port map( B1 => n44, B2 => regs(1245), C1 => n322, C2 => 
                           regs(2269), A => n1546, ZN => n1545);
   U1932 : INV_X1 port map( A => n1547, ZN => n1546);
   U1933 : AOI222_X1 port map( A1 => regs(221), A2 => n124, B1 => regs(1757), 
                           B2 => n182, C1 => regs(733), C2 => n257, ZN => n1547
                           );
   U1934 : INV_X1 port map( A => n1548, ZN => curr_proc_regs(733));
   U1935 : AOI221_X1 port map( B1 => n44, B2 => regs(1757), C1 => n322, C2 => 
                           regs(221), A => n1549, ZN => n1548);
   U1936 : INV_X1 port map( A => n1550, ZN => n1549);
   U1937 : AOI222_X1 port map( A1 => regs(733), A2 => n124, B1 => regs(2269), 
                           B2 => n182, C1 => regs(1245), C2 => n257, ZN => 
                           n1550);
   U1938 : INV_X1 port map( A => n1551, ZN => curr_proc_regs(220));
   U1939 : AOI221_X1 port map( B1 => n44, B2 => regs(1244), C1 => n322, C2 => 
                           regs(2268), A => n1552, ZN => n1551);
   U1940 : INV_X1 port map( A => n1553, ZN => n1552);
   U1941 : AOI222_X1 port map( A1 => regs(220), A2 => n124, B1 => regs(1756), 
                           B2 => n182, C1 => regs(732), C2 => n257, ZN => n1553
                           );
   U1942 : INV_X1 port map( A => n1554, ZN => curr_proc_regs(732));
   U1943 : AOI221_X1 port map( B1 => n44, B2 => regs(1756), C1 => n321, C2 => 
                           regs(220), A => n1555, ZN => n1554);
   U1944 : INV_X1 port map( A => n1556, ZN => n1555);
   U1945 : AOI222_X1 port map( A1 => regs(732), A2 => n124, B1 => regs(2268), 
                           B2 => n182, C1 => regs(1244), C2 => n257, ZN => 
                           n1556);
   U1946 : INV_X1 port map( A => n1557, ZN => curr_proc_regs(219));
   U1947 : AOI221_X1 port map( B1 => n44, B2 => regs(1243), C1 => n321, C2 => 
                           regs(2267), A => n1558, ZN => n1557);
   U1948 : INV_X1 port map( A => n1559, ZN => n1558);
   U1949 : AOI222_X1 port map( A1 => regs(219), A2 => n124, B1 => regs(1755), 
                           B2 => n182, C1 => regs(731), C2 => n257, ZN => n1559
                           );
   U1950 : INV_X1 port map( A => n1560, ZN => curr_proc_regs(731));
   U1951 : AOI221_X1 port map( B1 => n44, B2 => regs(1755), C1 => n321, C2 => 
                           regs(219), A => n1561, ZN => n1560);
   U1952 : INV_X1 port map( A => n1562, ZN => n1561);
   U1953 : AOI222_X1 port map( A1 => regs(731), A2 => n124, B1 => regs(2267), 
                           B2 => n182, C1 => regs(1243), C2 => n257, ZN => 
                           n1562);
   U1954 : INV_X1 port map( A => n1563, ZN => curr_proc_regs(218));
   U1955 : AOI221_X1 port map( B1 => n44, B2 => regs(1242), C1 => n321, C2 => 
                           regs(2266), A => n1564, ZN => n1563);
   U1956 : INV_X1 port map( A => n1565, ZN => n1564);
   U1957 : AOI222_X1 port map( A1 => regs(218), A2 => n124, B1 => regs(1754), 
                           B2 => n182, C1 => regs(730), C2 => n257, ZN => n1565
                           );
   U1958 : INV_X1 port map( A => n1566, ZN => curr_proc_regs(730));
   U1959 : AOI221_X1 port map( B1 => n44, B2 => regs(1754), C1 => n321, C2 => 
                           regs(218), A => n1567, ZN => n1566);
   U1960 : INV_X1 port map( A => n1568, ZN => n1567);
   U1961 : AOI222_X1 port map( A1 => regs(730), A2 => n124, B1 => regs(2266), 
                           B2 => n182, C1 => regs(1242), C2 => n257, ZN => 
                           n1568);
   U1962 : INV_X1 port map( A => n1569, ZN => curr_proc_regs(217));
   U1963 : AOI221_X1 port map( B1 => n44, B2 => regs(1241), C1 => n321, C2 => 
                           regs(2265), A => n1570, ZN => n1569);
   U1964 : INV_X1 port map( A => n1571, ZN => n1570);
   U1965 : AOI222_X1 port map( A1 => regs(217), A2 => n124, B1 => regs(1753), 
                           B2 => n181, C1 => regs(729), C2 => n256, ZN => n1571
                           );
   U1966 : INV_X1 port map( A => n1572, ZN => curr_proc_regs(729));
   U1967 : AOI221_X1 port map( B1 => n44, B2 => regs(1753), C1 => n321, C2 => 
                           regs(217), A => n1573, ZN => n1572);
   U1968 : INV_X1 port map( A => n1574, ZN => n1573);
   U1969 : AOI222_X1 port map( A1 => regs(729), A2 => n125, B1 => regs(2265), 
                           B2 => n181, C1 => regs(1241), C2 => n256, ZN => 
                           n1574);
   U1970 : INV_X1 port map( A => n1575, ZN => curr_proc_regs(216));
   U1971 : AOI221_X1 port map( B1 => n44, B2 => regs(1240), C1 => n321, C2 => 
                           regs(2264), A => n1576, ZN => n1575);
   U1972 : INV_X1 port map( A => n1577, ZN => n1576);
   U1973 : AOI222_X1 port map( A1 => regs(216), A2 => n125, B1 => regs(1752), 
                           B2 => n181, C1 => regs(728), C2 => n256, ZN => n1577
                           );
   U1974 : INV_X1 port map( A => n1578, ZN => curr_proc_regs(728));
   U1975 : AOI221_X1 port map( B1 => n45, B2 => regs(1752), C1 => n321, C2 => 
                           regs(216), A => n1579, ZN => n1578);
   U1976 : INV_X1 port map( A => n1580, ZN => n1579);
   U1977 : AOI222_X1 port map( A1 => regs(728), A2 => n125, B1 => regs(2264), 
                           B2 => n181, C1 => regs(1240), C2 => n256, ZN => 
                           n1580);
   U1978 : INV_X1 port map( A => n1581, ZN => curr_proc_regs(215));
   U1979 : AOI221_X1 port map( B1 => n45, B2 => regs(1239), C1 => n321, C2 => 
                           regs(2263), A => n1582, ZN => n1581);
   U1980 : INV_X1 port map( A => n1583, ZN => n1582);
   U1981 : AOI222_X1 port map( A1 => regs(215), A2 => n125, B1 => regs(1751), 
                           B2 => n181, C1 => regs(727), C2 => n256, ZN => n1583
                           );
   U1982 : INV_X1 port map( A => n1584, ZN => curr_proc_regs(727));
   U1983 : AOI221_X1 port map( B1 => n45, B2 => regs(1751), C1 => n321, C2 => 
                           regs(215), A => n1585, ZN => n1584);
   U1984 : INV_X1 port map( A => n1586, ZN => n1585);
   U1985 : AOI222_X1 port map( A1 => regs(727), A2 => n125, B1 => regs(2263), 
                           B2 => n181, C1 => regs(1239), C2 => n256, ZN => 
                           n1586);
   U1986 : INV_X1 port map( A => n1587, ZN => curr_proc_regs(214));
   U1987 : AOI221_X1 port map( B1 => n45, B2 => regs(1238), C1 => n321, C2 => 
                           regs(2262), A => n1588, ZN => n1587);
   U1988 : INV_X1 port map( A => n1589, ZN => n1588);
   U1989 : AOI222_X1 port map( A1 => regs(214), A2 => n125, B1 => regs(1750), 
                           B2 => n181, C1 => regs(726), C2 => n256, ZN => n1589
                           );
   U1990 : INV_X1 port map( A => n1590, ZN => curr_proc_regs(726));
   U1991 : AOI221_X1 port map( B1 => n45, B2 => regs(1750), C1 => n320, C2 => 
                           regs(214), A => n1591, ZN => n1590);
   U1992 : INV_X1 port map( A => n1592, ZN => n1591);
   U1993 : AOI222_X1 port map( A1 => regs(726), A2 => n125, B1 => regs(2262), 
                           B2 => n181, C1 => regs(1238), C2 => n256, ZN => 
                           n1592);
   U1994 : INV_X1 port map( A => n1593, ZN => curr_proc_regs(213));
   U1995 : AOI221_X1 port map( B1 => n45, B2 => regs(1237), C1 => n320, C2 => 
                           regs(2261), A => n1594, ZN => n1593);
   U1996 : INV_X1 port map( A => n1595, ZN => n1594);
   U1997 : AOI222_X1 port map( A1 => regs(213), A2 => n125, B1 => regs(1749), 
                           B2 => n181, C1 => regs(725), C2 => n256, ZN => n1595
                           );
   U1998 : INV_X1 port map( A => n1596, ZN => curr_proc_regs(725));
   U1999 : AOI221_X1 port map( B1 => n45, B2 => regs(1749), C1 => n320, C2 => 
                           regs(213), A => n1597, ZN => n1596);
   U2000 : INV_X1 port map( A => n1598, ZN => n1597);
   U2001 : AOI222_X1 port map( A1 => regs(725), A2 => n125, B1 => regs(2261), 
                           B2 => n181, C1 => regs(1237), C2 => n256, ZN => 
                           n1598);
   U2002 : INV_X1 port map( A => n1599, ZN => curr_proc_regs(212));
   U2003 : AOI221_X1 port map( B1 => n45, B2 => regs(1236), C1 => n320, C2 => 
                           regs(2260), A => n1600, ZN => n1599);
   U2004 : INV_X1 port map( A => n1601, ZN => n1600);
   U2005 : AOI222_X1 port map( A1 => regs(212), A2 => n125, B1 => regs(1748), 
                           B2 => n181, C1 => regs(724), C2 => n256, ZN => n1601
                           );
   U2006 : INV_X1 port map( A => n1602, ZN => curr_proc_regs(724));
   U2007 : AOI221_X1 port map( B1 => n45, B2 => regs(1748), C1 => n320, C2 => 
                           regs(212), A => n1603, ZN => n1602);
   U2008 : INV_X1 port map( A => n1604, ZN => n1603);
   U2009 : AOI222_X1 port map( A1 => regs(724), A2 => n125, B1 => regs(2260), 
                           B2 => n181, C1 => regs(1236), C2 => n256, ZN => 
                           n1604);
   U2010 : INV_X1 port map( A => n1605, ZN => curr_proc_regs(211));
   U2011 : AOI221_X1 port map( B1 => n45, B2 => regs(1235), C1 => n320, C2 => 
                           regs(2259), A => n1606, ZN => n1605);
   U2012 : INV_X1 port map( A => n1607, ZN => n1606);
   U2013 : AOI222_X1 port map( A1 => regs(211), A2 => n125, B1 => regs(1747), 
                           B2 => n180, C1 => regs(723), C2 => n255, ZN => n1607
                           );
   U2014 : INV_X1 port map( A => n1608, ZN => curr_proc_regs(723));
   U2015 : AOI221_X1 port map( B1 => n45, B2 => regs(1747), C1 => n320, C2 => 
                           regs(211), A => n1609, ZN => n1608);
   U2016 : INV_X1 port map( A => n1610, ZN => n1609);
   U2017 : AOI222_X1 port map( A1 => regs(723), A2 => n126, B1 => regs(2259), 
                           B2 => n180, C1 => regs(1235), C2 => n255, ZN => 
                           n1610);
   U2018 : INV_X1 port map( A => n1611, ZN => curr_proc_regs(210));
   U2019 : AOI221_X1 port map( B1 => n45, B2 => regs(1234), C1 => n320, C2 => 
                           regs(2258), A => n1612, ZN => n1611);
   U2020 : INV_X1 port map( A => n1613, ZN => n1612);
   U2021 : AOI222_X1 port map( A1 => regs(210), A2 => n126, B1 => regs(1746), 
                           B2 => n180, C1 => regs(722), C2 => n255, ZN => n1613
                           );
   U2022 : INV_X1 port map( A => n1614, ZN => curr_proc_regs(722));
   U2023 : AOI221_X1 port map( B1 => n46, B2 => regs(1746), C1 => n320, C2 => 
                           regs(210), A => n1615, ZN => n1614);
   U2024 : INV_X1 port map( A => n1616, ZN => n1615);
   U2025 : AOI222_X1 port map( A1 => regs(722), A2 => n126, B1 => regs(2258), 
                           B2 => n180, C1 => regs(1234), C2 => n255, ZN => 
                           n1616);
   U2026 : INV_X1 port map( A => n1617, ZN => curr_proc_regs(209));
   U2027 : AOI221_X1 port map( B1 => n46, B2 => regs(1233), C1 => n320, C2 => 
                           regs(2257), A => n1618, ZN => n1617);
   U2028 : INV_X1 port map( A => n1619, ZN => n1618);
   U2029 : AOI222_X1 port map( A1 => regs(209), A2 => n126, B1 => regs(1745), 
                           B2 => n180, C1 => regs(721), C2 => n255, ZN => n1619
                           );
   U2030 : INV_X1 port map( A => n1620, ZN => curr_proc_regs(721));
   U2031 : AOI221_X1 port map( B1 => n46, B2 => regs(1745), C1 => n320, C2 => 
                           regs(209), A => n1621, ZN => n1620);
   U2032 : INV_X1 port map( A => n1622, ZN => n1621);
   U2033 : AOI222_X1 port map( A1 => regs(721), A2 => n126, B1 => regs(2257), 
                           B2 => n180, C1 => regs(1233), C2 => n255, ZN => 
                           n1622);
   U2034 : INV_X1 port map( A => n1623, ZN => curr_proc_regs(208));
   U2035 : AOI221_X1 port map( B1 => n46, B2 => regs(1232), C1 => n320, C2 => 
                           regs(2256), A => n1624, ZN => n1623);
   U2036 : INV_X1 port map( A => n1625, ZN => n1624);
   U2037 : AOI222_X1 port map( A1 => regs(208), A2 => n126, B1 => regs(1744), 
                           B2 => n180, C1 => regs(720), C2 => n255, ZN => n1625
                           );
   U2038 : INV_X1 port map( A => n1626, ZN => curr_proc_regs(720));
   U2039 : AOI221_X1 port map( B1 => n46, B2 => regs(1744), C1 => n319, C2 => 
                           regs(208), A => n1627, ZN => n1626);
   U2040 : INV_X1 port map( A => n1628, ZN => n1627);
   U2041 : AOI222_X1 port map( A1 => regs(720), A2 => n126, B1 => regs(2256), 
                           B2 => n180, C1 => regs(1232), C2 => n255, ZN => 
                           n1628);
   U2042 : INV_X1 port map( A => n1629, ZN => curr_proc_regs(207));
   U2043 : AOI221_X1 port map( B1 => n46, B2 => regs(1231), C1 => n319, C2 => 
                           regs(2255), A => n1630, ZN => n1629);
   U2044 : INV_X1 port map( A => n1631, ZN => n1630);
   U2045 : AOI222_X1 port map( A1 => regs(207), A2 => n126, B1 => regs(1743), 
                           B2 => n180, C1 => regs(719), C2 => n255, ZN => n1631
                           );
   U2046 : INV_X1 port map( A => n1632, ZN => curr_proc_regs(719));
   U2047 : AOI221_X1 port map( B1 => n46, B2 => regs(1743), C1 => n319, C2 => 
                           regs(207), A => n1633, ZN => n1632);
   U2048 : INV_X1 port map( A => n1634, ZN => n1633);
   U2049 : AOI222_X1 port map( A1 => regs(719), A2 => n126, B1 => regs(2255), 
                           B2 => n180, C1 => regs(1231), C2 => n255, ZN => 
                           n1634);
   U2050 : INV_X1 port map( A => n1635, ZN => curr_proc_regs(206));
   U2051 : AOI221_X1 port map( B1 => n46, B2 => regs(1230), C1 => n319, C2 => 
                           regs(2254), A => n1636, ZN => n1635);
   U2052 : INV_X1 port map( A => n1637, ZN => n1636);
   U2053 : AOI222_X1 port map( A1 => regs(206), A2 => n126, B1 => regs(1742), 
                           B2 => n180, C1 => regs(718), C2 => n255, ZN => n1637
                           );
   U2054 : INV_X1 port map( A => n1638, ZN => curr_proc_regs(718));
   U2055 : AOI221_X1 port map( B1 => n46, B2 => regs(1742), C1 => n319, C2 => 
                           regs(206), A => n1639, ZN => n1638);
   U2056 : INV_X1 port map( A => n1640, ZN => n1639);
   U2057 : AOI222_X1 port map( A1 => regs(718), A2 => n126, B1 => regs(2254), 
                           B2 => n180, C1 => regs(1230), C2 => n255, ZN => 
                           n1640);
   U2058 : INV_X1 port map( A => n1641, ZN => curr_proc_regs(205));
   U2059 : AOI221_X1 port map( B1 => n46, B2 => regs(1229), C1 => n319, C2 => 
                           regs(2253), A => n1642, ZN => n1641);
   U2060 : INV_X1 port map( A => n1643, ZN => n1642);
   U2061 : AOI222_X1 port map( A1 => regs(205), A2 => n126, B1 => regs(1741), 
                           B2 => n179, C1 => regs(717), C2 => n254, ZN => n1643
                           );
   U2062 : INV_X1 port map( A => n1644, ZN => curr_proc_regs(717));
   U2063 : AOI221_X1 port map( B1 => n46, B2 => regs(1741), C1 => n319, C2 => 
                           regs(205), A => n1645, ZN => n1644);
   U2064 : INV_X1 port map( A => n1646, ZN => n1645);
   U2065 : AOI222_X1 port map( A1 => regs(717), A2 => n127, B1 => regs(2253), 
                           B2 => n179, C1 => regs(1229), C2 => n254, ZN => 
                           n1646);
   U2066 : INV_X1 port map( A => n1647, ZN => curr_proc_regs(204));
   U2067 : AOI221_X1 port map( B1 => n46, B2 => regs(1228), C1 => n319, C2 => 
                           regs(2252), A => n1648, ZN => n1647);
   U2068 : INV_X1 port map( A => n1649, ZN => n1648);
   U2069 : AOI222_X1 port map( A1 => regs(204), A2 => n127, B1 => regs(1740), 
                           B2 => n179, C1 => regs(716), C2 => n254, ZN => n1649
                           );
   U2070 : INV_X1 port map( A => n1650, ZN => curr_proc_regs(716));
   U2071 : AOI221_X1 port map( B1 => n47, B2 => regs(1740), C1 => n319, C2 => 
                           regs(204), A => n1651, ZN => n1650);
   U2072 : INV_X1 port map( A => n1652, ZN => n1651);
   U2073 : AOI222_X1 port map( A1 => regs(716), A2 => n127, B1 => regs(2252), 
                           B2 => n179, C1 => regs(1228), C2 => n254, ZN => 
                           n1652);
   U2074 : INV_X1 port map( A => n1653, ZN => curr_proc_regs(203));
   U2075 : AOI221_X1 port map( B1 => n47, B2 => regs(1227), C1 => n319, C2 => 
                           regs(2251), A => n1654, ZN => n1653);
   U2076 : INV_X1 port map( A => n1655, ZN => n1654);
   U2077 : AOI222_X1 port map( A1 => regs(203), A2 => n127, B1 => regs(1739), 
                           B2 => n179, C1 => regs(715), C2 => n254, ZN => n1655
                           );
   U2078 : INV_X1 port map( A => n1656, ZN => curr_proc_regs(715));
   U2079 : AOI221_X1 port map( B1 => n47, B2 => regs(1739), C1 => n319, C2 => 
                           regs(203), A => n1657, ZN => n1656);
   U2080 : INV_X1 port map( A => n1658, ZN => n1657);
   U2081 : AOI222_X1 port map( A1 => regs(715), A2 => n127, B1 => regs(2251), 
                           B2 => n179, C1 => regs(1227), C2 => n254, ZN => 
                           n1658);
   U2082 : INV_X1 port map( A => n1659, ZN => curr_proc_regs(202));
   U2083 : AOI221_X1 port map( B1 => n47, B2 => regs(1226), C1 => n319, C2 => 
                           regs(2250), A => n1660, ZN => n1659);
   U2084 : INV_X1 port map( A => n1661, ZN => n1660);
   U2085 : AOI222_X1 port map( A1 => regs(202), A2 => n127, B1 => regs(1738), 
                           B2 => n179, C1 => regs(714), C2 => n254, ZN => n1661
                           );
   U2086 : INV_X1 port map( A => n1662, ZN => curr_proc_regs(714));
   U2087 : AOI221_X1 port map( B1 => n47, B2 => regs(1738), C1 => n318, C2 => 
                           regs(202), A => n1663, ZN => n1662);
   U2088 : INV_X1 port map( A => n1664, ZN => n1663);
   U2089 : AOI222_X1 port map( A1 => regs(714), A2 => n127, B1 => regs(2250), 
                           B2 => n179, C1 => regs(1226), C2 => n254, ZN => 
                           n1664);
   U2090 : INV_X1 port map( A => n1665, ZN => curr_proc_regs(201));
   U2091 : AOI221_X1 port map( B1 => n47, B2 => regs(1225), C1 => n318, C2 => 
                           regs(2249), A => n1666, ZN => n1665);
   U2092 : INV_X1 port map( A => n1667, ZN => n1666);
   U2093 : AOI222_X1 port map( A1 => regs(201), A2 => n127, B1 => regs(1737), 
                           B2 => n179, C1 => regs(713), C2 => n254, ZN => n1667
                           );
   U2094 : INV_X1 port map( A => n1668, ZN => curr_proc_regs(713));
   U2095 : AOI221_X1 port map( B1 => n47, B2 => regs(1737), C1 => n318, C2 => 
                           regs(201), A => n1669, ZN => n1668);
   U2096 : INV_X1 port map( A => n1670, ZN => n1669);
   U2097 : AOI222_X1 port map( A1 => regs(713), A2 => n127, B1 => regs(2249), 
                           B2 => n179, C1 => regs(1225), C2 => n254, ZN => 
                           n1670);
   U2098 : INV_X1 port map( A => n1671, ZN => curr_proc_regs(200));
   U2099 : AOI221_X1 port map( B1 => n47, B2 => regs(1224), C1 => n318, C2 => 
                           regs(2248), A => n1672, ZN => n1671);
   U2100 : INV_X1 port map( A => n1673, ZN => n1672);
   U2101 : AOI222_X1 port map( A1 => regs(200), A2 => n127, B1 => regs(1736), 
                           B2 => n179, C1 => regs(712), C2 => n254, ZN => n1673
                           );
   U2102 : INV_X1 port map( A => n1674, ZN => curr_proc_regs(712));
   U2103 : AOI221_X1 port map( B1 => n47, B2 => regs(1736), C1 => n318, C2 => 
                           regs(200), A => n1675, ZN => n1674);
   U2104 : INV_X1 port map( A => n1676, ZN => n1675);
   U2105 : AOI222_X1 port map( A1 => regs(712), A2 => n127, B1 => regs(2248), 
                           B2 => n179, C1 => regs(1224), C2 => n254, ZN => 
                           n1676);
   U2106 : INV_X1 port map( A => n1677, ZN => curr_proc_regs(199));
   U2107 : AOI221_X1 port map( B1 => n47, B2 => regs(1223), C1 => n318, C2 => 
                           regs(2247), A => n1678, ZN => n1677);
   U2108 : INV_X1 port map( A => n1679, ZN => n1678);
   U2109 : AOI222_X1 port map( A1 => regs(199), A2 => n127, B1 => regs(1735), 
                           B2 => n178, C1 => regs(711), C2 => n253, ZN => n1679
                           );
   U2110 : INV_X1 port map( A => n1680, ZN => curr_proc_regs(711));
   U2111 : AOI221_X1 port map( B1 => n47, B2 => regs(1735), C1 => n318, C2 => 
                           regs(199), A => n1681, ZN => n1680);
   U2112 : INV_X1 port map( A => n1682, ZN => n1681);
   U2113 : AOI222_X1 port map( A1 => regs(711), A2 => n128, B1 => regs(2247), 
                           B2 => n178, C1 => regs(1223), C2 => n253, ZN => 
                           n1682);
   U2114 : INV_X1 port map( A => n1683, ZN => curr_proc_regs(198));
   U2115 : AOI221_X1 port map( B1 => n47, B2 => regs(1222), C1 => n318, C2 => 
                           regs(2246), A => n1684, ZN => n1683);
   U2116 : INV_X1 port map( A => n1685, ZN => n1684);
   U2117 : AOI222_X1 port map( A1 => regs(198), A2 => n128, B1 => regs(1734), 
                           B2 => n178, C1 => regs(710), C2 => n253, ZN => n1685
                           );
   U2118 : INV_X1 port map( A => n1686, ZN => curr_proc_regs(710));
   U2119 : AOI221_X1 port map( B1 => n48, B2 => regs(1734), C1 => n318, C2 => 
                           regs(198), A => n1687, ZN => n1686);
   U2120 : INV_X1 port map( A => n1688, ZN => n1687);
   U2121 : AOI222_X1 port map( A1 => regs(710), A2 => n128, B1 => regs(2246), 
                           B2 => n178, C1 => regs(1222), C2 => n253, ZN => 
                           n1688);
   U2122 : INV_X1 port map( A => n1689, ZN => curr_proc_regs(197));
   U2123 : AOI221_X1 port map( B1 => n48, B2 => regs(1221), C1 => n318, C2 => 
                           regs(2245), A => n1690, ZN => n1689);
   U2124 : INV_X1 port map( A => n1691, ZN => n1690);
   U2125 : AOI222_X1 port map( A1 => regs(197), A2 => n128, B1 => regs(1733), 
                           B2 => n178, C1 => regs(709), C2 => n253, ZN => n1691
                           );
   U2126 : INV_X1 port map( A => n1692, ZN => curr_proc_regs(709));
   U2127 : AOI221_X1 port map( B1 => n48, B2 => regs(1733), C1 => n318, C2 => 
                           regs(197), A => n1693, ZN => n1692);
   U2128 : INV_X1 port map( A => n1694, ZN => n1693);
   U2129 : AOI222_X1 port map( A1 => regs(709), A2 => n128, B1 => regs(2245), 
                           B2 => n178, C1 => regs(1221), C2 => n253, ZN => 
                           n1694);
   U2130 : INV_X1 port map( A => n1695, ZN => curr_proc_regs(196));
   U2131 : AOI221_X1 port map( B1 => n48, B2 => regs(1220), C1 => n318, C2 => 
                           regs(2244), A => n1696, ZN => n1695);
   U2132 : INV_X1 port map( A => n1697, ZN => n1696);
   U2133 : AOI222_X1 port map( A1 => regs(196), A2 => n128, B1 => regs(1732), 
                           B2 => n178, C1 => regs(708), C2 => n253, ZN => n1697
                           );
   U2134 : INV_X1 port map( A => n1698, ZN => curr_proc_regs(708));
   U2135 : AOI221_X1 port map( B1 => n48, B2 => regs(1732), C1 => n317, C2 => 
                           regs(196), A => n1699, ZN => n1698);
   U2136 : INV_X1 port map( A => n1700, ZN => n1699);
   U2137 : AOI222_X1 port map( A1 => regs(708), A2 => n128, B1 => regs(2244), 
                           B2 => n178, C1 => regs(1220), C2 => n253, ZN => 
                           n1700);
   U2138 : INV_X1 port map( A => n1701, ZN => curr_proc_regs(195));
   U2139 : AOI221_X1 port map( B1 => n48, B2 => regs(1219), C1 => n317, C2 => 
                           regs(2243), A => n1702, ZN => n1701);
   U2140 : INV_X1 port map( A => n1703, ZN => n1702);
   U2141 : AOI222_X1 port map( A1 => regs(195), A2 => n128, B1 => regs(1731), 
                           B2 => n178, C1 => regs(707), C2 => n253, ZN => n1703
                           );
   U2142 : INV_X1 port map( A => n1704, ZN => curr_proc_regs(707));
   U2143 : AOI221_X1 port map( B1 => n48, B2 => regs(1731), C1 => n317, C2 => 
                           regs(195), A => n1705, ZN => n1704);
   U2144 : INV_X1 port map( A => n1706, ZN => n1705);
   U2145 : AOI222_X1 port map( A1 => regs(707), A2 => n128, B1 => regs(2243), 
                           B2 => n178, C1 => regs(1219), C2 => n253, ZN => 
                           n1706);
   U2146 : INV_X1 port map( A => n1707, ZN => curr_proc_regs(194));
   U2147 : AOI221_X1 port map( B1 => n48, B2 => regs(1218), C1 => n317, C2 => 
                           regs(2242), A => n1708, ZN => n1707);
   U2148 : INV_X1 port map( A => n1709, ZN => n1708);
   U2149 : AOI222_X1 port map( A1 => regs(194), A2 => n128, B1 => regs(1730), 
                           B2 => n178, C1 => regs(706), C2 => n253, ZN => n1709
                           );
   U2150 : INV_X1 port map( A => n1710, ZN => curr_proc_regs(706));
   U2151 : AOI221_X1 port map( B1 => n48, B2 => regs(1730), C1 => n317, C2 => 
                           regs(194), A => n1711, ZN => n1710);
   U2152 : INV_X1 port map( A => n1712, ZN => n1711);
   U2153 : AOI222_X1 port map( A1 => regs(706), A2 => n128, B1 => regs(2242), 
                           B2 => n178, C1 => regs(1218), C2 => n253, ZN => 
                           n1712);
   U2154 : INV_X1 port map( A => n1713, ZN => curr_proc_regs(193));
   U2155 : AOI221_X1 port map( B1 => n48, B2 => regs(1217), C1 => n317, C2 => 
                           regs(2241), A => n1714, ZN => n1713);
   U2156 : INV_X1 port map( A => n1715, ZN => n1714);
   U2157 : AOI222_X1 port map( A1 => regs(193), A2 => n128, B1 => regs(1729), 
                           B2 => n177, C1 => regs(705), C2 => n252, ZN => n1715
                           );
   U2158 : INV_X1 port map( A => n1716, ZN => curr_proc_regs(705));
   U2159 : AOI221_X1 port map( B1 => n48, B2 => regs(1729), C1 => n317, C2 => 
                           regs(193), A => n1717, ZN => n1716);
   U2160 : INV_X1 port map( A => n1718, ZN => n1717);
   U2161 : AOI222_X1 port map( A1 => regs(705), A2 => n129, B1 => regs(2241), 
                           B2 => n177, C1 => regs(1217), C2 => n252, ZN => 
                           n1718);
   U2162 : INV_X1 port map( A => n1719, ZN => curr_proc_regs(192));
   U2163 : AOI221_X1 port map( B1 => n48, B2 => regs(1216), C1 => n317, C2 => 
                           regs(2240), A => n1720, ZN => n1719);
   U2164 : INV_X1 port map( A => n1721, ZN => n1720);
   U2165 : AOI222_X1 port map( A1 => regs(192), A2 => n129, B1 => regs(1728), 
                           B2 => n177, C1 => regs(704), C2 => n252, ZN => n1721
                           );
   U2166 : INV_X1 port map( A => n1722, ZN => curr_proc_regs(704));
   U2167 : AOI221_X1 port map( B1 => n49, B2 => regs(1728), C1 => n317, C2 => 
                           regs(192), A => n1723, ZN => n1722);
   U2168 : INV_X1 port map( A => n1724, ZN => n1723);
   U2169 : AOI222_X1 port map( A1 => regs(704), A2 => n129, B1 => regs(2240), 
                           B2 => n177, C1 => regs(1216), C2 => n252, ZN => 
                           n1724);
   U2170 : INV_X1 port map( A => n1725, ZN => curr_proc_regs(255));
   U2171 : AOI221_X1 port map( B1 => n49, B2 => regs(1279), C1 => n317, C2 => 
                           regs(2303), A => n1726, ZN => n1725);
   U2172 : INV_X1 port map( A => n1727, ZN => n1726);
   U2173 : AOI222_X1 port map( A1 => regs(255), A2 => n129, B1 => regs(1791), 
                           B2 => n177, C1 => regs(767), C2 => n252, ZN => n1727
                           );
   U2174 : INV_X1 port map( A => n1728, ZN => curr_proc_regs(767));
   U2175 : AOI221_X1 port map( B1 => n49, B2 => regs(1791), C1 => n317, C2 => 
                           regs(255), A => n1729, ZN => n1728);
   U2176 : INV_X1 port map( A => n1730, ZN => n1729);
   U2177 : AOI222_X1 port map( A1 => regs(767), A2 => n129, B1 => regs(2303), 
                           B2 => n177, C1 => regs(1279), C2 => n252, ZN => 
                           n1730);
   U2178 : INV_X1 port map( A => n1731, ZN => curr_proc_regs(254));
   U2179 : AOI221_X1 port map( B1 => n49, B2 => regs(1278), C1 => n316, C2 => 
                           regs(2302), A => n1732, ZN => n1731);
   U2180 : INV_X1 port map( A => n1733, ZN => n1732);
   U2181 : AOI222_X1 port map( A1 => regs(254), A2 => n129, B1 => regs(1790), 
                           B2 => n177, C1 => regs(766), C2 => n252, ZN => n1733
                           );
   U2182 : INV_X1 port map( A => n1734, ZN => curr_proc_regs(766));
   U2183 : AOI221_X1 port map( B1 => n49, B2 => regs(1790), C1 => n316, C2 => 
                           regs(254), A => n1735, ZN => n1734);
   U2184 : INV_X1 port map( A => n1736, ZN => n1735);
   U2185 : AOI222_X1 port map( A1 => regs(766), A2 => n129, B1 => regs(2302), 
                           B2 => n177, C1 => regs(1278), C2 => n252, ZN => 
                           n1736);
   U2186 : INV_X1 port map( A => n1737, ZN => curr_proc_regs(253));
   U2187 : AOI221_X1 port map( B1 => n49, B2 => regs(1277), C1 => n316, C2 => 
                           regs(2301), A => n1738, ZN => n1737);
   U2188 : INV_X1 port map( A => n1739, ZN => n1738);
   U2189 : AOI222_X1 port map( A1 => regs(253), A2 => n129, B1 => regs(1789), 
                           B2 => n177, C1 => regs(765), C2 => n252, ZN => n1739
                           );
   U2190 : INV_X1 port map( A => n1740, ZN => curr_proc_regs(765));
   U2191 : AOI221_X1 port map( B1 => n49, B2 => regs(1789), C1 => n316, C2 => 
                           regs(253), A => n1741, ZN => n1740);
   U2192 : INV_X1 port map( A => n1742, ZN => n1741);
   U2193 : AOI222_X1 port map( A1 => regs(765), A2 => n129, B1 => regs(2301), 
                           B2 => n177, C1 => regs(1277), C2 => n252, ZN => 
                           n1742);
   U2194 : INV_X1 port map( A => n1743, ZN => curr_proc_regs(252));
   U2195 : AOI221_X1 port map( B1 => n49, B2 => regs(1276), C1 => n316, C2 => 
                           regs(2300), A => n1744, ZN => n1743);
   U2196 : INV_X1 port map( A => n1745, ZN => n1744);
   U2197 : AOI222_X1 port map( A1 => regs(252), A2 => n129, B1 => regs(1788), 
                           B2 => n177, C1 => regs(764), C2 => n252, ZN => n1745
                           );
   U2198 : INV_X1 port map( A => n1746, ZN => curr_proc_regs(764));
   U2199 : AOI221_X1 port map( B1 => n49, B2 => regs(1788), C1 => n316, C2 => 
                           regs(252), A => n1747, ZN => n1746);
   U2200 : INV_X1 port map( A => n1748, ZN => n1747);
   U2201 : AOI222_X1 port map( A1 => regs(764), A2 => n129, B1 => regs(2300), 
                           B2 => n177, C1 => regs(1276), C2 => n252, ZN => 
                           n1748);
   U2202 : INV_X1 port map( A => n1749, ZN => curr_proc_regs(251));
   U2203 : AOI221_X1 port map( B1 => n49, B2 => regs(1275), C1 => n316, C2 => 
                           regs(2299), A => n1750, ZN => n1749);
   U2204 : INV_X1 port map( A => n1751, ZN => n1750);
   U2205 : AOI222_X1 port map( A1 => regs(251), A2 => n129, B1 => regs(1787), 
                           B2 => n176, C1 => regs(763), C2 => n251, ZN => n1751
                           );
   U2206 : INV_X1 port map( A => n1752, ZN => curr_proc_regs(763));
   U2207 : AOI221_X1 port map( B1 => n49, B2 => regs(1787), C1 => n316, C2 => 
                           regs(251), A => n1753, ZN => n1752);
   U2208 : INV_X1 port map( A => n1754, ZN => n1753);
   U2209 : AOI222_X1 port map( A1 => regs(763), A2 => n130, B1 => regs(2299), 
                           B2 => n176, C1 => regs(1275), C2 => n251, ZN => 
                           n1754);
   U2210 : INV_X1 port map( A => n1755, ZN => curr_proc_regs(250));
   U2211 : AOI221_X1 port map( B1 => n50, B2 => regs(1274), C1 => n316, C2 => 
                           regs(2298), A => n1756, ZN => n1755);
   U2212 : INV_X1 port map( A => n1757, ZN => n1756);
   U2213 : AOI222_X1 port map( A1 => regs(250), A2 => n130, B1 => regs(1786), 
                           B2 => n176, C1 => regs(762), C2 => n251, ZN => n1757
                           );
   U2214 : INV_X1 port map( A => n1758, ZN => curr_proc_regs(762));
   U2215 : AOI221_X1 port map( B1 => n50, B2 => regs(1786), C1 => n316, C2 => 
                           regs(250), A => n1759, ZN => n1758);
   U2216 : INV_X1 port map( A => n1760, ZN => n1759);
   U2217 : AOI222_X1 port map( A1 => regs(762), A2 => n130, B1 => regs(2298), 
                           B2 => n176, C1 => regs(1274), C2 => n251, ZN => 
                           n1760);
   U2218 : INV_X1 port map( A => n1761, ZN => curr_proc_regs(249));
   U2219 : AOI221_X1 port map( B1 => n50, B2 => regs(1273), C1 => n316, C2 => 
                           regs(2297), A => n1762, ZN => n1761);
   U2220 : INV_X1 port map( A => n1763, ZN => n1762);
   U2221 : AOI222_X1 port map( A1 => regs(249), A2 => n130, B1 => regs(1785), 
                           B2 => n176, C1 => regs(761), C2 => n251, ZN => n1763
                           );
   U2222 : INV_X1 port map( A => n1764, ZN => curr_proc_regs(761));
   U2223 : AOI221_X1 port map( B1 => n50, B2 => regs(1785), C1 => n316, C2 => 
                           regs(249), A => n1765, ZN => n1764);
   U2224 : INV_X1 port map( A => n1766, ZN => n1765);
   U2225 : AOI222_X1 port map( A1 => regs(761), A2 => n130, B1 => regs(2297), 
                           B2 => n176, C1 => regs(1273), C2 => n251, ZN => 
                           n1766);
   U2226 : INV_X1 port map( A => n1767, ZN => curr_proc_regs(248));
   U2227 : AOI221_X1 port map( B1 => n50, B2 => regs(1272), C1 => n315, C2 => 
                           regs(2296), A => n1768, ZN => n1767);
   U2228 : INV_X1 port map( A => n1769, ZN => n1768);
   U2229 : AOI222_X1 port map( A1 => regs(248), A2 => n130, B1 => regs(1784), 
                           B2 => n176, C1 => regs(760), C2 => n251, ZN => n1769
                           );
   U2230 : INV_X1 port map( A => n1770, ZN => curr_proc_regs(760));
   U2231 : AOI221_X1 port map( B1 => n50, B2 => regs(1784), C1 => n315, C2 => 
                           regs(248), A => n1771, ZN => n1770);
   U2232 : INV_X1 port map( A => n1772, ZN => n1771);
   U2233 : AOI222_X1 port map( A1 => regs(760), A2 => n130, B1 => regs(2296), 
                           B2 => n176, C1 => regs(1272), C2 => n251, ZN => 
                           n1772);
   U2234 : INV_X1 port map( A => n1773, ZN => curr_proc_regs(247));
   U2235 : AOI221_X1 port map( B1 => n50, B2 => regs(1271), C1 => n315, C2 => 
                           regs(2295), A => n1774, ZN => n1773);
   U2236 : INV_X1 port map( A => n1775, ZN => n1774);
   U2237 : AOI222_X1 port map( A1 => regs(247), A2 => n130, B1 => regs(1783), 
                           B2 => n176, C1 => regs(759), C2 => n251, ZN => n1775
                           );
   U2238 : INV_X1 port map( A => n1776, ZN => curr_proc_regs(759));
   U2239 : AOI221_X1 port map( B1 => n50, B2 => regs(1783), C1 => n315, C2 => 
                           regs(247), A => n1777, ZN => n1776);
   U2240 : INV_X1 port map( A => n1778, ZN => n1777);
   U2241 : AOI222_X1 port map( A1 => regs(759), A2 => n130, B1 => regs(2295), 
                           B2 => n176, C1 => regs(1271), C2 => n251, ZN => 
                           n1778);
   U2242 : INV_X1 port map( A => n1779, ZN => curr_proc_regs(246));
   U2243 : AOI221_X1 port map( B1 => n50, B2 => regs(1270), C1 => n315, C2 => 
                           regs(2294), A => n1780, ZN => n1779);
   U2244 : INV_X1 port map( A => n1781, ZN => n1780);
   U2245 : AOI222_X1 port map( A1 => regs(246), A2 => n130, B1 => regs(1782), 
                           B2 => n176, C1 => regs(758), C2 => n251, ZN => n1781
                           );
   U2246 : INV_X1 port map( A => n1782, ZN => curr_proc_regs(758));
   U2247 : AOI221_X1 port map( B1 => n50, B2 => regs(1782), C1 => n315, C2 => 
                           regs(246), A => n1783, ZN => n1782);
   U2248 : INV_X1 port map( A => n1784, ZN => n1783);
   U2249 : AOI222_X1 port map( A1 => regs(758), A2 => n130, B1 => regs(2294), 
                           B2 => n176, C1 => regs(1270), C2 => n251, ZN => 
                           n1784);
   U2250 : INV_X1 port map( A => n1785, ZN => curr_proc_regs(245));
   U2251 : AOI221_X1 port map( B1 => n50, B2 => regs(1269), C1 => n315, C2 => 
                           regs(2293), A => n1786, ZN => n1785);
   U2252 : INV_X1 port map( A => n1787, ZN => n1786);
   U2253 : AOI222_X1 port map( A1 => regs(245), A2 => n130, B1 => regs(1781), 
                           B2 => n175, C1 => regs(757), C2 => n250, ZN => n1787
                           );
   U2254 : INV_X1 port map( A => n1788, ZN => curr_proc_regs(757));
   U2255 : AOI221_X1 port map( B1 => n50, B2 => regs(1781), C1 => n315, C2 => 
                           regs(245), A => n1789, ZN => n1788);
   U2256 : INV_X1 port map( A => n1790, ZN => n1789);
   U2257 : AOI222_X1 port map( A1 => regs(757), A2 => n131, B1 => regs(2293), 
                           B2 => n175, C1 => regs(1269), C2 => n250, ZN => 
                           n1790);
   U2258 : INV_X1 port map( A => n1791, ZN => curr_proc_regs(244));
   U2259 : AOI221_X1 port map( B1 => n51, B2 => regs(1268), C1 => n315, C2 => 
                           regs(2292), A => n1792, ZN => n1791);
   U2260 : INV_X1 port map( A => n1793, ZN => n1792);
   U2261 : AOI222_X1 port map( A1 => regs(244), A2 => n131, B1 => regs(1780), 
                           B2 => n175, C1 => regs(756), C2 => n250, ZN => n1793
                           );
   U2262 : INV_X1 port map( A => n1794, ZN => curr_proc_regs(756));
   U2263 : AOI221_X1 port map( B1 => n51, B2 => regs(1780), C1 => n315, C2 => 
                           regs(244), A => n1795, ZN => n1794);
   U2264 : INV_X1 port map( A => n1796, ZN => n1795);
   U2265 : AOI222_X1 port map( A1 => regs(756), A2 => n131, B1 => regs(2292), 
                           B2 => n175, C1 => regs(1268), C2 => n250, ZN => 
                           n1796);
   U2266 : INV_X1 port map( A => n1797, ZN => curr_proc_regs(243));
   U2267 : AOI221_X1 port map( B1 => n51, B2 => regs(1267), C1 => n315, C2 => 
                           regs(2291), A => n1798, ZN => n1797);
   U2268 : INV_X1 port map( A => n1799, ZN => n1798);
   U2269 : AOI222_X1 port map( A1 => regs(243), A2 => n131, B1 => regs(1779), 
                           B2 => n175, C1 => regs(755), C2 => n250, ZN => n1799
                           );
   U2270 : INV_X1 port map( A => n1800, ZN => curr_proc_regs(755));
   U2271 : AOI221_X1 port map( B1 => n51, B2 => regs(1779), C1 => n315, C2 => 
                           regs(243), A => n1801, ZN => n1800);
   U2272 : INV_X1 port map( A => n1802, ZN => n1801);
   U2273 : AOI222_X1 port map( A1 => regs(755), A2 => n131, B1 => regs(2291), 
                           B2 => n175, C1 => regs(1267), C2 => n250, ZN => 
                           n1802);
   U2274 : INV_X1 port map( A => n1803, ZN => curr_proc_regs(242));
   U2275 : AOI221_X1 port map( B1 => n51, B2 => regs(1266), C1 => n314, C2 => 
                           regs(2290), A => n1804, ZN => n1803);
   U2276 : INV_X1 port map( A => n1805, ZN => n1804);
   U2277 : AOI222_X1 port map( A1 => regs(242), A2 => n131, B1 => regs(1778), 
                           B2 => n175, C1 => regs(754), C2 => n250, ZN => n1805
                           );
   U2278 : INV_X1 port map( A => n1806, ZN => curr_proc_regs(754));
   U2279 : AOI221_X1 port map( B1 => n51, B2 => regs(1778), C1 => n314, C2 => 
                           regs(242), A => n1807, ZN => n1806);
   U2280 : INV_X1 port map( A => n1808, ZN => n1807);
   U2281 : AOI222_X1 port map( A1 => regs(754), A2 => n131, B1 => regs(2290), 
                           B2 => n175, C1 => regs(1266), C2 => n250, ZN => 
                           n1808);
   U2282 : INV_X1 port map( A => n1809, ZN => curr_proc_regs(241));
   U2283 : AOI221_X1 port map( B1 => n51, B2 => regs(1265), C1 => n314, C2 => 
                           regs(2289), A => n1810, ZN => n1809);
   U2284 : INV_X1 port map( A => n1811, ZN => n1810);
   U2285 : AOI222_X1 port map( A1 => regs(241), A2 => n131, B1 => regs(1777), 
                           B2 => n175, C1 => regs(753), C2 => n250, ZN => n1811
                           );
   U2286 : INV_X1 port map( A => n1812, ZN => curr_proc_regs(753));
   U2287 : AOI221_X1 port map( B1 => n51, B2 => regs(1777), C1 => n314, C2 => 
                           regs(241), A => n1813, ZN => n1812);
   U2288 : INV_X1 port map( A => n1814, ZN => n1813);
   U2289 : AOI222_X1 port map( A1 => regs(753), A2 => n131, B1 => regs(2289), 
                           B2 => n175, C1 => regs(1265), C2 => n250, ZN => 
                           n1814);
   U2290 : INV_X1 port map( A => n1815, ZN => curr_proc_regs(240));
   U2291 : AOI221_X1 port map( B1 => n51, B2 => regs(1264), C1 => n314, C2 => 
                           regs(2288), A => n1816, ZN => n1815);
   U2292 : INV_X1 port map( A => n1817, ZN => n1816);
   U2293 : AOI222_X1 port map( A1 => regs(240), A2 => n131, B1 => regs(1776), 
                           B2 => n175, C1 => regs(752), C2 => n250, ZN => n1817
                           );
   U2294 : INV_X1 port map( A => n1818, ZN => curr_proc_regs(752));
   U2295 : AOI221_X1 port map( B1 => n51, B2 => regs(1776), C1 => n314, C2 => 
                           regs(240), A => n1819, ZN => n1818);
   U2296 : INV_X1 port map( A => n1820, ZN => n1819);
   U2297 : AOI222_X1 port map( A1 => regs(752), A2 => n131, B1 => regs(2288), 
                           B2 => n175, C1 => regs(1264), C2 => n250, ZN => 
                           n1820);
   U2298 : INV_X1 port map( A => n1821, ZN => curr_proc_regs(239));
   U2299 : AOI221_X1 port map( B1 => n51, B2 => regs(1263), C1 => n314, C2 => 
                           regs(2287), A => n1822, ZN => n1821);
   U2300 : INV_X1 port map( A => n1823, ZN => n1822);
   U2301 : AOI222_X1 port map( A1 => regs(239), A2 => n132, B1 => regs(1775), 
                           B2 => n174, C1 => regs(751), C2 => n249, ZN => n1823
                           );
   U2302 : INV_X1 port map( A => n1824, ZN => curr_proc_regs(751));
   U2303 : AOI221_X1 port map( B1 => n51, B2 => regs(1775), C1 => n314, C2 => 
                           regs(239), A => n1825, ZN => n1824);
   U2304 : INV_X1 port map( A => n1826, ZN => n1825);
   U2305 : AOI222_X1 port map( A1 => regs(751), A2 => n132, B1 => regs(2287), 
                           B2 => n174, C1 => regs(1263), C2 => n249, ZN => 
                           n1826);
   U2306 : INV_X1 port map( A => n1827, ZN => curr_proc_regs(238));
   U2307 : AOI221_X1 port map( B1 => n52, B2 => regs(1262), C1 => n314, C2 => 
                           regs(2286), A => n1828, ZN => n1827);
   U2308 : INV_X1 port map( A => n1829, ZN => n1828);
   U2309 : AOI222_X1 port map( A1 => regs(238), A2 => n132, B1 => regs(1774), 
                           B2 => n174, C1 => regs(750), C2 => n249, ZN => n1829
                           );
   U2310 : INV_X1 port map( A => n1830, ZN => curr_proc_regs(750));
   U2311 : AOI221_X1 port map( B1 => n52, B2 => regs(1774), C1 => n314, C2 => 
                           regs(238), A => n1831, ZN => n1830);
   U2312 : INV_X1 port map( A => n1832, ZN => n1831);
   U2313 : AOI222_X1 port map( A1 => regs(750), A2 => n132, B1 => regs(2286), 
                           B2 => n174, C1 => regs(1262), C2 => n249, ZN => 
                           n1832);
   U2314 : INV_X1 port map( A => n1833, ZN => curr_proc_regs(237));
   U2315 : AOI221_X1 port map( B1 => n52, B2 => regs(1261), C1 => n314, C2 => 
                           regs(2285), A => n1834, ZN => n1833);
   U2316 : INV_X1 port map( A => n1835, ZN => n1834);
   U2317 : AOI222_X1 port map( A1 => regs(237), A2 => n132, B1 => regs(1773), 
                           B2 => n174, C1 => regs(749), C2 => n249, ZN => n1835
                           );
   U2318 : INV_X1 port map( A => n1836, ZN => curr_proc_regs(749));
   U2319 : AOI221_X1 port map( B1 => n52, B2 => regs(1773), C1 => n314, C2 => 
                           regs(237), A => n1837, ZN => n1836);
   U2320 : INV_X1 port map( A => n1838, ZN => n1837);
   U2321 : AOI222_X1 port map( A1 => regs(749), A2 => n132, B1 => regs(2285), 
                           B2 => n174, C1 => regs(1261), C2 => n249, ZN => 
                           n1838);
   U2322 : INV_X1 port map( A => n1839, ZN => curr_proc_regs(236));
   U2323 : AOI221_X1 port map( B1 => n52, B2 => regs(1260), C1 => n313, C2 => 
                           regs(2284), A => n1840, ZN => n1839);
   U2324 : INV_X1 port map( A => n1841, ZN => n1840);
   U2325 : AOI222_X1 port map( A1 => regs(236), A2 => n132, B1 => regs(1772), 
                           B2 => n174, C1 => regs(748), C2 => n249, ZN => n1841
                           );
   U2326 : INV_X1 port map( A => n1842, ZN => curr_proc_regs(748));
   U2327 : AOI221_X1 port map( B1 => n52, B2 => regs(1772), C1 => n313, C2 => 
                           regs(236), A => n1843, ZN => n1842);
   U2328 : INV_X1 port map( A => n1844, ZN => n1843);
   U2329 : AOI222_X1 port map( A1 => regs(748), A2 => n132, B1 => regs(2284), 
                           B2 => n174, C1 => regs(1260), C2 => n249, ZN => 
                           n1844);
   U2330 : INV_X1 port map( A => n1845, ZN => curr_proc_regs(235));
   U2331 : AOI221_X1 port map( B1 => n52, B2 => regs(1259), C1 => n313, C2 => 
                           regs(2283), A => n1846, ZN => n1845);
   U2332 : INV_X1 port map( A => n1847, ZN => n1846);
   U2333 : AOI222_X1 port map( A1 => regs(235), A2 => n132, B1 => regs(1771), 
                           B2 => n174, C1 => regs(747), C2 => n249, ZN => n1847
                           );
   U2334 : INV_X1 port map( A => n1848, ZN => curr_proc_regs(747));
   U2335 : AOI221_X1 port map( B1 => n52, B2 => regs(1771), C1 => n313, C2 => 
                           regs(235), A => n1849, ZN => n1848);
   U2336 : INV_X1 port map( A => n1850, ZN => n1849);
   U2337 : AOI222_X1 port map( A1 => regs(747), A2 => n132, B1 => regs(2283), 
                           B2 => n174, C1 => regs(1259), C2 => n249, ZN => 
                           n1850);
   U2338 : INV_X1 port map( A => n1851, ZN => curr_proc_regs(234));
   U2339 : AOI221_X1 port map( B1 => n52, B2 => regs(1258), C1 => n313, C2 => 
                           regs(2282), A => n1852, ZN => n1851);
   U2340 : INV_X1 port map( A => n1853, ZN => n1852);
   U2341 : AOI222_X1 port map( A1 => regs(234), A2 => n132, B1 => regs(1770), 
                           B2 => n174, C1 => regs(746), C2 => n249, ZN => n1853
                           );
   U2342 : INV_X1 port map( A => n1854, ZN => curr_proc_regs(746));
   U2343 : AOI221_X1 port map( B1 => n52, B2 => regs(1770), C1 => n313, C2 => 
                           regs(234), A => n1855, ZN => n1854);
   U2344 : INV_X1 port map( A => n1856, ZN => n1855);
   U2345 : AOI222_X1 port map( A1 => regs(746), A2 => n132, B1 => regs(2282), 
                           B2 => n174, C1 => regs(1258), C2 => n249, ZN => 
                           n1856);
   U2346 : INV_X1 port map( A => n1857, ZN => curr_proc_regs(233));
   U2347 : AOI221_X1 port map( B1 => n52, B2 => regs(1257), C1 => n313, C2 => 
                           regs(2281), A => n1858, ZN => n1857);
   U2348 : INV_X1 port map( A => n1859, ZN => n1858);
   U2349 : AOI222_X1 port map( A1 => regs(233), A2 => n133, B1 => regs(1769), 
                           B2 => n173, C1 => regs(745), C2 => n248, ZN => n1859
                           );
   U2350 : INV_X1 port map( A => n1860, ZN => curr_proc_regs(745));
   U2351 : AOI221_X1 port map( B1 => n52, B2 => regs(1769), C1 => n313, C2 => 
                           regs(233), A => n1861, ZN => n1860);
   U2352 : INV_X1 port map( A => n1862, ZN => n1861);
   U2353 : AOI222_X1 port map( A1 => regs(745), A2 => n133, B1 => regs(2281), 
                           B2 => n173, C1 => regs(1257), C2 => n248, ZN => 
                           n1862);
   U2354 : INV_X1 port map( A => n1863, ZN => curr_proc_regs(232));
   U2355 : AOI221_X1 port map( B1 => n53, B2 => regs(1256), C1 => n313, C2 => 
                           regs(2280), A => n1864, ZN => n1863);
   U2356 : INV_X1 port map( A => n1865, ZN => n1864);
   U2357 : AOI222_X1 port map( A1 => regs(232), A2 => n133, B1 => regs(1768), 
                           B2 => n173, C1 => regs(744), C2 => n248, ZN => n1865
                           );
   U2358 : INV_X1 port map( A => n1866, ZN => curr_proc_regs(744));
   U2359 : AOI221_X1 port map( B1 => n53, B2 => regs(1768), C1 => n313, C2 => 
                           regs(232), A => n1867, ZN => n1866);
   U2360 : INV_X1 port map( A => n1868, ZN => n1867);
   U2361 : AOI222_X1 port map( A1 => regs(744), A2 => n133, B1 => regs(2280), 
                           B2 => n173, C1 => regs(1256), C2 => n248, ZN => 
                           n1868);
   U2362 : INV_X1 port map( A => n1869, ZN => curr_proc_regs(231));
   U2363 : AOI221_X1 port map( B1 => n53, B2 => regs(1255), C1 => n313, C2 => 
                           regs(2279), A => n1870, ZN => n1869);
   U2364 : INV_X1 port map( A => n1871, ZN => n1870);
   U2365 : AOI222_X1 port map( A1 => regs(231), A2 => n133, B1 => regs(1767), 
                           B2 => n173, C1 => regs(743), C2 => n248, ZN => n1871
                           );
   U2366 : INV_X1 port map( A => n1872, ZN => curr_proc_regs(743));
   U2367 : AOI221_X1 port map( B1 => n53, B2 => regs(1767), C1 => n313, C2 => 
                           regs(231), A => n1873, ZN => n1872);
   U2368 : INV_X1 port map( A => n1874, ZN => n1873);
   U2369 : AOI222_X1 port map( A1 => regs(743), A2 => n133, B1 => regs(2279), 
                           B2 => n173, C1 => regs(1255), C2 => n248, ZN => 
                           n1874);
   U2370 : INV_X1 port map( A => n1875, ZN => curr_proc_regs(230));
   U2371 : AOI221_X1 port map( B1 => n53, B2 => regs(1254), C1 => n312, C2 => 
                           regs(2278), A => n1876, ZN => n1875);
   U2372 : INV_X1 port map( A => n1877, ZN => n1876);
   U2373 : AOI222_X1 port map( A1 => regs(230), A2 => n133, B1 => regs(1766), 
                           B2 => n173, C1 => regs(742), C2 => n248, ZN => n1877
                           );
   U2374 : INV_X1 port map( A => n1878, ZN => curr_proc_regs(742));
   U2375 : AOI221_X1 port map( B1 => n53, B2 => regs(1766), C1 => n312, C2 => 
                           regs(230), A => n1879, ZN => n1878);
   U2376 : INV_X1 port map( A => n1880, ZN => n1879);
   U2377 : AOI222_X1 port map( A1 => regs(742), A2 => n133, B1 => regs(2278), 
                           B2 => n173, C1 => regs(1254), C2 => n248, ZN => 
                           n1880);
   U2378 : INV_X1 port map( A => n1881, ZN => curr_proc_regs(229));
   U2379 : AOI221_X1 port map( B1 => n53, B2 => regs(1253), C1 => n312, C2 => 
                           regs(2277), A => n1882, ZN => n1881);
   U2380 : INV_X1 port map( A => n1883, ZN => n1882);
   U2381 : AOI222_X1 port map( A1 => regs(229), A2 => n133, B1 => regs(1765), 
                           B2 => n173, C1 => regs(741), C2 => n248, ZN => n1883
                           );
   U2382 : INV_X1 port map( A => n1884, ZN => curr_proc_regs(741));
   U2383 : AOI221_X1 port map( B1 => n53, B2 => regs(1765), C1 => n312, C2 => 
                           regs(229), A => n1885, ZN => n1884);
   U2384 : INV_X1 port map( A => n1886, ZN => n1885);
   U2385 : AOI222_X1 port map( A1 => regs(741), A2 => n133, B1 => regs(2277), 
                           B2 => n173, C1 => regs(1253), C2 => n248, ZN => 
                           n1886);
   U2386 : INV_X1 port map( A => n1887, ZN => curr_proc_regs(228));
   U2387 : AOI221_X1 port map( B1 => n53, B2 => regs(1252), C1 => n312, C2 => 
                           regs(2276), A => n1888, ZN => n1887);
   U2388 : INV_X1 port map( A => n1889, ZN => n1888);
   U2389 : AOI222_X1 port map( A1 => regs(228), A2 => n133, B1 => regs(1764), 
                           B2 => n173, C1 => regs(740), C2 => n248, ZN => n1889
                           );
   U2390 : INV_X1 port map( A => n1890, ZN => curr_proc_regs(740));
   U2391 : AOI221_X1 port map( B1 => n53, B2 => regs(1764), C1 => n312, C2 => 
                           regs(228), A => n1891, ZN => n1890);
   U2392 : INV_X1 port map( A => n1892, ZN => n1891);
   U2393 : AOI222_X1 port map( A1 => regs(740), A2 => n133, B1 => regs(2276), 
                           B2 => n173, C1 => regs(1252), C2 => n248, ZN => 
                           n1892);
   U2394 : INV_X1 port map( A => n1893, ZN => curr_proc_regs(227));
   U2395 : AOI221_X1 port map( B1 => n53, B2 => regs(1251), C1 => n312, C2 => 
                           regs(2275), A => n1894, ZN => n1893);
   U2396 : INV_X1 port map( A => n1895, ZN => n1894);
   U2397 : AOI222_X1 port map( A1 => regs(227), A2 => n134, B1 => regs(1763), 
                           B2 => n172, C1 => regs(739), C2 => n247, ZN => n1895
                           );
   U2398 : INV_X1 port map( A => n1896, ZN => curr_proc_regs(739));
   U2399 : AOI221_X1 port map( B1 => n53, B2 => regs(1763), C1 => n312, C2 => 
                           regs(227), A => n1897, ZN => n1896);
   U2400 : INV_X1 port map( A => n1898, ZN => n1897);
   U2401 : AOI222_X1 port map( A1 => regs(739), A2 => n134, B1 => regs(2275), 
                           B2 => n172, C1 => regs(1251), C2 => n247, ZN => 
                           n1898);
   U2402 : INV_X1 port map( A => n1899, ZN => curr_proc_regs(226));
   U2403 : AOI221_X1 port map( B1 => n54, B2 => regs(1250), C1 => n312, C2 => 
                           regs(2274), A => n1900, ZN => n1899);
   U2404 : INV_X1 port map( A => n1901, ZN => n1900);
   U2405 : AOI222_X1 port map( A1 => regs(226), A2 => n134, B1 => regs(1762), 
                           B2 => n172, C1 => regs(738), C2 => n247, ZN => n1901
                           );
   U2406 : INV_X1 port map( A => n1902, ZN => curr_proc_regs(738));
   U2407 : AOI221_X1 port map( B1 => n54, B2 => regs(1762), C1 => n312, C2 => 
                           regs(226), A => n1903, ZN => n1902);
   U2408 : INV_X1 port map( A => n1904, ZN => n1903);
   U2409 : AOI222_X1 port map( A1 => regs(738), A2 => n134, B1 => regs(2274), 
                           B2 => n172, C1 => regs(1250), C2 => n247, ZN => 
                           n1904);
   U2410 : INV_X1 port map( A => n1905, ZN => curr_proc_regs(225));
   U2411 : AOI221_X1 port map( B1 => n54, B2 => regs(1249), C1 => n312, C2 => 
                           regs(2273), A => n1906, ZN => n1905);
   U2412 : INV_X1 port map( A => n1907, ZN => n1906);
   U2413 : AOI222_X1 port map( A1 => regs(225), A2 => n134, B1 => regs(1761), 
                           B2 => n172, C1 => regs(737), C2 => n247, ZN => n1907
                           );
   U2414 : INV_X1 port map( A => n1908, ZN => curr_proc_regs(737));
   U2415 : AOI221_X1 port map( B1 => n54, B2 => regs(1761), C1 => n312, C2 => 
                           regs(225), A => n1909, ZN => n1908);
   U2416 : INV_X1 port map( A => n1910, ZN => n1909);
   U2417 : AOI222_X1 port map( A1 => regs(737), A2 => n134, B1 => regs(2273), 
                           B2 => n172, C1 => regs(1249), C2 => n247, ZN => 
                           n1910);
   U2418 : INV_X1 port map( A => n1911, ZN => curr_proc_regs(224));
   U2419 : AOI221_X1 port map( B1 => n54, B2 => regs(1248), C1 => n311, C2 => 
                           regs(2272), A => n1912, ZN => n1911);
   U2420 : INV_X1 port map( A => n1913, ZN => n1912);
   U2421 : AOI222_X1 port map( A1 => regs(224), A2 => n134, B1 => regs(1760), 
                           B2 => n172, C1 => regs(736), C2 => n247, ZN => n1913
                           );
   U2422 : INV_X1 port map( A => n1914, ZN => curr_proc_regs(736));
   U2423 : AOI221_X1 port map( B1 => n22, B2 => regs(1760), C1 => n317, C2 => 
                           regs(224), A => n1915, ZN => n1914);
   U2424 : INV_X1 port map( A => n1916, ZN => n1915);
   U2425 : AOI222_X1 port map( A1 => regs(736), A2 => n134, B1 => regs(2272), 
                           B2 => n172, C1 => regs(1248), C2 => n247, ZN => 
                           n1916);
   U2426 : NAND2_X1 port map( A1 => n1917, A2 => n1918, ZN => 
                           curr_proc_regs(511));
   U2427 : AOI222_X1 port map( A1 => regs(511), A2 => n134, B1 => regs(2047), 
                           B2 => n172, C1 => regs(1023), C2 => n247, ZN => 
                           n1918);
   U2428 : AOI22_X1 port map( A1 => regs(1535), A2 => n1, B1 => regs(2559), B2 
                           => n343, ZN => n1917);
   U2429 : NAND2_X1 port map( A1 => n1919, A2 => n1920, ZN => 
                           curr_proc_regs(510));
   U2430 : AOI222_X1 port map( A1 => regs(510), A2 => n134, B1 => regs(2046), 
                           B2 => n172, C1 => regs(1022), C2 => n247, ZN => 
                           n1920);
   U2431 : AOI22_X1 port map( A1 => regs(1534), A2 => n11, B1 => regs(2558), B2
                           => n359, ZN => n1919);
   U2432 : NAND2_X1 port map( A1 => n1921, A2 => n1922, ZN => 
                           curr_proc_regs(509));
   U2433 : AOI222_X1 port map( A1 => regs(509), A2 => n134, B1 => regs(2045), 
                           B2 => n172, C1 => regs(1021), C2 => n247, ZN => 
                           n1922);
   U2434 : AOI22_X1 port map( A1 => regs(1533), A2 => n11, B1 => regs(2557), B2
                           => n354, ZN => n1921);
   U2435 : NAND2_X1 port map( A1 => n1923, A2 => n1924, ZN => 
                           curr_proc_regs(508));
   U2436 : AOI222_X1 port map( A1 => regs(508), A2 => n134, B1 => regs(2044), 
                           B2 => n172, C1 => regs(1020), C2 => n247, ZN => 
                           n1924);
   U2437 : AOI22_X1 port map( A1 => regs(1532), A2 => n11, B1 => regs(2556), B2
                           => n354, ZN => n1923);
   U2438 : NAND2_X1 port map( A1 => n1925, A2 => n1926, ZN => 
                           curr_proc_regs(507));
   U2439 : AOI222_X1 port map( A1 => regs(507), A2 => n135, B1 => regs(2043), 
                           B2 => n171, C1 => regs(1019), C2 => n246, ZN => 
                           n1926);
   U2440 : AOI22_X1 port map( A1 => regs(1531), A2 => n11, B1 => regs(2555), B2
                           => n354, ZN => n1925);
   U2441 : NAND2_X1 port map( A1 => n1927, A2 => n1928, ZN => 
                           curr_proc_regs(506));
   U2442 : AOI222_X1 port map( A1 => regs(506), A2 => n135, B1 => regs(2042), 
                           B2 => n171, C1 => regs(1018), C2 => n246, ZN => 
                           n1928);
   U2443 : AOI22_X1 port map( A1 => regs(1530), A2 => n11, B1 => regs(2554), B2
                           => n354, ZN => n1927);
   U2444 : NAND2_X1 port map( A1 => n1929, A2 => n1930, ZN => 
                           curr_proc_regs(505));
   U2445 : AOI222_X1 port map( A1 => regs(505), A2 => n135, B1 => regs(2041), 
                           B2 => n171, C1 => regs(1017), C2 => n246, ZN => 
                           n1930);
   U2446 : AOI22_X1 port map( A1 => regs(1529), A2 => n11, B1 => regs(2553), B2
                           => n354, ZN => n1929);
   U2447 : NAND2_X1 port map( A1 => n1931, A2 => n1932, ZN => 
                           curr_proc_regs(504));
   U2448 : AOI222_X1 port map( A1 => regs(504), A2 => n135, B1 => regs(2040), 
                           B2 => n171, C1 => regs(1016), C2 => n246, ZN => 
                           n1932);
   U2449 : AOI22_X1 port map( A1 => regs(1528), A2 => n11, B1 => regs(2552), B2
                           => n354, ZN => n1931);
   U2450 : NAND2_X1 port map( A1 => n1933, A2 => n1934, ZN => 
                           curr_proc_regs(503));
   U2451 : AOI222_X1 port map( A1 => regs(503), A2 => n135, B1 => regs(2039), 
                           B2 => n171, C1 => regs(1015), C2 => n246, ZN => 
                           n1934);
   U2452 : AOI22_X1 port map( A1 => regs(1527), A2 => n11, B1 => regs(2551), B2
                           => n355, ZN => n1933);
   U2453 : NAND2_X1 port map( A1 => n1935, A2 => n1936, ZN => 
                           curr_proc_regs(502));
   U2454 : AOI222_X1 port map( A1 => regs(502), A2 => n135, B1 => regs(2038), 
                           B2 => n171, C1 => regs(1014), C2 => n246, ZN => 
                           n1936);
   U2455 : AOI22_X1 port map( A1 => regs(1526), A2 => n10, B1 => regs(2550), B2
                           => n355, ZN => n1935);
   U2456 : NAND2_X1 port map( A1 => n1937, A2 => n1938, ZN => 
                           curr_proc_regs(501));
   U2457 : AOI222_X1 port map( A1 => regs(501), A2 => n135, B1 => regs(2037), 
                           B2 => n171, C1 => regs(1013), C2 => n246, ZN => 
                           n1938);
   U2458 : AOI22_X1 port map( A1 => regs(1525), A2 => n10, B1 => regs(2549), B2
                           => n355, ZN => n1937);
   U2459 : NAND2_X1 port map( A1 => n1939, A2 => n1940, ZN => 
                           curr_proc_regs(500));
   U2460 : AOI222_X1 port map( A1 => regs(500), A2 => n135, B1 => regs(2036), 
                           B2 => n171, C1 => regs(1012), C2 => n246, ZN => 
                           n1940);
   U2461 : AOI22_X1 port map( A1 => regs(1524), A2 => n10, B1 => regs(2548), B2
                           => n355, ZN => n1939);
   U2462 : NAND2_X1 port map( A1 => n1941, A2 => n1942, ZN => 
                           curr_proc_regs(499));
   U2463 : AOI222_X1 port map( A1 => regs(499), A2 => n135, B1 => regs(2035), 
                           B2 => n171, C1 => regs(1011), C2 => n246, ZN => 
                           n1942);
   U2464 : AOI22_X1 port map( A1 => regs(1523), A2 => n10, B1 => regs(2547), B2
                           => n355, ZN => n1941);
   U2465 : NAND2_X1 port map( A1 => n1943, A2 => n1944, ZN => 
                           curr_proc_regs(498));
   U2466 : AOI222_X1 port map( A1 => regs(498), A2 => n135, B1 => regs(2034), 
                           B2 => n171, C1 => regs(1010), C2 => n246, ZN => 
                           n1944);
   U2467 : AOI22_X1 port map( A1 => regs(1522), A2 => n10, B1 => regs(2546), B2
                           => n355, ZN => n1943);
   U2468 : NAND2_X1 port map( A1 => n1945, A2 => n1946, ZN => 
                           curr_proc_regs(497));
   U2469 : AOI222_X1 port map( A1 => regs(497), A2 => n135, B1 => regs(2033), 
                           B2 => n171, C1 => regs(1009), C2 => n246, ZN => 
                           n1946);
   U2470 : AOI22_X1 port map( A1 => regs(1521), A2 => n10, B1 => regs(2545), B2
                           => n355, ZN => n1945);
   U2471 : NAND2_X1 port map( A1 => n1947, A2 => n1948, ZN => 
                           curr_proc_regs(496));
   U2472 : AOI222_X1 port map( A1 => regs(496), A2 => n135, B1 => regs(2032), 
                           B2 => n171, C1 => regs(1008), C2 => n246, ZN => 
                           n1948);
   U2473 : AOI22_X1 port map( A1 => regs(1520), A2 => n10, B1 => regs(2544), B2
                           => n355, ZN => n1947);
   U2474 : NAND2_X1 port map( A1 => n1949, A2 => n1950, ZN => 
                           curr_proc_regs(495));
   U2475 : AOI222_X1 port map( A1 => regs(495), A2 => n136, B1 => regs(2031), 
                           B2 => n170, C1 => regs(1007), C2 => n245, ZN => 
                           n1950);
   U2476 : AOI22_X1 port map( A1 => regs(1519), A2 => n10, B1 => regs(2543), B2
                           => n355, ZN => n1949);
   U2477 : NAND2_X1 port map( A1 => n1951, A2 => n1952, ZN => 
                           curr_proc_regs(494));
   U2478 : AOI222_X1 port map( A1 => regs(494), A2 => n136, B1 => regs(2030), 
                           B2 => n170, C1 => regs(1006), C2 => n245, ZN => 
                           n1952);
   U2479 : AOI22_X1 port map( A1 => regs(1518), A2 => n10, B1 => regs(2542), B2
                           => n355, ZN => n1951);
   U2480 : NAND2_X1 port map( A1 => n1953, A2 => n1954, ZN => 
                           curr_proc_regs(493));
   U2481 : AOI222_X1 port map( A1 => regs(493), A2 => n136, B1 => regs(2029), 
                           B2 => n170, C1 => regs(1005), C2 => n245, ZN => 
                           n1954);
   U2482 : AOI22_X1 port map( A1 => regs(1517), A2 => n10, B1 => regs(2541), B2
                           => n355, ZN => n1953);
   U2483 : NAND2_X1 port map( A1 => n1955, A2 => n1956, ZN => 
                           curr_proc_regs(492));
   U2484 : AOI222_X1 port map( A1 => regs(492), A2 => n136, B1 => regs(2028), 
                           B2 => n170, C1 => regs(1004), C2 => n245, ZN => 
                           n1956);
   U2485 : AOI22_X1 port map( A1 => regs(1516), A2 => n10, B1 => regs(2540), B2
                           => n355, ZN => n1955);
   U2486 : NAND2_X1 port map( A1 => n1957, A2 => n1958, ZN => 
                           curr_proc_regs(491));
   U2487 : AOI222_X1 port map( A1 => regs(491), A2 => n136, B1 => regs(2027), 
                           B2 => n170, C1 => regs(1003), C2 => n245, ZN => 
                           n1958);
   U2488 : AOI22_X1 port map( A1 => regs(1515), A2 => n10, B1 => regs(2539), B2
                           => n356, ZN => n1957);
   U2489 : NAND2_X1 port map( A1 => n1959, A2 => n1960, ZN => 
                           curr_proc_regs(490));
   U2490 : AOI222_X1 port map( A1 => regs(490), A2 => n136, B1 => regs(2026), 
                           B2 => n170, C1 => regs(1002), C2 => n245, ZN => 
                           n1960);
   U2491 : AOI22_X1 port map( A1 => regs(1514), A2 => n9, B1 => regs(2538), B2 
                           => n356, ZN => n1959);
   U2492 : NAND2_X1 port map( A1 => n1961, A2 => n1962, ZN => 
                           curr_proc_regs(489));
   U2493 : AOI222_X1 port map( A1 => regs(489), A2 => n136, B1 => regs(2025), 
                           B2 => n170, C1 => regs(1001), C2 => n245, ZN => 
                           n1962);
   U2494 : AOI22_X1 port map( A1 => regs(1513), A2 => n9, B1 => regs(2537), B2 
                           => n356, ZN => n1961);
   U2495 : NAND2_X1 port map( A1 => n1963, A2 => n1964, ZN => 
                           curr_proc_regs(488));
   U2496 : AOI222_X1 port map( A1 => regs(488), A2 => n136, B1 => regs(2024), 
                           B2 => n170, C1 => regs(1000), C2 => n245, ZN => 
                           n1964);
   U2497 : AOI22_X1 port map( A1 => regs(1512), A2 => n9, B1 => regs(2536), B2 
                           => n356, ZN => n1963);
   U2498 : NAND2_X1 port map( A1 => n1965, A2 => n1966, ZN => 
                           curr_proc_regs(487));
   U2499 : AOI222_X1 port map( A1 => regs(487), A2 => n136, B1 => regs(2023), 
                           B2 => n170, C1 => regs(999), C2 => n245, ZN => n1966
                           );
   U2500 : AOI22_X1 port map( A1 => regs(1511), A2 => n9, B1 => regs(2535), B2 
                           => n356, ZN => n1965);
   U2501 : NAND2_X1 port map( A1 => n1967, A2 => n1968, ZN => 
                           curr_proc_regs(486));
   U2502 : AOI222_X1 port map( A1 => regs(486), A2 => n136, B1 => regs(2022), 
                           B2 => n170, C1 => regs(998), C2 => n245, ZN => n1968
                           );
   U2503 : AOI22_X1 port map( A1 => regs(1510), A2 => n9, B1 => regs(2534), B2 
                           => n356, ZN => n1967);
   U2504 : NAND2_X1 port map( A1 => n1969, A2 => n1970, ZN => 
                           curr_proc_regs(485));
   U2505 : AOI222_X1 port map( A1 => regs(485), A2 => n136, B1 => regs(2021), 
                           B2 => n170, C1 => regs(997), C2 => n245, ZN => n1970
                           );
   U2506 : AOI22_X1 port map( A1 => regs(1509), A2 => n9, B1 => regs(2533), B2 
                           => n356, ZN => n1969);
   U2507 : NAND2_X1 port map( A1 => n1971, A2 => n1972, ZN => 
                           curr_proc_regs(484));
   U2508 : AOI222_X1 port map( A1 => regs(484), A2 => n136, B1 => regs(2020), 
                           B2 => n170, C1 => regs(996), C2 => n245, ZN => n1972
                           );
   U2509 : AOI22_X1 port map( A1 => regs(1508), A2 => n9, B1 => regs(2532), B2 
                           => n356, ZN => n1971);
   U2510 : NAND2_X1 port map( A1 => n1973, A2 => n1974, ZN => 
                           curr_proc_regs(483));
   U2511 : AOI222_X1 port map( A1 => regs(483), A2 => n137, B1 => regs(2019), 
                           B2 => n169, C1 => regs(995), C2 => n244, ZN => n1974
                           );
   U2512 : AOI22_X1 port map( A1 => regs(1507), A2 => n9, B1 => regs(2531), B2 
                           => n356, ZN => n1973);
   U2513 : NAND2_X1 port map( A1 => n1975, A2 => n1976, ZN => 
                           curr_proc_regs(482));
   U2514 : AOI222_X1 port map( A1 => regs(482), A2 => n137, B1 => regs(2018), 
                           B2 => n169, C1 => regs(994), C2 => n244, ZN => n1976
                           );
   U2515 : AOI22_X1 port map( A1 => regs(1506), A2 => n9, B1 => regs(2530), B2 
                           => n356, ZN => n1975);
   U2516 : NAND2_X1 port map( A1 => n1977, A2 => n1978, ZN => 
                           curr_proc_regs(481));
   U2517 : AOI222_X1 port map( A1 => regs(481), A2 => n137, B1 => regs(2017), 
                           B2 => n169, C1 => regs(993), C2 => n244, ZN => n1978
                           );
   U2518 : AOI22_X1 port map( A1 => regs(1505), A2 => n9, B1 => regs(2529), B2 
                           => n356, ZN => n1977);
   U2519 : NAND2_X1 port map( A1 => n1979, A2 => n1980, ZN => 
                           curr_proc_regs(480));
   U2520 : AOI222_X1 port map( A1 => regs(480), A2 => n137, B1 => regs(2016), 
                           B2 => n169, C1 => regs(992), C2 => n244, ZN => n1980
                           );
   U2521 : AOI22_X1 port map( A1 => regs(1504), A2 => n9, B1 => regs(2528), B2 
                           => n356, ZN => n1979);
   U2522 : NAND2_X1 port map( A1 => n1981, A2 => n1982, ZN => 
                           curr_proc_regs(479));
   U2523 : AOI222_X1 port map( A1 => regs(479), A2 => n137, B1 => regs(2015), 
                           B2 => n169, C1 => regs(991), C2 => n244, ZN => n1982
                           );
   U2524 : AOI22_X1 port map( A1 => regs(1503), A2 => n9, B1 => regs(2527), B2 
                           => n357, ZN => n1981);
   U2525 : NAND2_X1 port map( A1 => n1983, A2 => n1984, ZN => 
                           curr_proc_regs(478));
   U2526 : AOI222_X1 port map( A1 => regs(478), A2 => n137, B1 => regs(2014), 
                           B2 => n169, C1 => regs(990), C2 => n244, ZN => n1984
                           );
   U2527 : AOI22_X1 port map( A1 => regs(1502), A2 => n8, B1 => regs(2526), B2 
                           => n357, ZN => n1983);
   U2528 : NAND2_X1 port map( A1 => n1985, A2 => n1986, ZN => 
                           curr_proc_regs(477));
   U2529 : AOI222_X1 port map( A1 => regs(477), A2 => n137, B1 => regs(2013), 
                           B2 => n169, C1 => regs(989), C2 => n244, ZN => n1986
                           );
   U2530 : AOI22_X1 port map( A1 => regs(1501), A2 => n8, B1 => regs(2525), B2 
                           => n357, ZN => n1985);
   U2531 : NAND2_X1 port map( A1 => n1987, A2 => n1988, ZN => 
                           curr_proc_regs(476));
   U2532 : AOI222_X1 port map( A1 => regs(476), A2 => n137, B1 => regs(2012), 
                           B2 => n169, C1 => regs(988), C2 => n244, ZN => n1988
                           );
   U2533 : AOI22_X1 port map( A1 => regs(1500), A2 => n8, B1 => regs(2524), B2 
                           => n357, ZN => n1987);
   U2534 : NAND2_X1 port map( A1 => n1989, A2 => n1990, ZN => 
                           curr_proc_regs(475));
   U2535 : AOI222_X1 port map( A1 => regs(475), A2 => n137, B1 => regs(2011), 
                           B2 => n169, C1 => regs(987), C2 => n244, ZN => n1990
                           );
   U2536 : AOI22_X1 port map( A1 => regs(1499), A2 => n8, B1 => regs(2523), B2 
                           => n357, ZN => n1989);
   U2537 : NAND2_X1 port map( A1 => n1991, A2 => n1992, ZN => 
                           curr_proc_regs(474));
   U2538 : AOI222_X1 port map( A1 => regs(474), A2 => n137, B1 => regs(2010), 
                           B2 => n169, C1 => regs(986), C2 => n244, ZN => n1992
                           );
   U2539 : AOI22_X1 port map( A1 => regs(1498), A2 => n8, B1 => regs(2522), B2 
                           => n357, ZN => n1991);
   U2540 : NAND2_X1 port map( A1 => n1993, A2 => n1994, ZN => 
                           curr_proc_regs(473));
   U2541 : AOI222_X1 port map( A1 => regs(473), A2 => n137, B1 => regs(2009), 
                           B2 => n169, C1 => regs(985), C2 => n244, ZN => n1994
                           );
   U2542 : AOI22_X1 port map( A1 => regs(1497), A2 => n8, B1 => regs(2521), B2 
                           => n357, ZN => n1993);
   U2543 : NAND2_X1 port map( A1 => n1995, A2 => n1996, ZN => 
                           curr_proc_regs(472));
   U2544 : AOI222_X1 port map( A1 => regs(472), A2 => n137, B1 => regs(2008), 
                           B2 => n169, C1 => regs(984), C2 => n244, ZN => n1996
                           );
   U2545 : AOI22_X1 port map( A1 => regs(1496), A2 => n8, B1 => regs(2520), B2 
                           => n357, ZN => n1995);
   U2546 : NAND2_X1 port map( A1 => n1997, A2 => n1998, ZN => 
                           curr_proc_regs(471));
   U2547 : AOI222_X1 port map( A1 => regs(471), A2 => n138, B1 => regs(2007), 
                           B2 => n168, C1 => regs(983), C2 => n243, ZN => n1998
                           );
   U2548 : AOI22_X1 port map( A1 => regs(1495), A2 => n8, B1 => regs(2519), B2 
                           => n357, ZN => n1997);
   U2549 : NAND2_X1 port map( A1 => n1999, A2 => n2000, ZN => 
                           curr_proc_regs(470));
   U2550 : AOI222_X1 port map( A1 => regs(470), A2 => n138, B1 => regs(2006), 
                           B2 => n168, C1 => regs(982), C2 => n243, ZN => n2000
                           );
   U2551 : AOI22_X1 port map( A1 => regs(1494), A2 => n8, B1 => regs(2518), B2 
                           => n357, ZN => n1999);
   U2552 : NAND2_X1 port map( A1 => n2001, A2 => n2002, ZN => 
                           curr_proc_regs(469));
   U2553 : AOI222_X1 port map( A1 => regs(469), A2 => n138, B1 => regs(2005), 
                           B2 => n168, C1 => regs(981), C2 => n243, ZN => n2002
                           );
   U2554 : AOI22_X1 port map( A1 => regs(1493), A2 => n8, B1 => regs(2517), B2 
                           => n357, ZN => n2001);
   U2555 : NAND2_X1 port map( A1 => n2003, A2 => n2004, ZN => 
                           curr_proc_regs(468));
   U2556 : AOI222_X1 port map( A1 => regs(468), A2 => n138, B1 => regs(2004), 
                           B2 => n168, C1 => regs(980), C2 => n243, ZN => n2004
                           );
   U2557 : AOI22_X1 port map( A1 => regs(1492), A2 => n8, B1 => regs(2516), B2 
                           => n357, ZN => n2003);
   U2558 : NAND2_X1 port map( A1 => n2005, A2 => n2006, ZN => 
                           curr_proc_regs(467));
   U2559 : AOI222_X1 port map( A1 => regs(467), A2 => n138, B1 => regs(2003), 
                           B2 => n168, C1 => regs(979), C2 => n243, ZN => n2006
                           );
   U2560 : AOI22_X1 port map( A1 => regs(1491), A2 => n8, B1 => regs(2515), B2 
                           => n358, ZN => n2005);
   U2561 : NAND2_X1 port map( A1 => n2007, A2 => n2008, ZN => 
                           curr_proc_regs(466));
   U2562 : AOI222_X1 port map( A1 => regs(466), A2 => n138, B1 => regs(2002), 
                           B2 => n168, C1 => regs(978), C2 => n243, ZN => n2008
                           );
   U2563 : AOI22_X1 port map( A1 => regs(1490), A2 => n7, B1 => regs(2514), B2 
                           => n358, ZN => n2007);
   U2564 : NAND2_X1 port map( A1 => n2009, A2 => n2010, ZN => 
                           curr_proc_regs(465));
   U2565 : AOI222_X1 port map( A1 => regs(465), A2 => n138, B1 => regs(2001), 
                           B2 => n168, C1 => regs(977), C2 => n243, ZN => n2010
                           );
   U2566 : AOI22_X1 port map( A1 => regs(1489), A2 => n7, B1 => regs(2513), B2 
                           => n358, ZN => n2009);
   U2567 : NAND2_X1 port map( A1 => n2011, A2 => n2012, ZN => 
                           curr_proc_regs(464));
   U2568 : AOI222_X1 port map( A1 => regs(464), A2 => n138, B1 => regs(2000), 
                           B2 => n168, C1 => regs(976), C2 => n243, ZN => n2012
                           );
   U2569 : AOI22_X1 port map( A1 => regs(1488), A2 => n7, B1 => regs(2512), B2 
                           => n358, ZN => n2011);
   U2570 : NAND2_X1 port map( A1 => n2013, A2 => n2014, ZN => 
                           curr_proc_regs(463));
   U2571 : AOI222_X1 port map( A1 => regs(463), A2 => n138, B1 => regs(1999), 
                           B2 => n168, C1 => regs(975), C2 => n243, ZN => n2014
                           );
   U2572 : AOI22_X1 port map( A1 => regs(1487), A2 => n7, B1 => regs(2511), B2 
                           => n358, ZN => n2013);
   U2573 : NAND2_X1 port map( A1 => n2015, A2 => n2016, ZN => 
                           curr_proc_regs(462));
   U2574 : AOI222_X1 port map( A1 => regs(462), A2 => n138, B1 => regs(1998), 
                           B2 => n168, C1 => regs(974), C2 => n243, ZN => n2016
                           );
   U2575 : AOI22_X1 port map( A1 => regs(1486), A2 => n7, B1 => regs(2510), B2 
                           => n358, ZN => n2015);
   U2576 : NAND2_X1 port map( A1 => n2017, A2 => n2018, ZN => 
                           curr_proc_regs(461));
   U2577 : AOI222_X1 port map( A1 => regs(461), A2 => n138, B1 => regs(1997), 
                           B2 => n168, C1 => regs(973), C2 => n243, ZN => n2018
                           );
   U2578 : AOI22_X1 port map( A1 => regs(1485), A2 => n7, B1 => regs(2509), B2 
                           => n358, ZN => n2017);
   U2579 : NAND2_X1 port map( A1 => n2019, A2 => n2020, ZN => 
                           curr_proc_regs(460));
   U2580 : AOI222_X1 port map( A1 => regs(460), A2 => n138, B1 => regs(1996), 
                           B2 => n168, C1 => regs(972), C2 => n243, ZN => n2020
                           );
   U2581 : AOI22_X1 port map( A1 => regs(1484), A2 => n7, B1 => regs(2508), B2 
                           => n358, ZN => n2019);
   U2582 : NAND2_X1 port map( A1 => n2021, A2 => n2022, ZN => 
                           curr_proc_regs(459));
   U2583 : AOI222_X1 port map( A1 => regs(459), A2 => n139, B1 => regs(1995), 
                           B2 => n167, C1 => regs(971), C2 => n242, ZN => n2022
                           );
   U2584 : AOI22_X1 port map( A1 => regs(1483), A2 => n7, B1 => regs(2507), B2 
                           => n358, ZN => n2021);
   U2585 : NAND2_X1 port map( A1 => n2023, A2 => n2024, ZN => 
                           curr_proc_regs(458));
   U2586 : AOI222_X1 port map( A1 => regs(458), A2 => n139, B1 => regs(1994), 
                           B2 => n167, C1 => regs(970), C2 => n242, ZN => n2024
                           );
   U2587 : AOI22_X1 port map( A1 => regs(1482), A2 => n7, B1 => regs(2506), B2 
                           => n358, ZN => n2023);
   U2588 : NAND2_X1 port map( A1 => n2025, A2 => n2026, ZN => 
                           curr_proc_regs(457));
   U2589 : AOI222_X1 port map( A1 => regs(457), A2 => n139, B1 => regs(1993), 
                           B2 => n167, C1 => regs(969), C2 => n242, ZN => n2026
                           );
   U2590 : AOI22_X1 port map( A1 => regs(1481), A2 => n7, B1 => regs(2505), B2 
                           => n358, ZN => n2025);
   U2591 : NAND2_X1 port map( A1 => n2027, A2 => n2028, ZN => 
                           curr_proc_regs(456));
   U2592 : AOI222_X1 port map( A1 => regs(456), A2 => n139, B1 => regs(1992), 
                           B2 => n167, C1 => regs(968), C2 => n242, ZN => n2028
                           );
   U2593 : AOI22_X1 port map( A1 => regs(1480), A2 => n7, B1 => regs(2504), B2 
                           => n358, ZN => n2027);
   U2594 : NAND2_X1 port map( A1 => n2029, A2 => n2030, ZN => 
                           curr_proc_regs(455));
   U2595 : AOI222_X1 port map( A1 => regs(455), A2 => n139, B1 => regs(1991), 
                           B2 => n167, C1 => regs(967), C2 => n242, ZN => n2030
                           );
   U2596 : AOI22_X1 port map( A1 => regs(1479), A2 => n7, B1 => regs(2503), B2 
                           => n359, ZN => n2029);
   U2597 : NAND2_X1 port map( A1 => n2031, A2 => n2032, ZN => 
                           curr_proc_regs(454));
   U2598 : AOI222_X1 port map( A1 => regs(454), A2 => n139, B1 => regs(1990), 
                           B2 => n167, C1 => regs(966), C2 => n242, ZN => n2032
                           );
   U2599 : AOI22_X1 port map( A1 => regs(1478), A2 => n6, B1 => regs(2502), B2 
                           => n359, ZN => n2031);
   U2600 : NAND2_X1 port map( A1 => n2033, A2 => n2034, ZN => 
                           curr_proc_regs(453));
   U2601 : AOI222_X1 port map( A1 => regs(453), A2 => n139, B1 => regs(1989), 
                           B2 => n167, C1 => regs(965), C2 => n242, ZN => n2034
                           );
   U2602 : AOI22_X1 port map( A1 => regs(1477), A2 => n6, B1 => regs(2501), B2 
                           => n359, ZN => n2033);
   U2603 : NAND2_X1 port map( A1 => n2035, A2 => n2036, ZN => 
                           curr_proc_regs(452));
   U2604 : AOI222_X1 port map( A1 => regs(452), A2 => n139, B1 => regs(1988), 
                           B2 => n167, C1 => regs(964), C2 => n242, ZN => n2036
                           );
   U2605 : AOI22_X1 port map( A1 => regs(1476), A2 => n6, B1 => regs(2500), B2 
                           => n359, ZN => n2035);
   U2606 : NAND2_X1 port map( A1 => n2037, A2 => n2038, ZN => 
                           curr_proc_regs(451));
   U2607 : AOI222_X1 port map( A1 => regs(451), A2 => n139, B1 => regs(1987), 
                           B2 => n167, C1 => regs(963), C2 => n242, ZN => n2038
                           );
   U2608 : AOI22_X1 port map( A1 => regs(1475), A2 => n6, B1 => regs(2499), B2 
                           => n359, ZN => n2037);
   U2609 : NAND2_X1 port map( A1 => n2039, A2 => n2040, ZN => 
                           curr_proc_regs(450));
   U2610 : AOI222_X1 port map( A1 => regs(450), A2 => n139, B1 => regs(1986), 
                           B2 => n167, C1 => regs(962), C2 => n242, ZN => n2040
                           );
   U2611 : AOI22_X1 port map( A1 => regs(1474), A2 => n6, B1 => regs(2498), B2 
                           => n359, ZN => n2039);
   U2612 : NAND2_X1 port map( A1 => n2041, A2 => n2042, ZN => 
                           curr_proc_regs(449));
   U2613 : AOI222_X1 port map( A1 => regs(449), A2 => n139, B1 => regs(1985), 
                           B2 => n167, C1 => regs(961), C2 => n242, ZN => n2042
                           );
   U2614 : AOI22_X1 port map( A1 => regs(1473), A2 => n6, B1 => regs(2497), B2 
                           => n359, ZN => n2041);
   U2615 : NAND2_X1 port map( A1 => n2043, A2 => n2044, ZN => 
                           curr_proc_regs(448));
   U2616 : AOI222_X1 port map( A1 => regs(448), A2 => n115, B1 => regs(1984), 
                           B2 => n167, C1 => regs(960), C2 => n242, ZN => n2044
                           );
   U2617 : AOI22_X1 port map( A1 => regs(1472), A2 => n6, B1 => regs(2496), B2 
                           => n359, ZN => n2043);
   U2618 : NAND2_X1 port map( A1 => n2045, A2 => n2046, ZN => 
                           curr_proc_regs(447));
   U2619 : AOI222_X1 port map( A1 => regs(447), A2 => n108, B1 => regs(1983), 
                           B2 => n166, C1 => regs(959), C2 => n241, ZN => n2046
                           );
   U2620 : AOI22_X1 port map( A1 => regs(1471), A2 => n6, B1 => regs(2495), B2 
                           => n359, ZN => n2045);
   U2621 : NAND2_X1 port map( A1 => n2047, A2 => n2048, ZN => 
                           curr_proc_regs(446));
   U2622 : AOI222_X1 port map( A1 => regs(446), A2 => n108, B1 => regs(1982), 
                           B2 => n166, C1 => regs(958), C2 => n241, ZN => n2048
                           );
   U2623 : AOI22_X1 port map( A1 => regs(1470), A2 => n6, B1 => regs(2494), B2 
                           => n359, ZN => n2047);
   U2624 : NAND2_X1 port map( A1 => n2049, A2 => n2050, ZN => 
                           curr_proc_regs(445));
   U2625 : AOI222_X1 port map( A1 => regs(445), A2 => n108, B1 => regs(1981), 
                           B2 => n166, C1 => regs(957), C2 => n241, ZN => n2050
                           );
   U2626 : AOI22_X1 port map( A1 => regs(1469), A2 => n6, B1 => regs(2493), B2 
                           => n359, ZN => n2049);
   U2627 : NAND2_X1 port map( A1 => n2051, A2 => n2052, ZN => 
                           curr_proc_regs(444));
   U2628 : AOI222_X1 port map( A1 => regs(444), A2 => n108, B1 => regs(1980), 
                           B2 => n166, C1 => regs(956), C2 => n241, ZN => n2052
                           );
   U2629 : AOI22_X1 port map( A1 => regs(1468), A2 => n6, B1 => regs(2492), B2 
                           => n360, ZN => n2051);
   U2630 : NAND2_X1 port map( A1 => n2053, A2 => n2054, ZN => 
                           curr_proc_regs(443));
   U2631 : AOI222_X1 port map( A1 => regs(443), A2 => n108, B1 => regs(1979), 
                           B2 => n166, C1 => regs(955), C2 => n241, ZN => n2054
                           );
   U2632 : AOI22_X1 port map( A1 => regs(1467), A2 => n5, B1 => regs(2491), B2 
                           => n360, ZN => n2053);
   U2633 : NAND2_X1 port map( A1 => n2055, A2 => n2056, ZN => 
                           curr_proc_regs(442));
   U2634 : AOI222_X1 port map( A1 => regs(442), A2 => n108, B1 => regs(1978), 
                           B2 => n166, C1 => regs(954), C2 => n241, ZN => n2056
                           );
   U2635 : AOI22_X1 port map( A1 => regs(1466), A2 => n5, B1 => regs(2490), B2 
                           => n360, ZN => n2055);
   U2636 : NAND2_X1 port map( A1 => n2057, A2 => n2058, ZN => 
                           curr_proc_regs(441));
   U2637 : AOI222_X1 port map( A1 => regs(441), A2 => n108, B1 => regs(1977), 
                           B2 => n166, C1 => regs(953), C2 => n241, ZN => n2058
                           );
   U2638 : AOI22_X1 port map( A1 => regs(1465), A2 => n5, B1 => regs(2489), B2 
                           => n360, ZN => n2057);
   U2639 : NAND2_X1 port map( A1 => n2059, A2 => n2060, ZN => 
                           curr_proc_regs(440));
   U2640 : AOI222_X1 port map( A1 => regs(440), A2 => n108, B1 => regs(1976), 
                           B2 => n166, C1 => regs(952), C2 => n241, ZN => n2060
                           );
   U2641 : AOI22_X1 port map( A1 => regs(1464), A2 => n5, B1 => regs(2488), B2 
                           => n360, ZN => n2059);
   U2642 : NAND2_X1 port map( A1 => n2061, A2 => n2062, ZN => 
                           curr_proc_regs(439));
   U2643 : AOI222_X1 port map( A1 => regs(439), A2 => n108, B1 => regs(1975), 
                           B2 => n166, C1 => regs(951), C2 => n241, ZN => n2062
                           );
   U2644 : AOI22_X1 port map( A1 => regs(1463), A2 => n5, B1 => regs(2487), B2 
                           => n360, ZN => n2061);
   U2645 : NAND2_X1 port map( A1 => n2063, A2 => n2064, ZN => 
                           curr_proc_regs(438));
   U2646 : AOI222_X1 port map( A1 => regs(438), A2 => n108, B1 => regs(1974), 
                           B2 => n166, C1 => regs(950), C2 => n241, ZN => n2064
                           );
   U2647 : AOI22_X1 port map( A1 => regs(1462), A2 => n5, B1 => regs(2486), B2 
                           => n360, ZN => n2063);
   U2648 : NAND2_X1 port map( A1 => n2065, A2 => n2066, ZN => 
                           curr_proc_regs(437));
   U2649 : AOI222_X1 port map( A1 => regs(437), A2 => n108, B1 => regs(1973), 
                           B2 => n166, C1 => regs(949), C2 => n241, ZN => n2066
                           );
   U2650 : AOI22_X1 port map( A1 => regs(1461), A2 => n5, B1 => regs(2485), B2 
                           => n360, ZN => n2065);
   U2651 : NAND2_X1 port map( A1 => n2067, A2 => n2068, ZN => 
                           curr_proc_regs(436));
   U2652 : AOI222_X1 port map( A1 => regs(436), A2 => n108, B1 => regs(1972), 
                           B2 => n166, C1 => regs(948), C2 => n241, ZN => n2068
                           );
   U2653 : AOI22_X1 port map( A1 => regs(1460), A2 => n5, B1 => regs(2484), B2 
                           => n360, ZN => n2067);
   U2654 : NAND2_X1 port map( A1 => n2069, A2 => n2070, ZN => 
                           curr_proc_regs(435));
   U2655 : AOI222_X1 port map( A1 => regs(435), A2 => n109, B1 => regs(1971), 
                           B2 => n165, C1 => regs(947), C2 => n240, ZN => n2070
                           );
   U2656 : AOI22_X1 port map( A1 => regs(1459), A2 => n5, B1 => regs(2483), B2 
                           => n360, ZN => n2069);
   U2657 : NAND2_X1 port map( A1 => n2071, A2 => n2072, ZN => 
                           curr_proc_regs(434));
   U2658 : AOI222_X1 port map( A1 => regs(434), A2 => n109, B1 => regs(1970), 
                           B2 => n165, C1 => regs(946), C2 => n240, ZN => n2072
                           );
   U2659 : AOI22_X1 port map( A1 => regs(1458), A2 => n5, B1 => regs(2482), B2 
                           => n360, ZN => n2071);
   U2660 : NAND2_X1 port map( A1 => n2073, A2 => n2074, ZN => 
                           curr_proc_regs(433));
   U2661 : AOI222_X1 port map( A1 => regs(433), A2 => n109, B1 => regs(1969), 
                           B2 => n165, C1 => regs(945), C2 => n240, ZN => n2074
                           );
   U2662 : AOI22_X1 port map( A1 => regs(1457), A2 => n5, B1 => regs(2481), B2 
                           => n360, ZN => n2073);
   U2663 : NAND2_X1 port map( A1 => n2075, A2 => n2076, ZN => 
                           curr_proc_regs(432));
   U2664 : AOI222_X1 port map( A1 => regs(432), A2 => n109, B1 => regs(1968), 
                           B2 => n165, C1 => regs(944), C2 => n240, ZN => n2076
                           );
   U2665 : AOI22_X1 port map( A1 => regs(1456), A2 => n5, B1 => regs(2480), B2 
                           => n361, ZN => n2075);
   U2666 : NAND2_X1 port map( A1 => n2077, A2 => n2078, ZN => 
                           curr_proc_regs(431));
   U2667 : AOI222_X1 port map( A1 => regs(431), A2 => n109, B1 => regs(1967), 
                           B2 => n165, C1 => regs(943), C2 => n240, ZN => n2078
                           );
   U2668 : AOI22_X1 port map( A1 => regs(1455), A2 => n4, B1 => regs(2479), B2 
                           => n361, ZN => n2077);
   U2669 : NAND2_X1 port map( A1 => n2079, A2 => n2080, ZN => 
                           curr_proc_regs(430));
   U2670 : AOI222_X1 port map( A1 => regs(430), A2 => n109, B1 => regs(1966), 
                           B2 => n165, C1 => regs(942), C2 => n240, ZN => n2080
                           );
   U2671 : AOI22_X1 port map( A1 => regs(1454), A2 => n4, B1 => regs(2478), B2 
                           => n361, ZN => n2079);
   U2672 : NAND2_X1 port map( A1 => n2081, A2 => n2082, ZN => 
                           curr_proc_regs(429));
   U2673 : AOI222_X1 port map( A1 => regs(429), A2 => n109, B1 => regs(1965), 
                           B2 => n165, C1 => regs(941), C2 => n240, ZN => n2082
                           );
   U2674 : AOI22_X1 port map( A1 => regs(1453), A2 => n4, B1 => regs(2477), B2 
                           => n361, ZN => n2081);
   U2675 : NAND2_X1 port map( A1 => n2083, A2 => n2084, ZN => 
                           curr_proc_regs(428));
   U2676 : AOI222_X1 port map( A1 => regs(428), A2 => n109, B1 => regs(1964), 
                           B2 => n165, C1 => regs(940), C2 => n240, ZN => n2084
                           );
   U2677 : AOI22_X1 port map( A1 => regs(1452), A2 => n4, B1 => regs(2476), B2 
                           => n361, ZN => n2083);
   U2678 : NAND2_X1 port map( A1 => n2085, A2 => n2086, ZN => 
                           curr_proc_regs(427));
   U2679 : AOI222_X1 port map( A1 => regs(427), A2 => n109, B1 => regs(1963), 
                           B2 => n165, C1 => regs(939), C2 => n240, ZN => n2086
                           );
   U2680 : AOI22_X1 port map( A1 => regs(1451), A2 => n4, B1 => regs(2475), B2 
                           => n361, ZN => n2085);
   U2681 : NAND2_X1 port map( A1 => n2087, A2 => n2088, ZN => 
                           curr_proc_regs(426));
   U2682 : AOI222_X1 port map( A1 => regs(426), A2 => n109, B1 => regs(1962), 
                           B2 => n165, C1 => regs(938), C2 => n240, ZN => n2088
                           );
   U2683 : AOI22_X1 port map( A1 => regs(1450), A2 => n4, B1 => regs(2474), B2 
                           => n361, ZN => n2087);
   U2684 : NAND2_X1 port map( A1 => n2089, A2 => n2090, ZN => 
                           curr_proc_regs(425));
   U2685 : AOI222_X1 port map( A1 => regs(425), A2 => n109, B1 => regs(1961), 
                           B2 => n165, C1 => regs(937), C2 => n240, ZN => n2090
                           );
   U2686 : AOI22_X1 port map( A1 => regs(1449), A2 => n4, B1 => regs(2473), B2 
                           => n361, ZN => n2089);
   U2687 : NAND2_X1 port map( A1 => n2091, A2 => n2092, ZN => 
                           curr_proc_regs(424));
   U2688 : AOI222_X1 port map( A1 => regs(424), A2 => n109, B1 => regs(1960), 
                           B2 => n165, C1 => regs(936), C2 => n240, ZN => n2092
                           );
   U2689 : AOI22_X1 port map( A1 => regs(1448), A2 => n4, B1 => regs(2472), B2 
                           => n361, ZN => n2091);
   U2690 : NAND2_X1 port map( A1 => n2093, A2 => n2094, ZN => 
                           curr_proc_regs(423));
   U2691 : AOI222_X1 port map( A1 => regs(423), A2 => n110, B1 => regs(1959), 
                           B2 => n164, C1 => regs(935), C2 => n239, ZN => n2094
                           );
   U2692 : AOI22_X1 port map( A1 => regs(1447), A2 => n4, B1 => regs(2471), B2 
                           => n361, ZN => n2093);
   U2693 : NAND2_X1 port map( A1 => n2095, A2 => n2096, ZN => 
                           curr_proc_regs(422));
   U2694 : AOI222_X1 port map( A1 => regs(422), A2 => n110, B1 => regs(1958), 
                           B2 => n164, C1 => regs(934), C2 => n239, ZN => n2096
                           );
   U2695 : AOI22_X1 port map( A1 => regs(1446), A2 => n4, B1 => regs(2470), B2 
                           => n361, ZN => n2095);
   U2696 : NAND2_X1 port map( A1 => n2097, A2 => n2098, ZN => 
                           curr_proc_regs(421));
   U2697 : AOI222_X1 port map( A1 => regs(421), A2 => n110, B1 => regs(1957), 
                           B2 => n164, C1 => regs(933), C2 => n239, ZN => n2098
                           );
   U2698 : AOI22_X1 port map( A1 => regs(1445), A2 => n4, B1 => regs(2469), B2 
                           => n361, ZN => n2097);
   U2699 : NAND2_X1 port map( A1 => n2099, A2 => n2100, ZN => 
                           curr_proc_regs(420));
   U2700 : AOI222_X1 port map( A1 => regs(420), A2 => n110, B1 => regs(1956), 
                           B2 => n164, C1 => regs(932), C2 => n239, ZN => n2100
                           );
   U2701 : AOI22_X1 port map( A1 => regs(1444), A2 => n4, B1 => regs(2468), B2 
                           => n362, ZN => n2099);
   U2702 : NAND2_X1 port map( A1 => n2101, A2 => n2102, ZN => 
                           curr_proc_regs(419));
   U2703 : AOI222_X1 port map( A1 => regs(419), A2 => n110, B1 => regs(1955), 
                           B2 => n164, C1 => regs(931), C2 => n239, ZN => n2102
                           );
   U2704 : AOI22_X1 port map( A1 => regs(1443), A2 => n3, B1 => regs(2467), B2 
                           => n362, ZN => n2101);
   U2705 : NAND2_X1 port map( A1 => n2103, A2 => n2104, ZN => 
                           curr_proc_regs(418));
   U2706 : AOI222_X1 port map( A1 => regs(418), A2 => n110, B1 => regs(1954), 
                           B2 => n164, C1 => regs(930), C2 => n239, ZN => n2104
                           );
   U2707 : AOI22_X1 port map( A1 => regs(1442), A2 => n3, B1 => regs(2466), B2 
                           => n362, ZN => n2103);
   U2708 : NAND2_X1 port map( A1 => n2105, A2 => n2106, ZN => 
                           curr_proc_regs(417));
   U2709 : AOI222_X1 port map( A1 => regs(417), A2 => n110, B1 => regs(1953), 
                           B2 => n164, C1 => regs(929), C2 => n239, ZN => n2106
                           );
   U2710 : AOI22_X1 port map( A1 => regs(1441), A2 => n3, B1 => regs(2465), B2 
                           => n362, ZN => n2105);
   U2711 : NAND2_X1 port map( A1 => n2107, A2 => n2108, ZN => 
                           curr_proc_regs(416));
   U2712 : AOI222_X1 port map( A1 => regs(416), A2 => n110, B1 => regs(1952), 
                           B2 => n164, C1 => regs(928), C2 => n239, ZN => n2108
                           );
   U2713 : AOI22_X1 port map( A1 => regs(1440), A2 => n3, B1 => regs(2464), B2 
                           => n362, ZN => n2107);
   U2714 : NAND2_X1 port map( A1 => n2109, A2 => n2110, ZN => 
                           curr_proc_regs(415));
   U2715 : AOI222_X1 port map( A1 => regs(415), A2 => n110, B1 => regs(1951), 
                           B2 => n164, C1 => regs(927), C2 => n239, ZN => n2110
                           );
   U2716 : AOI22_X1 port map( A1 => regs(1439), A2 => n3, B1 => regs(2463), B2 
                           => n362, ZN => n2109);
   U2717 : NAND2_X1 port map( A1 => n2111, A2 => n2112, ZN => 
                           curr_proc_regs(414));
   U2718 : AOI222_X1 port map( A1 => regs(414), A2 => n110, B1 => regs(1950), 
                           B2 => n164, C1 => regs(926), C2 => n239, ZN => n2112
                           );
   U2719 : AOI22_X1 port map( A1 => regs(1438), A2 => n3, B1 => regs(2462), B2 
                           => n362, ZN => n2111);
   U2720 : NAND2_X1 port map( A1 => n2113, A2 => n2114, ZN => 
                           curr_proc_regs(413));
   U2721 : AOI222_X1 port map( A1 => regs(413), A2 => n110, B1 => regs(1949), 
                           B2 => n164, C1 => regs(925), C2 => n239, ZN => n2114
                           );
   U2722 : AOI22_X1 port map( A1 => regs(1437), A2 => n3, B1 => regs(2461), B2 
                           => n362, ZN => n2113);
   U2723 : NAND2_X1 port map( A1 => n2115, A2 => n2116, ZN => 
                           curr_proc_regs(412));
   U2724 : AOI222_X1 port map( A1 => regs(412), A2 => n110, B1 => regs(1948), 
                           B2 => n164, C1 => regs(924), C2 => n239, ZN => n2116
                           );
   U2725 : AOI22_X1 port map( A1 => regs(1436), A2 => n3, B1 => regs(2460), B2 
                           => n362, ZN => n2115);
   U2726 : NAND2_X1 port map( A1 => n2117, A2 => n2118, ZN => 
                           curr_proc_regs(411));
   U2727 : AOI222_X1 port map( A1 => regs(411), A2 => n111, B1 => regs(1947), 
                           B2 => n163, C1 => regs(923), C2 => n238, ZN => n2118
                           );
   U2728 : AOI22_X1 port map( A1 => regs(1435), A2 => n3, B1 => regs(2459), B2 
                           => n362, ZN => n2117);
   U2729 : NAND2_X1 port map( A1 => n2119, A2 => n2120, ZN => 
                           curr_proc_regs(410));
   U2730 : AOI222_X1 port map( A1 => regs(410), A2 => n111, B1 => regs(1946), 
                           B2 => n163, C1 => regs(922), C2 => n238, ZN => n2120
                           );
   U2731 : AOI22_X1 port map( A1 => regs(1434), A2 => n3, B1 => regs(2458), B2 
                           => n362, ZN => n2119);
   U2732 : NAND2_X1 port map( A1 => n2121, A2 => n2122, ZN => 
                           curr_proc_regs(409));
   U2733 : AOI222_X1 port map( A1 => regs(409), A2 => n111, B1 => regs(1945), 
                           B2 => n163, C1 => regs(921), C2 => n238, ZN => n2122
                           );
   U2734 : AOI22_X1 port map( A1 => regs(1433), A2 => n3, B1 => regs(2457), B2 
                           => n362, ZN => n2121);
   U2735 : NAND2_X1 port map( A1 => n2123, A2 => n2124, ZN => 
                           curr_proc_regs(408));
   U2736 : AOI222_X1 port map( A1 => regs(408), A2 => n111, B1 => regs(1944), 
                           B2 => n163, C1 => regs(920), C2 => n238, ZN => n2124
                           );
   U2737 : AOI22_X1 port map( A1 => regs(1432), A2 => n3, B1 => regs(2456), B2 
                           => n363, ZN => n2123);
   U2738 : NAND2_X1 port map( A1 => n2125, A2 => n2126, ZN => 
                           curr_proc_regs(407));
   U2739 : AOI222_X1 port map( A1 => regs(407), A2 => n111, B1 => regs(1943), 
                           B2 => n163, C1 => regs(919), C2 => n238, ZN => n2126
                           );
   U2740 : AOI22_X1 port map( A1 => regs(1431), A2 => n2, B1 => regs(2455), B2 
                           => n363, ZN => n2125);
   U2741 : NAND2_X1 port map( A1 => n2127, A2 => n2128, ZN => 
                           curr_proc_regs(406));
   U2742 : AOI222_X1 port map( A1 => regs(406), A2 => n111, B1 => regs(1942), 
                           B2 => n163, C1 => regs(918), C2 => n238, ZN => n2128
                           );
   U2743 : AOI22_X1 port map( A1 => regs(1430), A2 => n2, B1 => regs(2454), B2 
                           => n363, ZN => n2127);
   U2744 : NAND2_X1 port map( A1 => n2129, A2 => n2130, ZN => 
                           curr_proc_regs(405));
   U2745 : AOI222_X1 port map( A1 => regs(405), A2 => n111, B1 => regs(1941), 
                           B2 => n163, C1 => regs(917), C2 => n238, ZN => n2130
                           );
   U2746 : AOI22_X1 port map( A1 => regs(1429), A2 => n2, B1 => regs(2453), B2 
                           => n363, ZN => n2129);
   U2747 : NAND2_X1 port map( A1 => n2131, A2 => n2132, ZN => 
                           curr_proc_regs(404));
   U2748 : AOI222_X1 port map( A1 => regs(404), A2 => n111, B1 => regs(1940), 
                           B2 => n163, C1 => regs(916), C2 => n238, ZN => n2132
                           );
   U2749 : AOI22_X1 port map( A1 => regs(1428), A2 => n2, B1 => regs(2452), B2 
                           => n363, ZN => n2131);
   U2750 : NAND2_X1 port map( A1 => n2133, A2 => n2134, ZN => 
                           curr_proc_regs(403));
   U2751 : AOI222_X1 port map( A1 => regs(403), A2 => n111, B1 => regs(1939), 
                           B2 => n163, C1 => regs(915), C2 => n238, ZN => n2134
                           );
   U2752 : AOI22_X1 port map( A1 => regs(1427), A2 => n2, B1 => regs(2451), B2 
                           => n363, ZN => n2133);
   U2753 : NAND2_X1 port map( A1 => n2135, A2 => n2136, ZN => 
                           curr_proc_regs(402));
   U2754 : AOI222_X1 port map( A1 => regs(402), A2 => n111, B1 => regs(1938), 
                           B2 => n163, C1 => regs(914), C2 => n238, ZN => n2136
                           );
   U2755 : AOI22_X1 port map( A1 => regs(1426), A2 => n2, B1 => regs(2450), B2 
                           => n363, ZN => n2135);
   U2756 : NAND2_X1 port map( A1 => n2137, A2 => n2138, ZN => 
                           curr_proc_regs(401));
   U2757 : AOI222_X1 port map( A1 => regs(401), A2 => n111, B1 => regs(1937), 
                           B2 => n163, C1 => regs(913), C2 => n238, ZN => n2138
                           );
   U2758 : AOI22_X1 port map( A1 => regs(1425), A2 => n2, B1 => regs(2449), B2 
                           => n363, ZN => n2137);
   U2759 : NAND2_X1 port map( A1 => n2139, A2 => n2140, ZN => 
                           curr_proc_regs(400));
   U2760 : AOI222_X1 port map( A1 => regs(400), A2 => n111, B1 => regs(1936), 
                           B2 => n163, C1 => regs(912), C2 => n238, ZN => n2140
                           );
   U2761 : AOI22_X1 port map( A1 => regs(1424), A2 => n2, B1 => regs(2448), B2 
                           => n363, ZN => n2139);
   U2762 : NAND2_X1 port map( A1 => n2141, A2 => n2142, ZN => 
                           curr_proc_regs(399));
   U2763 : AOI222_X1 port map( A1 => regs(399), A2 => n112, B1 => regs(1935), 
                           B2 => n162, C1 => regs(911), C2 => n237, ZN => n2142
                           );
   U2764 : AOI22_X1 port map( A1 => regs(1423), A2 => n2, B1 => regs(2447), B2 
                           => n363, ZN => n2141);
   U2765 : NAND2_X1 port map( A1 => n2143, A2 => n2144, ZN => 
                           curr_proc_regs(398));
   U2766 : AOI222_X1 port map( A1 => regs(398), A2 => n112, B1 => regs(1934), 
                           B2 => n162, C1 => regs(910), C2 => n237, ZN => n2144
                           );
   U2767 : AOI22_X1 port map( A1 => regs(1422), A2 => n2, B1 => regs(2446), B2 
                           => n363, ZN => n2143);
   U2768 : NAND2_X1 port map( A1 => n2145, A2 => n2146, ZN => 
                           curr_proc_regs(397));
   U2769 : AOI222_X1 port map( A1 => regs(397), A2 => n112, B1 => regs(1933), 
                           B2 => n162, C1 => regs(909), C2 => n237, ZN => n2146
                           );
   U2770 : AOI22_X1 port map( A1 => regs(1421), A2 => n2, B1 => regs(2445), B2 
                           => n363, ZN => n2145);
   U2771 : NAND2_X1 port map( A1 => n2147, A2 => n2148, ZN => 
                           curr_proc_regs(396));
   U2772 : AOI222_X1 port map( A1 => regs(396), A2 => n112, B1 => regs(1932), 
                           B2 => n162, C1 => regs(908), C2 => n237, ZN => n2148
                           );
   U2773 : AOI22_X1 port map( A1 => regs(1420), A2 => n2, B1 => regs(2444), B2 
                           => n364, ZN => n2147);
   U2774 : NAND2_X1 port map( A1 => n2149, A2 => n2150, ZN => 
                           curr_proc_regs(395));
   U2775 : AOI222_X1 port map( A1 => regs(395), A2 => n112, B1 => regs(1931), 
                           B2 => n162, C1 => regs(907), C2 => n237, ZN => n2150
                           );
   U2776 : AOI22_X1 port map( A1 => regs(1419), A2 => n1, B1 => regs(2443), B2 
                           => n364, ZN => n2149);
   U2777 : NAND2_X1 port map( A1 => n2151, A2 => n2152, ZN => 
                           curr_proc_regs(394));
   U2778 : AOI222_X1 port map( A1 => regs(394), A2 => n112, B1 => regs(1930), 
                           B2 => n162, C1 => regs(906), C2 => n237, ZN => n2152
                           );
   U2779 : AOI22_X1 port map( A1 => regs(1418), A2 => n1, B1 => regs(2442), B2 
                           => n364, ZN => n2151);
   U2780 : NAND2_X1 port map( A1 => n2153, A2 => n2154, ZN => 
                           curr_proc_regs(393));
   U2781 : AOI222_X1 port map( A1 => regs(393), A2 => n112, B1 => regs(1929), 
                           B2 => n162, C1 => regs(905), C2 => n237, ZN => n2154
                           );
   U2782 : AOI22_X1 port map( A1 => regs(1417), A2 => n1, B1 => regs(2441), B2 
                           => n364, ZN => n2153);
   U2783 : NAND2_X1 port map( A1 => n2155, A2 => n2156, ZN => 
                           curr_proc_regs(392));
   U2784 : AOI222_X1 port map( A1 => regs(392), A2 => n112, B1 => regs(1928), 
                           B2 => n162, C1 => regs(904), C2 => n237, ZN => n2156
                           );
   U2785 : AOI22_X1 port map( A1 => regs(1416), A2 => n1, B1 => regs(2440), B2 
                           => n364, ZN => n2155);
   U2786 : NAND2_X1 port map( A1 => n2157, A2 => n2158, ZN => 
                           curr_proc_regs(391));
   U2787 : AOI222_X1 port map( A1 => regs(391), A2 => n112, B1 => regs(1927), 
                           B2 => n162, C1 => regs(903), C2 => n237, ZN => n2158
                           );
   U2788 : AOI22_X1 port map( A1 => regs(1415), A2 => n1, B1 => regs(2439), B2 
                           => n364, ZN => n2157);
   U2789 : NAND2_X1 port map( A1 => n2159, A2 => n2160, ZN => 
                           curr_proc_regs(390));
   U2790 : AOI222_X1 port map( A1 => regs(390), A2 => n112, B1 => regs(1926), 
                           B2 => n162, C1 => regs(902), C2 => n237, ZN => n2160
                           );
   U2791 : AOI22_X1 port map( A1 => regs(1414), A2 => n1, B1 => regs(2438), B2 
                           => n364, ZN => n2159);
   U2792 : NAND2_X1 port map( A1 => n2161, A2 => n2162, ZN => 
                           curr_proc_regs(389));
   U2793 : AOI222_X1 port map( A1 => regs(389), A2 => n112, B1 => regs(1925), 
                           B2 => n162, C1 => regs(901), C2 => n237, ZN => n2162
                           );
   U2794 : AOI22_X1 port map( A1 => regs(1413), A2 => n1, B1 => regs(2437), B2 
                           => n364, ZN => n2161);
   U2795 : NAND2_X1 port map( A1 => n2163, A2 => n2164, ZN => 
                           curr_proc_regs(388));
   U2796 : AOI222_X1 port map( A1 => regs(388), A2 => n112, B1 => regs(1924), 
                           B2 => n162, C1 => regs(900), C2 => n237, ZN => n2164
                           );
   U2797 : AOI22_X1 port map( A1 => regs(1412), A2 => n1, B1 => regs(2436), B2 
                           => n364, ZN => n2163);
   U2798 : NAND2_X1 port map( A1 => n2165, A2 => n2166, ZN => 
                           curr_proc_regs(387));
   U2799 : AOI222_X1 port map( A1 => regs(387), A2 => n113, B1 => regs(1923), 
                           B2 => n161, C1 => regs(899), C2 => n236, ZN => n2166
                           );
   U2800 : AOI22_X1 port map( A1 => regs(1411), A2 => n1, B1 => regs(2435), B2 
                           => n364, ZN => n2165);
   U2801 : NAND2_X1 port map( A1 => n2167, A2 => n2168, ZN => 
                           curr_proc_regs(386));
   U2802 : AOI222_X1 port map( A1 => regs(386), A2 => n113, B1 => regs(1922), 
                           B2 => n161, C1 => regs(898), C2 => n236, ZN => n2168
                           );
   U2803 : AOI22_X1 port map( A1 => regs(1410), A2 => n1, B1 => regs(2434), B2 
                           => n364, ZN => n2167);
   U2804 : NAND2_X1 port map( A1 => n2169, A2 => n2170, ZN => 
                           curr_proc_regs(385));
   U2805 : AOI222_X1 port map( A1 => regs(385), A2 => n113, B1 => regs(1921), 
                           B2 => n161, C1 => regs(897), C2 => n236, ZN => n2170
                           );
   U2806 : AOI22_X1 port map( A1 => regs(1409), A2 => n1, B1 => regs(2433), B2 
                           => n364, ZN => n2169);
   U2807 : NAND2_X1 port map( A1 => n2171, A2 => n2172, ZN => 
                           curr_proc_regs(384));
   U2808 : AOI222_X1 port map( A1 => regs(384), A2 => n113, B1 => regs(1920), 
                           B2 => n161, C1 => regs(896), C2 => n236, ZN => n2172
                           );
   U2809 : AOI22_X1 port map( A1 => regs(1408), A2 => n6, B1 => regs(2432), B2 
                           => n365, ZN => n2171);
   U2810 : NAND2_X1 port map( A1 => n2173, A2 => n2174, ZN => 
                           curr_proc_regs(383));
   U2811 : AOI222_X1 port map( A1 => regs(383), A2 => n113, B1 => regs(1919), 
                           B2 => n161, C1 => regs(895), C2 => n236, ZN => n2174
                           );
   U2812 : AOI22_X1 port map( A1 => regs(1407), A2 => n17, B1 => regs(2431), B2
                           => n365, ZN => n2173);
   U2813 : NAND2_X1 port map( A1 => n2175, A2 => n2176, ZN => 
                           curr_proc_regs(382));
   U2814 : AOI222_X1 port map( A1 => regs(382), A2 => n113, B1 => regs(1918), 
                           B2 => n161, C1 => regs(894), C2 => n236, ZN => n2176
                           );
   U2815 : AOI22_X1 port map( A1 => regs(1406), A2 => n17, B1 => regs(2430), B2
                           => n354, ZN => n2175);
   U2816 : NAND2_X1 port map( A1 => n2177, A2 => n2178, ZN => 
                           curr_proc_regs(381));
   U2817 : AOI222_X1 port map( A1 => regs(381), A2 => n113, B1 => regs(1917), 
                           B2 => n161, C1 => regs(893), C2 => n236, ZN => n2178
                           );
   U2818 : AOI22_X1 port map( A1 => regs(1405), A2 => n17, B1 => regs(2429), B2
                           => n349, ZN => n2177);
   U2819 : NAND2_X1 port map( A1 => n2179, A2 => n2180, ZN => 
                           curr_proc_regs(380));
   U2820 : AOI222_X1 port map( A1 => regs(380), A2 => n113, B1 => regs(1916), 
                           B2 => n161, C1 => regs(892), C2 => n236, ZN => n2180
                           );
   U2821 : AOI22_X1 port map( A1 => regs(1404), A2 => n17, B1 => regs(2428), B2
                           => n348, ZN => n2179);
   U2822 : NAND2_X1 port map( A1 => n2181, A2 => n2182, ZN => 
                           curr_proc_regs(379));
   U2823 : AOI222_X1 port map( A1 => regs(379), A2 => n113, B1 => regs(1915), 
                           B2 => n161, C1 => regs(891), C2 => n236, ZN => n2182
                           );
   U2824 : AOI22_X1 port map( A1 => regs(1403), A2 => n17, B1 => regs(2427), B2
                           => n348, ZN => n2181);
   U2825 : NAND2_X1 port map( A1 => n2183, A2 => n2184, ZN => 
                           curr_proc_regs(378));
   U2826 : AOI222_X1 port map( A1 => regs(378), A2 => n113, B1 => regs(1914), 
                           B2 => n161, C1 => regs(890), C2 => n236, ZN => n2184
                           );
   U2827 : AOI22_X1 port map( A1 => regs(1402), A2 => n17, B1 => regs(2426), B2
                           => n348, ZN => n2183);
   U2828 : NAND2_X1 port map( A1 => n2185, A2 => n2186, ZN => 
                           curr_proc_regs(377));
   U2829 : AOI222_X1 port map( A1 => regs(377), A2 => n113, B1 => regs(1913), 
                           B2 => n161, C1 => regs(889), C2 => n236, ZN => n2186
                           );
   U2830 : AOI22_X1 port map( A1 => regs(1401), A2 => n17, B1 => regs(2425), B2
                           => n348, ZN => n2185);
   U2831 : NAND2_X1 port map( A1 => n2187, A2 => n2188, ZN => 
                           curr_proc_regs(376));
   U2832 : AOI222_X1 port map( A1 => regs(376), A2 => n113, B1 => regs(1912), 
                           B2 => n161, C1 => regs(888), C2 => n236, ZN => n2188
                           );
   U2833 : AOI22_X1 port map( A1 => regs(1400), A2 => n17, B1 => regs(2424), B2
                           => n348, ZN => n2187);
   U2834 : NAND2_X1 port map( A1 => n2189, A2 => n2190, ZN => 
                           curr_proc_regs(375));
   U2835 : AOI222_X1 port map( A1 => regs(375), A2 => n114, B1 => regs(1911), 
                           B2 => n160, C1 => regs(887), C2 => n235, ZN => n2190
                           );
   U2836 : AOI22_X1 port map( A1 => regs(1399), A2 => n17, B1 => regs(2423), B2
                           => n348, ZN => n2189);
   U2837 : NAND2_X1 port map( A1 => n2191, A2 => n2192, ZN => 
                           curr_proc_regs(374));
   U2838 : AOI222_X1 port map( A1 => regs(374), A2 => n114, B1 => regs(1910), 
                           B2 => n160, C1 => regs(886), C2 => n235, ZN => n2192
                           );
   U2839 : AOI22_X1 port map( A1 => regs(1398), A2 => n17, B1 => regs(2422), B2
                           => n348, ZN => n2191);
   U2840 : NAND2_X1 port map( A1 => n2193, A2 => n2194, ZN => 
                           curr_proc_regs(373));
   U2841 : AOI222_X1 port map( A1 => regs(373), A2 => n114, B1 => regs(1909), 
                           B2 => n160, C1 => regs(885), C2 => n235, ZN => n2194
                           );
   U2842 : AOI22_X1 port map( A1 => regs(1397), A2 => n17, B1 => regs(2421), B2
                           => n348, ZN => n2193);
   U2843 : NAND2_X1 port map( A1 => n2195, A2 => n2196, ZN => 
                           curr_proc_regs(372));
   U2844 : AOI222_X1 port map( A1 => regs(372), A2 => n114, B1 => regs(1908), 
                           B2 => n160, C1 => regs(884), C2 => n235, ZN => n2196
                           );
   U2845 : AOI22_X1 port map( A1 => regs(1396), A2 => n17, B1 => regs(2420), B2
                           => n348, ZN => n2195);
   U2846 : NAND2_X1 port map( A1 => n2197, A2 => n2198, ZN => 
                           curr_proc_regs(371));
   U2847 : AOI222_X1 port map( A1 => regs(371), A2 => n114, B1 => regs(1907), 
                           B2 => n160, C1 => regs(883), C2 => n235, ZN => n2198
                           );
   U2848 : AOI22_X1 port map( A1 => regs(1395), A2 => n18, B1 => regs(2419), B2
                           => n348, ZN => n2197);
   U2849 : NAND2_X1 port map( A1 => n2199, A2 => n2200, ZN => 
                           curr_proc_regs(370));
   U2850 : AOI222_X1 port map( A1 => regs(370), A2 => n114, B1 => regs(1906), 
                           B2 => n160, C1 => regs(882), C2 => n235, ZN => n2200
                           );
   U2851 : AOI22_X1 port map( A1 => regs(1394), A2 => n18, B1 => regs(2418), B2
                           => n348, ZN => n2199);
   U2852 : NAND2_X1 port map( A1 => n2201, A2 => n2202, ZN => 
                           curr_proc_regs(369));
   U2853 : AOI222_X1 port map( A1 => regs(369), A2 => n114, B1 => regs(1905), 
                           B2 => n160, C1 => regs(881), C2 => n235, ZN => n2202
                           );
   U2854 : AOI22_X1 port map( A1 => regs(1393), A2 => n18, B1 => regs(2417), B2
                           => n348, ZN => n2201);
   U2855 : NAND2_X1 port map( A1 => n2203, A2 => n2204, ZN => 
                           curr_proc_regs(368));
   U2856 : AOI222_X1 port map( A1 => regs(368), A2 => n114, B1 => regs(1904), 
                           B2 => n160, C1 => regs(880), C2 => n235, ZN => n2204
                           );
   U2857 : AOI22_X1 port map( A1 => regs(1392), A2 => n18, B1 => regs(2416), B2
                           => n347, ZN => n2203);
   U2858 : NAND2_X1 port map( A1 => n2205, A2 => n2206, ZN => 
                           curr_proc_regs(367));
   U2859 : AOI222_X1 port map( A1 => regs(367), A2 => n114, B1 => regs(1903), 
                           B2 => n160, C1 => regs(879), C2 => n235, ZN => n2206
                           );
   U2860 : AOI22_X1 port map( A1 => regs(1391), A2 => n18, B1 => regs(2415), B2
                           => n347, ZN => n2205);
   U2861 : NAND2_X1 port map( A1 => n2207, A2 => n2208, ZN => 
                           curr_proc_regs(366));
   U2862 : AOI222_X1 port map( A1 => regs(366), A2 => n114, B1 => regs(1902), 
                           B2 => n160, C1 => regs(878), C2 => n235, ZN => n2208
                           );
   U2863 : AOI22_X1 port map( A1 => regs(1390), A2 => n18, B1 => regs(2414), B2
                           => n347, ZN => n2207);
   U2864 : NAND2_X1 port map( A1 => n2209, A2 => n2210, ZN => 
                           curr_proc_regs(365));
   U2865 : AOI222_X1 port map( A1 => regs(365), A2 => n114, B1 => regs(1901), 
                           B2 => n160, C1 => regs(877), C2 => n235, ZN => n2210
                           );
   U2866 : AOI22_X1 port map( A1 => regs(1389), A2 => n18, B1 => regs(2413), B2
                           => n347, ZN => n2209);
   U2867 : NAND2_X1 port map( A1 => n2211, A2 => n2212, ZN => 
                           curr_proc_regs(364));
   U2868 : AOI222_X1 port map( A1 => regs(364), A2 => n114, B1 => regs(1900), 
                           B2 => n160, C1 => regs(876), C2 => n235, ZN => n2212
                           );
   U2869 : AOI22_X1 port map( A1 => regs(1388), A2 => n18, B1 => regs(2412), B2
                           => n347, ZN => n2211);
   U2870 : NAND2_X1 port map( A1 => n2213, A2 => n2214, ZN => 
                           curr_proc_regs(363));
   U2871 : AOI222_X1 port map( A1 => regs(363), A2 => n115, B1 => regs(1899), 
                           B2 => n159, C1 => regs(875), C2 => n234, ZN => n2214
                           );
   U2872 : AOI22_X1 port map( A1 => regs(1387), A2 => n18, B1 => regs(2411), B2
                           => n347, ZN => n2213);
   U2873 : NAND2_X1 port map( A1 => n2215, A2 => n2216, ZN => 
                           curr_proc_regs(362));
   U2874 : AOI222_X1 port map( A1 => regs(362), A2 => n115, B1 => regs(1898), 
                           B2 => n159, C1 => regs(874), C2 => n234, ZN => n2216
                           );
   U2875 : AOI22_X1 port map( A1 => regs(1386), A2 => n18, B1 => regs(2410), B2
                           => n347, ZN => n2215);
   U2876 : NAND2_X1 port map( A1 => n2217, A2 => n2218, ZN => 
                           curr_proc_regs(361));
   U2877 : AOI222_X1 port map( A1 => regs(361), A2 => n115, B1 => regs(1897), 
                           B2 => n159, C1 => regs(873), C2 => n234, ZN => n2218
                           );
   U2878 : AOI22_X1 port map( A1 => regs(1385), A2 => n18, B1 => regs(2409), B2
                           => n347, ZN => n2217);
   U2879 : NAND2_X1 port map( A1 => n2219, A2 => n2220, ZN => 
                           curr_proc_regs(360));
   U2880 : AOI222_X1 port map( A1 => regs(360), A2 => n115, B1 => regs(1896), 
                           B2 => n159, C1 => regs(872), C2 => n234, ZN => n2220
                           );
   U2881 : AOI22_X1 port map( A1 => regs(1384), A2 => n18, B1 => regs(2408), B2
                           => n347, ZN => n2219);
   U2882 : NAND2_X1 port map( A1 => n2221, A2 => n2222, ZN => 
                           curr_proc_regs(359));
   U2883 : AOI222_X1 port map( A1 => regs(359), A2 => n115, B1 => regs(1895), 
                           B2 => n159, C1 => regs(871), C2 => n234, ZN => n2222
                           );
   U2884 : AOI22_X1 port map( A1 => regs(1383), A2 => n19, B1 => regs(2407), B2
                           => n347, ZN => n2221);
   U2885 : NAND2_X1 port map( A1 => n2223, A2 => n2224, ZN => 
                           curr_proc_regs(358));
   U2886 : AOI222_X1 port map( A1 => regs(358), A2 => n115, B1 => regs(1894), 
                           B2 => n159, C1 => regs(870), C2 => n234, ZN => n2224
                           );
   U2887 : AOI22_X1 port map( A1 => regs(1382), A2 => n19, B1 => regs(2406), B2
                           => n347, ZN => n2223);
   U2888 : NAND2_X1 port map( A1 => n2225, A2 => n2226, ZN => 
                           curr_proc_regs(357));
   U2889 : AOI222_X1 port map( A1 => regs(357), A2 => n115, B1 => regs(1893), 
                           B2 => n159, C1 => regs(869), C2 => n234, ZN => n2226
                           );
   U2890 : AOI22_X1 port map( A1 => regs(1381), A2 => n19, B1 => regs(2405), B2
                           => n347, ZN => n2225);
   U2891 : NAND2_X1 port map( A1 => n2227, A2 => n2228, ZN => 
                           curr_proc_regs(356));
   U2892 : AOI222_X1 port map( A1 => regs(356), A2 => n115, B1 => regs(1892), 
                           B2 => n159, C1 => regs(868), C2 => n234, ZN => n2228
                           );
   U2893 : AOI22_X1 port map( A1 => regs(1380), A2 => n19, B1 => regs(2404), B2
                           => n346, ZN => n2227);
   U2894 : NAND2_X1 port map( A1 => n2229, A2 => n2230, ZN => 
                           curr_proc_regs(355));
   U2895 : AOI222_X1 port map( A1 => regs(355), A2 => n115, B1 => regs(1891), 
                           B2 => n159, C1 => regs(867), C2 => n234, ZN => n2230
                           );
   U2896 : AOI22_X1 port map( A1 => regs(1379), A2 => n19, B1 => regs(2403), B2
                           => n346, ZN => n2229);
   U2897 : NAND2_X1 port map( A1 => n2231, A2 => n2232, ZN => 
                           curr_proc_regs(354));
   U2898 : AOI222_X1 port map( A1 => regs(354), A2 => n115, B1 => regs(1890), 
                           B2 => n159, C1 => regs(866), C2 => n234, ZN => n2232
                           );
   U2899 : AOI22_X1 port map( A1 => regs(1378), A2 => n19, B1 => regs(2402), B2
                           => n346, ZN => n2231);
   U2900 : NAND2_X1 port map( A1 => n2233, A2 => n2234, ZN => 
                           curr_proc_regs(353));
   U2901 : AOI222_X1 port map( A1 => regs(353), A2 => n115, B1 => regs(1889), 
                           B2 => n159, C1 => regs(865), C2 => n234, ZN => n2234
                           );
   U2902 : AOI22_X1 port map( A1 => regs(1377), A2 => n19, B1 => regs(2401), B2
                           => n346, ZN => n2233);
   U2903 : NAND2_X1 port map( A1 => n2235, A2 => n2236, ZN => 
                           curr_proc_regs(352));
   U2904 : AOI222_X1 port map( A1 => regs(352), A2 => n116, B1 => regs(1888), 
                           B2 => n159, C1 => regs(864), C2 => n234, ZN => n2236
                           );
   U2905 : AOI22_X1 port map( A1 => regs(1376), A2 => n19, B1 => regs(2400), B2
                           => n346, ZN => n2235);
   U2906 : NAND2_X1 port map( A1 => n2237, A2 => n2238, ZN => 
                           curr_proc_regs(351));
   U2907 : AOI222_X1 port map( A1 => regs(351), A2 => n116, B1 => regs(1887), 
                           B2 => n158, C1 => regs(863), C2 => n233, ZN => n2238
                           );
   U2908 : AOI22_X1 port map( A1 => regs(1375), A2 => n19, B1 => regs(2399), B2
                           => n346, ZN => n2237);
   U2909 : NAND2_X1 port map( A1 => n2239, A2 => n2240, ZN => 
                           curr_proc_regs(350));
   U2910 : AOI222_X1 port map( A1 => regs(350), A2 => n116, B1 => regs(1886), 
                           B2 => n158, C1 => regs(862), C2 => n233, ZN => n2240
                           );
   U2911 : AOI22_X1 port map( A1 => regs(1374), A2 => n19, B1 => regs(2398), B2
                           => n346, ZN => n2239);
   U2912 : NAND2_X1 port map( A1 => n2241, A2 => n2242, ZN => 
                           curr_proc_regs(349));
   U2913 : AOI222_X1 port map( A1 => regs(349), A2 => n116, B1 => regs(1885), 
                           B2 => n158, C1 => regs(861), C2 => n233, ZN => n2242
                           );
   U2914 : AOI22_X1 port map( A1 => regs(1373), A2 => n19, B1 => regs(2397), B2
                           => n346, ZN => n2241);
   U2915 : NAND2_X1 port map( A1 => n2243, A2 => n2244, ZN => 
                           curr_proc_regs(348));
   U2916 : AOI222_X1 port map( A1 => regs(348), A2 => n116, B1 => regs(1884), 
                           B2 => n158, C1 => regs(860), C2 => n233, ZN => n2244
                           );
   U2917 : AOI22_X1 port map( A1 => regs(1372), A2 => n20, B1 => regs(2396), B2
                           => n346, ZN => n2243);
   U2918 : NAND2_X1 port map( A1 => n2245, A2 => n2246, ZN => 
                           curr_proc_regs(347));
   U2919 : AOI222_X1 port map( A1 => regs(347), A2 => n116, B1 => regs(1883), 
                           B2 => n158, C1 => regs(859), C2 => n233, ZN => n2246
                           );
   U2920 : AOI22_X1 port map( A1 => regs(1371), A2 => n20, B1 => regs(2395), B2
                           => n346, ZN => n2245);
   U2921 : NAND2_X1 port map( A1 => n2247, A2 => n2248, ZN => 
                           curr_proc_regs(346));
   U2922 : AOI222_X1 port map( A1 => regs(346), A2 => n116, B1 => regs(1882), 
                           B2 => n158, C1 => regs(858), C2 => n233, ZN => n2248
                           );
   U2923 : AOI22_X1 port map( A1 => regs(1370), A2 => n20, B1 => regs(2394), B2
                           => n346, ZN => n2247);
   U2924 : NAND2_X1 port map( A1 => n2249, A2 => n2250, ZN => 
                           curr_proc_regs(345));
   U2925 : AOI222_X1 port map( A1 => regs(345), A2 => n116, B1 => regs(1881), 
                           B2 => n158, C1 => regs(857), C2 => n233, ZN => n2250
                           );
   U2926 : AOI22_X1 port map( A1 => regs(1369), A2 => n20, B1 => regs(2393), B2
                           => n345, ZN => n2249);
   U2927 : NAND2_X1 port map( A1 => n2251, A2 => n2252, ZN => 
                           curr_proc_regs(344));
   U2928 : AOI222_X1 port map( A1 => regs(344), A2 => n116, B1 => regs(1880), 
                           B2 => n158, C1 => regs(856), C2 => n233, ZN => n2252
                           );
   U2929 : AOI22_X1 port map( A1 => regs(1368), A2 => n20, B1 => regs(2392), B2
                           => n345, ZN => n2251);
   U2930 : NAND2_X1 port map( A1 => n2253, A2 => n2254, ZN => 
                           curr_proc_regs(343));
   U2931 : AOI222_X1 port map( A1 => regs(343), A2 => n116, B1 => regs(1879), 
                           B2 => n158, C1 => regs(855), C2 => n233, ZN => n2254
                           );
   U2932 : AOI22_X1 port map( A1 => regs(1367), A2 => n20, B1 => regs(2391), B2
                           => n345, ZN => n2253);
   U2933 : NAND2_X1 port map( A1 => n2255, A2 => n2256, ZN => 
                           curr_proc_regs(342));
   U2934 : AOI222_X1 port map( A1 => regs(342), A2 => n116, B1 => regs(1878), 
                           B2 => n158, C1 => regs(854), C2 => n233, ZN => n2256
                           );
   U2935 : AOI22_X1 port map( A1 => regs(1366), A2 => n20, B1 => regs(2390), B2
                           => n345, ZN => n2255);
   U2936 : NAND2_X1 port map( A1 => n2257, A2 => n2258, ZN => 
                           curr_proc_regs(341));
   U2937 : AOI222_X1 port map( A1 => regs(341), A2 => n116, B1 => regs(1877), 
                           B2 => n158, C1 => regs(853), C2 => n233, ZN => n2258
                           );
   U2938 : AOI22_X1 port map( A1 => regs(1365), A2 => n20, B1 => regs(2389), B2
                           => n345, ZN => n2257);
   U2939 : NAND2_X1 port map( A1 => n2259, A2 => n2260, ZN => 
                           curr_proc_regs(340));
   U2940 : AOI222_X1 port map( A1 => regs(340), A2 => n117, B1 => regs(1876), 
                           B2 => n158, C1 => regs(852), C2 => n233, ZN => n2260
                           );
   U2941 : AOI22_X1 port map( A1 => regs(1364), A2 => n20, B1 => regs(2388), B2
                           => n345, ZN => n2259);
   U2942 : NAND2_X1 port map( A1 => n2261, A2 => n2262, ZN => 
                           curr_proc_regs(339));
   U2943 : AOI222_X1 port map( A1 => regs(339), A2 => n117, B1 => regs(1875), 
                           B2 => n157, C1 => regs(851), C2 => n232, ZN => n2262
                           );
   U2944 : AOI22_X1 port map( A1 => regs(1363), A2 => n20, B1 => regs(2387), B2
                           => n345, ZN => n2261);
   U2945 : NAND2_X1 port map( A1 => n2263, A2 => n2264, ZN => 
                           curr_proc_regs(338));
   U2946 : AOI222_X1 port map( A1 => regs(338), A2 => n117, B1 => regs(1874), 
                           B2 => n157, C1 => regs(850), C2 => n232, ZN => n2264
                           );
   U2947 : AOI22_X1 port map( A1 => regs(1362), A2 => n20, B1 => regs(2386), B2
                           => n345, ZN => n2263);
   U2948 : NAND2_X1 port map( A1 => n2265, A2 => n2266, ZN => 
                           curr_proc_regs(337));
   U2949 : AOI222_X1 port map( A1 => regs(337), A2 => n117, B1 => regs(1873), 
                           B2 => n157, C1 => regs(849), C2 => n232, ZN => n2266
                           );
   U2950 : AOI22_X1 port map( A1 => regs(1361), A2 => n20, B1 => regs(2385), B2
                           => n345, ZN => n2265);
   U2951 : NAND2_X1 port map( A1 => n2267, A2 => n2268, ZN => 
                           curr_proc_regs(336));
   U2952 : AOI222_X1 port map( A1 => regs(336), A2 => n117, B1 => regs(1872), 
                           B2 => n157, C1 => regs(848), C2 => n232, ZN => n2268
                           );
   U2953 : AOI22_X1 port map( A1 => regs(1360), A2 => n21, B1 => regs(2384), B2
                           => n345, ZN => n2267);
   U2954 : NAND2_X1 port map( A1 => n2269, A2 => n2270, ZN => 
                           curr_proc_regs(335));
   U2955 : AOI222_X1 port map( A1 => regs(335), A2 => n117, B1 => regs(1871), 
                           B2 => n157, C1 => regs(847), C2 => n232, ZN => n2270
                           );
   U2956 : AOI22_X1 port map( A1 => regs(1359), A2 => n21, B1 => regs(2383), B2
                           => n345, ZN => n2269);
   U2957 : NAND2_X1 port map( A1 => n2271, A2 => n2272, ZN => 
                           curr_proc_regs(334));
   U2958 : AOI222_X1 port map( A1 => regs(334), A2 => n117, B1 => regs(1870), 
                           B2 => n157, C1 => regs(846), C2 => n232, ZN => n2272
                           );
   U2959 : AOI22_X1 port map( A1 => regs(1358), A2 => n21, B1 => regs(2382), B2
                           => n345, ZN => n2271);
   U2960 : NAND2_X1 port map( A1 => n2273, A2 => n2274, ZN => 
                           curr_proc_regs(333));
   U2961 : AOI222_X1 port map( A1 => regs(333), A2 => n117, B1 => regs(1869), 
                           B2 => n157, C1 => regs(845), C2 => n232, ZN => n2274
                           );
   U2962 : AOI22_X1 port map( A1 => regs(1357), A2 => n21, B1 => regs(2381), B2
                           => n344, ZN => n2273);
   U2963 : NAND2_X1 port map( A1 => n2275, A2 => n2276, ZN => 
                           curr_proc_regs(332));
   U2964 : AOI222_X1 port map( A1 => regs(332), A2 => n117, B1 => regs(1868), 
                           B2 => n157, C1 => regs(844), C2 => n232, ZN => n2276
                           );
   U2965 : AOI22_X1 port map( A1 => regs(1356), A2 => n21, B1 => regs(2380), B2
                           => n344, ZN => n2275);
   U2966 : NAND2_X1 port map( A1 => n2277, A2 => n2278, ZN => 
                           curr_proc_regs(331));
   U2967 : AOI222_X1 port map( A1 => regs(331), A2 => n117, B1 => regs(1867), 
                           B2 => n157, C1 => regs(843), C2 => n232, ZN => n2278
                           );
   U2968 : AOI22_X1 port map( A1 => regs(1355), A2 => n21, B1 => regs(2379), B2
                           => n344, ZN => n2277);
   U2969 : NAND2_X1 port map( A1 => n2279, A2 => n2280, ZN => 
                           curr_proc_regs(330));
   U2970 : AOI222_X1 port map( A1 => regs(330), A2 => n117, B1 => regs(1866), 
                           B2 => n157, C1 => regs(842), C2 => n232, ZN => n2280
                           );
   U2971 : AOI22_X1 port map( A1 => regs(1354), A2 => n21, B1 => regs(2378), B2
                           => n344, ZN => n2279);
   U2972 : NAND2_X1 port map( A1 => n2281, A2 => n2282, ZN => 
                           curr_proc_regs(329));
   U2973 : AOI222_X1 port map( A1 => regs(329), A2 => n117, B1 => regs(1865), 
                           B2 => n157, C1 => regs(841), C2 => n232, ZN => n2282
                           );
   U2974 : AOI22_X1 port map( A1 => regs(1353), A2 => n21, B1 => regs(2377), B2
                           => n344, ZN => n2281);
   U2975 : NAND2_X1 port map( A1 => n2283, A2 => n2284, ZN => 
                           curr_proc_regs(328));
   U2976 : AOI222_X1 port map( A1 => regs(328), A2 => n118, B1 => regs(1864), 
                           B2 => n157, C1 => regs(840), C2 => n232, ZN => n2284
                           );
   U2977 : AOI22_X1 port map( A1 => regs(1352), A2 => n21, B1 => regs(2376), B2
                           => n344, ZN => n2283);
   U2978 : NAND2_X1 port map( A1 => n2285, A2 => n2286, ZN => 
                           curr_proc_regs(327));
   U2979 : AOI222_X1 port map( A1 => regs(327), A2 => n118, B1 => regs(1863), 
                           B2 => n156, C1 => regs(839), C2 => n231, ZN => n2286
                           );
   U2980 : AOI22_X1 port map( A1 => regs(1351), A2 => n21, B1 => regs(2375), B2
                           => n344, ZN => n2285);
   U2981 : NAND2_X1 port map( A1 => n2287, A2 => n2288, ZN => 
                           curr_proc_regs(326));
   U2982 : AOI222_X1 port map( A1 => regs(326), A2 => n118, B1 => regs(1862), 
                           B2 => n156, C1 => regs(838), C2 => n231, ZN => n2288
                           );
   U2983 : AOI22_X1 port map( A1 => regs(1350), A2 => n21, B1 => regs(2374), B2
                           => n344, ZN => n2287);
   U2984 : NAND2_X1 port map( A1 => n2289, A2 => n2290, ZN => 
                           curr_proc_regs(325));
   U2985 : AOI222_X1 port map( A1 => regs(325), A2 => n118, B1 => regs(1861), 
                           B2 => n156, C1 => regs(837), C2 => n231, ZN => n2290
                           );
   U2986 : AOI22_X1 port map( A1 => regs(1349), A2 => n21, B1 => regs(2373), B2
                           => n344, ZN => n2289);
   U2987 : NAND2_X1 port map( A1 => n2291, A2 => n2292, ZN => 
                           curr_proc_regs(324));
   U2988 : AOI222_X1 port map( A1 => regs(324), A2 => n118, B1 => regs(1860), 
                           B2 => n156, C1 => regs(836), C2 => n231, ZN => n2292
                           );
   U2989 : AOI22_X1 port map( A1 => regs(1348), A2 => n22, B1 => regs(2372), B2
                           => n344, ZN => n2291);
   U2990 : NAND2_X1 port map( A1 => n2293, A2 => n2294, ZN => 
                           curr_proc_regs(323));
   U2991 : AOI222_X1 port map( A1 => regs(323), A2 => n118, B1 => regs(1859), 
                           B2 => n156, C1 => regs(835), C2 => n231, ZN => n2294
                           );
   U2992 : AOI22_X1 port map( A1 => regs(1347), A2 => n22, B1 => regs(2371), B2
                           => n344, ZN => n2293);
   U2993 : NAND2_X1 port map( A1 => n2295, A2 => n2296, ZN => 
                           curr_proc_regs(322));
   U2994 : AOI222_X1 port map( A1 => regs(322), A2 => n118, B1 => regs(1858), 
                           B2 => n156, C1 => regs(834), C2 => n231, ZN => n2296
                           );
   U2995 : AOI22_X1 port map( A1 => regs(1346), A2 => n22, B1 => regs(2370), B2
                           => n344, ZN => n2295);
   U2996 : NAND2_X1 port map( A1 => n2297, A2 => n2298, ZN => 
                           curr_proc_regs(321));
   U2997 : AOI222_X1 port map( A1 => regs(321), A2 => n118, B1 => regs(1857), 
                           B2 => n156, C1 => regs(833), C2 => n231, ZN => n2298
                           );
   U2998 : AOI22_X1 port map( A1 => regs(1345), A2 => n22, B1 => regs(2369), B2
                           => n343, ZN => n2297);
   U2999 : NAND2_X1 port map( A1 => n2299, A2 => n2300, ZN => 
                           curr_proc_regs(320));
   U3000 : AOI222_X1 port map( A1 => regs(320), A2 => n118, B1 => regs(1856), 
                           B2 => n156, C1 => regs(832), C2 => n231, ZN => n2300
                           );
   U3001 : AOI22_X1 port map( A1 => regs(1344), A2 => n16, B1 => regs(2368), B2
                           => n349, ZN => n2299);
   U3002 : NAND2_X1 port map( A1 => n2301, A2 => n2302, ZN => 
                           curr_proc_regs(319));
   U3003 : AOI222_X1 port map( A1 => regs(319), A2 => n118, B1 => regs(1855), 
                           B2 => n156, C1 => regs(831), C2 => n231, ZN => n2302
                           );
   U3004 : AOI22_X1 port map( A1 => regs(1343), A2 => n16, B1 => regs(2367), B2
                           => n346, ZN => n2301);
   U3005 : NAND2_X1 port map( A1 => n2303, A2 => n2304, ZN => 
                           curr_proc_regs(318));
   U3006 : AOI222_X1 port map( A1 => regs(318), A2 => n118, B1 => regs(1854), 
                           B2 => n156, C1 => regs(830), C2 => n231, ZN => n2304
                           );
   U3007 : AOI22_X1 port map( A1 => regs(1342), A2 => n16, B1 => regs(2366), B2
                           => n349, ZN => n2303);
   U3008 : NAND2_X1 port map( A1 => n2305, A2 => n2306, ZN => 
                           curr_proc_regs(317));
   U3009 : AOI222_X1 port map( A1 => regs(317), A2 => n118, B1 => regs(1853), 
                           B2 => n156, C1 => regs(829), C2 => n231, ZN => n2306
                           );
   U3010 : AOI22_X1 port map( A1 => regs(1341), A2 => n16, B1 => regs(2365), B2
                           => n349, ZN => n2305);
   U3011 : NAND2_X1 port map( A1 => n2307, A2 => n2308, ZN => 
                           curr_proc_regs(316));
   U3012 : AOI222_X1 port map( A1 => regs(316), A2 => n119, B1 => regs(1852), 
                           B2 => n156, C1 => regs(828), C2 => n231, ZN => n2308
                           );
   U3013 : AOI22_X1 port map( A1 => regs(1340), A2 => n16, B1 => regs(2364), B2
                           => n349, ZN => n2307);
   U3014 : NAND2_X1 port map( A1 => n2309, A2 => n2310, ZN => 
                           curr_proc_regs(315));
   U3015 : AOI222_X1 port map( A1 => regs(315), A2 => n119, B1 => regs(1851), 
                           B2 => n155, C1 => regs(827), C2 => n230, ZN => n2310
                           );
   U3016 : AOI22_X1 port map( A1 => regs(1339), A2 => n16, B1 => regs(2363), B2
                           => n349, ZN => n2309);
   U3017 : NAND2_X1 port map( A1 => n2311, A2 => n2312, ZN => 
                           curr_proc_regs(314));
   U3018 : AOI222_X1 port map( A1 => regs(314), A2 => n119, B1 => regs(1850), 
                           B2 => n155, C1 => regs(826), C2 => n230, ZN => n2312
                           );
   U3019 : AOI22_X1 port map( A1 => regs(1338), A2 => n16, B1 => regs(2362), B2
                           => n349, ZN => n2311);
   U3020 : NAND2_X1 port map( A1 => n2313, A2 => n2314, ZN => 
                           curr_proc_regs(313));
   U3021 : AOI222_X1 port map( A1 => regs(313), A2 => n119, B1 => regs(1849), 
                           B2 => n155, C1 => regs(825), C2 => n230, ZN => n2314
                           );
   U3022 : AOI22_X1 port map( A1 => regs(1337), A2 => n16, B1 => regs(2361), B2
                           => n349, ZN => n2313);
   U3023 : NAND2_X1 port map( A1 => n2315, A2 => n2316, ZN => 
                           curr_proc_regs(312));
   U3024 : AOI222_X1 port map( A1 => regs(312), A2 => n119, B1 => regs(1848), 
                           B2 => n155, C1 => regs(824), C2 => n230, ZN => n2316
                           );
   U3025 : AOI22_X1 port map( A1 => regs(1336), A2 => n16, B1 => regs(2360), B2
                           => n349, ZN => n2315);
   U3026 : NAND2_X1 port map( A1 => n2317, A2 => n2318, ZN => 
                           curr_proc_regs(311));
   U3027 : AOI222_X1 port map( A1 => regs(311), A2 => n119, B1 => regs(1847), 
                           B2 => n155, C1 => regs(823), C2 => n230, ZN => n2318
                           );
   U3028 : AOI22_X1 port map( A1 => regs(1335), A2 => n16, B1 => regs(2359), B2
                           => n349, ZN => n2317);
   U3029 : NAND2_X1 port map( A1 => n2319, A2 => n2320, ZN => 
                           curr_proc_regs(310));
   U3030 : AOI222_X1 port map( A1 => regs(310), A2 => n119, B1 => regs(1846), 
                           B2 => n155, C1 => regs(822), C2 => n230, ZN => n2320
                           );
   U3031 : AOI22_X1 port map( A1 => regs(1334), A2 => n16, B1 => regs(2358), B2
                           => n349, ZN => n2319);
   U3032 : NAND2_X1 port map( A1 => n2321, A2 => n2322, ZN => 
                           curr_proc_regs(309));
   U3033 : AOI222_X1 port map( A1 => regs(309), A2 => n119, B1 => regs(1845), 
                           B2 => n155, C1 => regs(821), C2 => n230, ZN => n2322
                           );
   U3034 : AOI22_X1 port map( A1 => regs(1333), A2 => n16, B1 => regs(2357), B2
                           => n349, ZN => n2321);
   U3035 : NAND2_X1 port map( A1 => n2323, A2 => n2324, ZN => 
                           curr_proc_regs(308));
   U3036 : AOI222_X1 port map( A1 => regs(308), A2 => n119, B1 => regs(1844), 
                           B2 => n155, C1 => regs(820), C2 => n230, ZN => n2324
                           );
   U3037 : AOI22_X1 port map( A1 => regs(1332), A2 => n15, B1 => regs(2356), B2
                           => n350, ZN => n2323);
   U3038 : NAND2_X1 port map( A1 => n2325, A2 => n2326, ZN => 
                           curr_proc_regs(307));
   U3039 : AOI222_X1 port map( A1 => regs(307), A2 => n119, B1 => regs(1843), 
                           B2 => n155, C1 => regs(819), C2 => n230, ZN => n2326
                           );
   U3040 : AOI22_X1 port map( A1 => regs(1331), A2 => n15, B1 => regs(2355), B2
                           => n350, ZN => n2325);
   U3041 : NAND2_X1 port map( A1 => n2327, A2 => n2328, ZN => 
                           curr_proc_regs(306));
   U3042 : AOI222_X1 port map( A1 => regs(306), A2 => n119, B1 => regs(1842), 
                           B2 => n155, C1 => regs(818), C2 => n230, ZN => n2328
                           );
   U3043 : AOI22_X1 port map( A1 => regs(1330), A2 => n15, B1 => regs(2354), B2
                           => n350, ZN => n2327);
   U3044 : NAND2_X1 port map( A1 => n2329, A2 => n2330, ZN => 
                           curr_proc_regs(305));
   U3045 : AOI222_X1 port map( A1 => regs(305), A2 => n119, B1 => regs(1841), 
                           B2 => n155, C1 => regs(817), C2 => n230, ZN => n2330
                           );
   U3046 : AOI22_X1 port map( A1 => regs(1329), A2 => n15, B1 => regs(2353), B2
                           => n350, ZN => n2329);
   U3047 : NAND2_X1 port map( A1 => n2331, A2 => n2332, ZN => 
                           curr_proc_regs(304));
   U3048 : AOI222_X1 port map( A1 => regs(304), A2 => n120, B1 => regs(1840), 
                           B2 => n155, C1 => regs(816), C2 => n230, ZN => n2332
                           );
   U3049 : AOI22_X1 port map( A1 => regs(1328), A2 => n15, B1 => regs(2352), B2
                           => n350, ZN => n2331);
   U3050 : NAND2_X1 port map( A1 => n2333, A2 => n2334, ZN => 
                           curr_proc_regs(303));
   U3051 : AOI222_X1 port map( A1 => regs(303), A2 => n120, B1 => regs(1839), 
                           B2 => n154, C1 => regs(815), C2 => n229, ZN => n2334
                           );
   U3052 : AOI22_X1 port map( A1 => regs(1327), A2 => n15, B1 => regs(2351), B2
                           => n350, ZN => n2333);
   U3053 : NAND2_X1 port map( A1 => n2335, A2 => n2336, ZN => 
                           curr_proc_regs(302));
   U3054 : AOI222_X1 port map( A1 => regs(302), A2 => n120, B1 => regs(1838), 
                           B2 => n154, C1 => regs(814), C2 => n229, ZN => n2336
                           );
   U3055 : AOI22_X1 port map( A1 => regs(1326), A2 => n15, B1 => regs(2350), B2
                           => n350, ZN => n2335);
   U3056 : NAND2_X1 port map( A1 => n2337, A2 => n2338, ZN => 
                           curr_proc_regs(301));
   U3057 : AOI222_X1 port map( A1 => regs(301), A2 => n120, B1 => regs(1837), 
                           B2 => n154, C1 => regs(813), C2 => n229, ZN => n2338
                           );
   U3058 : AOI22_X1 port map( A1 => regs(1325), A2 => n15, B1 => regs(2349), B2
                           => n350, ZN => n2337);
   U3059 : NAND2_X1 port map( A1 => n2339, A2 => n2340, ZN => 
                           curr_proc_regs(300));
   U3060 : AOI222_X1 port map( A1 => regs(300), A2 => n120, B1 => regs(1836), 
                           B2 => n154, C1 => regs(812), C2 => n229, ZN => n2340
                           );
   U3061 : AOI22_X1 port map( A1 => regs(1324), A2 => n15, B1 => regs(2348), B2
                           => n350, ZN => n2339);
   U3062 : NAND2_X1 port map( A1 => n2341, A2 => n2342, ZN => 
                           curr_proc_regs(299));
   U3063 : AOI222_X1 port map( A1 => regs(299), A2 => n120, B1 => regs(1835), 
                           B2 => n154, C1 => regs(811), C2 => n229, ZN => n2342
                           );
   U3064 : AOI22_X1 port map( A1 => regs(1323), A2 => n15, B1 => regs(2347), B2
                           => n350, ZN => n2341);
   U3065 : NAND2_X1 port map( A1 => n2343, A2 => n2344, ZN => 
                           curr_proc_regs(298));
   U3066 : AOI222_X1 port map( A1 => regs(298), A2 => n120, B1 => regs(1834), 
                           B2 => n154, C1 => regs(810), C2 => n229, ZN => n2344
                           );
   U3067 : AOI22_X1 port map( A1 => regs(1322), A2 => n15, B1 => regs(2346), B2
                           => n350, ZN => n2343);
   U3068 : NAND2_X1 port map( A1 => n2345, A2 => n2346, ZN => 
                           curr_proc_regs(297));
   U3069 : AOI222_X1 port map( A1 => regs(297), A2 => n120, B1 => regs(1833), 
                           B2 => n154, C1 => regs(809), C2 => n229, ZN => n2346
                           );
   U3070 : AOI22_X1 port map( A1 => regs(1321), A2 => n15, B1 => regs(2345), B2
                           => n350, ZN => n2345);
   U3071 : NAND2_X1 port map( A1 => n2347, A2 => n2348, ZN => 
                           curr_proc_regs(296));
   U3072 : AOI222_X1 port map( A1 => regs(296), A2 => n120, B1 => regs(1832), 
                           B2 => n154, C1 => regs(808), C2 => n229, ZN => n2348
                           );
   U3073 : AOI22_X1 port map( A1 => regs(1320), A2 => n14, B1 => regs(2344), B2
                           => n351, ZN => n2347);
   U3074 : NAND2_X1 port map( A1 => n2349, A2 => n2350, ZN => 
                           curr_proc_regs(295));
   U3075 : AOI222_X1 port map( A1 => regs(295), A2 => n120, B1 => regs(1831), 
                           B2 => n154, C1 => regs(807), C2 => n229, ZN => n2350
                           );
   U3076 : AOI22_X1 port map( A1 => regs(1319), A2 => n14, B1 => regs(2343), B2
                           => n351, ZN => n2349);
   U3077 : NAND2_X1 port map( A1 => n2351, A2 => n2352, ZN => 
                           curr_proc_regs(294));
   U3078 : AOI222_X1 port map( A1 => regs(294), A2 => n120, B1 => regs(1830), 
                           B2 => n154, C1 => regs(806), C2 => n229, ZN => n2352
                           );
   U3079 : AOI22_X1 port map( A1 => regs(1318), A2 => n14, B1 => regs(2342), B2
                           => n351, ZN => n2351);
   U3080 : NAND2_X1 port map( A1 => n2353, A2 => n2354, ZN => 
                           curr_proc_regs(293));
   U3081 : AOI222_X1 port map( A1 => regs(293), A2 => n120, B1 => regs(1829), 
                           B2 => n154, C1 => regs(805), C2 => n229, ZN => n2354
                           );
   U3082 : AOI22_X1 port map( A1 => regs(1317), A2 => n14, B1 => regs(2341), B2
                           => n351, ZN => n2353);
   U3083 : NAND2_X1 port map( A1 => n2355, A2 => n2356, ZN => 
                           curr_proc_regs(292));
   U3084 : AOI222_X1 port map( A1 => regs(292), A2 => n121, B1 => regs(1828), 
                           B2 => n154, C1 => regs(804), C2 => n229, ZN => n2356
                           );
   U3085 : AOI22_X1 port map( A1 => regs(1316), A2 => n14, B1 => regs(2340), B2
                           => n351, ZN => n2355);
   U3086 : NAND2_X1 port map( A1 => n2357, A2 => n2358, ZN => 
                           curr_proc_regs(291));
   U3087 : AOI222_X1 port map( A1 => regs(291), A2 => n121, B1 => regs(1827), 
                           B2 => n153, C1 => regs(803), C2 => n228, ZN => n2358
                           );
   U3088 : AOI22_X1 port map( A1 => regs(1315), A2 => n14, B1 => regs(2339), B2
                           => n351, ZN => n2357);
   U3089 : NAND2_X1 port map( A1 => n2359, A2 => n2360, ZN => 
                           curr_proc_regs(290));
   U3090 : AOI222_X1 port map( A1 => regs(290), A2 => n121, B1 => regs(1826), 
                           B2 => n153, C1 => regs(802), C2 => n228, ZN => n2360
                           );
   U3091 : AOI22_X1 port map( A1 => regs(1314), A2 => n14, B1 => regs(2338), B2
                           => n351, ZN => n2359);
   U3092 : NAND2_X1 port map( A1 => n2361, A2 => n2362, ZN => 
                           curr_proc_regs(289));
   U3093 : AOI222_X1 port map( A1 => regs(289), A2 => n121, B1 => regs(1825), 
                           B2 => n153, C1 => regs(801), C2 => n228, ZN => n2362
                           );
   U3094 : AOI22_X1 port map( A1 => regs(1313), A2 => n14, B1 => regs(2337), B2
                           => n351, ZN => n2361);
   U3095 : NAND2_X1 port map( A1 => n2363, A2 => n2364, ZN => 
                           curr_proc_regs(288));
   U3096 : AOI222_X1 port map( A1 => regs(288), A2 => n121, B1 => regs(1824), 
                           B2 => n153, C1 => regs(800), C2 => n228, ZN => n2364
                           );
   U3097 : AOI22_X1 port map( A1 => regs(1312), A2 => n14, B1 => regs(2336), B2
                           => n351, ZN => n2363);
   U3098 : NAND2_X1 port map( A1 => n2365, A2 => n2366, ZN => 
                           curr_proc_regs(287));
   U3099 : AOI222_X1 port map( A1 => regs(287), A2 => n121, B1 => regs(1823), 
                           B2 => n153, C1 => regs(799), C2 => n228, ZN => n2366
                           );
   U3100 : AOI22_X1 port map( A1 => regs(1311), A2 => n14, B1 => regs(2335), B2
                           => n351, ZN => n2365);
   U3101 : NAND2_X1 port map( A1 => n2367, A2 => n2368, ZN => 
                           curr_proc_regs(286));
   U3102 : AOI222_X1 port map( A1 => regs(286), A2 => n121, B1 => regs(1822), 
                           B2 => n153, C1 => regs(798), C2 => n228, ZN => n2368
                           );
   U3103 : AOI22_X1 port map( A1 => regs(1310), A2 => n14, B1 => regs(2334), B2
                           => n351, ZN => n2367);
   U3104 : NAND2_X1 port map( A1 => n2369, A2 => n2370, ZN => 
                           curr_proc_regs(285));
   U3105 : AOI222_X1 port map( A1 => regs(285), A2 => n121, B1 => regs(1821), 
                           B2 => n153, C1 => regs(797), C2 => n228, ZN => n2370
                           );
   U3106 : AOI22_X1 port map( A1 => regs(1309), A2 => n14, B1 => regs(2333), B2
                           => n351, ZN => n2369);
   U3107 : NAND2_X1 port map( A1 => n2371, A2 => n2372, ZN => 
                           curr_proc_regs(284));
   U3108 : AOI222_X1 port map( A1 => regs(284), A2 => n121, B1 => regs(1820), 
                           B2 => n153, C1 => regs(796), C2 => n228, ZN => n2372
                           );
   U3109 : AOI22_X1 port map( A1 => regs(1308), A2 => n13, B1 => regs(2332), B2
                           => n352, ZN => n2371);
   U3110 : NAND2_X1 port map( A1 => n2373, A2 => n2374, ZN => 
                           curr_proc_regs(283));
   U3111 : AOI222_X1 port map( A1 => regs(283), A2 => n121, B1 => regs(1819), 
                           B2 => n153, C1 => regs(795), C2 => n228, ZN => n2374
                           );
   U3112 : AOI22_X1 port map( A1 => regs(1307), A2 => n13, B1 => regs(2331), B2
                           => n352, ZN => n2373);
   U3113 : NAND2_X1 port map( A1 => n2375, A2 => n2376, ZN => 
                           curr_proc_regs(282));
   U3114 : AOI222_X1 port map( A1 => regs(282), A2 => n121, B1 => regs(1818), 
                           B2 => n153, C1 => regs(794), C2 => n228, ZN => n2376
                           );
   U3115 : AOI22_X1 port map( A1 => regs(1306), A2 => n13, B1 => regs(2330), B2
                           => n352, ZN => n2375);
   U3116 : NAND2_X1 port map( A1 => n2377, A2 => n2378, ZN => 
                           curr_proc_regs(281));
   U3117 : AOI222_X1 port map( A1 => regs(281), A2 => n121, B1 => regs(1817), 
                           B2 => n153, C1 => regs(793), C2 => n228, ZN => n2378
                           );
   U3118 : AOI22_X1 port map( A1 => regs(1305), A2 => n13, B1 => regs(2329), B2
                           => n352, ZN => n2377);
   U3119 : NAND2_X1 port map( A1 => n2379, A2 => n2380, ZN => 
                           curr_proc_regs(280));
   U3120 : AOI222_X1 port map( A1 => regs(280), A2 => n122, B1 => regs(1816), 
                           B2 => n153, C1 => regs(792), C2 => n228, ZN => n2380
                           );
   U3121 : AOI22_X1 port map( A1 => regs(1304), A2 => n13, B1 => regs(2328), B2
                           => n352, ZN => n2379);
   U3122 : NAND2_X1 port map( A1 => n2381, A2 => n2382, ZN => 
                           curr_proc_regs(279));
   U3123 : AOI222_X1 port map( A1 => regs(279), A2 => n122, B1 => regs(1815), 
                           B2 => n152, C1 => regs(791), C2 => n227, ZN => n2382
                           );
   U3124 : AOI22_X1 port map( A1 => regs(1303), A2 => n13, B1 => regs(2327), B2
                           => n352, ZN => n2381);
   U3125 : NAND2_X1 port map( A1 => n2383, A2 => n2384, ZN => 
                           curr_proc_regs(278));
   U3126 : AOI222_X1 port map( A1 => regs(278), A2 => n122, B1 => regs(1814), 
                           B2 => n152, C1 => regs(790), C2 => n227, ZN => n2384
                           );
   U3127 : AOI22_X1 port map( A1 => regs(1302), A2 => n13, B1 => regs(2326), B2
                           => n352, ZN => n2383);
   U3128 : NAND2_X1 port map( A1 => n2385, A2 => n2386, ZN => 
                           curr_proc_regs(277));
   U3129 : AOI222_X1 port map( A1 => regs(277), A2 => n122, B1 => regs(1813), 
                           B2 => n152, C1 => regs(789), C2 => n227, ZN => n2386
                           );
   U3130 : AOI22_X1 port map( A1 => regs(1301), A2 => n13, B1 => regs(2325), B2
                           => n352, ZN => n2385);
   U3131 : NAND2_X1 port map( A1 => n2387, A2 => n2388, ZN => 
                           curr_proc_regs(276));
   U3132 : AOI222_X1 port map( A1 => regs(276), A2 => n122, B1 => regs(1812), 
                           B2 => n152, C1 => regs(788), C2 => n227, ZN => n2388
                           );
   U3133 : AOI22_X1 port map( A1 => regs(1300), A2 => n13, B1 => regs(2324), B2
                           => n352, ZN => n2387);
   U3134 : NAND2_X1 port map( A1 => n2389, A2 => n2390, ZN => 
                           curr_proc_regs(275));
   U3135 : AOI222_X1 port map( A1 => regs(275), A2 => n122, B1 => regs(1811), 
                           B2 => n152, C1 => regs(787), C2 => n227, ZN => n2390
                           );
   U3136 : AOI22_X1 port map( A1 => regs(1299), A2 => n13, B1 => regs(2323), B2
                           => n352, ZN => n2389);
   U3137 : NAND2_X1 port map( A1 => n2391, A2 => n2392, ZN => 
                           curr_proc_regs(274));
   U3138 : AOI222_X1 port map( A1 => regs(274), A2 => n122, B1 => regs(1810), 
                           B2 => n152, C1 => regs(786), C2 => n227, ZN => n2392
                           );
   U3139 : AOI22_X1 port map( A1 => regs(1298), A2 => n13, B1 => regs(2322), B2
                           => n352, ZN => n2391);
   U3140 : NAND2_X1 port map( A1 => n2393, A2 => n2394, ZN => 
                           curr_proc_regs(273));
   U3141 : AOI222_X1 port map( A1 => regs(273), A2 => n122, B1 => regs(1809), 
                           B2 => n152, C1 => regs(785), C2 => n227, ZN => n2394
                           );
   U3142 : AOI22_X1 port map( A1 => regs(1297), A2 => n13, B1 => regs(2321), B2
                           => n352, ZN => n2393);
   U3143 : NAND2_X1 port map( A1 => n2395, A2 => n2396, ZN => 
                           curr_proc_regs(272));
   U3144 : AOI222_X1 port map( A1 => regs(272), A2 => n122, B1 => regs(1808), 
                           B2 => n152, C1 => regs(784), C2 => n227, ZN => n2396
                           );
   U3145 : AOI22_X1 port map( A1 => regs(1296), A2 => n12, B1 => regs(2320), B2
                           => n353, ZN => n2395);
   U3146 : NAND2_X1 port map( A1 => n2397, A2 => n2398, ZN => 
                           curr_proc_regs(271));
   U3147 : AOI222_X1 port map( A1 => regs(271), A2 => n122, B1 => regs(1807), 
                           B2 => n152, C1 => regs(783), C2 => n227, ZN => n2398
                           );
   U3148 : AOI22_X1 port map( A1 => regs(1295), A2 => n12, B1 => regs(2319), B2
                           => n353, ZN => n2397);
   U3149 : NAND2_X1 port map( A1 => n2399, A2 => n2400, ZN => 
                           curr_proc_regs(270));
   U3150 : AOI222_X1 port map( A1 => regs(270), A2 => n122, B1 => regs(1806), 
                           B2 => n152, C1 => regs(782), C2 => n227, ZN => n2400
                           );
   U3151 : AOI22_X1 port map( A1 => regs(1294), A2 => n12, B1 => regs(2318), B2
                           => n353, ZN => n2399);
   U3152 : NAND2_X1 port map( A1 => n2401, A2 => n2402, ZN => 
                           curr_proc_regs(269));
   U3153 : AOI222_X1 port map( A1 => regs(269), A2 => n122, B1 => regs(1805), 
                           B2 => n152, C1 => regs(781), C2 => n227, ZN => n2402
                           );
   U3154 : AOI22_X1 port map( A1 => regs(1293), A2 => n12, B1 => regs(2317), B2
                           => n353, ZN => n2401);
   U3155 : NAND2_X1 port map( A1 => n2403, A2 => n2404, ZN => 
                           curr_proc_regs(268));
   U3156 : AOI222_X1 port map( A1 => regs(268), A2 => n123, B1 => regs(1804), 
                           B2 => n152, C1 => regs(780), C2 => n227, ZN => n2404
                           );
   U3157 : AOI22_X1 port map( A1 => regs(1292), A2 => n12, B1 => regs(2316), B2
                           => n353, ZN => n2403);
   U3158 : NAND2_X1 port map( A1 => n2405, A2 => n2406, ZN => 
                           curr_proc_regs(267));
   U3159 : AOI222_X1 port map( A1 => regs(267), A2 => n123, B1 => regs(1803), 
                           B2 => n151, C1 => regs(779), C2 => n226, ZN => n2406
                           );
   U3160 : AOI22_X1 port map( A1 => regs(1291), A2 => n12, B1 => regs(2315), B2
                           => n353, ZN => n2405);
   U3161 : NAND2_X1 port map( A1 => n2407, A2 => n2408, ZN => 
                           curr_proc_regs(266));
   U3162 : AOI222_X1 port map( A1 => regs(266), A2 => n123, B1 => regs(1802), 
                           B2 => n151, C1 => regs(778), C2 => n226, ZN => n2408
                           );
   U3163 : AOI22_X1 port map( A1 => regs(1290), A2 => n12, B1 => regs(2314), B2
                           => n353, ZN => n2407);
   U3164 : NAND2_X1 port map( A1 => n2409, A2 => n2410, ZN => 
                           curr_proc_regs(265));
   U3165 : AOI222_X1 port map( A1 => regs(265), A2 => n123, B1 => regs(1801), 
                           B2 => n151, C1 => regs(777), C2 => n226, ZN => n2410
                           );
   U3166 : AOI22_X1 port map( A1 => regs(1289), A2 => n12, B1 => regs(2313), B2
                           => n353, ZN => n2409);
   U3167 : NAND2_X1 port map( A1 => n2411, A2 => n2412, ZN => 
                           curr_proc_regs(264));
   U3168 : AOI222_X1 port map( A1 => regs(264), A2 => n123, B1 => regs(1800), 
                           B2 => n151, C1 => regs(776), C2 => n226, ZN => n2412
                           );
   U3169 : AOI22_X1 port map( A1 => regs(1288), A2 => n12, B1 => regs(2312), B2
                           => n353, ZN => n2411);
   U3170 : NAND2_X1 port map( A1 => n2413, A2 => n2414, ZN => 
                           curr_proc_regs(263));
   U3171 : AOI222_X1 port map( A1 => regs(263), A2 => n123, B1 => regs(1799), 
                           B2 => n151, C1 => regs(775), C2 => n226, ZN => n2414
                           );
   U3172 : AOI22_X1 port map( A1 => regs(1287), A2 => n12, B1 => regs(2311), B2
                           => n353, ZN => n2413);
   U3173 : NAND2_X1 port map( A1 => n2415, A2 => n2416, ZN => 
                           curr_proc_regs(262));
   U3174 : AOI222_X1 port map( A1 => regs(262), A2 => n123, B1 => regs(1798), 
                           B2 => n151, C1 => regs(774), C2 => n226, ZN => n2416
                           );
   U3175 : AOI22_X1 port map( A1 => regs(1286), A2 => n12, B1 => regs(2310), B2
                           => n353, ZN => n2415);
   U3176 : NAND2_X1 port map( A1 => n2417, A2 => n2418, ZN => 
                           curr_proc_regs(261));
   U3177 : AOI222_X1 port map( A1 => regs(261), A2 => n123, B1 => regs(1797), 
                           B2 => n151, C1 => regs(773), C2 => n226, ZN => n2418
                           );
   U3178 : AOI22_X1 port map( A1 => regs(1285), A2 => n12, B1 => regs(2309), B2
                           => n353, ZN => n2417);
   U3179 : NAND2_X1 port map( A1 => n2419, A2 => n2420, ZN => 
                           curr_proc_regs(260));
   U3180 : AOI222_X1 port map( A1 => regs(260), A2 => n123, B1 => regs(1796), 
                           B2 => n151, C1 => regs(772), C2 => n226, ZN => n2420
                           );
   U3181 : AOI22_X1 port map( A1 => regs(1284), A2 => n11, B1 => regs(2308), B2
                           => n354, ZN => n2419);
   U3182 : NAND2_X1 port map( A1 => n2421, A2 => n2422, ZN => 
                           curr_proc_regs(259));
   U3183 : AOI222_X1 port map( A1 => regs(259), A2 => n123, B1 => regs(1795), 
                           B2 => n151, C1 => regs(771), C2 => n226, ZN => n2422
                           );
   U3184 : AOI22_X1 port map( A1 => regs(1283), A2 => n11, B1 => regs(2307), B2
                           => n354, ZN => n2421);
   U3185 : NAND2_X1 port map( A1 => n2423, A2 => n2424, ZN => 
                           curr_proc_regs(258));
   U3186 : AOI222_X1 port map( A1 => regs(258), A2 => n123, B1 => regs(1794), 
                           B2 => n151, C1 => regs(770), C2 => n226, ZN => n2424
                           );
   U3187 : AOI22_X1 port map( A1 => regs(1282), A2 => n11, B1 => regs(2306), B2
                           => n354, ZN => n2423);
   U3188 : NAND2_X1 port map( A1 => n2425, A2 => n2426, ZN => 
                           curr_proc_regs(257));
   U3189 : AOI222_X1 port map( A1 => regs(257), A2 => n123, B1 => regs(1793), 
                           B2 => n151, C1 => regs(769), C2 => n226, ZN => n2426
                           );
   U3190 : AOI22_X1 port map( A1 => regs(1281), A2 => n11, B1 => regs(2305), B2
                           => n354, ZN => n2425);
   U3191 : NAND2_X1 port map( A1 => n2427, A2 => n2428, ZN => 
                           curr_proc_regs(256));
   U3192 : AOI222_X1 port map( A1 => regs(256), A2 => n76, B1 => regs(1792), B2
                           => n151, C1 => regs(768), C2 => n226, ZN => n2428);
   U3193 : AND3_X1 port map( A1 => n2429, A2 => n2430, A3 => win(1), ZN => n383
                           );
   U3194 : NOR2_X1 port map( A1 => n2431, A2 => n301, ZN => n382);
   U3195 : INV_X1 port map( A => win(3), ZN => n2431);
   U3196 : AND4_X1 port map( A1 => win(0), A2 => n2429, A3 => n2432, A4 => 
                           n2430, ZN => n381);
   U3197 : INV_X1 port map( A => win(2), ZN => n2430);
   U3198 : INV_X1 port map( A => win(1), ZN => n2432);
   U3199 : AOI22_X1 port map( A1 => regs(1280), A2 => n19, B1 => regs(2304), B2
                           => n354, ZN => n2427);
   U3200 : AND2_X1 port map( A1 => win(2), A2 => n2429, ZN => n378);
   U3201 : NOR2_X1 port map( A1 => win(3), A2 => n301, ZN => n2429);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity reg_generic_N5_RSTVAL1_0 is

   port( D : in std_logic_vector (4 downto 0);  Q : out std_logic_vector (4 
         downto 0);  Clk, Rst, Enable : in std_logic);

end reg_generic_N5_RSTVAL1_0;

architecture SYN_Behavioural of reg_generic_N5_RSTVAL1_0 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n14, n1, n2, n3, n4
      , n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n_1001 : 
      std_logic;

begin
   Q <= ( Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_4_inst : DFF_X1 port map( D => n17, CK => Clk, Q => Q_4_port, QN => 
                           n12);
   Q_reg_3_inst : DFF_X1 port map( D => n16, CK => Clk, Q => Q_3_port, QN => 
                           n11);
   Q_reg_2_inst : DFF_X1 port map( D => n15, CK => Clk, Q => Q_2_port, QN => 
                           n10);
   Q_reg_1_inst : DFF_X1 port map( D => n13, CK => Clk, Q => Q_1_port, QN => n9
                           );
   Q_reg_0_inst : DFF_X1 port map( D => n14, CK => Clk, Q => Q_0_port, QN => 
                           n_1001);
   U3 : OAI22_X1 port map( A1 => n9, A2 => n1, B1 => n2, B2 => n3, ZN => n13);
   U4 : INV_X1 port map( A => D(1), ZN => n3);
   U5 : OAI22_X1 port map( A1 => n10, A2 => n1, B1 => n2, B2 => n4, ZN => n15);
   U6 : INV_X1 port map( A => D(2), ZN => n4);
   U7 : OAI22_X1 port map( A1 => n11, A2 => n1, B1 => n2, B2 => n5, ZN => n16);
   U8 : INV_X1 port map( A => D(3), ZN => n5);
   U9 : OAI22_X1 port map( A1 => n12, A2 => n1, B1 => n2, B2 => n6, ZN => n17);
   U10 : INV_X1 port map( A => D(4), ZN => n6);
   U11 : OR2_X1 port map( A1 => n7, A2 => Rst, ZN => n2);
   U12 : MUX2_X1 port map( A => Q_0_port, B => n8, S => n1, Z => n14);
   U13 : INV_X1 port map( A => n7, ZN => n1);
   U14 : NOR2_X1 port map( A1 => Rst, A2 => Enable, ZN => n7);
   U15 : OR2_X1 port map( A1 => D(0), A2 => Rst, ZN => n8);

end SYN_Behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity nwin_calc_F5_0 is

   port( c_win : in std_logic_vector (4 downto 0);  sel : in std_logic_vector 
         (1 downto 0);  n_win : out std_logic_vector (4 downto 0));

end nwin_calc_F5_0;

architecture SYN_struct of nwin_calc_F5_0 is

   component mux_N5_M2_0
      port( S : in std_logic_vector (1 downto 0);  Q : in std_logic_vector (19 
            downto 0);  Y : out std_logic_vector (4 downto 0));
   end component;

begin
   
   MUX_SEL : mux_N5_M2_0 port map( S(1) => sel(1), S(0) => sel(0), Q(19) => 
                           c_win(4), Q(18) => c_win(3), Q(17) => c_win(2), 
                           Q(16) => c_win(1), Q(15) => c_win(0), Q(14) => 
                           c_win(0), Q(13) => c_win(4), Q(12) => c_win(3), 
                           Q(11) => c_win(2), Q(10) => c_win(1), Q(9) => 
                           c_win(3), Q(8) => c_win(2), Q(7) => c_win(1), Q(6) 
                           => c_win(0), Q(5) => c_win(4), Q(4) => c_win(4), 
                           Q(3) => c_win(3), Q(2) => c_win(2), Q(1) => c_win(1)
                           , Q(0) => c_win(0), Y(4) => n_win(4), Y(3) => 
                           n_win(3), Y(2) => n_win(2), Y(1) => n_win(1), Y(0) 
                           => n_win(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5.all;

entity windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0);  CALL, RET : in std_logic;  FILL, SPILL : out std_logic;  
         BUS_TOMEM : out std_logic_vector (31 downto 0);  BUS_FROMEM : in 
         std_logic_vector (31 downto 0));

end windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5;

architecture SYN_mix of windowing_rf_NBIT_DATA32_NBIT_ADD5_M8_N8_F5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component address_generator_N16_1
      port( clk, rst, enable : in std_logic;  done, working : out std_logic;  
            addr : out std_logic_vector (15 downto 0));
   end component;
   
   component equal_check_N5_1
      port( A, B : in std_logic_vector (4 downto 0);  EQUAL : out std_logic);
   end component;
   
   component mux_N32_M4
      port( S : in std_logic_vector (3 downto 0);  Q : in std_logic_vector (511
            downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component addr_encoder_N4
      port( Q : in std_logic_vector (15 downto 0);  Y : out std_logic_vector (3
            downto 0));
   end component;
   
   component address_generator_N16_0
      port( clk, rst, enable : in std_logic;  done, working : out std_logic;  
            addr : out std_logic_vector (15 downto 0));
   end component;
   
   component in_loc_selblock_NBIT_DATA32_N8_F5
      port( regs : in std_logic_vector (2559 downto 0);  win : in 
            std_logic_vector (4 downto 0);  curr_proc_regs : out 
            std_logic_vector (511 downto 0));
   end component;
   
   component equal_check_N5_0
      port( A, B : in std_logic_vector (4 downto 0);  EQUAL : out std_logic);
   end component;
   
   component reg_generic_N5_RSTVAL1_1
      port( D : in std_logic_vector (4 downto 0);  Q : out std_logic_vector (4 
            downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component nwin_calc_F5_1
      port( c_win : in std_logic_vector (4 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  n_win : out std_logic_vector (4 
            downto 0));
   end component;
   
   component connection_mtx_M8_N8_F5
      port( dec : in std_logic_vector (31 downto 0);  addr_pop : in 
            std_logic_vector (15 downto 0);  win, swp : in std_logic_vector (4 
            downto 0);  sel : out std_logic_vector (87 downto 0));
   end component;
   
   component decoder_N5
      port( Q : in std_logic_vector (4 downto 0);  Y : out std_logic_vector (31
            downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_1
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_2
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_1
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_3
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_4
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_2
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_5
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_6
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_3
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_7
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_8
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_4
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_9
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_10
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_5
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_11
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_12
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_6
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_13
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_14
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_7
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_15
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_16
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_8
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_17
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_18
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_9
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_19
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_20
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_10
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_21
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_22
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_11
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_23
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_24
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_12
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_25
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_26
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_13
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_27
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_28
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_14
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_29
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_30
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_15
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_31
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_32
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_16
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_33
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_34
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_17
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_35
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_36
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_18
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_37
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_38
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_19
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_39
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_40
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_20
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_41
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_42
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_21
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_43
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_44
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_22
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_45
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_46
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_23
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_47
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_48
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_24
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_49
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_50
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_25
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_51
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_52
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_26
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_53
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_54
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_27
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_55
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_56
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_28
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_57
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_58
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_29
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_59
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_60
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_30
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_61
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_62
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_31
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_63
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_64
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_32
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_65
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_66
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_33
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_67
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_68
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_34
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_69
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_70
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_35
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_71
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_72
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_36
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_73
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_74
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_37
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_75
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_76
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_38
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_77
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_78
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_39
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_79
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_80
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M1_0
      port( S : in std_logic;  Q : in std_logic_vector (63 downto 0);  Y : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_81
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_82
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_83
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_84
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_85
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_86
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_87
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_88
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component reg_generic_N32_RSTVAL0_89
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M5_1
      port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector 
            (1023 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component reg_generic_N32_RSTVAL0_0
      port( D : in std_logic_vector (31 downto 0);  Q : out std_logic_vector 
            (31 downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component mux_N32_M5_0
      port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector 
            (1023 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component select_block_NBIT_DATA32_N8_F5
      port( regs : in std_logic_vector (2559 downto 0);  win : in 
            std_logic_vector (4 downto 0);  curr_proc_regs : out 
            std_logic_vector (767 downto 0));
   end component;
   
   component reg_generic_N5_RSTVAL1_0
      port( D : in std_logic_vector (4 downto 0);  Q : out std_logic_vector (4 
            downto 0);  Clk, Rst, Enable : in std_logic);
   end component;
   
   component nwin_calc_F5_0
      port( c_win : in std_logic_vector (4 downto 0);  sel : in 
            std_logic_vector (1 downto 0);  n_win : out std_logic_vector (4 
            downto 0));
   end component;
   
   signal X_Logic1_port, int_RD1, int_RD2, filleq, spilleq, c_win_4_port, 
      c_win_3_port, c_win_2_port, c_win_1_port, c_win_0_port, next_cwp_4_port, 
      next_cwp_3_port, next_cwp_2_port, next_cwp_1_port, next_cwp_0_port, 
      bus_reg_dataout_2559_port, bus_reg_dataout_2558_port, 
      bus_reg_dataout_2557_port, bus_reg_dataout_2556_port, 
      bus_reg_dataout_2555_port, bus_reg_dataout_2554_port, 
      bus_reg_dataout_2553_port, bus_reg_dataout_2552_port, 
      bus_reg_dataout_2551_port, bus_reg_dataout_2550_port, 
      bus_reg_dataout_2549_port, bus_reg_dataout_2548_port, 
      bus_reg_dataout_2547_port, bus_reg_dataout_2546_port, 
      bus_reg_dataout_2545_port, bus_reg_dataout_2544_port, 
      bus_reg_dataout_2543_port, bus_reg_dataout_2542_port, 
      bus_reg_dataout_2541_port, bus_reg_dataout_2540_port, 
      bus_reg_dataout_2539_port, bus_reg_dataout_2538_port, 
      bus_reg_dataout_2537_port, bus_reg_dataout_2536_port, 
      bus_reg_dataout_2535_port, bus_reg_dataout_2534_port, 
      bus_reg_dataout_2533_port, bus_reg_dataout_2532_port, 
      bus_reg_dataout_2531_port, bus_reg_dataout_2530_port, 
      bus_reg_dataout_2529_port, bus_reg_dataout_2528_port, 
      bus_reg_dataout_2527_port, bus_reg_dataout_2526_port, 
      bus_reg_dataout_2525_port, bus_reg_dataout_2524_port, 
      bus_reg_dataout_2523_port, bus_reg_dataout_2522_port, 
      bus_reg_dataout_2521_port, bus_reg_dataout_2520_port, 
      bus_reg_dataout_2519_port, bus_reg_dataout_2518_port, 
      bus_reg_dataout_2517_port, bus_reg_dataout_2516_port, 
      bus_reg_dataout_2515_port, bus_reg_dataout_2514_port, 
      bus_reg_dataout_2513_port, bus_reg_dataout_2512_port, 
      bus_reg_dataout_2511_port, bus_reg_dataout_2510_port, 
      bus_reg_dataout_2509_port, bus_reg_dataout_2508_port, 
      bus_reg_dataout_2507_port, bus_reg_dataout_2506_port, 
      bus_reg_dataout_2505_port, bus_reg_dataout_2504_port, 
      bus_reg_dataout_2503_port, bus_reg_dataout_2502_port, 
      bus_reg_dataout_2501_port, bus_reg_dataout_2500_port, 
      bus_reg_dataout_2499_port, bus_reg_dataout_2498_port, 
      bus_reg_dataout_2497_port, bus_reg_dataout_2496_port, 
      bus_reg_dataout_2495_port, bus_reg_dataout_2494_port, 
      bus_reg_dataout_2493_port, bus_reg_dataout_2492_port, 
      bus_reg_dataout_2491_port, bus_reg_dataout_2490_port, 
      bus_reg_dataout_2489_port, bus_reg_dataout_2488_port, 
      bus_reg_dataout_2487_port, bus_reg_dataout_2486_port, 
      bus_reg_dataout_2485_port, bus_reg_dataout_2484_port, 
      bus_reg_dataout_2483_port, bus_reg_dataout_2482_port, 
      bus_reg_dataout_2481_port, bus_reg_dataout_2480_port, 
      bus_reg_dataout_2479_port, bus_reg_dataout_2478_port, 
      bus_reg_dataout_2477_port, bus_reg_dataout_2476_port, 
      bus_reg_dataout_2475_port, bus_reg_dataout_2474_port, 
      bus_reg_dataout_2473_port, bus_reg_dataout_2472_port, 
      bus_reg_dataout_2471_port, bus_reg_dataout_2470_port, 
      bus_reg_dataout_2469_port, bus_reg_dataout_2468_port, 
      bus_reg_dataout_2467_port, bus_reg_dataout_2466_port, 
      bus_reg_dataout_2465_port, bus_reg_dataout_2464_port, 
      bus_reg_dataout_2463_port, bus_reg_dataout_2462_port, 
      bus_reg_dataout_2461_port, bus_reg_dataout_2460_port, 
      bus_reg_dataout_2459_port, bus_reg_dataout_2458_port, 
      bus_reg_dataout_2457_port, bus_reg_dataout_2456_port, 
      bus_reg_dataout_2455_port, bus_reg_dataout_2454_port, 
      bus_reg_dataout_2453_port, bus_reg_dataout_2452_port, 
      bus_reg_dataout_2451_port, bus_reg_dataout_2450_port, 
      bus_reg_dataout_2449_port, bus_reg_dataout_2448_port, 
      bus_reg_dataout_2447_port, bus_reg_dataout_2446_port, 
      bus_reg_dataout_2445_port, bus_reg_dataout_2444_port, 
      bus_reg_dataout_2443_port, bus_reg_dataout_2442_port, 
      bus_reg_dataout_2441_port, bus_reg_dataout_2440_port, 
      bus_reg_dataout_2439_port, bus_reg_dataout_2438_port, 
      bus_reg_dataout_2437_port, bus_reg_dataout_2436_port, 
      bus_reg_dataout_2435_port, bus_reg_dataout_2434_port, 
      bus_reg_dataout_2433_port, bus_reg_dataout_2432_port, 
      bus_reg_dataout_2431_port, bus_reg_dataout_2430_port, 
      bus_reg_dataout_2429_port, bus_reg_dataout_2428_port, 
      bus_reg_dataout_2427_port, bus_reg_dataout_2426_port, 
      bus_reg_dataout_2425_port, bus_reg_dataout_2424_port, 
      bus_reg_dataout_2423_port, bus_reg_dataout_2422_port, 
      bus_reg_dataout_2421_port, bus_reg_dataout_2420_port, 
      bus_reg_dataout_2419_port, bus_reg_dataout_2418_port, 
      bus_reg_dataout_2417_port, bus_reg_dataout_2416_port, 
      bus_reg_dataout_2415_port, bus_reg_dataout_2414_port, 
      bus_reg_dataout_2413_port, bus_reg_dataout_2412_port, 
      bus_reg_dataout_2411_port, bus_reg_dataout_2410_port, 
      bus_reg_dataout_2409_port, bus_reg_dataout_2408_port, 
      bus_reg_dataout_2407_port, bus_reg_dataout_2406_port, 
      bus_reg_dataout_2405_port, bus_reg_dataout_2404_port, 
      bus_reg_dataout_2403_port, bus_reg_dataout_2402_port, 
      bus_reg_dataout_2401_port, bus_reg_dataout_2400_port, 
      bus_reg_dataout_2399_port, bus_reg_dataout_2398_port, 
      bus_reg_dataout_2397_port, bus_reg_dataout_2396_port, 
      bus_reg_dataout_2395_port, bus_reg_dataout_2394_port, 
      bus_reg_dataout_2393_port, bus_reg_dataout_2392_port, 
      bus_reg_dataout_2391_port, bus_reg_dataout_2390_port, 
      bus_reg_dataout_2389_port, bus_reg_dataout_2388_port, 
      bus_reg_dataout_2387_port, bus_reg_dataout_2386_port, 
      bus_reg_dataout_2385_port, bus_reg_dataout_2384_port, 
      bus_reg_dataout_2383_port, bus_reg_dataout_2382_port, 
      bus_reg_dataout_2381_port, bus_reg_dataout_2380_port, 
      bus_reg_dataout_2379_port, bus_reg_dataout_2378_port, 
      bus_reg_dataout_2377_port, bus_reg_dataout_2376_port, 
      bus_reg_dataout_2375_port, bus_reg_dataout_2374_port, 
      bus_reg_dataout_2373_port, bus_reg_dataout_2372_port, 
      bus_reg_dataout_2371_port, bus_reg_dataout_2370_port, 
      bus_reg_dataout_2369_port, bus_reg_dataout_2368_port, 
      bus_reg_dataout_2367_port, bus_reg_dataout_2366_port, 
      bus_reg_dataout_2365_port, bus_reg_dataout_2364_port, 
      bus_reg_dataout_2363_port, bus_reg_dataout_2362_port, 
      bus_reg_dataout_2361_port, bus_reg_dataout_2360_port, 
      bus_reg_dataout_2359_port, bus_reg_dataout_2358_port, 
      bus_reg_dataout_2357_port, bus_reg_dataout_2356_port, 
      bus_reg_dataout_2355_port, bus_reg_dataout_2354_port, 
      bus_reg_dataout_2353_port, bus_reg_dataout_2352_port, 
      bus_reg_dataout_2351_port, bus_reg_dataout_2350_port, 
      bus_reg_dataout_2349_port, bus_reg_dataout_2348_port, 
      bus_reg_dataout_2347_port, bus_reg_dataout_2346_port, 
      bus_reg_dataout_2345_port, bus_reg_dataout_2344_port, 
      bus_reg_dataout_2343_port, bus_reg_dataout_2342_port, 
      bus_reg_dataout_2341_port, bus_reg_dataout_2340_port, 
      bus_reg_dataout_2339_port, bus_reg_dataout_2338_port, 
      bus_reg_dataout_2337_port, bus_reg_dataout_2336_port, 
      bus_reg_dataout_2335_port, bus_reg_dataout_2334_port, 
      bus_reg_dataout_2333_port, bus_reg_dataout_2332_port, 
      bus_reg_dataout_2331_port, bus_reg_dataout_2330_port, 
      bus_reg_dataout_2329_port, bus_reg_dataout_2328_port, 
      bus_reg_dataout_2327_port, bus_reg_dataout_2326_port, 
      bus_reg_dataout_2325_port, bus_reg_dataout_2324_port, 
      bus_reg_dataout_2323_port, bus_reg_dataout_2322_port, 
      bus_reg_dataout_2321_port, bus_reg_dataout_2320_port, 
      bus_reg_dataout_2319_port, bus_reg_dataout_2318_port, 
      bus_reg_dataout_2317_port, bus_reg_dataout_2316_port, 
      bus_reg_dataout_2315_port, bus_reg_dataout_2314_port, 
      bus_reg_dataout_2313_port, bus_reg_dataout_2312_port, 
      bus_reg_dataout_2311_port, bus_reg_dataout_2310_port, 
      bus_reg_dataout_2309_port, bus_reg_dataout_2308_port, 
      bus_reg_dataout_2307_port, bus_reg_dataout_2306_port, 
      bus_reg_dataout_2305_port, bus_reg_dataout_2304_port, 
      bus_reg_dataout_2303_port, bus_reg_dataout_2302_port, 
      bus_reg_dataout_2301_port, bus_reg_dataout_2300_port, 
      bus_reg_dataout_2299_port, bus_reg_dataout_2298_port, 
      bus_reg_dataout_2297_port, bus_reg_dataout_2296_port, 
      bus_reg_dataout_2295_port, bus_reg_dataout_2294_port, 
      bus_reg_dataout_2293_port, bus_reg_dataout_2292_port, 
      bus_reg_dataout_2291_port, bus_reg_dataout_2290_port, 
      bus_reg_dataout_2289_port, bus_reg_dataout_2288_port, 
      bus_reg_dataout_2287_port, bus_reg_dataout_2286_port, 
      bus_reg_dataout_2285_port, bus_reg_dataout_2284_port, 
      bus_reg_dataout_2283_port, bus_reg_dataout_2282_port, 
      bus_reg_dataout_2281_port, bus_reg_dataout_2280_port, 
      bus_reg_dataout_2279_port, bus_reg_dataout_2278_port, 
      bus_reg_dataout_2277_port, bus_reg_dataout_2276_port, 
      bus_reg_dataout_2275_port, bus_reg_dataout_2274_port, 
      bus_reg_dataout_2273_port, bus_reg_dataout_2272_port, 
      bus_reg_dataout_2271_port, bus_reg_dataout_2270_port, 
      bus_reg_dataout_2269_port, bus_reg_dataout_2268_port, 
      bus_reg_dataout_2267_port, bus_reg_dataout_2266_port, 
      bus_reg_dataout_2265_port, bus_reg_dataout_2264_port, 
      bus_reg_dataout_2263_port, bus_reg_dataout_2262_port, 
      bus_reg_dataout_2261_port, bus_reg_dataout_2260_port, 
      bus_reg_dataout_2259_port, bus_reg_dataout_2258_port, 
      bus_reg_dataout_2257_port, bus_reg_dataout_2256_port, 
      bus_reg_dataout_2255_port, bus_reg_dataout_2254_port, 
      bus_reg_dataout_2253_port, bus_reg_dataout_2252_port, 
      bus_reg_dataout_2251_port, bus_reg_dataout_2250_port, 
      bus_reg_dataout_2249_port, bus_reg_dataout_2248_port, 
      bus_reg_dataout_2247_port, bus_reg_dataout_2246_port, 
      bus_reg_dataout_2245_port, bus_reg_dataout_2244_port, 
      bus_reg_dataout_2243_port, bus_reg_dataout_2242_port, 
      bus_reg_dataout_2241_port, bus_reg_dataout_2240_port, 
      bus_reg_dataout_2239_port, bus_reg_dataout_2238_port, 
      bus_reg_dataout_2237_port, bus_reg_dataout_2236_port, 
      bus_reg_dataout_2235_port, bus_reg_dataout_2234_port, 
      bus_reg_dataout_2233_port, bus_reg_dataout_2232_port, 
      bus_reg_dataout_2231_port, bus_reg_dataout_2230_port, 
      bus_reg_dataout_2229_port, bus_reg_dataout_2228_port, 
      bus_reg_dataout_2227_port, bus_reg_dataout_2226_port, 
      bus_reg_dataout_2225_port, bus_reg_dataout_2224_port, 
      bus_reg_dataout_2223_port, bus_reg_dataout_2222_port, 
      bus_reg_dataout_2221_port, bus_reg_dataout_2220_port, 
      bus_reg_dataout_2219_port, bus_reg_dataout_2218_port, 
      bus_reg_dataout_2217_port, bus_reg_dataout_2216_port, 
      bus_reg_dataout_2215_port, bus_reg_dataout_2214_port, 
      bus_reg_dataout_2213_port, bus_reg_dataout_2212_port, 
      bus_reg_dataout_2211_port, bus_reg_dataout_2210_port, 
      bus_reg_dataout_2209_port, bus_reg_dataout_2208_port, 
      bus_reg_dataout_2207_port, bus_reg_dataout_2206_port, 
      bus_reg_dataout_2205_port, bus_reg_dataout_2204_port, 
      bus_reg_dataout_2203_port, bus_reg_dataout_2202_port, 
      bus_reg_dataout_2201_port, bus_reg_dataout_2200_port, 
      bus_reg_dataout_2199_port, bus_reg_dataout_2198_port, 
      bus_reg_dataout_2197_port, bus_reg_dataout_2196_port, 
      bus_reg_dataout_2195_port, bus_reg_dataout_2194_port, 
      bus_reg_dataout_2193_port, bus_reg_dataout_2192_port, 
      bus_reg_dataout_2191_port, bus_reg_dataout_2190_port, 
      bus_reg_dataout_2189_port, bus_reg_dataout_2188_port, 
      bus_reg_dataout_2187_port, bus_reg_dataout_2186_port, 
      bus_reg_dataout_2185_port, bus_reg_dataout_2184_port, 
      bus_reg_dataout_2183_port, bus_reg_dataout_2182_port, 
      bus_reg_dataout_2181_port, bus_reg_dataout_2180_port, 
      bus_reg_dataout_2179_port, bus_reg_dataout_2178_port, 
      bus_reg_dataout_2177_port, bus_reg_dataout_2176_port, 
      bus_reg_dataout_2175_port, bus_reg_dataout_2174_port, 
      bus_reg_dataout_2173_port, bus_reg_dataout_2172_port, 
      bus_reg_dataout_2171_port, bus_reg_dataout_2170_port, 
      bus_reg_dataout_2169_port, bus_reg_dataout_2168_port, 
      bus_reg_dataout_2167_port, bus_reg_dataout_2166_port, 
      bus_reg_dataout_2165_port, bus_reg_dataout_2164_port, 
      bus_reg_dataout_2163_port, bus_reg_dataout_2162_port, 
      bus_reg_dataout_2161_port, bus_reg_dataout_2160_port, 
      bus_reg_dataout_2159_port, bus_reg_dataout_2158_port, 
      bus_reg_dataout_2157_port, bus_reg_dataout_2156_port, 
      bus_reg_dataout_2155_port, bus_reg_dataout_2154_port, 
      bus_reg_dataout_2153_port, bus_reg_dataout_2152_port, 
      bus_reg_dataout_2151_port, bus_reg_dataout_2150_port, 
      bus_reg_dataout_2149_port, bus_reg_dataout_2148_port, 
      bus_reg_dataout_2147_port, bus_reg_dataout_2146_port, 
      bus_reg_dataout_2145_port, bus_reg_dataout_2144_port, 
      bus_reg_dataout_2143_port, bus_reg_dataout_2142_port, 
      bus_reg_dataout_2141_port, bus_reg_dataout_2140_port, 
      bus_reg_dataout_2139_port, bus_reg_dataout_2138_port, 
      bus_reg_dataout_2137_port, bus_reg_dataout_2136_port, 
      bus_reg_dataout_2135_port, bus_reg_dataout_2134_port, 
      bus_reg_dataout_2133_port, bus_reg_dataout_2132_port, 
      bus_reg_dataout_2131_port, bus_reg_dataout_2130_port, 
      bus_reg_dataout_2129_port, bus_reg_dataout_2128_port, 
      bus_reg_dataout_2127_port, bus_reg_dataout_2126_port, 
      bus_reg_dataout_2125_port, bus_reg_dataout_2124_port, 
      bus_reg_dataout_2123_port, bus_reg_dataout_2122_port, 
      bus_reg_dataout_2121_port, bus_reg_dataout_2120_port, 
      bus_reg_dataout_2119_port, bus_reg_dataout_2118_port, 
      bus_reg_dataout_2117_port, bus_reg_dataout_2116_port, 
      bus_reg_dataout_2115_port, bus_reg_dataout_2114_port, 
      bus_reg_dataout_2113_port, bus_reg_dataout_2112_port, 
      bus_reg_dataout_2111_port, bus_reg_dataout_2110_port, 
      bus_reg_dataout_2109_port, bus_reg_dataout_2108_port, 
      bus_reg_dataout_2107_port, bus_reg_dataout_2106_port, 
      bus_reg_dataout_2105_port, bus_reg_dataout_2104_port, 
      bus_reg_dataout_2103_port, bus_reg_dataout_2102_port, 
      bus_reg_dataout_2101_port, bus_reg_dataout_2100_port, 
      bus_reg_dataout_2099_port, bus_reg_dataout_2098_port, 
      bus_reg_dataout_2097_port, bus_reg_dataout_2096_port, 
      bus_reg_dataout_2095_port, bus_reg_dataout_2094_port, 
      bus_reg_dataout_2093_port, bus_reg_dataout_2092_port, 
      bus_reg_dataout_2091_port, bus_reg_dataout_2090_port, 
      bus_reg_dataout_2089_port, bus_reg_dataout_2088_port, 
      bus_reg_dataout_2087_port, bus_reg_dataout_2086_port, 
      bus_reg_dataout_2085_port, bus_reg_dataout_2084_port, 
      bus_reg_dataout_2083_port, bus_reg_dataout_2082_port, 
      bus_reg_dataout_2081_port, bus_reg_dataout_2080_port, 
      bus_reg_dataout_2079_port, bus_reg_dataout_2078_port, 
      bus_reg_dataout_2077_port, bus_reg_dataout_2076_port, 
      bus_reg_dataout_2075_port, bus_reg_dataout_2074_port, 
      bus_reg_dataout_2073_port, bus_reg_dataout_2072_port, 
      bus_reg_dataout_2071_port, bus_reg_dataout_2070_port, 
      bus_reg_dataout_2069_port, bus_reg_dataout_2068_port, 
      bus_reg_dataout_2067_port, bus_reg_dataout_2066_port, 
      bus_reg_dataout_2065_port, bus_reg_dataout_2064_port, 
      bus_reg_dataout_2063_port, bus_reg_dataout_2062_port, 
      bus_reg_dataout_2061_port, bus_reg_dataout_2060_port, 
      bus_reg_dataout_2059_port, bus_reg_dataout_2058_port, 
      bus_reg_dataout_2057_port, bus_reg_dataout_2056_port, 
      bus_reg_dataout_2055_port, bus_reg_dataout_2054_port, 
      bus_reg_dataout_2053_port, bus_reg_dataout_2052_port, 
      bus_reg_dataout_2051_port, bus_reg_dataout_2050_port, 
      bus_reg_dataout_2049_port, bus_reg_dataout_2048_port, 
      bus_reg_dataout_2047_port, bus_reg_dataout_2046_port, 
      bus_reg_dataout_2045_port, bus_reg_dataout_2044_port, 
      bus_reg_dataout_2043_port, bus_reg_dataout_2042_port, 
      bus_reg_dataout_2041_port, bus_reg_dataout_2040_port, 
      bus_reg_dataout_2039_port, bus_reg_dataout_2038_port, 
      bus_reg_dataout_2037_port, bus_reg_dataout_2036_port, 
      bus_reg_dataout_2035_port, bus_reg_dataout_2034_port, 
      bus_reg_dataout_2033_port, bus_reg_dataout_2032_port, 
      bus_reg_dataout_2031_port, bus_reg_dataout_2030_port, 
      bus_reg_dataout_2029_port, bus_reg_dataout_2028_port, 
      bus_reg_dataout_2027_port, bus_reg_dataout_2026_port, 
      bus_reg_dataout_2025_port, bus_reg_dataout_2024_port, 
      bus_reg_dataout_2023_port, bus_reg_dataout_2022_port, 
      bus_reg_dataout_2021_port, bus_reg_dataout_2020_port, 
      bus_reg_dataout_2019_port, bus_reg_dataout_2018_port, 
      bus_reg_dataout_2017_port, bus_reg_dataout_2016_port, 
      bus_reg_dataout_2015_port, bus_reg_dataout_2014_port, 
      bus_reg_dataout_2013_port, bus_reg_dataout_2012_port, 
      bus_reg_dataout_2011_port, bus_reg_dataout_2010_port, 
      bus_reg_dataout_2009_port, bus_reg_dataout_2008_port, 
      bus_reg_dataout_2007_port, bus_reg_dataout_2006_port, 
      bus_reg_dataout_2005_port, bus_reg_dataout_2004_port, 
      bus_reg_dataout_2003_port, bus_reg_dataout_2002_port, 
      bus_reg_dataout_2001_port, bus_reg_dataout_2000_port, 
      bus_reg_dataout_1999_port, bus_reg_dataout_1998_port, 
      bus_reg_dataout_1997_port, bus_reg_dataout_1996_port, 
      bus_reg_dataout_1995_port, bus_reg_dataout_1994_port, 
      bus_reg_dataout_1993_port, bus_reg_dataout_1992_port, 
      bus_reg_dataout_1991_port, bus_reg_dataout_1990_port, 
      bus_reg_dataout_1989_port, bus_reg_dataout_1988_port, 
      bus_reg_dataout_1987_port, bus_reg_dataout_1986_port, 
      bus_reg_dataout_1985_port, bus_reg_dataout_1984_port, 
      bus_reg_dataout_1983_port, bus_reg_dataout_1982_port, 
      bus_reg_dataout_1981_port, bus_reg_dataout_1980_port, 
      bus_reg_dataout_1979_port, bus_reg_dataout_1978_port, 
      bus_reg_dataout_1977_port, bus_reg_dataout_1976_port, 
      bus_reg_dataout_1975_port, bus_reg_dataout_1974_port, 
      bus_reg_dataout_1973_port, bus_reg_dataout_1972_port, 
      bus_reg_dataout_1971_port, bus_reg_dataout_1970_port, 
      bus_reg_dataout_1969_port, bus_reg_dataout_1968_port, 
      bus_reg_dataout_1967_port, bus_reg_dataout_1966_port, 
      bus_reg_dataout_1965_port, bus_reg_dataout_1964_port, 
      bus_reg_dataout_1963_port, bus_reg_dataout_1962_port, 
      bus_reg_dataout_1961_port, bus_reg_dataout_1960_port, 
      bus_reg_dataout_1959_port, bus_reg_dataout_1958_port, 
      bus_reg_dataout_1957_port, bus_reg_dataout_1956_port, 
      bus_reg_dataout_1955_port, bus_reg_dataout_1954_port, 
      bus_reg_dataout_1953_port, bus_reg_dataout_1952_port, 
      bus_reg_dataout_1951_port, bus_reg_dataout_1950_port, 
      bus_reg_dataout_1949_port, bus_reg_dataout_1948_port, 
      bus_reg_dataout_1947_port, bus_reg_dataout_1946_port, 
      bus_reg_dataout_1945_port, bus_reg_dataout_1944_port, 
      bus_reg_dataout_1943_port, bus_reg_dataout_1942_port, 
      bus_reg_dataout_1941_port, bus_reg_dataout_1940_port, 
      bus_reg_dataout_1939_port, bus_reg_dataout_1938_port, 
      bus_reg_dataout_1937_port, bus_reg_dataout_1936_port, 
      bus_reg_dataout_1935_port, bus_reg_dataout_1934_port, 
      bus_reg_dataout_1933_port, bus_reg_dataout_1932_port, 
      bus_reg_dataout_1931_port, bus_reg_dataout_1930_port, 
      bus_reg_dataout_1929_port, bus_reg_dataout_1928_port, 
      bus_reg_dataout_1927_port, bus_reg_dataout_1926_port, 
      bus_reg_dataout_1925_port, bus_reg_dataout_1924_port, 
      bus_reg_dataout_1923_port, bus_reg_dataout_1922_port, 
      bus_reg_dataout_1921_port, bus_reg_dataout_1920_port, 
      bus_reg_dataout_1919_port, bus_reg_dataout_1918_port, 
      bus_reg_dataout_1917_port, bus_reg_dataout_1916_port, 
      bus_reg_dataout_1915_port, bus_reg_dataout_1914_port, 
      bus_reg_dataout_1913_port, bus_reg_dataout_1912_port, 
      bus_reg_dataout_1911_port, bus_reg_dataout_1910_port, 
      bus_reg_dataout_1909_port, bus_reg_dataout_1908_port, 
      bus_reg_dataout_1907_port, bus_reg_dataout_1906_port, 
      bus_reg_dataout_1905_port, bus_reg_dataout_1904_port, 
      bus_reg_dataout_1903_port, bus_reg_dataout_1902_port, 
      bus_reg_dataout_1901_port, bus_reg_dataout_1900_port, 
      bus_reg_dataout_1899_port, bus_reg_dataout_1898_port, 
      bus_reg_dataout_1897_port, bus_reg_dataout_1896_port, 
      bus_reg_dataout_1895_port, bus_reg_dataout_1894_port, 
      bus_reg_dataout_1893_port, bus_reg_dataout_1892_port, 
      bus_reg_dataout_1891_port, bus_reg_dataout_1890_port, 
      bus_reg_dataout_1889_port, bus_reg_dataout_1888_port, 
      bus_reg_dataout_1887_port, bus_reg_dataout_1886_port, 
      bus_reg_dataout_1885_port, bus_reg_dataout_1884_port, 
      bus_reg_dataout_1883_port, bus_reg_dataout_1882_port, 
      bus_reg_dataout_1881_port, bus_reg_dataout_1880_port, 
      bus_reg_dataout_1879_port, bus_reg_dataout_1878_port, 
      bus_reg_dataout_1877_port, bus_reg_dataout_1876_port, 
      bus_reg_dataout_1875_port, bus_reg_dataout_1874_port, 
      bus_reg_dataout_1873_port, bus_reg_dataout_1872_port, 
      bus_reg_dataout_1871_port, bus_reg_dataout_1870_port, 
      bus_reg_dataout_1869_port, bus_reg_dataout_1868_port, 
      bus_reg_dataout_1867_port, bus_reg_dataout_1866_port, 
      bus_reg_dataout_1865_port, bus_reg_dataout_1864_port, 
      bus_reg_dataout_1863_port, bus_reg_dataout_1862_port, 
      bus_reg_dataout_1861_port, bus_reg_dataout_1860_port, 
      bus_reg_dataout_1859_port, bus_reg_dataout_1858_port, 
      bus_reg_dataout_1857_port, bus_reg_dataout_1856_port, 
      bus_reg_dataout_1855_port, bus_reg_dataout_1854_port, 
      bus_reg_dataout_1853_port, bus_reg_dataout_1852_port, 
      bus_reg_dataout_1851_port, bus_reg_dataout_1850_port, 
      bus_reg_dataout_1849_port, bus_reg_dataout_1848_port, 
      bus_reg_dataout_1847_port, bus_reg_dataout_1846_port, 
      bus_reg_dataout_1845_port, bus_reg_dataout_1844_port, 
      bus_reg_dataout_1843_port, bus_reg_dataout_1842_port, 
      bus_reg_dataout_1841_port, bus_reg_dataout_1840_port, 
      bus_reg_dataout_1839_port, bus_reg_dataout_1838_port, 
      bus_reg_dataout_1837_port, bus_reg_dataout_1836_port, 
      bus_reg_dataout_1835_port, bus_reg_dataout_1834_port, 
      bus_reg_dataout_1833_port, bus_reg_dataout_1832_port, 
      bus_reg_dataout_1831_port, bus_reg_dataout_1830_port, 
      bus_reg_dataout_1829_port, bus_reg_dataout_1828_port, 
      bus_reg_dataout_1827_port, bus_reg_dataout_1826_port, 
      bus_reg_dataout_1825_port, bus_reg_dataout_1824_port, 
      bus_reg_dataout_1823_port, bus_reg_dataout_1822_port, 
      bus_reg_dataout_1821_port, bus_reg_dataout_1820_port, 
      bus_reg_dataout_1819_port, bus_reg_dataout_1818_port, 
      bus_reg_dataout_1817_port, bus_reg_dataout_1816_port, 
      bus_reg_dataout_1815_port, bus_reg_dataout_1814_port, 
      bus_reg_dataout_1813_port, bus_reg_dataout_1812_port, 
      bus_reg_dataout_1811_port, bus_reg_dataout_1810_port, 
      bus_reg_dataout_1809_port, bus_reg_dataout_1808_port, 
      bus_reg_dataout_1807_port, bus_reg_dataout_1806_port, 
      bus_reg_dataout_1805_port, bus_reg_dataout_1804_port, 
      bus_reg_dataout_1803_port, bus_reg_dataout_1802_port, 
      bus_reg_dataout_1801_port, bus_reg_dataout_1800_port, 
      bus_reg_dataout_1799_port, bus_reg_dataout_1798_port, 
      bus_reg_dataout_1797_port, bus_reg_dataout_1796_port, 
      bus_reg_dataout_1795_port, bus_reg_dataout_1794_port, 
      bus_reg_dataout_1793_port, bus_reg_dataout_1792_port, 
      bus_reg_dataout_1791_port, bus_reg_dataout_1790_port, 
      bus_reg_dataout_1789_port, bus_reg_dataout_1788_port, 
      bus_reg_dataout_1787_port, bus_reg_dataout_1786_port, 
      bus_reg_dataout_1785_port, bus_reg_dataout_1784_port, 
      bus_reg_dataout_1783_port, bus_reg_dataout_1782_port, 
      bus_reg_dataout_1781_port, bus_reg_dataout_1780_port, 
      bus_reg_dataout_1779_port, bus_reg_dataout_1778_port, 
      bus_reg_dataout_1777_port, bus_reg_dataout_1776_port, 
      bus_reg_dataout_1775_port, bus_reg_dataout_1774_port, 
      bus_reg_dataout_1773_port, bus_reg_dataout_1772_port, 
      bus_reg_dataout_1771_port, bus_reg_dataout_1770_port, 
      bus_reg_dataout_1769_port, bus_reg_dataout_1768_port, 
      bus_reg_dataout_1767_port, bus_reg_dataout_1766_port, 
      bus_reg_dataout_1765_port, bus_reg_dataout_1764_port, 
      bus_reg_dataout_1763_port, bus_reg_dataout_1762_port, 
      bus_reg_dataout_1761_port, bus_reg_dataout_1760_port, 
      bus_reg_dataout_1759_port, bus_reg_dataout_1758_port, 
      bus_reg_dataout_1757_port, bus_reg_dataout_1756_port, 
      bus_reg_dataout_1755_port, bus_reg_dataout_1754_port, 
      bus_reg_dataout_1753_port, bus_reg_dataout_1752_port, 
      bus_reg_dataout_1751_port, bus_reg_dataout_1750_port, 
      bus_reg_dataout_1749_port, bus_reg_dataout_1748_port, 
      bus_reg_dataout_1747_port, bus_reg_dataout_1746_port, 
      bus_reg_dataout_1745_port, bus_reg_dataout_1744_port, 
      bus_reg_dataout_1743_port, bus_reg_dataout_1742_port, 
      bus_reg_dataout_1741_port, bus_reg_dataout_1740_port, 
      bus_reg_dataout_1739_port, bus_reg_dataout_1738_port, 
      bus_reg_dataout_1737_port, bus_reg_dataout_1736_port, 
      bus_reg_dataout_1735_port, bus_reg_dataout_1734_port, 
      bus_reg_dataout_1733_port, bus_reg_dataout_1732_port, 
      bus_reg_dataout_1731_port, bus_reg_dataout_1730_port, 
      bus_reg_dataout_1729_port, bus_reg_dataout_1728_port, 
      bus_reg_dataout_1727_port, bus_reg_dataout_1726_port, 
      bus_reg_dataout_1725_port, bus_reg_dataout_1724_port, 
      bus_reg_dataout_1723_port, bus_reg_dataout_1722_port, 
      bus_reg_dataout_1721_port, bus_reg_dataout_1720_port, 
      bus_reg_dataout_1719_port, bus_reg_dataout_1718_port, 
      bus_reg_dataout_1717_port, bus_reg_dataout_1716_port, 
      bus_reg_dataout_1715_port, bus_reg_dataout_1714_port, 
      bus_reg_dataout_1713_port, bus_reg_dataout_1712_port, 
      bus_reg_dataout_1711_port, bus_reg_dataout_1710_port, 
      bus_reg_dataout_1709_port, bus_reg_dataout_1708_port, 
      bus_reg_dataout_1707_port, bus_reg_dataout_1706_port, 
      bus_reg_dataout_1705_port, bus_reg_dataout_1704_port, 
      bus_reg_dataout_1703_port, bus_reg_dataout_1702_port, 
      bus_reg_dataout_1701_port, bus_reg_dataout_1700_port, 
      bus_reg_dataout_1699_port, bus_reg_dataout_1698_port, 
      bus_reg_dataout_1697_port, bus_reg_dataout_1696_port, 
      bus_reg_dataout_1695_port, bus_reg_dataout_1694_port, 
      bus_reg_dataout_1693_port, bus_reg_dataout_1692_port, 
      bus_reg_dataout_1691_port, bus_reg_dataout_1690_port, 
      bus_reg_dataout_1689_port, bus_reg_dataout_1688_port, 
      bus_reg_dataout_1687_port, bus_reg_dataout_1686_port, 
      bus_reg_dataout_1685_port, bus_reg_dataout_1684_port, 
      bus_reg_dataout_1683_port, bus_reg_dataout_1682_port, 
      bus_reg_dataout_1681_port, bus_reg_dataout_1680_port, 
      bus_reg_dataout_1679_port, bus_reg_dataout_1678_port, 
      bus_reg_dataout_1677_port, bus_reg_dataout_1676_port, 
      bus_reg_dataout_1675_port, bus_reg_dataout_1674_port, 
      bus_reg_dataout_1673_port, bus_reg_dataout_1672_port, 
      bus_reg_dataout_1671_port, bus_reg_dataout_1670_port, 
      bus_reg_dataout_1669_port, bus_reg_dataout_1668_port, 
      bus_reg_dataout_1667_port, bus_reg_dataout_1666_port, 
      bus_reg_dataout_1665_port, bus_reg_dataout_1664_port, 
      bus_reg_dataout_1663_port, bus_reg_dataout_1662_port, 
      bus_reg_dataout_1661_port, bus_reg_dataout_1660_port, 
      bus_reg_dataout_1659_port, bus_reg_dataout_1658_port, 
      bus_reg_dataout_1657_port, bus_reg_dataout_1656_port, 
      bus_reg_dataout_1655_port, bus_reg_dataout_1654_port, 
      bus_reg_dataout_1653_port, bus_reg_dataout_1652_port, 
      bus_reg_dataout_1651_port, bus_reg_dataout_1650_port, 
      bus_reg_dataout_1649_port, bus_reg_dataout_1648_port, 
      bus_reg_dataout_1647_port, bus_reg_dataout_1646_port, 
      bus_reg_dataout_1645_port, bus_reg_dataout_1644_port, 
      bus_reg_dataout_1643_port, bus_reg_dataout_1642_port, 
      bus_reg_dataout_1641_port, bus_reg_dataout_1640_port, 
      bus_reg_dataout_1639_port, bus_reg_dataout_1638_port, 
      bus_reg_dataout_1637_port, bus_reg_dataout_1636_port, 
      bus_reg_dataout_1635_port, bus_reg_dataout_1634_port, 
      bus_reg_dataout_1633_port, bus_reg_dataout_1632_port, 
      bus_reg_dataout_1631_port, bus_reg_dataout_1630_port, 
      bus_reg_dataout_1629_port, bus_reg_dataout_1628_port, 
      bus_reg_dataout_1627_port, bus_reg_dataout_1626_port, 
      bus_reg_dataout_1625_port, bus_reg_dataout_1624_port, 
      bus_reg_dataout_1623_port, bus_reg_dataout_1622_port, 
      bus_reg_dataout_1621_port, bus_reg_dataout_1620_port, 
      bus_reg_dataout_1619_port, bus_reg_dataout_1618_port, 
      bus_reg_dataout_1617_port, bus_reg_dataout_1616_port, 
      bus_reg_dataout_1615_port, bus_reg_dataout_1614_port, 
      bus_reg_dataout_1613_port, bus_reg_dataout_1612_port, 
      bus_reg_dataout_1611_port, bus_reg_dataout_1610_port, 
      bus_reg_dataout_1609_port, bus_reg_dataout_1608_port, 
      bus_reg_dataout_1607_port, bus_reg_dataout_1606_port, 
      bus_reg_dataout_1605_port, bus_reg_dataout_1604_port, 
      bus_reg_dataout_1603_port, bus_reg_dataout_1602_port, 
      bus_reg_dataout_1601_port, bus_reg_dataout_1600_port, 
      bus_reg_dataout_1599_port, bus_reg_dataout_1598_port, 
      bus_reg_dataout_1597_port, bus_reg_dataout_1596_port, 
      bus_reg_dataout_1595_port, bus_reg_dataout_1594_port, 
      bus_reg_dataout_1593_port, bus_reg_dataout_1592_port, 
      bus_reg_dataout_1591_port, bus_reg_dataout_1590_port, 
      bus_reg_dataout_1589_port, bus_reg_dataout_1588_port, 
      bus_reg_dataout_1587_port, bus_reg_dataout_1586_port, 
      bus_reg_dataout_1585_port, bus_reg_dataout_1584_port, 
      bus_reg_dataout_1583_port, bus_reg_dataout_1582_port, 
      bus_reg_dataout_1581_port, bus_reg_dataout_1580_port, 
      bus_reg_dataout_1579_port, bus_reg_dataout_1578_port, 
      bus_reg_dataout_1577_port, bus_reg_dataout_1576_port, 
      bus_reg_dataout_1575_port, bus_reg_dataout_1574_port, 
      bus_reg_dataout_1573_port, bus_reg_dataout_1572_port, 
      bus_reg_dataout_1571_port, bus_reg_dataout_1570_port, 
      bus_reg_dataout_1569_port, bus_reg_dataout_1568_port, 
      bus_reg_dataout_1567_port, bus_reg_dataout_1566_port, 
      bus_reg_dataout_1565_port, bus_reg_dataout_1564_port, 
      bus_reg_dataout_1563_port, bus_reg_dataout_1562_port, 
      bus_reg_dataout_1561_port, bus_reg_dataout_1560_port, 
      bus_reg_dataout_1559_port, bus_reg_dataout_1558_port, 
      bus_reg_dataout_1557_port, bus_reg_dataout_1556_port, 
      bus_reg_dataout_1555_port, bus_reg_dataout_1554_port, 
      bus_reg_dataout_1553_port, bus_reg_dataout_1552_port, 
      bus_reg_dataout_1551_port, bus_reg_dataout_1550_port, 
      bus_reg_dataout_1549_port, bus_reg_dataout_1548_port, 
      bus_reg_dataout_1547_port, bus_reg_dataout_1546_port, 
      bus_reg_dataout_1545_port, bus_reg_dataout_1544_port, 
      bus_reg_dataout_1543_port, bus_reg_dataout_1542_port, 
      bus_reg_dataout_1541_port, bus_reg_dataout_1540_port, 
      bus_reg_dataout_1539_port, bus_reg_dataout_1538_port, 
      bus_reg_dataout_1537_port, bus_reg_dataout_1536_port, 
      bus_reg_dataout_1535_port, bus_reg_dataout_1534_port, 
      bus_reg_dataout_1533_port, bus_reg_dataout_1532_port, 
      bus_reg_dataout_1531_port, bus_reg_dataout_1530_port, 
      bus_reg_dataout_1529_port, bus_reg_dataout_1528_port, 
      bus_reg_dataout_1527_port, bus_reg_dataout_1526_port, 
      bus_reg_dataout_1525_port, bus_reg_dataout_1524_port, 
      bus_reg_dataout_1523_port, bus_reg_dataout_1522_port, 
      bus_reg_dataout_1521_port, bus_reg_dataout_1520_port, 
      bus_reg_dataout_1519_port, bus_reg_dataout_1518_port, 
      bus_reg_dataout_1517_port, bus_reg_dataout_1516_port, 
      bus_reg_dataout_1515_port, bus_reg_dataout_1514_port, 
      bus_reg_dataout_1513_port, bus_reg_dataout_1512_port, 
      bus_reg_dataout_1511_port, bus_reg_dataout_1510_port, 
      bus_reg_dataout_1509_port, bus_reg_dataout_1508_port, 
      bus_reg_dataout_1507_port, bus_reg_dataout_1506_port, 
      bus_reg_dataout_1505_port, bus_reg_dataout_1504_port, 
      bus_reg_dataout_1503_port, bus_reg_dataout_1502_port, 
      bus_reg_dataout_1501_port, bus_reg_dataout_1500_port, 
      bus_reg_dataout_1499_port, bus_reg_dataout_1498_port, 
      bus_reg_dataout_1497_port, bus_reg_dataout_1496_port, 
      bus_reg_dataout_1495_port, bus_reg_dataout_1494_port, 
      bus_reg_dataout_1493_port, bus_reg_dataout_1492_port, 
      bus_reg_dataout_1491_port, bus_reg_dataout_1490_port, 
      bus_reg_dataout_1489_port, bus_reg_dataout_1488_port, 
      bus_reg_dataout_1487_port, bus_reg_dataout_1486_port, 
      bus_reg_dataout_1485_port, bus_reg_dataout_1484_port, 
      bus_reg_dataout_1483_port, bus_reg_dataout_1482_port, 
      bus_reg_dataout_1481_port, bus_reg_dataout_1480_port, 
      bus_reg_dataout_1479_port, bus_reg_dataout_1478_port, 
      bus_reg_dataout_1477_port, bus_reg_dataout_1476_port, 
      bus_reg_dataout_1475_port, bus_reg_dataout_1474_port, 
      bus_reg_dataout_1473_port, bus_reg_dataout_1472_port, 
      bus_reg_dataout_1471_port, bus_reg_dataout_1470_port, 
      bus_reg_dataout_1469_port, bus_reg_dataout_1468_port, 
      bus_reg_dataout_1467_port, bus_reg_dataout_1466_port, 
      bus_reg_dataout_1465_port, bus_reg_dataout_1464_port, 
      bus_reg_dataout_1463_port, bus_reg_dataout_1462_port, 
      bus_reg_dataout_1461_port, bus_reg_dataout_1460_port, 
      bus_reg_dataout_1459_port, bus_reg_dataout_1458_port, 
      bus_reg_dataout_1457_port, bus_reg_dataout_1456_port, 
      bus_reg_dataout_1455_port, bus_reg_dataout_1454_port, 
      bus_reg_dataout_1453_port, bus_reg_dataout_1452_port, 
      bus_reg_dataout_1451_port, bus_reg_dataout_1450_port, 
      bus_reg_dataout_1449_port, bus_reg_dataout_1448_port, 
      bus_reg_dataout_1447_port, bus_reg_dataout_1446_port, 
      bus_reg_dataout_1445_port, bus_reg_dataout_1444_port, 
      bus_reg_dataout_1443_port, bus_reg_dataout_1442_port, 
      bus_reg_dataout_1441_port, bus_reg_dataout_1440_port, 
      bus_reg_dataout_1439_port, bus_reg_dataout_1438_port, 
      bus_reg_dataout_1437_port, bus_reg_dataout_1436_port, 
      bus_reg_dataout_1435_port, bus_reg_dataout_1434_port, 
      bus_reg_dataout_1433_port, bus_reg_dataout_1432_port, 
      bus_reg_dataout_1431_port, bus_reg_dataout_1430_port, 
      bus_reg_dataout_1429_port, bus_reg_dataout_1428_port, 
      bus_reg_dataout_1427_port, bus_reg_dataout_1426_port, 
      bus_reg_dataout_1425_port, bus_reg_dataout_1424_port, 
      bus_reg_dataout_1423_port, bus_reg_dataout_1422_port, 
      bus_reg_dataout_1421_port, bus_reg_dataout_1420_port, 
      bus_reg_dataout_1419_port, bus_reg_dataout_1418_port, 
      bus_reg_dataout_1417_port, bus_reg_dataout_1416_port, 
      bus_reg_dataout_1415_port, bus_reg_dataout_1414_port, 
      bus_reg_dataout_1413_port, bus_reg_dataout_1412_port, 
      bus_reg_dataout_1411_port, bus_reg_dataout_1410_port, 
      bus_reg_dataout_1409_port, bus_reg_dataout_1408_port, 
      bus_reg_dataout_1407_port, bus_reg_dataout_1406_port, 
      bus_reg_dataout_1405_port, bus_reg_dataout_1404_port, 
      bus_reg_dataout_1403_port, bus_reg_dataout_1402_port, 
      bus_reg_dataout_1401_port, bus_reg_dataout_1400_port, 
      bus_reg_dataout_1399_port, bus_reg_dataout_1398_port, 
      bus_reg_dataout_1397_port, bus_reg_dataout_1396_port, 
      bus_reg_dataout_1395_port, bus_reg_dataout_1394_port, 
      bus_reg_dataout_1393_port, bus_reg_dataout_1392_port, 
      bus_reg_dataout_1391_port, bus_reg_dataout_1390_port, 
      bus_reg_dataout_1389_port, bus_reg_dataout_1388_port, 
      bus_reg_dataout_1387_port, bus_reg_dataout_1386_port, 
      bus_reg_dataout_1385_port, bus_reg_dataout_1384_port, 
      bus_reg_dataout_1383_port, bus_reg_dataout_1382_port, 
      bus_reg_dataout_1381_port, bus_reg_dataout_1380_port, 
      bus_reg_dataout_1379_port, bus_reg_dataout_1378_port, 
      bus_reg_dataout_1377_port, bus_reg_dataout_1376_port, 
      bus_reg_dataout_1375_port, bus_reg_dataout_1374_port, 
      bus_reg_dataout_1373_port, bus_reg_dataout_1372_port, 
      bus_reg_dataout_1371_port, bus_reg_dataout_1370_port, 
      bus_reg_dataout_1369_port, bus_reg_dataout_1368_port, 
      bus_reg_dataout_1367_port, bus_reg_dataout_1366_port, 
      bus_reg_dataout_1365_port, bus_reg_dataout_1364_port, 
      bus_reg_dataout_1363_port, bus_reg_dataout_1362_port, 
      bus_reg_dataout_1361_port, bus_reg_dataout_1360_port, 
      bus_reg_dataout_1359_port, bus_reg_dataout_1358_port, 
      bus_reg_dataout_1357_port, bus_reg_dataout_1356_port, 
      bus_reg_dataout_1355_port, bus_reg_dataout_1354_port, 
      bus_reg_dataout_1353_port, bus_reg_dataout_1352_port, 
      bus_reg_dataout_1351_port, bus_reg_dataout_1350_port, 
      bus_reg_dataout_1349_port, bus_reg_dataout_1348_port, 
      bus_reg_dataout_1347_port, bus_reg_dataout_1346_port, 
      bus_reg_dataout_1345_port, bus_reg_dataout_1344_port, 
      bus_reg_dataout_1343_port, bus_reg_dataout_1342_port, 
      bus_reg_dataout_1341_port, bus_reg_dataout_1340_port, 
      bus_reg_dataout_1339_port, bus_reg_dataout_1338_port, 
      bus_reg_dataout_1337_port, bus_reg_dataout_1336_port, 
      bus_reg_dataout_1335_port, bus_reg_dataout_1334_port, 
      bus_reg_dataout_1333_port, bus_reg_dataout_1332_port, 
      bus_reg_dataout_1331_port, bus_reg_dataout_1330_port, 
      bus_reg_dataout_1329_port, bus_reg_dataout_1328_port, 
      bus_reg_dataout_1327_port, bus_reg_dataout_1326_port, 
      bus_reg_dataout_1325_port, bus_reg_dataout_1324_port, 
      bus_reg_dataout_1323_port, bus_reg_dataout_1322_port, 
      bus_reg_dataout_1321_port, bus_reg_dataout_1320_port, 
      bus_reg_dataout_1319_port, bus_reg_dataout_1318_port, 
      bus_reg_dataout_1317_port, bus_reg_dataout_1316_port, 
      bus_reg_dataout_1315_port, bus_reg_dataout_1314_port, 
      bus_reg_dataout_1313_port, bus_reg_dataout_1312_port, 
      bus_reg_dataout_1311_port, bus_reg_dataout_1310_port, 
      bus_reg_dataout_1309_port, bus_reg_dataout_1308_port, 
      bus_reg_dataout_1307_port, bus_reg_dataout_1306_port, 
      bus_reg_dataout_1305_port, bus_reg_dataout_1304_port, 
      bus_reg_dataout_1303_port, bus_reg_dataout_1302_port, 
      bus_reg_dataout_1301_port, bus_reg_dataout_1300_port, 
      bus_reg_dataout_1299_port, bus_reg_dataout_1298_port, 
      bus_reg_dataout_1297_port, bus_reg_dataout_1296_port, 
      bus_reg_dataout_1295_port, bus_reg_dataout_1294_port, 
      bus_reg_dataout_1293_port, bus_reg_dataout_1292_port, 
      bus_reg_dataout_1291_port, bus_reg_dataout_1290_port, 
      bus_reg_dataout_1289_port, bus_reg_dataout_1288_port, 
      bus_reg_dataout_1287_port, bus_reg_dataout_1286_port, 
      bus_reg_dataout_1285_port, bus_reg_dataout_1284_port, 
      bus_reg_dataout_1283_port, bus_reg_dataout_1282_port, 
      bus_reg_dataout_1281_port, bus_reg_dataout_1280_port, 
      bus_reg_dataout_1279_port, bus_reg_dataout_1278_port, 
      bus_reg_dataout_1277_port, bus_reg_dataout_1276_port, 
      bus_reg_dataout_1275_port, bus_reg_dataout_1274_port, 
      bus_reg_dataout_1273_port, bus_reg_dataout_1272_port, 
      bus_reg_dataout_1271_port, bus_reg_dataout_1270_port, 
      bus_reg_dataout_1269_port, bus_reg_dataout_1268_port, 
      bus_reg_dataout_1267_port, bus_reg_dataout_1266_port, 
      bus_reg_dataout_1265_port, bus_reg_dataout_1264_port, 
      bus_reg_dataout_1263_port, bus_reg_dataout_1262_port, 
      bus_reg_dataout_1261_port, bus_reg_dataout_1260_port, 
      bus_reg_dataout_1259_port, bus_reg_dataout_1258_port, 
      bus_reg_dataout_1257_port, bus_reg_dataout_1256_port, 
      bus_reg_dataout_1255_port, bus_reg_dataout_1254_port, 
      bus_reg_dataout_1253_port, bus_reg_dataout_1252_port, 
      bus_reg_dataout_1251_port, bus_reg_dataout_1250_port, 
      bus_reg_dataout_1249_port, bus_reg_dataout_1248_port, 
      bus_reg_dataout_1247_port, bus_reg_dataout_1246_port, 
      bus_reg_dataout_1245_port, bus_reg_dataout_1244_port, 
      bus_reg_dataout_1243_port, bus_reg_dataout_1242_port, 
      bus_reg_dataout_1241_port, bus_reg_dataout_1240_port, 
      bus_reg_dataout_1239_port, bus_reg_dataout_1238_port, 
      bus_reg_dataout_1237_port, bus_reg_dataout_1236_port, 
      bus_reg_dataout_1235_port, bus_reg_dataout_1234_port, 
      bus_reg_dataout_1233_port, bus_reg_dataout_1232_port, 
      bus_reg_dataout_1231_port, bus_reg_dataout_1230_port, 
      bus_reg_dataout_1229_port, bus_reg_dataout_1228_port, 
      bus_reg_dataout_1227_port, bus_reg_dataout_1226_port, 
      bus_reg_dataout_1225_port, bus_reg_dataout_1224_port, 
      bus_reg_dataout_1223_port, bus_reg_dataout_1222_port, 
      bus_reg_dataout_1221_port, bus_reg_dataout_1220_port, 
      bus_reg_dataout_1219_port, bus_reg_dataout_1218_port, 
      bus_reg_dataout_1217_port, bus_reg_dataout_1216_port, 
      bus_reg_dataout_1215_port, bus_reg_dataout_1214_port, 
      bus_reg_dataout_1213_port, bus_reg_dataout_1212_port, 
      bus_reg_dataout_1211_port, bus_reg_dataout_1210_port, 
      bus_reg_dataout_1209_port, bus_reg_dataout_1208_port, 
      bus_reg_dataout_1207_port, bus_reg_dataout_1206_port, 
      bus_reg_dataout_1205_port, bus_reg_dataout_1204_port, 
      bus_reg_dataout_1203_port, bus_reg_dataout_1202_port, 
      bus_reg_dataout_1201_port, bus_reg_dataout_1200_port, 
      bus_reg_dataout_1199_port, bus_reg_dataout_1198_port, 
      bus_reg_dataout_1197_port, bus_reg_dataout_1196_port, 
      bus_reg_dataout_1195_port, bus_reg_dataout_1194_port, 
      bus_reg_dataout_1193_port, bus_reg_dataout_1192_port, 
      bus_reg_dataout_1191_port, bus_reg_dataout_1190_port, 
      bus_reg_dataout_1189_port, bus_reg_dataout_1188_port, 
      bus_reg_dataout_1187_port, bus_reg_dataout_1186_port, 
      bus_reg_dataout_1185_port, bus_reg_dataout_1184_port, 
      bus_reg_dataout_1183_port, bus_reg_dataout_1182_port, 
      bus_reg_dataout_1181_port, bus_reg_dataout_1180_port, 
      bus_reg_dataout_1179_port, bus_reg_dataout_1178_port, 
      bus_reg_dataout_1177_port, bus_reg_dataout_1176_port, 
      bus_reg_dataout_1175_port, bus_reg_dataout_1174_port, 
      bus_reg_dataout_1173_port, bus_reg_dataout_1172_port, 
      bus_reg_dataout_1171_port, bus_reg_dataout_1170_port, 
      bus_reg_dataout_1169_port, bus_reg_dataout_1168_port, 
      bus_reg_dataout_1167_port, bus_reg_dataout_1166_port, 
      bus_reg_dataout_1165_port, bus_reg_dataout_1164_port, 
      bus_reg_dataout_1163_port, bus_reg_dataout_1162_port, 
      bus_reg_dataout_1161_port, bus_reg_dataout_1160_port, 
      bus_reg_dataout_1159_port, bus_reg_dataout_1158_port, 
      bus_reg_dataout_1157_port, bus_reg_dataout_1156_port, 
      bus_reg_dataout_1155_port, bus_reg_dataout_1154_port, 
      bus_reg_dataout_1153_port, bus_reg_dataout_1152_port, 
      bus_reg_dataout_1151_port, bus_reg_dataout_1150_port, 
      bus_reg_dataout_1149_port, bus_reg_dataout_1148_port, 
      bus_reg_dataout_1147_port, bus_reg_dataout_1146_port, 
      bus_reg_dataout_1145_port, bus_reg_dataout_1144_port, 
      bus_reg_dataout_1143_port, bus_reg_dataout_1142_port, 
      bus_reg_dataout_1141_port, bus_reg_dataout_1140_port, 
      bus_reg_dataout_1139_port, bus_reg_dataout_1138_port, 
      bus_reg_dataout_1137_port, bus_reg_dataout_1136_port, 
      bus_reg_dataout_1135_port, bus_reg_dataout_1134_port, 
      bus_reg_dataout_1133_port, bus_reg_dataout_1132_port, 
      bus_reg_dataout_1131_port, bus_reg_dataout_1130_port, 
      bus_reg_dataout_1129_port, bus_reg_dataout_1128_port, 
      bus_reg_dataout_1127_port, bus_reg_dataout_1126_port, 
      bus_reg_dataout_1125_port, bus_reg_dataout_1124_port, 
      bus_reg_dataout_1123_port, bus_reg_dataout_1122_port, 
      bus_reg_dataout_1121_port, bus_reg_dataout_1120_port, 
      bus_reg_dataout_1119_port, bus_reg_dataout_1118_port, 
      bus_reg_dataout_1117_port, bus_reg_dataout_1116_port, 
      bus_reg_dataout_1115_port, bus_reg_dataout_1114_port, 
      bus_reg_dataout_1113_port, bus_reg_dataout_1112_port, 
      bus_reg_dataout_1111_port, bus_reg_dataout_1110_port, 
      bus_reg_dataout_1109_port, bus_reg_dataout_1108_port, 
      bus_reg_dataout_1107_port, bus_reg_dataout_1106_port, 
      bus_reg_dataout_1105_port, bus_reg_dataout_1104_port, 
      bus_reg_dataout_1103_port, bus_reg_dataout_1102_port, 
      bus_reg_dataout_1101_port, bus_reg_dataout_1100_port, 
      bus_reg_dataout_1099_port, bus_reg_dataout_1098_port, 
      bus_reg_dataout_1097_port, bus_reg_dataout_1096_port, 
      bus_reg_dataout_1095_port, bus_reg_dataout_1094_port, 
      bus_reg_dataout_1093_port, bus_reg_dataout_1092_port, 
      bus_reg_dataout_1091_port, bus_reg_dataout_1090_port, 
      bus_reg_dataout_1089_port, bus_reg_dataout_1088_port, 
      bus_reg_dataout_1087_port, bus_reg_dataout_1086_port, 
      bus_reg_dataout_1085_port, bus_reg_dataout_1084_port, 
      bus_reg_dataout_1083_port, bus_reg_dataout_1082_port, 
      bus_reg_dataout_1081_port, bus_reg_dataout_1080_port, 
      bus_reg_dataout_1079_port, bus_reg_dataout_1078_port, 
      bus_reg_dataout_1077_port, bus_reg_dataout_1076_port, 
      bus_reg_dataout_1075_port, bus_reg_dataout_1074_port, 
      bus_reg_dataout_1073_port, bus_reg_dataout_1072_port, 
      bus_reg_dataout_1071_port, bus_reg_dataout_1070_port, 
      bus_reg_dataout_1069_port, bus_reg_dataout_1068_port, 
      bus_reg_dataout_1067_port, bus_reg_dataout_1066_port, 
      bus_reg_dataout_1065_port, bus_reg_dataout_1064_port, 
      bus_reg_dataout_1063_port, bus_reg_dataout_1062_port, 
      bus_reg_dataout_1061_port, bus_reg_dataout_1060_port, 
      bus_reg_dataout_1059_port, bus_reg_dataout_1058_port, 
      bus_reg_dataout_1057_port, bus_reg_dataout_1056_port, 
      bus_reg_dataout_1055_port, bus_reg_dataout_1054_port, 
      bus_reg_dataout_1053_port, bus_reg_dataout_1052_port, 
      bus_reg_dataout_1051_port, bus_reg_dataout_1050_port, 
      bus_reg_dataout_1049_port, bus_reg_dataout_1048_port, 
      bus_reg_dataout_1047_port, bus_reg_dataout_1046_port, 
      bus_reg_dataout_1045_port, bus_reg_dataout_1044_port, 
      bus_reg_dataout_1043_port, bus_reg_dataout_1042_port, 
      bus_reg_dataout_1041_port, bus_reg_dataout_1040_port, 
      bus_reg_dataout_1039_port, bus_reg_dataout_1038_port, 
      bus_reg_dataout_1037_port, bus_reg_dataout_1036_port, 
      bus_reg_dataout_1035_port, bus_reg_dataout_1034_port, 
      bus_reg_dataout_1033_port, bus_reg_dataout_1032_port, 
      bus_reg_dataout_1031_port, bus_reg_dataout_1030_port, 
      bus_reg_dataout_1029_port, bus_reg_dataout_1028_port, 
      bus_reg_dataout_1027_port, bus_reg_dataout_1026_port, 
      bus_reg_dataout_1025_port, bus_reg_dataout_1024_port, 
      bus_reg_dataout_1023_port, bus_reg_dataout_1022_port, 
      bus_reg_dataout_1021_port, bus_reg_dataout_1020_port, 
      bus_reg_dataout_1019_port, bus_reg_dataout_1018_port, 
      bus_reg_dataout_1017_port, bus_reg_dataout_1016_port, 
      bus_reg_dataout_1015_port, bus_reg_dataout_1014_port, 
      bus_reg_dataout_1013_port, bus_reg_dataout_1012_port, 
      bus_reg_dataout_1011_port, bus_reg_dataout_1010_port, 
      bus_reg_dataout_1009_port, bus_reg_dataout_1008_port, 
      bus_reg_dataout_1007_port, bus_reg_dataout_1006_port, 
      bus_reg_dataout_1005_port, bus_reg_dataout_1004_port, 
      bus_reg_dataout_1003_port, bus_reg_dataout_1002_port, 
      bus_reg_dataout_1001_port, bus_reg_dataout_1000_port, 
      bus_reg_dataout_999_port, bus_reg_dataout_998_port, 
      bus_reg_dataout_997_port, bus_reg_dataout_996_port, 
      bus_reg_dataout_995_port, bus_reg_dataout_994_port, 
      bus_reg_dataout_993_port, bus_reg_dataout_992_port, 
      bus_reg_dataout_991_port, bus_reg_dataout_990_port, 
      bus_reg_dataout_989_port, bus_reg_dataout_988_port, 
      bus_reg_dataout_987_port, bus_reg_dataout_986_port, 
      bus_reg_dataout_985_port, bus_reg_dataout_984_port, 
      bus_reg_dataout_983_port, bus_reg_dataout_982_port, 
      bus_reg_dataout_981_port, bus_reg_dataout_980_port, 
      bus_reg_dataout_979_port, bus_reg_dataout_978_port, 
      bus_reg_dataout_977_port, bus_reg_dataout_976_port, 
      bus_reg_dataout_975_port, bus_reg_dataout_974_port, 
      bus_reg_dataout_973_port, bus_reg_dataout_972_port, 
      bus_reg_dataout_971_port, bus_reg_dataout_970_port, 
      bus_reg_dataout_969_port, bus_reg_dataout_968_port, 
      bus_reg_dataout_967_port, bus_reg_dataout_966_port, 
      bus_reg_dataout_965_port, bus_reg_dataout_964_port, 
      bus_reg_dataout_963_port, bus_reg_dataout_962_port, 
      bus_reg_dataout_961_port, bus_reg_dataout_960_port, 
      bus_reg_dataout_959_port, bus_reg_dataout_958_port, 
      bus_reg_dataout_957_port, bus_reg_dataout_956_port, 
      bus_reg_dataout_955_port, bus_reg_dataout_954_port, 
      bus_reg_dataout_953_port, bus_reg_dataout_952_port, 
      bus_reg_dataout_951_port, bus_reg_dataout_950_port, 
      bus_reg_dataout_949_port, bus_reg_dataout_948_port, 
      bus_reg_dataout_947_port, bus_reg_dataout_946_port, 
      bus_reg_dataout_945_port, bus_reg_dataout_944_port, 
      bus_reg_dataout_943_port, bus_reg_dataout_942_port, 
      bus_reg_dataout_941_port, bus_reg_dataout_940_port, 
      bus_reg_dataout_939_port, bus_reg_dataout_938_port, 
      bus_reg_dataout_937_port, bus_reg_dataout_936_port, 
      bus_reg_dataout_935_port, bus_reg_dataout_934_port, 
      bus_reg_dataout_933_port, bus_reg_dataout_932_port, 
      bus_reg_dataout_931_port, bus_reg_dataout_930_port, 
      bus_reg_dataout_929_port, bus_reg_dataout_928_port, 
      bus_reg_dataout_927_port, bus_reg_dataout_926_port, 
      bus_reg_dataout_925_port, bus_reg_dataout_924_port, 
      bus_reg_dataout_923_port, bus_reg_dataout_922_port, 
      bus_reg_dataout_921_port, bus_reg_dataout_920_port, 
      bus_reg_dataout_919_port, bus_reg_dataout_918_port, 
      bus_reg_dataout_917_port, bus_reg_dataout_916_port, 
      bus_reg_dataout_915_port, bus_reg_dataout_914_port, 
      bus_reg_dataout_913_port, bus_reg_dataout_912_port, 
      bus_reg_dataout_911_port, bus_reg_dataout_910_port, 
      bus_reg_dataout_909_port, bus_reg_dataout_908_port, 
      bus_reg_dataout_907_port, bus_reg_dataout_906_port, 
      bus_reg_dataout_905_port, bus_reg_dataout_904_port, 
      bus_reg_dataout_903_port, bus_reg_dataout_902_port, 
      bus_reg_dataout_901_port, bus_reg_dataout_900_port, 
      bus_reg_dataout_899_port, bus_reg_dataout_898_port, 
      bus_reg_dataout_897_port, bus_reg_dataout_896_port, 
      bus_reg_dataout_895_port, bus_reg_dataout_894_port, 
      bus_reg_dataout_893_port, bus_reg_dataout_892_port, 
      bus_reg_dataout_891_port, bus_reg_dataout_890_port, 
      bus_reg_dataout_889_port, bus_reg_dataout_888_port, 
      bus_reg_dataout_887_port, bus_reg_dataout_886_port, 
      bus_reg_dataout_885_port, bus_reg_dataout_884_port, 
      bus_reg_dataout_883_port, bus_reg_dataout_882_port, 
      bus_reg_dataout_881_port, bus_reg_dataout_880_port, 
      bus_reg_dataout_879_port, bus_reg_dataout_878_port, 
      bus_reg_dataout_877_port, bus_reg_dataout_876_port, 
      bus_reg_dataout_875_port, bus_reg_dataout_874_port, 
      bus_reg_dataout_873_port, bus_reg_dataout_872_port, 
      bus_reg_dataout_871_port, bus_reg_dataout_870_port, 
      bus_reg_dataout_869_port, bus_reg_dataout_868_port, 
      bus_reg_dataout_867_port, bus_reg_dataout_866_port, 
      bus_reg_dataout_865_port, bus_reg_dataout_864_port, 
      bus_reg_dataout_863_port, bus_reg_dataout_862_port, 
      bus_reg_dataout_861_port, bus_reg_dataout_860_port, 
      bus_reg_dataout_859_port, bus_reg_dataout_858_port, 
      bus_reg_dataout_857_port, bus_reg_dataout_856_port, 
      bus_reg_dataout_855_port, bus_reg_dataout_854_port, 
      bus_reg_dataout_853_port, bus_reg_dataout_852_port, 
      bus_reg_dataout_851_port, bus_reg_dataout_850_port, 
      bus_reg_dataout_849_port, bus_reg_dataout_848_port, 
      bus_reg_dataout_847_port, bus_reg_dataout_846_port, 
      bus_reg_dataout_845_port, bus_reg_dataout_844_port, 
      bus_reg_dataout_843_port, bus_reg_dataout_842_port, 
      bus_reg_dataout_841_port, bus_reg_dataout_840_port, 
      bus_reg_dataout_839_port, bus_reg_dataout_838_port, 
      bus_reg_dataout_837_port, bus_reg_dataout_836_port, 
      bus_reg_dataout_835_port, bus_reg_dataout_834_port, 
      bus_reg_dataout_833_port, bus_reg_dataout_832_port, 
      bus_reg_dataout_831_port, bus_reg_dataout_830_port, 
      bus_reg_dataout_829_port, bus_reg_dataout_828_port, 
      bus_reg_dataout_827_port, bus_reg_dataout_826_port, 
      bus_reg_dataout_825_port, bus_reg_dataout_824_port, 
      bus_reg_dataout_823_port, bus_reg_dataout_822_port, 
      bus_reg_dataout_821_port, bus_reg_dataout_820_port, 
      bus_reg_dataout_819_port, bus_reg_dataout_818_port, 
      bus_reg_dataout_817_port, bus_reg_dataout_816_port, 
      bus_reg_dataout_815_port, bus_reg_dataout_814_port, 
      bus_reg_dataout_813_port, bus_reg_dataout_812_port, 
      bus_reg_dataout_811_port, bus_reg_dataout_810_port, 
      bus_reg_dataout_809_port, bus_reg_dataout_808_port, 
      bus_reg_dataout_807_port, bus_reg_dataout_806_port, 
      bus_reg_dataout_805_port, bus_reg_dataout_804_port, 
      bus_reg_dataout_803_port, bus_reg_dataout_802_port, 
      bus_reg_dataout_801_port, bus_reg_dataout_800_port, 
      bus_reg_dataout_799_port, bus_reg_dataout_798_port, 
      bus_reg_dataout_797_port, bus_reg_dataout_796_port, 
      bus_reg_dataout_795_port, bus_reg_dataout_794_port, 
      bus_reg_dataout_793_port, bus_reg_dataout_792_port, 
      bus_reg_dataout_791_port, bus_reg_dataout_790_port, 
      bus_reg_dataout_789_port, bus_reg_dataout_788_port, 
      bus_reg_dataout_787_port, bus_reg_dataout_786_port, 
      bus_reg_dataout_785_port, bus_reg_dataout_784_port, 
      bus_reg_dataout_783_port, bus_reg_dataout_782_port, 
      bus_reg_dataout_781_port, bus_reg_dataout_780_port, 
      bus_reg_dataout_779_port, bus_reg_dataout_778_port, 
      bus_reg_dataout_777_port, bus_reg_dataout_776_port, 
      bus_reg_dataout_775_port, bus_reg_dataout_774_port, 
      bus_reg_dataout_773_port, bus_reg_dataout_772_port, 
      bus_reg_dataout_771_port, bus_reg_dataout_770_port, 
      bus_reg_dataout_769_port, bus_reg_dataout_768_port, 
      bus_reg_dataout_767_port, bus_reg_dataout_766_port, 
      bus_reg_dataout_765_port, bus_reg_dataout_764_port, 
      bus_reg_dataout_763_port, bus_reg_dataout_762_port, 
      bus_reg_dataout_761_port, bus_reg_dataout_760_port, 
      bus_reg_dataout_759_port, bus_reg_dataout_758_port, 
      bus_reg_dataout_757_port, bus_reg_dataout_756_port, 
      bus_reg_dataout_755_port, bus_reg_dataout_754_port, 
      bus_reg_dataout_753_port, bus_reg_dataout_752_port, 
      bus_reg_dataout_751_port, bus_reg_dataout_750_port, 
      bus_reg_dataout_749_port, bus_reg_dataout_748_port, 
      bus_reg_dataout_747_port, bus_reg_dataout_746_port, 
      bus_reg_dataout_745_port, bus_reg_dataout_744_port, 
      bus_reg_dataout_743_port, bus_reg_dataout_742_port, 
      bus_reg_dataout_741_port, bus_reg_dataout_740_port, 
      bus_reg_dataout_739_port, bus_reg_dataout_738_port, 
      bus_reg_dataout_737_port, bus_reg_dataout_736_port, 
      bus_reg_dataout_735_port, bus_reg_dataout_734_port, 
      bus_reg_dataout_733_port, bus_reg_dataout_732_port, 
      bus_reg_dataout_731_port, bus_reg_dataout_730_port, 
      bus_reg_dataout_729_port, bus_reg_dataout_728_port, 
      bus_reg_dataout_727_port, bus_reg_dataout_726_port, 
      bus_reg_dataout_725_port, bus_reg_dataout_724_port, 
      bus_reg_dataout_723_port, bus_reg_dataout_722_port, 
      bus_reg_dataout_721_port, bus_reg_dataout_720_port, 
      bus_reg_dataout_719_port, bus_reg_dataout_718_port, 
      bus_reg_dataout_717_port, bus_reg_dataout_716_port, 
      bus_reg_dataout_715_port, bus_reg_dataout_714_port, 
      bus_reg_dataout_713_port, bus_reg_dataout_712_port, 
      bus_reg_dataout_711_port, bus_reg_dataout_710_port, 
      bus_reg_dataout_709_port, bus_reg_dataout_708_port, 
      bus_reg_dataout_707_port, bus_reg_dataout_706_port, 
      bus_reg_dataout_705_port, bus_reg_dataout_704_port, 
      bus_reg_dataout_703_port, bus_reg_dataout_702_port, 
      bus_reg_dataout_701_port, bus_reg_dataout_700_port, 
      bus_reg_dataout_699_port, bus_reg_dataout_698_port, 
      bus_reg_dataout_697_port, bus_reg_dataout_696_port, 
      bus_reg_dataout_695_port, bus_reg_dataout_694_port, 
      bus_reg_dataout_693_port, bus_reg_dataout_692_port, 
      bus_reg_dataout_691_port, bus_reg_dataout_690_port, 
      bus_reg_dataout_689_port, bus_reg_dataout_688_port, 
      bus_reg_dataout_687_port, bus_reg_dataout_686_port, 
      bus_reg_dataout_685_port, bus_reg_dataout_684_port, 
      bus_reg_dataout_683_port, bus_reg_dataout_682_port, 
      bus_reg_dataout_681_port, bus_reg_dataout_680_port, 
      bus_reg_dataout_679_port, bus_reg_dataout_678_port, 
      bus_reg_dataout_677_port, bus_reg_dataout_676_port, 
      bus_reg_dataout_675_port, bus_reg_dataout_674_port, 
      bus_reg_dataout_673_port, bus_reg_dataout_672_port, 
      bus_reg_dataout_671_port, bus_reg_dataout_670_port, 
      bus_reg_dataout_669_port, bus_reg_dataout_668_port, 
      bus_reg_dataout_667_port, bus_reg_dataout_666_port, 
      bus_reg_dataout_665_port, bus_reg_dataout_664_port, 
      bus_reg_dataout_663_port, bus_reg_dataout_662_port, 
      bus_reg_dataout_661_port, bus_reg_dataout_660_port, 
      bus_reg_dataout_659_port, bus_reg_dataout_658_port, 
      bus_reg_dataout_657_port, bus_reg_dataout_656_port, 
      bus_reg_dataout_655_port, bus_reg_dataout_654_port, 
      bus_reg_dataout_653_port, bus_reg_dataout_652_port, 
      bus_reg_dataout_651_port, bus_reg_dataout_650_port, 
      bus_reg_dataout_649_port, bus_reg_dataout_648_port, 
      bus_reg_dataout_647_port, bus_reg_dataout_646_port, 
      bus_reg_dataout_645_port, bus_reg_dataout_644_port, 
      bus_reg_dataout_643_port, bus_reg_dataout_642_port, 
      bus_reg_dataout_641_port, bus_reg_dataout_640_port, 
      bus_reg_dataout_639_port, bus_reg_dataout_638_port, 
      bus_reg_dataout_637_port, bus_reg_dataout_636_port, 
      bus_reg_dataout_635_port, bus_reg_dataout_634_port, 
      bus_reg_dataout_633_port, bus_reg_dataout_632_port, 
      bus_reg_dataout_631_port, bus_reg_dataout_630_port, 
      bus_reg_dataout_629_port, bus_reg_dataout_628_port, 
      bus_reg_dataout_627_port, bus_reg_dataout_626_port, 
      bus_reg_dataout_625_port, bus_reg_dataout_624_port, 
      bus_reg_dataout_623_port, bus_reg_dataout_622_port, 
      bus_reg_dataout_621_port, bus_reg_dataout_620_port, 
      bus_reg_dataout_619_port, bus_reg_dataout_618_port, 
      bus_reg_dataout_617_port, bus_reg_dataout_616_port, 
      bus_reg_dataout_615_port, bus_reg_dataout_614_port, 
      bus_reg_dataout_613_port, bus_reg_dataout_612_port, 
      bus_reg_dataout_611_port, bus_reg_dataout_610_port, 
      bus_reg_dataout_609_port, bus_reg_dataout_608_port, 
      bus_reg_dataout_607_port, bus_reg_dataout_606_port, 
      bus_reg_dataout_605_port, bus_reg_dataout_604_port, 
      bus_reg_dataout_603_port, bus_reg_dataout_602_port, 
      bus_reg_dataout_601_port, bus_reg_dataout_600_port, 
      bus_reg_dataout_599_port, bus_reg_dataout_598_port, 
      bus_reg_dataout_597_port, bus_reg_dataout_596_port, 
      bus_reg_dataout_595_port, bus_reg_dataout_594_port, 
      bus_reg_dataout_593_port, bus_reg_dataout_592_port, 
      bus_reg_dataout_591_port, bus_reg_dataout_590_port, 
      bus_reg_dataout_589_port, bus_reg_dataout_588_port, 
      bus_reg_dataout_587_port, bus_reg_dataout_586_port, 
      bus_reg_dataout_585_port, bus_reg_dataout_584_port, 
      bus_reg_dataout_583_port, bus_reg_dataout_582_port, 
      bus_reg_dataout_581_port, bus_reg_dataout_580_port, 
      bus_reg_dataout_579_port, bus_reg_dataout_578_port, 
      bus_reg_dataout_577_port, bus_reg_dataout_576_port, 
      bus_reg_dataout_575_port, bus_reg_dataout_574_port, 
      bus_reg_dataout_573_port, bus_reg_dataout_572_port, 
      bus_reg_dataout_571_port, bus_reg_dataout_570_port, 
      bus_reg_dataout_569_port, bus_reg_dataout_568_port, 
      bus_reg_dataout_567_port, bus_reg_dataout_566_port, 
      bus_reg_dataout_565_port, bus_reg_dataout_564_port, 
      bus_reg_dataout_563_port, bus_reg_dataout_562_port, 
      bus_reg_dataout_561_port, bus_reg_dataout_560_port, 
      bus_reg_dataout_559_port, bus_reg_dataout_558_port, 
      bus_reg_dataout_557_port, bus_reg_dataout_556_port, 
      bus_reg_dataout_555_port, bus_reg_dataout_554_port, 
      bus_reg_dataout_553_port, bus_reg_dataout_552_port, 
      bus_reg_dataout_551_port, bus_reg_dataout_550_port, 
      bus_reg_dataout_549_port, bus_reg_dataout_548_port, 
      bus_reg_dataout_547_port, bus_reg_dataout_546_port, 
      bus_reg_dataout_545_port, bus_reg_dataout_544_port, 
      bus_reg_dataout_543_port, bus_reg_dataout_542_port, 
      bus_reg_dataout_541_port, bus_reg_dataout_540_port, 
      bus_reg_dataout_539_port, bus_reg_dataout_538_port, 
      bus_reg_dataout_537_port, bus_reg_dataout_536_port, 
      bus_reg_dataout_535_port, bus_reg_dataout_534_port, 
      bus_reg_dataout_533_port, bus_reg_dataout_532_port, 
      bus_reg_dataout_531_port, bus_reg_dataout_530_port, 
      bus_reg_dataout_529_port, bus_reg_dataout_528_port, 
      bus_reg_dataout_527_port, bus_reg_dataout_526_port, 
      bus_reg_dataout_525_port, bus_reg_dataout_524_port, 
      bus_reg_dataout_523_port, bus_reg_dataout_522_port, 
      bus_reg_dataout_521_port, bus_reg_dataout_520_port, 
      bus_reg_dataout_519_port, bus_reg_dataout_518_port, 
      bus_reg_dataout_517_port, bus_reg_dataout_516_port, 
      bus_reg_dataout_515_port, bus_reg_dataout_514_port, 
      bus_reg_dataout_513_port, bus_reg_dataout_512_port, 
      bus_reg_dataout_511_port, bus_reg_dataout_510_port, 
      bus_reg_dataout_509_port, bus_reg_dataout_508_port, 
      bus_reg_dataout_507_port, bus_reg_dataout_506_port, 
      bus_reg_dataout_505_port, bus_reg_dataout_504_port, 
      bus_reg_dataout_503_port, bus_reg_dataout_502_port, 
      bus_reg_dataout_501_port, bus_reg_dataout_500_port, 
      bus_reg_dataout_499_port, bus_reg_dataout_498_port, 
      bus_reg_dataout_497_port, bus_reg_dataout_496_port, 
      bus_reg_dataout_495_port, bus_reg_dataout_494_port, 
      bus_reg_dataout_493_port, bus_reg_dataout_492_port, 
      bus_reg_dataout_491_port, bus_reg_dataout_490_port, 
      bus_reg_dataout_489_port, bus_reg_dataout_488_port, 
      bus_reg_dataout_487_port, bus_reg_dataout_486_port, 
      bus_reg_dataout_485_port, bus_reg_dataout_484_port, 
      bus_reg_dataout_483_port, bus_reg_dataout_482_port, 
      bus_reg_dataout_481_port, bus_reg_dataout_480_port, 
      bus_reg_dataout_479_port, bus_reg_dataout_478_port, 
      bus_reg_dataout_477_port, bus_reg_dataout_476_port, 
      bus_reg_dataout_475_port, bus_reg_dataout_474_port, 
      bus_reg_dataout_473_port, bus_reg_dataout_472_port, 
      bus_reg_dataout_471_port, bus_reg_dataout_470_port, 
      bus_reg_dataout_469_port, bus_reg_dataout_468_port, 
      bus_reg_dataout_467_port, bus_reg_dataout_466_port, 
      bus_reg_dataout_465_port, bus_reg_dataout_464_port, 
      bus_reg_dataout_463_port, bus_reg_dataout_462_port, 
      bus_reg_dataout_461_port, bus_reg_dataout_460_port, 
      bus_reg_dataout_459_port, bus_reg_dataout_458_port, 
      bus_reg_dataout_457_port, bus_reg_dataout_456_port, 
      bus_reg_dataout_455_port, bus_reg_dataout_454_port, 
      bus_reg_dataout_453_port, bus_reg_dataout_452_port, 
      bus_reg_dataout_451_port, bus_reg_dataout_450_port, 
      bus_reg_dataout_449_port, bus_reg_dataout_448_port, 
      bus_reg_dataout_447_port, bus_reg_dataout_446_port, 
      bus_reg_dataout_445_port, bus_reg_dataout_444_port, 
      bus_reg_dataout_443_port, bus_reg_dataout_442_port, 
      bus_reg_dataout_441_port, bus_reg_dataout_440_port, 
      bus_reg_dataout_439_port, bus_reg_dataout_438_port, 
      bus_reg_dataout_437_port, bus_reg_dataout_436_port, 
      bus_reg_dataout_435_port, bus_reg_dataout_434_port, 
      bus_reg_dataout_433_port, bus_reg_dataout_432_port, 
      bus_reg_dataout_431_port, bus_reg_dataout_430_port, 
      bus_reg_dataout_429_port, bus_reg_dataout_428_port, 
      bus_reg_dataout_427_port, bus_reg_dataout_426_port, 
      bus_reg_dataout_425_port, bus_reg_dataout_424_port, 
      bus_reg_dataout_423_port, bus_reg_dataout_422_port, 
      bus_reg_dataout_421_port, bus_reg_dataout_420_port, 
      bus_reg_dataout_419_port, bus_reg_dataout_418_port, 
      bus_reg_dataout_417_port, bus_reg_dataout_416_port, 
      bus_reg_dataout_415_port, bus_reg_dataout_414_port, 
      bus_reg_dataout_413_port, bus_reg_dataout_412_port, 
      bus_reg_dataout_411_port, bus_reg_dataout_410_port, 
      bus_reg_dataout_409_port, bus_reg_dataout_408_port, 
      bus_reg_dataout_407_port, bus_reg_dataout_406_port, 
      bus_reg_dataout_405_port, bus_reg_dataout_404_port, 
      bus_reg_dataout_403_port, bus_reg_dataout_402_port, 
      bus_reg_dataout_401_port, bus_reg_dataout_400_port, 
      bus_reg_dataout_399_port, bus_reg_dataout_398_port, 
      bus_reg_dataout_397_port, bus_reg_dataout_396_port, 
      bus_reg_dataout_395_port, bus_reg_dataout_394_port, 
      bus_reg_dataout_393_port, bus_reg_dataout_392_port, 
      bus_reg_dataout_391_port, bus_reg_dataout_390_port, 
      bus_reg_dataout_389_port, bus_reg_dataout_388_port, 
      bus_reg_dataout_387_port, bus_reg_dataout_386_port, 
      bus_reg_dataout_385_port, bus_reg_dataout_384_port, 
      bus_reg_dataout_383_port, bus_reg_dataout_382_port, 
      bus_reg_dataout_381_port, bus_reg_dataout_380_port, 
      bus_reg_dataout_379_port, bus_reg_dataout_378_port, 
      bus_reg_dataout_377_port, bus_reg_dataout_376_port, 
      bus_reg_dataout_375_port, bus_reg_dataout_374_port, 
      bus_reg_dataout_373_port, bus_reg_dataout_372_port, 
      bus_reg_dataout_371_port, bus_reg_dataout_370_port, 
      bus_reg_dataout_369_port, bus_reg_dataout_368_port, 
      bus_reg_dataout_367_port, bus_reg_dataout_366_port, 
      bus_reg_dataout_365_port, bus_reg_dataout_364_port, 
      bus_reg_dataout_363_port, bus_reg_dataout_362_port, 
      bus_reg_dataout_361_port, bus_reg_dataout_360_port, 
      bus_reg_dataout_359_port, bus_reg_dataout_358_port, 
      bus_reg_dataout_357_port, bus_reg_dataout_356_port, 
      bus_reg_dataout_355_port, bus_reg_dataout_354_port, 
      bus_reg_dataout_353_port, bus_reg_dataout_352_port, 
      bus_reg_dataout_351_port, bus_reg_dataout_350_port, 
      bus_reg_dataout_349_port, bus_reg_dataout_348_port, 
      bus_reg_dataout_347_port, bus_reg_dataout_346_port, 
      bus_reg_dataout_345_port, bus_reg_dataout_344_port, 
      bus_reg_dataout_343_port, bus_reg_dataout_342_port, 
      bus_reg_dataout_341_port, bus_reg_dataout_340_port, 
      bus_reg_dataout_339_port, bus_reg_dataout_338_port, 
      bus_reg_dataout_337_port, bus_reg_dataout_336_port, 
      bus_reg_dataout_335_port, bus_reg_dataout_334_port, 
      bus_reg_dataout_333_port, bus_reg_dataout_332_port, 
      bus_reg_dataout_331_port, bus_reg_dataout_330_port, 
      bus_reg_dataout_329_port, bus_reg_dataout_328_port, 
      bus_reg_dataout_327_port, bus_reg_dataout_326_port, 
      bus_reg_dataout_325_port, bus_reg_dataout_324_port, 
      bus_reg_dataout_323_port, bus_reg_dataout_322_port, 
      bus_reg_dataout_321_port, bus_reg_dataout_320_port, 
      bus_reg_dataout_319_port, bus_reg_dataout_318_port, 
      bus_reg_dataout_317_port, bus_reg_dataout_316_port, 
      bus_reg_dataout_315_port, bus_reg_dataout_314_port, 
      bus_reg_dataout_313_port, bus_reg_dataout_312_port, 
      bus_reg_dataout_311_port, bus_reg_dataout_310_port, 
      bus_reg_dataout_309_port, bus_reg_dataout_308_port, 
      bus_reg_dataout_307_port, bus_reg_dataout_306_port, 
      bus_reg_dataout_305_port, bus_reg_dataout_304_port, 
      bus_reg_dataout_303_port, bus_reg_dataout_302_port, 
      bus_reg_dataout_301_port, bus_reg_dataout_300_port, 
      bus_reg_dataout_299_port, bus_reg_dataout_298_port, 
      bus_reg_dataout_297_port, bus_reg_dataout_296_port, 
      bus_reg_dataout_295_port, bus_reg_dataout_294_port, 
      bus_reg_dataout_293_port, bus_reg_dataout_292_port, 
      bus_reg_dataout_291_port, bus_reg_dataout_290_port, 
      bus_reg_dataout_289_port, bus_reg_dataout_288_port, 
      bus_reg_dataout_287_port, bus_reg_dataout_286_port, 
      bus_reg_dataout_285_port, bus_reg_dataout_284_port, 
      bus_reg_dataout_283_port, bus_reg_dataout_282_port, 
      bus_reg_dataout_281_port, bus_reg_dataout_280_port, 
      bus_reg_dataout_279_port, bus_reg_dataout_278_port, 
      bus_reg_dataout_277_port, bus_reg_dataout_276_port, 
      bus_reg_dataout_275_port, bus_reg_dataout_274_port, 
      bus_reg_dataout_273_port, bus_reg_dataout_272_port, 
      bus_reg_dataout_271_port, bus_reg_dataout_270_port, 
      bus_reg_dataout_269_port, bus_reg_dataout_268_port, 
      bus_reg_dataout_267_port, bus_reg_dataout_266_port, 
      bus_reg_dataout_265_port, bus_reg_dataout_264_port, 
      bus_reg_dataout_263_port, bus_reg_dataout_262_port, 
      bus_reg_dataout_261_port, bus_reg_dataout_260_port, 
      bus_reg_dataout_259_port, bus_reg_dataout_258_port, 
      bus_reg_dataout_257_port, bus_reg_dataout_256_port, 
      bus_reg_dataout_255_port, bus_reg_dataout_254_port, 
      bus_reg_dataout_253_port, bus_reg_dataout_252_port, 
      bus_reg_dataout_251_port, bus_reg_dataout_250_port, 
      bus_reg_dataout_249_port, bus_reg_dataout_248_port, 
      bus_reg_dataout_247_port, bus_reg_dataout_246_port, 
      bus_reg_dataout_245_port, bus_reg_dataout_244_port, 
      bus_reg_dataout_243_port, bus_reg_dataout_242_port, 
      bus_reg_dataout_241_port, bus_reg_dataout_240_port, 
      bus_reg_dataout_239_port, bus_reg_dataout_238_port, 
      bus_reg_dataout_237_port, bus_reg_dataout_236_port, 
      bus_reg_dataout_235_port, bus_reg_dataout_234_port, 
      bus_reg_dataout_233_port, bus_reg_dataout_232_port, 
      bus_reg_dataout_231_port, bus_reg_dataout_230_port, 
      bus_reg_dataout_229_port, bus_reg_dataout_228_port, 
      bus_reg_dataout_227_port, bus_reg_dataout_226_port, 
      bus_reg_dataout_225_port, bus_reg_dataout_224_port, 
      bus_reg_dataout_223_port, bus_reg_dataout_222_port, 
      bus_reg_dataout_221_port, bus_reg_dataout_220_port, 
      bus_reg_dataout_219_port, bus_reg_dataout_218_port, 
      bus_reg_dataout_217_port, bus_reg_dataout_216_port, 
      bus_reg_dataout_215_port, bus_reg_dataout_214_port, 
      bus_reg_dataout_213_port, bus_reg_dataout_212_port, 
      bus_reg_dataout_211_port, bus_reg_dataout_210_port, 
      bus_reg_dataout_209_port, bus_reg_dataout_208_port, 
      bus_reg_dataout_207_port, bus_reg_dataout_206_port, 
      bus_reg_dataout_205_port, bus_reg_dataout_204_port, 
      bus_reg_dataout_203_port, bus_reg_dataout_202_port, 
      bus_reg_dataout_201_port, bus_reg_dataout_200_port, 
      bus_reg_dataout_199_port, bus_reg_dataout_198_port, 
      bus_reg_dataout_197_port, bus_reg_dataout_196_port, 
      bus_reg_dataout_195_port, bus_reg_dataout_194_port, 
      bus_reg_dataout_193_port, bus_reg_dataout_192_port, 
      bus_reg_dataout_191_port, bus_reg_dataout_190_port, 
      bus_reg_dataout_189_port, bus_reg_dataout_188_port, 
      bus_reg_dataout_187_port, bus_reg_dataout_186_port, 
      bus_reg_dataout_185_port, bus_reg_dataout_184_port, 
      bus_reg_dataout_183_port, bus_reg_dataout_182_port, 
      bus_reg_dataout_181_port, bus_reg_dataout_180_port, 
      bus_reg_dataout_179_port, bus_reg_dataout_178_port, 
      bus_reg_dataout_177_port, bus_reg_dataout_176_port, 
      bus_reg_dataout_175_port, bus_reg_dataout_174_port, 
      bus_reg_dataout_173_port, bus_reg_dataout_172_port, 
      bus_reg_dataout_171_port, bus_reg_dataout_170_port, 
      bus_reg_dataout_169_port, bus_reg_dataout_168_port, 
      bus_reg_dataout_167_port, bus_reg_dataout_166_port, 
      bus_reg_dataout_165_port, bus_reg_dataout_164_port, 
      bus_reg_dataout_163_port, bus_reg_dataout_162_port, 
      bus_reg_dataout_161_port, bus_reg_dataout_160_port, 
      bus_reg_dataout_159_port, bus_reg_dataout_158_port, 
      bus_reg_dataout_157_port, bus_reg_dataout_156_port, 
      bus_reg_dataout_155_port, bus_reg_dataout_154_port, 
      bus_reg_dataout_153_port, bus_reg_dataout_152_port, 
      bus_reg_dataout_151_port, bus_reg_dataout_150_port, 
      bus_reg_dataout_149_port, bus_reg_dataout_148_port, 
      bus_reg_dataout_147_port, bus_reg_dataout_146_port, 
      bus_reg_dataout_145_port, bus_reg_dataout_144_port, 
      bus_reg_dataout_143_port, bus_reg_dataout_142_port, 
      bus_reg_dataout_141_port, bus_reg_dataout_140_port, 
      bus_reg_dataout_139_port, bus_reg_dataout_138_port, 
      bus_reg_dataout_137_port, bus_reg_dataout_136_port, 
      bus_reg_dataout_135_port, bus_reg_dataout_134_port, 
      bus_reg_dataout_133_port, bus_reg_dataout_132_port, 
      bus_reg_dataout_131_port, bus_reg_dataout_130_port, 
      bus_reg_dataout_129_port, bus_reg_dataout_128_port, 
      bus_reg_dataout_127_port, bus_reg_dataout_126_port, 
      bus_reg_dataout_125_port, bus_reg_dataout_124_port, 
      bus_reg_dataout_123_port, bus_reg_dataout_122_port, 
      bus_reg_dataout_121_port, bus_reg_dataout_120_port, 
      bus_reg_dataout_119_port, bus_reg_dataout_118_port, 
      bus_reg_dataout_117_port, bus_reg_dataout_116_port, 
      bus_reg_dataout_115_port, bus_reg_dataout_114_port, 
      bus_reg_dataout_113_port, bus_reg_dataout_112_port, 
      bus_reg_dataout_111_port, bus_reg_dataout_110_port, 
      bus_reg_dataout_109_port, bus_reg_dataout_108_port, 
      bus_reg_dataout_107_port, bus_reg_dataout_106_port, 
      bus_reg_dataout_105_port, bus_reg_dataout_104_port, 
      bus_reg_dataout_103_port, bus_reg_dataout_102_port, 
      bus_reg_dataout_101_port, bus_reg_dataout_100_port, 
      bus_reg_dataout_99_port, bus_reg_dataout_98_port, bus_reg_dataout_97_port
      , bus_reg_dataout_96_port, bus_reg_dataout_95_port, 
      bus_reg_dataout_94_port, bus_reg_dataout_93_port, bus_reg_dataout_92_port
      , bus_reg_dataout_91_port, bus_reg_dataout_90_port, 
      bus_reg_dataout_89_port, bus_reg_dataout_88_port, bus_reg_dataout_87_port
      , bus_reg_dataout_86_port, bus_reg_dataout_85_port, 
      bus_reg_dataout_84_port, bus_reg_dataout_83_port, bus_reg_dataout_82_port
      , bus_reg_dataout_81_port, bus_reg_dataout_80_port, 
      bus_reg_dataout_79_port, bus_reg_dataout_78_port, bus_reg_dataout_77_port
      , bus_reg_dataout_76_port, bus_reg_dataout_75_port, 
      bus_reg_dataout_74_port, bus_reg_dataout_73_port, bus_reg_dataout_72_port
      , bus_reg_dataout_71_port, bus_reg_dataout_70_port, 
      bus_reg_dataout_69_port, bus_reg_dataout_68_port, bus_reg_dataout_67_port
      , bus_reg_dataout_66_port, bus_reg_dataout_65_port, 
      bus_reg_dataout_64_port, bus_reg_dataout_63_port, bus_reg_dataout_62_port
      , bus_reg_dataout_61_port, bus_reg_dataout_60_port, 
      bus_reg_dataout_59_port, bus_reg_dataout_58_port, bus_reg_dataout_57_port
      , bus_reg_dataout_56_port, bus_reg_dataout_55_port, 
      bus_reg_dataout_54_port, bus_reg_dataout_53_port, bus_reg_dataout_52_port
      , bus_reg_dataout_51_port, bus_reg_dataout_50_port, 
      bus_reg_dataout_49_port, bus_reg_dataout_48_port, bus_reg_dataout_47_port
      , bus_reg_dataout_46_port, bus_reg_dataout_45_port, 
      bus_reg_dataout_44_port, bus_reg_dataout_43_port, bus_reg_dataout_42_port
      , bus_reg_dataout_41_port, bus_reg_dataout_40_port, 
      bus_reg_dataout_39_port, bus_reg_dataout_38_port, bus_reg_dataout_37_port
      , bus_reg_dataout_36_port, bus_reg_dataout_35_port, 
      bus_reg_dataout_34_port, bus_reg_dataout_33_port, bus_reg_dataout_32_port
      , bus_reg_dataout_31_port, bus_reg_dataout_30_port, 
      bus_reg_dataout_29_port, bus_reg_dataout_28_port, bus_reg_dataout_27_port
      , bus_reg_dataout_26_port, bus_reg_dataout_25_port, 
      bus_reg_dataout_24_port, bus_reg_dataout_23_port, bus_reg_dataout_22_port
      , bus_reg_dataout_21_port, bus_reg_dataout_20_port, 
      bus_reg_dataout_19_port, bus_reg_dataout_18_port, bus_reg_dataout_17_port
      , bus_reg_dataout_16_port, bus_reg_dataout_15_port, 
      bus_reg_dataout_14_port, bus_reg_dataout_13_port, bus_reg_dataout_12_port
      , bus_reg_dataout_11_port, bus_reg_dataout_10_port, 
      bus_reg_dataout_9_port, bus_reg_dataout_8_port, bus_reg_dataout_7_port, 
      bus_reg_dataout_6_port, bus_reg_dataout_5_port, bus_reg_dataout_4_port, 
      bus_reg_dataout_3_port, bus_reg_dataout_2_port, bus_reg_dataout_1_port, 
      bus_reg_dataout_0_port, bus_selected_win_data_767_port, 
      bus_selected_win_data_766_port, bus_selected_win_data_765_port, 
      bus_selected_win_data_764_port, bus_selected_win_data_763_port, 
      bus_selected_win_data_762_port, bus_selected_win_data_761_port, 
      bus_selected_win_data_760_port, bus_selected_win_data_759_port, 
      bus_selected_win_data_758_port, bus_selected_win_data_757_port, 
      bus_selected_win_data_756_port, bus_selected_win_data_755_port, 
      bus_selected_win_data_754_port, bus_selected_win_data_753_port, 
      bus_selected_win_data_752_port, bus_selected_win_data_751_port, 
      bus_selected_win_data_750_port, bus_selected_win_data_749_port, 
      bus_selected_win_data_748_port, bus_selected_win_data_747_port, 
      bus_selected_win_data_746_port, bus_selected_win_data_745_port, 
      bus_selected_win_data_744_port, bus_selected_win_data_743_port, 
      bus_selected_win_data_742_port, bus_selected_win_data_741_port, 
      bus_selected_win_data_740_port, bus_selected_win_data_739_port, 
      bus_selected_win_data_738_port, bus_selected_win_data_737_port, 
      bus_selected_win_data_736_port, bus_selected_win_data_735_port, 
      bus_selected_win_data_734_port, bus_selected_win_data_733_port, 
      bus_selected_win_data_732_port, bus_selected_win_data_731_port, 
      bus_selected_win_data_730_port, bus_selected_win_data_729_port, 
      bus_selected_win_data_728_port, bus_selected_win_data_727_port, 
      bus_selected_win_data_726_port, bus_selected_win_data_725_port, 
      bus_selected_win_data_724_port, bus_selected_win_data_723_port, 
      bus_selected_win_data_722_port, bus_selected_win_data_721_port, 
      bus_selected_win_data_720_port, bus_selected_win_data_719_port, 
      bus_selected_win_data_718_port, bus_selected_win_data_717_port, 
      bus_selected_win_data_716_port, bus_selected_win_data_715_port, 
      bus_selected_win_data_714_port, bus_selected_win_data_713_port, 
      bus_selected_win_data_712_port, bus_selected_win_data_711_port, 
      bus_selected_win_data_710_port, bus_selected_win_data_709_port, 
      bus_selected_win_data_708_port, bus_selected_win_data_707_port, 
      bus_selected_win_data_706_port, bus_selected_win_data_705_port, 
      bus_selected_win_data_704_port, bus_selected_win_data_703_port, 
      bus_selected_win_data_702_port, bus_selected_win_data_701_port, 
      bus_selected_win_data_700_port, bus_selected_win_data_699_port, 
      bus_selected_win_data_698_port, bus_selected_win_data_697_port, 
      bus_selected_win_data_696_port, bus_selected_win_data_695_port, 
      bus_selected_win_data_694_port, bus_selected_win_data_693_port, 
      bus_selected_win_data_692_port, bus_selected_win_data_691_port, 
      bus_selected_win_data_690_port, bus_selected_win_data_689_port, 
      bus_selected_win_data_688_port, bus_selected_win_data_687_port, 
      bus_selected_win_data_686_port, bus_selected_win_data_685_port, 
      bus_selected_win_data_684_port, bus_selected_win_data_683_port, 
      bus_selected_win_data_682_port, bus_selected_win_data_681_port, 
      bus_selected_win_data_680_port, bus_selected_win_data_679_port, 
      bus_selected_win_data_678_port, bus_selected_win_data_677_port, 
      bus_selected_win_data_676_port, bus_selected_win_data_675_port, 
      bus_selected_win_data_674_port, bus_selected_win_data_673_port, 
      bus_selected_win_data_672_port, bus_selected_win_data_671_port, 
      bus_selected_win_data_670_port, bus_selected_win_data_669_port, 
      bus_selected_win_data_668_port, bus_selected_win_data_667_port, 
      bus_selected_win_data_666_port, bus_selected_win_data_665_port, 
      bus_selected_win_data_664_port, bus_selected_win_data_663_port, 
      bus_selected_win_data_662_port, bus_selected_win_data_661_port, 
      bus_selected_win_data_660_port, bus_selected_win_data_659_port, 
      bus_selected_win_data_658_port, bus_selected_win_data_657_port, 
      bus_selected_win_data_656_port, bus_selected_win_data_655_port, 
      bus_selected_win_data_654_port, bus_selected_win_data_653_port, 
      bus_selected_win_data_652_port, bus_selected_win_data_651_port, 
      bus_selected_win_data_650_port, bus_selected_win_data_649_port, 
      bus_selected_win_data_648_port, bus_selected_win_data_647_port, 
      bus_selected_win_data_646_port, bus_selected_win_data_645_port, 
      bus_selected_win_data_644_port, bus_selected_win_data_643_port, 
      bus_selected_win_data_642_port, bus_selected_win_data_641_port, 
      bus_selected_win_data_640_port, bus_selected_win_data_639_port, 
      bus_selected_win_data_638_port, bus_selected_win_data_637_port, 
      bus_selected_win_data_636_port, bus_selected_win_data_635_port, 
      bus_selected_win_data_634_port, bus_selected_win_data_633_port, 
      bus_selected_win_data_632_port, bus_selected_win_data_631_port, 
      bus_selected_win_data_630_port, bus_selected_win_data_629_port, 
      bus_selected_win_data_628_port, bus_selected_win_data_627_port, 
      bus_selected_win_data_626_port, bus_selected_win_data_625_port, 
      bus_selected_win_data_624_port, bus_selected_win_data_623_port, 
      bus_selected_win_data_622_port, bus_selected_win_data_621_port, 
      bus_selected_win_data_620_port, bus_selected_win_data_619_port, 
      bus_selected_win_data_618_port, bus_selected_win_data_617_port, 
      bus_selected_win_data_616_port, bus_selected_win_data_615_port, 
      bus_selected_win_data_614_port, bus_selected_win_data_613_port, 
      bus_selected_win_data_612_port, bus_selected_win_data_611_port, 
      bus_selected_win_data_610_port, bus_selected_win_data_609_port, 
      bus_selected_win_data_608_port, bus_selected_win_data_607_port, 
      bus_selected_win_data_606_port, bus_selected_win_data_605_port, 
      bus_selected_win_data_604_port, bus_selected_win_data_603_port, 
      bus_selected_win_data_602_port, bus_selected_win_data_601_port, 
      bus_selected_win_data_600_port, bus_selected_win_data_599_port, 
      bus_selected_win_data_598_port, bus_selected_win_data_597_port, 
      bus_selected_win_data_596_port, bus_selected_win_data_595_port, 
      bus_selected_win_data_594_port, bus_selected_win_data_593_port, 
      bus_selected_win_data_592_port, bus_selected_win_data_591_port, 
      bus_selected_win_data_590_port, bus_selected_win_data_589_port, 
      bus_selected_win_data_588_port, bus_selected_win_data_587_port, 
      bus_selected_win_data_586_port, bus_selected_win_data_585_port, 
      bus_selected_win_data_584_port, bus_selected_win_data_583_port, 
      bus_selected_win_data_582_port, bus_selected_win_data_581_port, 
      bus_selected_win_data_580_port, bus_selected_win_data_579_port, 
      bus_selected_win_data_578_port, bus_selected_win_data_577_port, 
      bus_selected_win_data_576_port, bus_selected_win_data_575_port, 
      bus_selected_win_data_574_port, bus_selected_win_data_573_port, 
      bus_selected_win_data_572_port, bus_selected_win_data_571_port, 
      bus_selected_win_data_570_port, bus_selected_win_data_569_port, 
      bus_selected_win_data_568_port, bus_selected_win_data_567_port, 
      bus_selected_win_data_566_port, bus_selected_win_data_565_port, 
      bus_selected_win_data_564_port, bus_selected_win_data_563_port, 
      bus_selected_win_data_562_port, bus_selected_win_data_561_port, 
      bus_selected_win_data_560_port, bus_selected_win_data_559_port, 
      bus_selected_win_data_558_port, bus_selected_win_data_557_port, 
      bus_selected_win_data_556_port, bus_selected_win_data_555_port, 
      bus_selected_win_data_554_port, bus_selected_win_data_553_port, 
      bus_selected_win_data_552_port, bus_selected_win_data_551_port, 
      bus_selected_win_data_550_port, bus_selected_win_data_549_port, 
      bus_selected_win_data_548_port, bus_selected_win_data_547_port, 
      bus_selected_win_data_546_port, bus_selected_win_data_545_port, 
      bus_selected_win_data_544_port, bus_selected_win_data_543_port, 
      bus_selected_win_data_542_port, bus_selected_win_data_541_port, 
      bus_selected_win_data_540_port, bus_selected_win_data_539_port, 
      bus_selected_win_data_538_port, bus_selected_win_data_537_port, 
      bus_selected_win_data_536_port, bus_selected_win_data_535_port, 
      bus_selected_win_data_534_port, bus_selected_win_data_533_port, 
      bus_selected_win_data_532_port, bus_selected_win_data_531_port, 
      bus_selected_win_data_530_port, bus_selected_win_data_529_port, 
      bus_selected_win_data_528_port, bus_selected_win_data_527_port, 
      bus_selected_win_data_526_port, bus_selected_win_data_525_port, 
      bus_selected_win_data_524_port, bus_selected_win_data_523_port, 
      bus_selected_win_data_522_port, bus_selected_win_data_521_port, 
      bus_selected_win_data_520_port, bus_selected_win_data_519_port, 
      bus_selected_win_data_518_port, bus_selected_win_data_517_port, 
      bus_selected_win_data_516_port, bus_selected_win_data_515_port, 
      bus_selected_win_data_514_port, bus_selected_win_data_513_port, 
      bus_selected_win_data_512_port, bus_selected_win_data_511_port, 
      bus_selected_win_data_510_port, bus_selected_win_data_509_port, 
      bus_selected_win_data_508_port, bus_selected_win_data_507_port, 
      bus_selected_win_data_506_port, bus_selected_win_data_505_port, 
      bus_selected_win_data_504_port, bus_selected_win_data_503_port, 
      bus_selected_win_data_502_port, bus_selected_win_data_501_port, 
      bus_selected_win_data_500_port, bus_selected_win_data_499_port, 
      bus_selected_win_data_498_port, bus_selected_win_data_497_port, 
      bus_selected_win_data_496_port, bus_selected_win_data_495_port, 
      bus_selected_win_data_494_port, bus_selected_win_data_493_port, 
      bus_selected_win_data_492_port, bus_selected_win_data_491_port, 
      bus_selected_win_data_490_port, bus_selected_win_data_489_port, 
      bus_selected_win_data_488_port, bus_selected_win_data_487_port, 
      bus_selected_win_data_486_port, bus_selected_win_data_485_port, 
      bus_selected_win_data_484_port, bus_selected_win_data_483_port, 
      bus_selected_win_data_482_port, bus_selected_win_data_481_port, 
      bus_selected_win_data_480_port, bus_selected_win_data_479_port, 
      bus_selected_win_data_478_port, bus_selected_win_data_477_port, 
      bus_selected_win_data_476_port, bus_selected_win_data_475_port, 
      bus_selected_win_data_474_port, bus_selected_win_data_473_port, 
      bus_selected_win_data_472_port, bus_selected_win_data_471_port, 
      bus_selected_win_data_470_port, bus_selected_win_data_469_port, 
      bus_selected_win_data_468_port, bus_selected_win_data_467_port, 
      bus_selected_win_data_466_port, bus_selected_win_data_465_port, 
      bus_selected_win_data_464_port, bus_selected_win_data_463_port, 
      bus_selected_win_data_462_port, bus_selected_win_data_461_port, 
      bus_selected_win_data_460_port, bus_selected_win_data_459_port, 
      bus_selected_win_data_458_port, bus_selected_win_data_457_port, 
      bus_selected_win_data_456_port, bus_selected_win_data_455_port, 
      bus_selected_win_data_454_port, bus_selected_win_data_453_port, 
      bus_selected_win_data_452_port, bus_selected_win_data_451_port, 
      bus_selected_win_data_450_port, bus_selected_win_data_449_port, 
      bus_selected_win_data_448_port, bus_selected_win_data_447_port, 
      bus_selected_win_data_446_port, bus_selected_win_data_445_port, 
      bus_selected_win_data_444_port, bus_selected_win_data_443_port, 
      bus_selected_win_data_442_port, bus_selected_win_data_441_port, 
      bus_selected_win_data_440_port, bus_selected_win_data_439_port, 
      bus_selected_win_data_438_port, bus_selected_win_data_437_port, 
      bus_selected_win_data_436_port, bus_selected_win_data_435_port, 
      bus_selected_win_data_434_port, bus_selected_win_data_433_port, 
      bus_selected_win_data_432_port, bus_selected_win_data_431_port, 
      bus_selected_win_data_430_port, bus_selected_win_data_429_port, 
      bus_selected_win_data_428_port, bus_selected_win_data_427_port, 
      bus_selected_win_data_426_port, bus_selected_win_data_425_port, 
      bus_selected_win_data_424_port, bus_selected_win_data_423_port, 
      bus_selected_win_data_422_port, bus_selected_win_data_421_port, 
      bus_selected_win_data_420_port, bus_selected_win_data_419_port, 
      bus_selected_win_data_418_port, bus_selected_win_data_417_port, 
      bus_selected_win_data_416_port, bus_selected_win_data_415_port, 
      bus_selected_win_data_414_port, bus_selected_win_data_413_port, 
      bus_selected_win_data_412_port, bus_selected_win_data_411_port, 
      bus_selected_win_data_410_port, bus_selected_win_data_409_port, 
      bus_selected_win_data_408_port, bus_selected_win_data_407_port, 
      bus_selected_win_data_406_port, bus_selected_win_data_405_port, 
      bus_selected_win_data_404_port, bus_selected_win_data_403_port, 
      bus_selected_win_data_402_port, bus_selected_win_data_401_port, 
      bus_selected_win_data_400_port, bus_selected_win_data_399_port, 
      bus_selected_win_data_398_port, bus_selected_win_data_397_port, 
      bus_selected_win_data_396_port, bus_selected_win_data_395_port, 
      bus_selected_win_data_394_port, bus_selected_win_data_393_port, 
      bus_selected_win_data_392_port, bus_selected_win_data_391_port, 
      bus_selected_win_data_390_port, bus_selected_win_data_389_port, 
      bus_selected_win_data_388_port, bus_selected_win_data_387_port, 
      bus_selected_win_data_386_port, bus_selected_win_data_385_port, 
      bus_selected_win_data_384_port, bus_selected_win_data_383_port, 
      bus_selected_win_data_382_port, bus_selected_win_data_381_port, 
      bus_selected_win_data_380_port, bus_selected_win_data_379_port, 
      bus_selected_win_data_378_port, bus_selected_win_data_377_port, 
      bus_selected_win_data_376_port, bus_selected_win_data_375_port, 
      bus_selected_win_data_374_port, bus_selected_win_data_373_port, 
      bus_selected_win_data_372_port, bus_selected_win_data_371_port, 
      bus_selected_win_data_370_port, bus_selected_win_data_369_port, 
      bus_selected_win_data_368_port, bus_selected_win_data_367_port, 
      bus_selected_win_data_366_port, bus_selected_win_data_365_port, 
      bus_selected_win_data_364_port, bus_selected_win_data_363_port, 
      bus_selected_win_data_362_port, bus_selected_win_data_361_port, 
      bus_selected_win_data_360_port, bus_selected_win_data_359_port, 
      bus_selected_win_data_358_port, bus_selected_win_data_357_port, 
      bus_selected_win_data_356_port, bus_selected_win_data_355_port, 
      bus_selected_win_data_354_port, bus_selected_win_data_353_port, 
      bus_selected_win_data_352_port, bus_selected_win_data_351_port, 
      bus_selected_win_data_350_port, bus_selected_win_data_349_port, 
      bus_selected_win_data_348_port, bus_selected_win_data_347_port, 
      bus_selected_win_data_346_port, bus_selected_win_data_345_port, 
      bus_selected_win_data_344_port, bus_selected_win_data_343_port, 
      bus_selected_win_data_342_port, bus_selected_win_data_341_port, 
      bus_selected_win_data_340_port, bus_selected_win_data_339_port, 
      bus_selected_win_data_338_port, bus_selected_win_data_337_port, 
      bus_selected_win_data_336_port, bus_selected_win_data_335_port, 
      bus_selected_win_data_334_port, bus_selected_win_data_333_port, 
      bus_selected_win_data_332_port, bus_selected_win_data_331_port, 
      bus_selected_win_data_330_port, bus_selected_win_data_329_port, 
      bus_selected_win_data_328_port, bus_selected_win_data_327_port, 
      bus_selected_win_data_326_port, bus_selected_win_data_325_port, 
      bus_selected_win_data_324_port, bus_selected_win_data_323_port, 
      bus_selected_win_data_322_port, bus_selected_win_data_321_port, 
      bus_selected_win_data_320_port, bus_selected_win_data_319_port, 
      bus_selected_win_data_318_port, bus_selected_win_data_317_port, 
      bus_selected_win_data_316_port, bus_selected_win_data_315_port, 
      bus_selected_win_data_314_port, bus_selected_win_data_313_port, 
      bus_selected_win_data_312_port, bus_selected_win_data_311_port, 
      bus_selected_win_data_310_port, bus_selected_win_data_309_port, 
      bus_selected_win_data_308_port, bus_selected_win_data_307_port, 
      bus_selected_win_data_306_port, bus_selected_win_data_305_port, 
      bus_selected_win_data_304_port, bus_selected_win_data_303_port, 
      bus_selected_win_data_302_port, bus_selected_win_data_301_port, 
      bus_selected_win_data_300_port, bus_selected_win_data_299_port, 
      bus_selected_win_data_298_port, bus_selected_win_data_297_port, 
      bus_selected_win_data_296_port, bus_selected_win_data_295_port, 
      bus_selected_win_data_294_port, bus_selected_win_data_293_port, 
      bus_selected_win_data_292_port, bus_selected_win_data_291_port, 
      bus_selected_win_data_290_port, bus_selected_win_data_289_port, 
      bus_selected_win_data_288_port, bus_selected_win_data_287_port, 
      bus_selected_win_data_286_port, bus_selected_win_data_285_port, 
      bus_selected_win_data_284_port, bus_selected_win_data_283_port, 
      bus_selected_win_data_282_port, bus_selected_win_data_281_port, 
      bus_selected_win_data_280_port, bus_selected_win_data_279_port, 
      bus_selected_win_data_278_port, bus_selected_win_data_277_port, 
      bus_selected_win_data_276_port, bus_selected_win_data_275_port, 
      bus_selected_win_data_274_port, bus_selected_win_data_273_port, 
      bus_selected_win_data_272_port, bus_selected_win_data_271_port, 
      bus_selected_win_data_270_port, bus_selected_win_data_269_port, 
      bus_selected_win_data_268_port, bus_selected_win_data_267_port, 
      bus_selected_win_data_266_port, bus_selected_win_data_265_port, 
      bus_selected_win_data_264_port, bus_selected_win_data_263_port, 
      bus_selected_win_data_262_port, bus_selected_win_data_261_port, 
      bus_selected_win_data_260_port, bus_selected_win_data_259_port, 
      bus_selected_win_data_258_port, bus_selected_win_data_257_port, 
      bus_selected_win_data_256_port, bus_selected_win_data_255_port, 
      bus_selected_win_data_254_port, bus_selected_win_data_253_port, 
      bus_selected_win_data_252_port, bus_selected_win_data_251_port, 
      bus_selected_win_data_250_port, bus_selected_win_data_249_port, 
      bus_selected_win_data_248_port, bus_selected_win_data_247_port, 
      bus_selected_win_data_246_port, bus_selected_win_data_245_port, 
      bus_selected_win_data_244_port, bus_selected_win_data_243_port, 
      bus_selected_win_data_242_port, bus_selected_win_data_241_port, 
      bus_selected_win_data_240_port, bus_selected_win_data_239_port, 
      bus_selected_win_data_238_port, bus_selected_win_data_237_port, 
      bus_selected_win_data_236_port, bus_selected_win_data_235_port, 
      bus_selected_win_data_234_port, bus_selected_win_data_233_port, 
      bus_selected_win_data_232_port, bus_selected_win_data_231_port, 
      bus_selected_win_data_230_port, bus_selected_win_data_229_port, 
      bus_selected_win_data_228_port, bus_selected_win_data_227_port, 
      bus_selected_win_data_226_port, bus_selected_win_data_225_port, 
      bus_selected_win_data_224_port, bus_selected_win_data_223_port, 
      bus_selected_win_data_222_port, bus_selected_win_data_221_port, 
      bus_selected_win_data_220_port, bus_selected_win_data_219_port, 
      bus_selected_win_data_218_port, bus_selected_win_data_217_port, 
      bus_selected_win_data_216_port, bus_selected_win_data_215_port, 
      bus_selected_win_data_214_port, bus_selected_win_data_213_port, 
      bus_selected_win_data_212_port, bus_selected_win_data_211_port, 
      bus_selected_win_data_210_port, bus_selected_win_data_209_port, 
      bus_selected_win_data_208_port, bus_selected_win_data_207_port, 
      bus_selected_win_data_206_port, bus_selected_win_data_205_port, 
      bus_selected_win_data_204_port, bus_selected_win_data_203_port, 
      bus_selected_win_data_202_port, bus_selected_win_data_201_port, 
      bus_selected_win_data_200_port, bus_selected_win_data_199_port, 
      bus_selected_win_data_198_port, bus_selected_win_data_197_port, 
      bus_selected_win_data_196_port, bus_selected_win_data_195_port, 
      bus_selected_win_data_194_port, bus_selected_win_data_193_port, 
      bus_selected_win_data_192_port, bus_selected_win_data_191_port, 
      bus_selected_win_data_190_port, bus_selected_win_data_189_port, 
      bus_selected_win_data_188_port, bus_selected_win_data_187_port, 
      bus_selected_win_data_186_port, bus_selected_win_data_185_port, 
      bus_selected_win_data_184_port, bus_selected_win_data_183_port, 
      bus_selected_win_data_182_port, bus_selected_win_data_181_port, 
      bus_selected_win_data_180_port, bus_selected_win_data_179_port, 
      bus_selected_win_data_178_port, bus_selected_win_data_177_port, 
      bus_selected_win_data_176_port, bus_selected_win_data_175_port, 
      bus_selected_win_data_174_port, bus_selected_win_data_173_port, 
      bus_selected_win_data_172_port, bus_selected_win_data_171_port, 
      bus_selected_win_data_170_port, bus_selected_win_data_169_port, 
      bus_selected_win_data_168_port, bus_selected_win_data_167_port, 
      bus_selected_win_data_166_port, bus_selected_win_data_165_port, 
      bus_selected_win_data_164_port, bus_selected_win_data_163_port, 
      bus_selected_win_data_162_port, bus_selected_win_data_161_port, 
      bus_selected_win_data_160_port, bus_selected_win_data_159_port, 
      bus_selected_win_data_158_port, bus_selected_win_data_157_port, 
      bus_selected_win_data_156_port, bus_selected_win_data_155_port, 
      bus_selected_win_data_154_port, bus_selected_win_data_153_port, 
      bus_selected_win_data_152_port, bus_selected_win_data_151_port, 
      bus_selected_win_data_150_port, bus_selected_win_data_149_port, 
      bus_selected_win_data_148_port, bus_selected_win_data_147_port, 
      bus_selected_win_data_146_port, bus_selected_win_data_145_port, 
      bus_selected_win_data_144_port, bus_selected_win_data_143_port, 
      bus_selected_win_data_142_port, bus_selected_win_data_141_port, 
      bus_selected_win_data_140_port, bus_selected_win_data_139_port, 
      bus_selected_win_data_138_port, bus_selected_win_data_137_port, 
      bus_selected_win_data_136_port, bus_selected_win_data_135_port, 
      bus_selected_win_data_134_port, bus_selected_win_data_133_port, 
      bus_selected_win_data_132_port, bus_selected_win_data_131_port, 
      bus_selected_win_data_130_port, bus_selected_win_data_129_port, 
      bus_selected_win_data_128_port, bus_selected_win_data_127_port, 
      bus_selected_win_data_126_port, bus_selected_win_data_125_port, 
      bus_selected_win_data_124_port, bus_selected_win_data_123_port, 
      bus_selected_win_data_122_port, bus_selected_win_data_121_port, 
      bus_selected_win_data_120_port, bus_selected_win_data_119_port, 
      bus_selected_win_data_118_port, bus_selected_win_data_117_port, 
      bus_selected_win_data_116_port, bus_selected_win_data_115_port, 
      bus_selected_win_data_114_port, bus_selected_win_data_113_port, 
      bus_selected_win_data_112_port, bus_selected_win_data_111_port, 
      bus_selected_win_data_110_port, bus_selected_win_data_109_port, 
      bus_selected_win_data_108_port, bus_selected_win_data_107_port, 
      bus_selected_win_data_106_port, bus_selected_win_data_105_port, 
      bus_selected_win_data_104_port, bus_selected_win_data_103_port, 
      bus_selected_win_data_102_port, bus_selected_win_data_101_port, 
      bus_selected_win_data_100_port, bus_selected_win_data_99_port, 
      bus_selected_win_data_98_port, bus_selected_win_data_97_port, 
      bus_selected_win_data_96_port, bus_selected_win_data_95_port, 
      bus_selected_win_data_94_port, bus_selected_win_data_93_port, 
      bus_selected_win_data_92_port, bus_selected_win_data_91_port, 
      bus_selected_win_data_90_port, bus_selected_win_data_89_port, 
      bus_selected_win_data_88_port, bus_selected_win_data_87_port, 
      bus_selected_win_data_86_port, bus_selected_win_data_85_port, 
      bus_selected_win_data_84_port, bus_selected_win_data_83_port, 
      bus_selected_win_data_82_port, bus_selected_win_data_81_port, 
      bus_selected_win_data_80_port, bus_selected_win_data_79_port, 
      bus_selected_win_data_78_port, bus_selected_win_data_77_port, 
      bus_selected_win_data_76_port, bus_selected_win_data_75_port, 
      bus_selected_win_data_74_port, bus_selected_win_data_73_port, 
      bus_selected_win_data_72_port, bus_selected_win_data_71_port, 
      bus_selected_win_data_70_port, bus_selected_win_data_69_port, 
      bus_selected_win_data_68_port, bus_selected_win_data_67_port, 
      bus_selected_win_data_66_port, bus_selected_win_data_65_port, 
      bus_selected_win_data_64_port, bus_selected_win_data_63_port, 
      bus_selected_win_data_62_port, bus_selected_win_data_61_port, 
      bus_selected_win_data_60_port, bus_selected_win_data_59_port, 
      bus_selected_win_data_58_port, bus_selected_win_data_57_port, 
      bus_selected_win_data_56_port, bus_selected_win_data_55_port, 
      bus_selected_win_data_54_port, bus_selected_win_data_53_port, 
      bus_selected_win_data_52_port, bus_selected_win_data_51_port, 
      bus_selected_win_data_50_port, bus_selected_win_data_49_port, 
      bus_selected_win_data_48_port, bus_selected_win_data_47_port, 
      bus_selected_win_data_46_port, bus_selected_win_data_45_port, 
      bus_selected_win_data_44_port, bus_selected_win_data_43_port, 
      bus_selected_win_data_42_port, bus_selected_win_data_41_port, 
      bus_selected_win_data_40_port, bus_selected_win_data_39_port, 
      bus_selected_win_data_38_port, bus_selected_win_data_37_port, 
      bus_selected_win_data_36_port, bus_selected_win_data_35_port, 
      bus_selected_win_data_34_port, bus_selected_win_data_33_port, 
      bus_selected_win_data_32_port, bus_selected_win_data_31_port, 
      bus_selected_win_data_30_port, bus_selected_win_data_29_port, 
      bus_selected_win_data_28_port, bus_selected_win_data_27_port, 
      bus_selected_win_data_26_port, bus_selected_win_data_25_port, 
      bus_selected_win_data_24_port, bus_selected_win_data_23_port, 
      bus_selected_win_data_22_port, bus_selected_win_data_21_port, 
      bus_selected_win_data_20_port, bus_selected_win_data_19_port, 
      bus_selected_win_data_18_port, bus_selected_win_data_17_port, 
      bus_selected_win_data_16_port, bus_selected_win_data_15_port, 
      bus_selected_win_data_14_port, bus_selected_win_data_13_port, 
      bus_selected_win_data_12_port, bus_selected_win_data_11_port, 
      bus_selected_win_data_10_port, bus_selected_win_data_9_port, 
      bus_selected_win_data_8_port, bus_selected_win_data_7_port, 
      bus_selected_win_data_6_port, bus_selected_win_data_5_port, 
      bus_selected_win_data_4_port, bus_selected_win_data_3_port, 
      bus_selected_win_data_2_port, bus_selected_win_data_1_port, 
      bus_selected_win_data_0_port, bus_complete_win_data_255_port, 
      bus_complete_win_data_254_port, bus_complete_win_data_253_port, 
      bus_complete_win_data_252_port, bus_complete_win_data_251_port, 
      bus_complete_win_data_250_port, bus_complete_win_data_249_port, 
      bus_complete_win_data_248_port, bus_complete_win_data_247_port, 
      bus_complete_win_data_246_port, bus_complete_win_data_245_port, 
      bus_complete_win_data_244_port, bus_complete_win_data_243_port, 
      bus_complete_win_data_242_port, bus_complete_win_data_241_port, 
      bus_complete_win_data_240_port, bus_complete_win_data_239_port, 
      bus_complete_win_data_238_port, bus_complete_win_data_237_port, 
      bus_complete_win_data_236_port, bus_complete_win_data_235_port, 
      bus_complete_win_data_234_port, bus_complete_win_data_233_port, 
      bus_complete_win_data_232_port, bus_complete_win_data_231_port, 
      bus_complete_win_data_230_port, bus_complete_win_data_229_port, 
      bus_complete_win_data_228_port, bus_complete_win_data_227_port, 
      bus_complete_win_data_226_port, bus_complete_win_data_225_port, 
      bus_complete_win_data_224_port, bus_complete_win_data_223_port, 
      bus_complete_win_data_222_port, bus_complete_win_data_221_port, 
      bus_complete_win_data_220_port, bus_complete_win_data_219_port, 
      bus_complete_win_data_218_port, bus_complete_win_data_217_port, 
      bus_complete_win_data_216_port, bus_complete_win_data_215_port, 
      bus_complete_win_data_214_port, bus_complete_win_data_213_port, 
      bus_complete_win_data_212_port, bus_complete_win_data_211_port, 
      bus_complete_win_data_210_port, bus_complete_win_data_209_port, 
      bus_complete_win_data_208_port, bus_complete_win_data_207_port, 
      bus_complete_win_data_206_port, bus_complete_win_data_205_port, 
      bus_complete_win_data_204_port, bus_complete_win_data_203_port, 
      bus_complete_win_data_202_port, bus_complete_win_data_201_port, 
      bus_complete_win_data_200_port, bus_complete_win_data_199_port, 
      bus_complete_win_data_198_port, bus_complete_win_data_197_port, 
      bus_complete_win_data_196_port, bus_complete_win_data_195_port, 
      bus_complete_win_data_194_port, bus_complete_win_data_193_port, 
      bus_complete_win_data_192_port, bus_complete_win_data_191_port, 
      bus_complete_win_data_190_port, bus_complete_win_data_189_port, 
      bus_complete_win_data_188_port, bus_complete_win_data_187_port, 
      bus_complete_win_data_186_port, bus_complete_win_data_185_port, 
      bus_complete_win_data_184_port, bus_complete_win_data_183_port, 
      bus_complete_win_data_182_port, bus_complete_win_data_181_port, 
      bus_complete_win_data_180_port, bus_complete_win_data_179_port, 
      bus_complete_win_data_178_port, bus_complete_win_data_177_port, 
      bus_complete_win_data_176_port, bus_complete_win_data_175_port, 
      bus_complete_win_data_174_port, bus_complete_win_data_173_port, 
      bus_complete_win_data_172_port, bus_complete_win_data_171_port, 
      bus_complete_win_data_170_port, bus_complete_win_data_169_port, 
      bus_complete_win_data_168_port, bus_complete_win_data_167_port, 
      bus_complete_win_data_166_port, bus_complete_win_data_165_port, 
      bus_complete_win_data_164_port, bus_complete_win_data_163_port, 
      bus_complete_win_data_162_port, bus_complete_win_data_161_port, 
      bus_complete_win_data_160_port, bus_complete_win_data_159_port, 
      bus_complete_win_data_158_port, bus_complete_win_data_157_port, 
      bus_complete_win_data_156_port, bus_complete_win_data_155_port, 
      bus_complete_win_data_154_port, bus_complete_win_data_153_port, 
      bus_complete_win_data_152_port, bus_complete_win_data_151_port, 
      bus_complete_win_data_150_port, bus_complete_win_data_149_port, 
      bus_complete_win_data_148_port, bus_complete_win_data_147_port, 
      bus_complete_win_data_146_port, bus_complete_win_data_145_port, 
      bus_complete_win_data_144_port, bus_complete_win_data_143_port, 
      bus_complete_win_data_142_port, bus_complete_win_data_141_port, 
      bus_complete_win_data_140_port, bus_complete_win_data_139_port, 
      bus_complete_win_data_138_port, bus_complete_win_data_137_port, 
      bus_complete_win_data_136_port, bus_complete_win_data_135_port, 
      bus_complete_win_data_134_port, bus_complete_win_data_133_port, 
      bus_complete_win_data_132_port, bus_complete_win_data_131_port, 
      bus_complete_win_data_130_port, bus_complete_win_data_129_port, 
      bus_complete_win_data_128_port, bus_complete_win_data_127_port, 
      bus_complete_win_data_126_port, bus_complete_win_data_125_port, 
      bus_complete_win_data_124_port, bus_complete_win_data_123_port, 
      bus_complete_win_data_122_port, bus_complete_win_data_121_port, 
      bus_complete_win_data_120_port, bus_complete_win_data_119_port, 
      bus_complete_win_data_118_port, bus_complete_win_data_117_port, 
      bus_complete_win_data_116_port, bus_complete_win_data_115_port, 
      bus_complete_win_data_114_port, bus_complete_win_data_113_port, 
      bus_complete_win_data_112_port, bus_complete_win_data_111_port, 
      bus_complete_win_data_110_port, bus_complete_win_data_109_port, 
      bus_complete_win_data_108_port, bus_complete_win_data_107_port, 
      bus_complete_win_data_106_port, bus_complete_win_data_105_port, 
      bus_complete_win_data_104_port, bus_complete_win_data_103_port, 
      bus_complete_win_data_102_port, bus_complete_win_data_101_port, 
      bus_complete_win_data_100_port, bus_complete_win_data_99_port, 
      bus_complete_win_data_98_port, bus_complete_win_data_97_port, 
      bus_complete_win_data_96_port, bus_complete_win_data_95_port, 
      bus_complete_win_data_94_port, bus_complete_win_data_93_port, 
      bus_complete_win_data_92_port, bus_complete_win_data_91_port, 
      bus_complete_win_data_90_port, bus_complete_win_data_89_port, 
      bus_complete_win_data_88_port, bus_complete_win_data_87_port, 
      bus_complete_win_data_86_port, bus_complete_win_data_85_port, 
      bus_complete_win_data_84_port, bus_complete_win_data_83_port, 
      bus_complete_win_data_82_port, bus_complete_win_data_81_port, 
      bus_complete_win_data_80_port, bus_complete_win_data_79_port, 
      bus_complete_win_data_78_port, bus_complete_win_data_77_port, 
      bus_complete_win_data_76_port, bus_complete_win_data_75_port, 
      bus_complete_win_data_74_port, bus_complete_win_data_73_port, 
      bus_complete_win_data_72_port, bus_complete_win_data_71_port, 
      bus_complete_win_data_70_port, bus_complete_win_data_69_port, 
      bus_complete_win_data_68_port, bus_complete_win_data_67_port, 
      bus_complete_win_data_66_port, bus_complete_win_data_65_port, 
      bus_complete_win_data_64_port, bus_complete_win_data_63_port, 
      bus_complete_win_data_62_port, bus_complete_win_data_61_port, 
      bus_complete_win_data_60_port, bus_complete_win_data_59_port, 
      bus_complete_win_data_58_port, bus_complete_win_data_57_port, 
      bus_complete_win_data_56_port, bus_complete_win_data_55_port, 
      bus_complete_win_data_54_port, bus_complete_win_data_53_port, 
      bus_complete_win_data_52_port, bus_complete_win_data_51_port, 
      bus_complete_win_data_50_port, bus_complete_win_data_49_port, 
      bus_complete_win_data_48_port, bus_complete_win_data_47_port, 
      bus_complete_win_data_46_port, bus_complete_win_data_45_port, 
      bus_complete_win_data_44_port, bus_complete_win_data_43_port, 
      bus_complete_win_data_42_port, bus_complete_win_data_41_port, 
      bus_complete_win_data_40_port, bus_complete_win_data_39_port, 
      bus_complete_win_data_38_port, bus_complete_win_data_37_port, 
      bus_complete_win_data_36_port, bus_complete_win_data_35_port, 
      bus_complete_win_data_34_port, bus_complete_win_data_33_port, 
      bus_complete_win_data_32_port, bus_complete_win_data_31_port, 
      bus_complete_win_data_30_port, bus_complete_win_data_29_port, 
      bus_complete_win_data_28_port, bus_complete_win_data_27_port, 
      bus_complete_win_data_26_port, bus_complete_win_data_25_port, 
      bus_complete_win_data_24_port, bus_complete_win_data_23_port, 
      bus_complete_win_data_22_port, bus_complete_win_data_21_port, 
      bus_complete_win_data_20_port, bus_complete_win_data_19_port, 
      bus_complete_win_data_18_port, bus_complete_win_data_17_port, 
      bus_complete_win_data_16_port, bus_complete_win_data_15_port, 
      bus_complete_win_data_14_port, bus_complete_win_data_13_port, 
      bus_complete_win_data_12_port, bus_complete_win_data_11_port, 
      bus_complete_win_data_10_port, bus_complete_win_data_9_port, 
      bus_complete_win_data_8_port, bus_complete_win_data_7_port, 
      bus_complete_win_data_6_port, bus_complete_win_data_5_port, 
      bus_complete_win_data_4_port, bus_complete_win_data_3_port, 
      bus_complete_win_data_2_port, bus_complete_win_data_1_port, 
      bus_complete_win_data_0_port, internal_out1_31_port, 
      internal_out1_30_port, internal_out1_29_port, internal_out1_28_port, 
      internal_out1_27_port, internal_out1_26_port, internal_out1_25_port, 
      internal_out1_24_port, internal_out1_23_port, internal_out1_22_port, 
      internal_out1_21_port, internal_out1_20_port, internal_out1_19_port, 
      internal_out1_18_port, internal_out1_17_port, internal_out1_16_port, 
      internal_out1_15_port, internal_out1_14_port, internal_out1_13_port, 
      internal_out1_12_port, internal_out1_11_port, internal_out1_10_port, 
      internal_out1_9_port, internal_out1_8_port, internal_out1_7_port, 
      internal_out1_6_port, internal_out1_5_port, internal_out1_4_port, 
      internal_out1_3_port, internal_out1_2_port, internal_out1_1_port, 
      internal_out1_0_port, internal_out2_31_port, internal_out2_30_port, 
      internal_out2_29_port, internal_out2_28_port, internal_out2_27_port, 
      internal_out2_26_port, internal_out2_25_port, internal_out2_24_port, 
      internal_out2_23_port, internal_out2_22_port, internal_out2_21_port, 
      internal_out2_20_port, internal_out2_19_port, internal_out2_18_port, 
      internal_out2_17_port, internal_out2_16_port, internal_out2_15_port, 
      internal_out2_14_port, internal_out2_13_port, internal_out2_12_port, 
      internal_out2_11_port, internal_out2_10_port, internal_out2_9_port, 
      internal_out2_8_port, internal_out2_7_port, internal_out2_6_port, 
      internal_out2_5_port, internal_out2_4_port, internal_out2_3_port, 
      internal_out2_2_port, internal_out2_1_port, internal_out2_0_port, 
      en_regi_87_port, en_regi_86_port, en_regi_85_port, en_regi_84_port, 
      en_regi_83_port, en_regi_82_port, en_regi_81_port, en_regi_80_port, 
      en_regi_79_port, en_regi_78_port, en_regi_77_port, en_regi_76_port, 
      en_regi_75_port, en_regi_74_port, en_regi_73_port, en_regi_72_port, 
      en_regi_71_port, en_regi_70_port, en_regi_69_port, en_regi_68_port, 
      en_regi_67_port, en_regi_66_port, en_regi_65_port, en_regi_64_port, 
      en_regi_63_port, en_regi_62_port, en_regi_61_port, en_regi_60_port, 
      en_regi_59_port, en_regi_58_port, en_regi_57_port, en_regi_56_port, 
      en_regi_55_port, en_regi_54_port, en_regi_53_port, en_regi_52_port, 
      en_regi_51_port, en_regi_50_port, en_regi_49_port, en_regi_48_port, 
      en_regi_47_port, en_regi_46_port, en_regi_45_port, en_regi_44_port, 
      en_regi_43_port, en_regi_42_port, en_regi_41_port, en_regi_40_port, 
      en_regi_39_port, en_regi_38_port, en_regi_37_port, en_regi_36_port, 
      en_regi_35_port, en_regi_34_port, en_regi_33_port, en_regi_32_port, 
      en_regi_31_port, en_regi_30_port, en_regi_29_port, en_regi_28_port, 
      en_regi_27_port, en_regi_26_port, en_regi_25_port, en_regi_24_port, 
      en_regi_23_port, en_regi_22_port, en_regi_21_port, en_regi_20_port, 
      en_regi_19_port, en_regi_18_port, en_regi_17_port, en_regi_16_port, 
      en_regi_15_port, en_regi_14_port, en_regi_13_port, en_regi_12_port, 
      en_regi_11_port, en_regi_10_port, en_regi_9_port, en_regi_8_port, 
      en_regi_7_port, en_regi_6_port, en_regi_5_port, en_regi_4_port, 
      en_regi_3_port, en_regi_2_port, en_regi_1_port, en_regi_0_port, 
      c_swin_masked_1bit_0_0_port, c_swin_masked_1bit_1_0_port, 
      c_swin_masked_1bit_2_0_port, c_swin_masked_1bit_3_0_port, 
      c_swin_masked_1bit_4_0_port, internal_inloc_data_0_31_port, 
      internal_inloc_data_0_30_port, internal_inloc_data_0_29_port, 
      internal_inloc_data_0_28_port, internal_inloc_data_0_27_port, 
      internal_inloc_data_0_26_port, internal_inloc_data_0_25_port, 
      internal_inloc_data_0_24_port, internal_inloc_data_0_23_port, 
      internal_inloc_data_0_22_port, internal_inloc_data_0_21_port, 
      internal_inloc_data_0_20_port, internal_inloc_data_0_19_port, 
      internal_inloc_data_0_18_port, internal_inloc_data_0_17_port, 
      internal_inloc_data_0_16_port, internal_inloc_data_0_15_port, 
      internal_inloc_data_0_14_port, internal_inloc_data_0_13_port, 
      internal_inloc_data_0_12_port, internal_inloc_data_0_11_port, 
      internal_inloc_data_0_10_port, internal_inloc_data_0_9_port, 
      internal_inloc_data_0_8_port, internal_inloc_data_0_7_port, 
      internal_inloc_data_0_6_port, internal_inloc_data_0_5_port, 
      internal_inloc_data_0_4_port, internal_inloc_data_0_3_port, 
      internal_inloc_data_0_2_port, internal_inloc_data_0_1_port, 
      internal_inloc_data_0_0_port, internal_inloc_data_1_31_port, 
      internal_inloc_data_1_30_port, internal_inloc_data_1_29_port, 
      internal_inloc_data_1_28_port, internal_inloc_data_1_27_port, 
      internal_inloc_data_1_26_port, internal_inloc_data_1_25_port, 
      internal_inloc_data_1_24_port, internal_inloc_data_1_23_port, 
      internal_inloc_data_1_22_port, internal_inloc_data_1_21_port, 
      internal_inloc_data_1_20_port, internal_inloc_data_1_19_port, 
      internal_inloc_data_1_18_port, internal_inloc_data_1_17_port, 
      internal_inloc_data_1_16_port, internal_inloc_data_1_15_port, 
      internal_inloc_data_1_14_port, internal_inloc_data_1_13_port, 
      internal_inloc_data_1_12_port, internal_inloc_data_1_11_port, 
      internal_inloc_data_1_10_port, internal_inloc_data_1_9_port, 
      internal_inloc_data_1_8_port, internal_inloc_data_1_7_port, 
      internal_inloc_data_1_6_port, internal_inloc_data_1_5_port, 
      internal_inloc_data_1_4_port, internal_inloc_data_1_3_port, 
      internal_inloc_data_1_2_port, internal_inloc_data_1_1_port, 
      internal_inloc_data_1_0_port, internal_inloc_data_2_31_port, 
      internal_inloc_data_2_30_port, internal_inloc_data_2_29_port, 
      internal_inloc_data_2_28_port, internal_inloc_data_2_27_port, 
      internal_inloc_data_2_26_port, internal_inloc_data_2_25_port, 
      internal_inloc_data_2_24_port, internal_inloc_data_2_23_port, 
      internal_inloc_data_2_22_port, internal_inloc_data_2_21_port, 
      internal_inloc_data_2_20_port, internal_inloc_data_2_19_port, 
      internal_inloc_data_2_18_port, internal_inloc_data_2_17_port, 
      internal_inloc_data_2_16_port, internal_inloc_data_2_15_port, 
      internal_inloc_data_2_14_port, internal_inloc_data_2_13_port, 
      internal_inloc_data_2_12_port, internal_inloc_data_2_11_port, 
      internal_inloc_data_2_10_port, internal_inloc_data_2_9_port, 
      internal_inloc_data_2_8_port, internal_inloc_data_2_7_port, 
      internal_inloc_data_2_6_port, internal_inloc_data_2_5_port, 
      internal_inloc_data_2_4_port, internal_inloc_data_2_3_port, 
      internal_inloc_data_2_2_port, internal_inloc_data_2_1_port, 
      internal_inloc_data_2_0_port, internal_inloc_data_3_31_port, 
      internal_inloc_data_3_30_port, internal_inloc_data_3_29_port, 
      internal_inloc_data_3_28_port, internal_inloc_data_3_27_port, 
      internal_inloc_data_3_26_port, internal_inloc_data_3_25_port, 
      internal_inloc_data_3_24_port, internal_inloc_data_3_23_port, 
      internal_inloc_data_3_22_port, internal_inloc_data_3_21_port, 
      internal_inloc_data_3_20_port, internal_inloc_data_3_19_port, 
      internal_inloc_data_3_18_port, internal_inloc_data_3_17_port, 
      internal_inloc_data_3_16_port, internal_inloc_data_3_15_port, 
      internal_inloc_data_3_14_port, internal_inloc_data_3_13_port, 
      internal_inloc_data_3_12_port, internal_inloc_data_3_11_port, 
      internal_inloc_data_3_10_port, internal_inloc_data_3_9_port, 
      internal_inloc_data_3_8_port, internal_inloc_data_3_7_port, 
      internal_inloc_data_3_6_port, internal_inloc_data_3_5_port, 
      internal_inloc_data_3_4_port, internal_inloc_data_3_3_port, 
      internal_inloc_data_3_2_port, internal_inloc_data_3_1_port, 
      internal_inloc_data_3_0_port, internal_inloc_data_4_31_port, 
      internal_inloc_data_4_30_port, internal_inloc_data_4_29_port, 
      internal_inloc_data_4_28_port, internal_inloc_data_4_27_port, 
      internal_inloc_data_4_26_port, internal_inloc_data_4_25_port, 
      internal_inloc_data_4_24_port, internal_inloc_data_4_23_port, 
      internal_inloc_data_4_22_port, internal_inloc_data_4_21_port, 
      internal_inloc_data_4_20_port, internal_inloc_data_4_19_port, 
      internal_inloc_data_4_18_port, internal_inloc_data_4_17_port, 
      internal_inloc_data_4_16_port, internal_inloc_data_4_15_port, 
      internal_inloc_data_4_14_port, internal_inloc_data_4_13_port, 
      internal_inloc_data_4_12_port, internal_inloc_data_4_11_port, 
      internal_inloc_data_4_10_port, internal_inloc_data_4_9_port, 
      internal_inloc_data_4_8_port, internal_inloc_data_4_7_port, 
      internal_inloc_data_4_6_port, internal_inloc_data_4_5_port, 
      internal_inloc_data_4_4_port, internal_inloc_data_4_3_port, 
      internal_inloc_data_4_2_port, internal_inloc_data_4_1_port, 
      internal_inloc_data_4_0_port, dec_output_31_port, dec_output_30_port, 
      dec_output_29_port, dec_output_28_port, dec_output_27_port, 
      dec_output_26_port, dec_output_25_port, dec_output_24_port, 
      dec_output_23_port, dec_output_22_port, dec_output_21_port, 
      dec_output_20_port, dec_output_19_port, dec_output_18_port, 
      dec_output_17_port, dec_output_16_port, dec_output_15_port, 
      dec_output_14_port, dec_output_13_port, dec_output_12_port, 
      dec_output_11_port, dec_output_10_port, dec_output_9_port, 
      dec_output_8_port, dec_output_7_port, dec_output_6_port, 
      dec_output_5_port, dec_output_4_port, dec_output_3_port, 
      dec_output_2_port, dec_output_1_port, dec_output_0_port, 
      dec_out_with_wen_31_port, dec_out_with_wen_30_port, 
      dec_out_with_wen_29_port, dec_out_with_wen_28_port, 
      dec_out_with_wen_27_port, dec_out_with_wen_26_port, 
      dec_out_with_wen_25_port, dec_out_with_wen_24_port, 
      dec_out_with_wen_23_port, dec_out_with_wen_22_port, 
      dec_out_with_wen_21_port, dec_out_with_wen_20_port, 
      dec_out_with_wen_19_port, dec_out_with_wen_18_port, 
      dec_out_with_wen_17_port, dec_out_with_wen_16_port, 
      dec_out_with_wen_15_port, dec_out_with_wen_14_port, 
      dec_out_with_wen_13_port, dec_out_with_wen_12_port, 
      dec_out_with_wen_11_port, dec_out_with_wen_10_port, 
      dec_out_with_wen_9_port, dec_out_with_wen_8_port, dec_out_with_wen_7_port
      , dec_out_with_wen_6_port, dec_out_with_wen_5_port, 
      dec_out_with_wen_4_port, dec_out_with_wen_3_port, dec_out_with_wen_2_port
      , dec_out_with_wen_1_port, dec_out_with_wen_0_port, 
      fill_address_ext_15_port, fill_address_ext_14_port, 
      fill_address_ext_13_port, fill_address_ext_12_port, 
      fill_address_ext_11_port, fill_address_ext_10_port, 
      fill_address_ext_9_port, fill_address_ext_8_port, fill_address_ext_7_port
      , fill_address_ext_6_port, fill_address_ext_5_port, 
      fill_address_ext_4_port, fill_address_ext_3_port, fill_address_ext_2_port
      , fill_address_ext_1_port, fill_address_ext_0_port, 
      donespill_donefill_encoding_1_port, donespill_donefill_encoding_0_port, 
      c_swin_4_port, c_swin_3_port, c_swin_2_port, c_swin_1_port, c_swin_0_port
      , next_swp_4_port, next_swp_3_port, next_swp_2_port, next_swp_1_port, 
      next_swp_0_port, working_PUSH, bus_sel_savedwin_data_511_port, 
      bus_sel_savedwin_data_510_port, bus_sel_savedwin_data_509_port, 
      bus_sel_savedwin_data_508_port, bus_sel_savedwin_data_507_port, 
      bus_sel_savedwin_data_506_port, bus_sel_savedwin_data_505_port, 
      bus_sel_savedwin_data_504_port, bus_sel_savedwin_data_503_port, 
      bus_sel_savedwin_data_502_port, bus_sel_savedwin_data_501_port, 
      bus_sel_savedwin_data_500_port, bus_sel_savedwin_data_499_port, 
      bus_sel_savedwin_data_498_port, bus_sel_savedwin_data_497_port, 
      bus_sel_savedwin_data_496_port, bus_sel_savedwin_data_495_port, 
      bus_sel_savedwin_data_494_port, bus_sel_savedwin_data_493_port, 
      bus_sel_savedwin_data_492_port, bus_sel_savedwin_data_491_port, 
      bus_sel_savedwin_data_490_port, bus_sel_savedwin_data_489_port, 
      bus_sel_savedwin_data_488_port, bus_sel_savedwin_data_487_port, 
      bus_sel_savedwin_data_486_port, bus_sel_savedwin_data_485_port, 
      bus_sel_savedwin_data_484_port, bus_sel_savedwin_data_483_port, 
      bus_sel_savedwin_data_482_port, bus_sel_savedwin_data_481_port, 
      bus_sel_savedwin_data_480_port, bus_sel_savedwin_data_479_port, 
      bus_sel_savedwin_data_478_port, bus_sel_savedwin_data_477_port, 
      bus_sel_savedwin_data_476_port, bus_sel_savedwin_data_475_port, 
      bus_sel_savedwin_data_474_port, bus_sel_savedwin_data_473_port, 
      bus_sel_savedwin_data_472_port, bus_sel_savedwin_data_471_port, 
      bus_sel_savedwin_data_470_port, bus_sel_savedwin_data_469_port, 
      bus_sel_savedwin_data_468_port, bus_sel_savedwin_data_467_port, 
      bus_sel_savedwin_data_466_port, bus_sel_savedwin_data_465_port, 
      bus_sel_savedwin_data_464_port, bus_sel_savedwin_data_463_port, 
      bus_sel_savedwin_data_462_port, bus_sel_savedwin_data_461_port, 
      bus_sel_savedwin_data_460_port, bus_sel_savedwin_data_459_port, 
      bus_sel_savedwin_data_458_port, bus_sel_savedwin_data_457_port, 
      bus_sel_savedwin_data_456_port, bus_sel_savedwin_data_455_port, 
      bus_sel_savedwin_data_454_port, bus_sel_savedwin_data_453_port, 
      bus_sel_savedwin_data_452_port, bus_sel_savedwin_data_451_port, 
      bus_sel_savedwin_data_450_port, bus_sel_savedwin_data_449_port, 
      bus_sel_savedwin_data_448_port, bus_sel_savedwin_data_447_port, 
      bus_sel_savedwin_data_446_port, bus_sel_savedwin_data_445_port, 
      bus_sel_savedwin_data_444_port, bus_sel_savedwin_data_443_port, 
      bus_sel_savedwin_data_442_port, bus_sel_savedwin_data_441_port, 
      bus_sel_savedwin_data_440_port, bus_sel_savedwin_data_439_port, 
      bus_sel_savedwin_data_438_port, bus_sel_savedwin_data_437_port, 
      bus_sel_savedwin_data_436_port, bus_sel_savedwin_data_435_port, 
      bus_sel_savedwin_data_434_port, bus_sel_savedwin_data_433_port, 
      bus_sel_savedwin_data_432_port, bus_sel_savedwin_data_431_port, 
      bus_sel_savedwin_data_430_port, bus_sel_savedwin_data_429_port, 
      bus_sel_savedwin_data_428_port, bus_sel_savedwin_data_427_port, 
      bus_sel_savedwin_data_426_port, bus_sel_savedwin_data_425_port, 
      bus_sel_savedwin_data_424_port, bus_sel_savedwin_data_423_port, 
      bus_sel_savedwin_data_422_port, bus_sel_savedwin_data_421_port, 
      bus_sel_savedwin_data_420_port, bus_sel_savedwin_data_419_port, 
      bus_sel_savedwin_data_418_port, bus_sel_savedwin_data_417_port, 
      bus_sel_savedwin_data_416_port, bus_sel_savedwin_data_415_port, 
      bus_sel_savedwin_data_414_port, bus_sel_savedwin_data_413_port, 
      bus_sel_savedwin_data_412_port, bus_sel_savedwin_data_411_port, 
      bus_sel_savedwin_data_410_port, bus_sel_savedwin_data_409_port, 
      bus_sel_savedwin_data_408_port, bus_sel_savedwin_data_407_port, 
      bus_sel_savedwin_data_406_port, bus_sel_savedwin_data_405_port, 
      bus_sel_savedwin_data_404_port, bus_sel_savedwin_data_403_port, 
      bus_sel_savedwin_data_402_port, bus_sel_savedwin_data_401_port, 
      bus_sel_savedwin_data_400_port, bus_sel_savedwin_data_399_port, 
      bus_sel_savedwin_data_398_port, bus_sel_savedwin_data_397_port, 
      bus_sel_savedwin_data_396_port, bus_sel_savedwin_data_395_port, 
      bus_sel_savedwin_data_394_port, bus_sel_savedwin_data_393_port, 
      bus_sel_savedwin_data_392_port, bus_sel_savedwin_data_391_port, 
      bus_sel_savedwin_data_390_port, bus_sel_savedwin_data_389_port, 
      bus_sel_savedwin_data_388_port, bus_sel_savedwin_data_387_port, 
      bus_sel_savedwin_data_386_port, bus_sel_savedwin_data_385_port, 
      bus_sel_savedwin_data_384_port, bus_sel_savedwin_data_383_port, 
      bus_sel_savedwin_data_382_port, bus_sel_savedwin_data_381_port, 
      bus_sel_savedwin_data_380_port, bus_sel_savedwin_data_379_port, 
      bus_sel_savedwin_data_378_port, bus_sel_savedwin_data_377_port, 
      bus_sel_savedwin_data_376_port, bus_sel_savedwin_data_375_port, 
      bus_sel_savedwin_data_374_port, bus_sel_savedwin_data_373_port, 
      bus_sel_savedwin_data_372_port, bus_sel_savedwin_data_371_port, 
      bus_sel_savedwin_data_370_port, bus_sel_savedwin_data_369_port, 
      bus_sel_savedwin_data_368_port, bus_sel_savedwin_data_367_port, 
      bus_sel_savedwin_data_366_port, bus_sel_savedwin_data_365_port, 
      bus_sel_savedwin_data_364_port, bus_sel_savedwin_data_363_port, 
      bus_sel_savedwin_data_362_port, bus_sel_savedwin_data_361_port, 
      bus_sel_savedwin_data_360_port, bus_sel_savedwin_data_359_port, 
      bus_sel_savedwin_data_358_port, bus_sel_savedwin_data_357_port, 
      bus_sel_savedwin_data_356_port, bus_sel_savedwin_data_355_port, 
      bus_sel_savedwin_data_354_port, bus_sel_savedwin_data_353_port, 
      bus_sel_savedwin_data_352_port, bus_sel_savedwin_data_351_port, 
      bus_sel_savedwin_data_350_port, bus_sel_savedwin_data_349_port, 
      bus_sel_savedwin_data_348_port, bus_sel_savedwin_data_347_port, 
      bus_sel_savedwin_data_346_port, bus_sel_savedwin_data_345_port, 
      bus_sel_savedwin_data_344_port, bus_sel_savedwin_data_343_port, 
      bus_sel_savedwin_data_342_port, bus_sel_savedwin_data_341_port, 
      bus_sel_savedwin_data_340_port, bus_sel_savedwin_data_339_port, 
      bus_sel_savedwin_data_338_port, bus_sel_savedwin_data_337_port, 
      bus_sel_savedwin_data_336_port, bus_sel_savedwin_data_335_port, 
      bus_sel_savedwin_data_334_port, bus_sel_savedwin_data_333_port, 
      bus_sel_savedwin_data_332_port, bus_sel_savedwin_data_331_port, 
      bus_sel_savedwin_data_330_port, bus_sel_savedwin_data_329_port, 
      bus_sel_savedwin_data_328_port, bus_sel_savedwin_data_327_port, 
      bus_sel_savedwin_data_326_port, bus_sel_savedwin_data_325_port, 
      bus_sel_savedwin_data_324_port, bus_sel_savedwin_data_323_port, 
      bus_sel_savedwin_data_322_port, bus_sel_savedwin_data_321_port, 
      bus_sel_savedwin_data_320_port, bus_sel_savedwin_data_319_port, 
      bus_sel_savedwin_data_318_port, bus_sel_savedwin_data_317_port, 
      bus_sel_savedwin_data_316_port, bus_sel_savedwin_data_315_port, 
      bus_sel_savedwin_data_314_port, bus_sel_savedwin_data_313_port, 
      bus_sel_savedwin_data_312_port, bus_sel_savedwin_data_311_port, 
      bus_sel_savedwin_data_310_port, bus_sel_savedwin_data_309_port, 
      bus_sel_savedwin_data_308_port, bus_sel_savedwin_data_307_port, 
      bus_sel_savedwin_data_306_port, bus_sel_savedwin_data_305_port, 
      bus_sel_savedwin_data_304_port, bus_sel_savedwin_data_303_port, 
      bus_sel_savedwin_data_302_port, bus_sel_savedwin_data_301_port, 
      bus_sel_savedwin_data_300_port, bus_sel_savedwin_data_299_port, 
      bus_sel_savedwin_data_298_port, bus_sel_savedwin_data_297_port, 
      bus_sel_savedwin_data_296_port, bus_sel_savedwin_data_295_port, 
      bus_sel_savedwin_data_294_port, bus_sel_savedwin_data_293_port, 
      bus_sel_savedwin_data_292_port, bus_sel_savedwin_data_291_port, 
      bus_sel_savedwin_data_290_port, bus_sel_savedwin_data_289_port, 
      bus_sel_savedwin_data_288_port, bus_sel_savedwin_data_287_port, 
      bus_sel_savedwin_data_286_port, bus_sel_savedwin_data_285_port, 
      bus_sel_savedwin_data_284_port, bus_sel_savedwin_data_283_port, 
      bus_sel_savedwin_data_282_port, bus_sel_savedwin_data_281_port, 
      bus_sel_savedwin_data_280_port, bus_sel_savedwin_data_279_port, 
      bus_sel_savedwin_data_278_port, bus_sel_savedwin_data_277_port, 
      bus_sel_savedwin_data_276_port, bus_sel_savedwin_data_275_port, 
      bus_sel_savedwin_data_274_port, bus_sel_savedwin_data_273_port, 
      bus_sel_savedwin_data_272_port, bus_sel_savedwin_data_271_port, 
      bus_sel_savedwin_data_270_port, bus_sel_savedwin_data_269_port, 
      bus_sel_savedwin_data_268_port, bus_sel_savedwin_data_267_port, 
      bus_sel_savedwin_data_266_port, bus_sel_savedwin_data_265_port, 
      bus_sel_savedwin_data_264_port, bus_sel_savedwin_data_263_port, 
      bus_sel_savedwin_data_262_port, bus_sel_savedwin_data_261_port, 
      bus_sel_savedwin_data_260_port, bus_sel_savedwin_data_259_port, 
      bus_sel_savedwin_data_258_port, bus_sel_savedwin_data_257_port, 
      bus_sel_savedwin_data_256_port, bus_sel_savedwin_data_255_port, 
      bus_sel_savedwin_data_254_port, bus_sel_savedwin_data_253_port, 
      bus_sel_savedwin_data_252_port, bus_sel_savedwin_data_251_port, 
      bus_sel_savedwin_data_250_port, bus_sel_savedwin_data_249_port, 
      bus_sel_savedwin_data_248_port, bus_sel_savedwin_data_247_port, 
      bus_sel_savedwin_data_246_port, bus_sel_savedwin_data_245_port, 
      bus_sel_savedwin_data_244_port, bus_sel_savedwin_data_243_port, 
      bus_sel_savedwin_data_242_port, bus_sel_savedwin_data_241_port, 
      bus_sel_savedwin_data_240_port, bus_sel_savedwin_data_239_port, 
      bus_sel_savedwin_data_238_port, bus_sel_savedwin_data_237_port, 
      bus_sel_savedwin_data_236_port, bus_sel_savedwin_data_235_port, 
      bus_sel_savedwin_data_234_port, bus_sel_savedwin_data_233_port, 
      bus_sel_savedwin_data_232_port, bus_sel_savedwin_data_231_port, 
      bus_sel_savedwin_data_230_port, bus_sel_savedwin_data_229_port, 
      bus_sel_savedwin_data_228_port, bus_sel_savedwin_data_227_port, 
      bus_sel_savedwin_data_226_port, bus_sel_savedwin_data_225_port, 
      bus_sel_savedwin_data_224_port, bus_sel_savedwin_data_223_port, 
      bus_sel_savedwin_data_222_port, bus_sel_savedwin_data_221_port, 
      bus_sel_savedwin_data_220_port, bus_sel_savedwin_data_219_port, 
      bus_sel_savedwin_data_218_port, bus_sel_savedwin_data_217_port, 
      bus_sel_savedwin_data_216_port, bus_sel_savedwin_data_215_port, 
      bus_sel_savedwin_data_214_port, bus_sel_savedwin_data_213_port, 
      bus_sel_savedwin_data_212_port, bus_sel_savedwin_data_211_port, 
      bus_sel_savedwin_data_210_port, bus_sel_savedwin_data_209_port, 
      bus_sel_savedwin_data_208_port, bus_sel_savedwin_data_207_port, 
      bus_sel_savedwin_data_206_port, bus_sel_savedwin_data_205_port, 
      bus_sel_savedwin_data_204_port, bus_sel_savedwin_data_203_port, 
      bus_sel_savedwin_data_202_port, bus_sel_savedwin_data_201_port, 
      bus_sel_savedwin_data_200_port, bus_sel_savedwin_data_199_port, 
      bus_sel_savedwin_data_198_port, bus_sel_savedwin_data_197_port, 
      bus_sel_savedwin_data_196_port, bus_sel_savedwin_data_195_port, 
      bus_sel_savedwin_data_194_port, bus_sel_savedwin_data_193_port, 
      bus_sel_savedwin_data_192_port, bus_sel_savedwin_data_191_port, 
      bus_sel_savedwin_data_190_port, bus_sel_savedwin_data_189_port, 
      bus_sel_savedwin_data_188_port, bus_sel_savedwin_data_187_port, 
      bus_sel_savedwin_data_186_port, bus_sel_savedwin_data_185_port, 
      bus_sel_savedwin_data_184_port, bus_sel_savedwin_data_183_port, 
      bus_sel_savedwin_data_182_port, bus_sel_savedwin_data_181_port, 
      bus_sel_savedwin_data_180_port, bus_sel_savedwin_data_179_port, 
      bus_sel_savedwin_data_178_port, bus_sel_savedwin_data_177_port, 
      bus_sel_savedwin_data_176_port, bus_sel_savedwin_data_175_port, 
      bus_sel_savedwin_data_174_port, bus_sel_savedwin_data_173_port, 
      bus_sel_savedwin_data_172_port, bus_sel_savedwin_data_171_port, 
      bus_sel_savedwin_data_170_port, bus_sel_savedwin_data_169_port, 
      bus_sel_savedwin_data_168_port, bus_sel_savedwin_data_167_port, 
      bus_sel_savedwin_data_166_port, bus_sel_savedwin_data_165_port, 
      bus_sel_savedwin_data_164_port, bus_sel_savedwin_data_163_port, 
      bus_sel_savedwin_data_162_port, bus_sel_savedwin_data_161_port, 
      bus_sel_savedwin_data_160_port, bus_sel_savedwin_data_159_port, 
      bus_sel_savedwin_data_158_port, bus_sel_savedwin_data_157_port, 
      bus_sel_savedwin_data_156_port, bus_sel_savedwin_data_155_port, 
      bus_sel_savedwin_data_154_port, bus_sel_savedwin_data_153_port, 
      bus_sel_savedwin_data_152_port, bus_sel_savedwin_data_151_port, 
      bus_sel_savedwin_data_150_port, bus_sel_savedwin_data_149_port, 
      bus_sel_savedwin_data_148_port, bus_sel_savedwin_data_147_port, 
      bus_sel_savedwin_data_146_port, bus_sel_savedwin_data_145_port, 
      bus_sel_savedwin_data_144_port, bus_sel_savedwin_data_143_port, 
      bus_sel_savedwin_data_142_port, bus_sel_savedwin_data_141_port, 
      bus_sel_savedwin_data_140_port, bus_sel_savedwin_data_139_port, 
      bus_sel_savedwin_data_138_port, bus_sel_savedwin_data_137_port, 
      bus_sel_savedwin_data_136_port, bus_sel_savedwin_data_135_port, 
      bus_sel_savedwin_data_134_port, bus_sel_savedwin_data_133_port, 
      bus_sel_savedwin_data_132_port, bus_sel_savedwin_data_131_port, 
      bus_sel_savedwin_data_130_port, bus_sel_savedwin_data_129_port, 
      bus_sel_savedwin_data_128_port, bus_sel_savedwin_data_127_port, 
      bus_sel_savedwin_data_126_port, bus_sel_savedwin_data_125_port, 
      bus_sel_savedwin_data_124_port, bus_sel_savedwin_data_123_port, 
      bus_sel_savedwin_data_122_port, bus_sel_savedwin_data_121_port, 
      bus_sel_savedwin_data_120_port, bus_sel_savedwin_data_119_port, 
      bus_sel_savedwin_data_118_port, bus_sel_savedwin_data_117_port, 
      bus_sel_savedwin_data_116_port, bus_sel_savedwin_data_115_port, 
      bus_sel_savedwin_data_114_port, bus_sel_savedwin_data_113_port, 
      bus_sel_savedwin_data_112_port, bus_sel_savedwin_data_111_port, 
      bus_sel_savedwin_data_110_port, bus_sel_savedwin_data_109_port, 
      bus_sel_savedwin_data_108_port, bus_sel_savedwin_data_107_port, 
      bus_sel_savedwin_data_106_port, bus_sel_savedwin_data_105_port, 
      bus_sel_savedwin_data_104_port, bus_sel_savedwin_data_103_port, 
      bus_sel_savedwin_data_102_port, bus_sel_savedwin_data_101_port, 
      bus_sel_savedwin_data_100_port, bus_sel_savedwin_data_99_port, 
      bus_sel_savedwin_data_98_port, bus_sel_savedwin_data_97_port, 
      bus_sel_savedwin_data_96_port, bus_sel_savedwin_data_95_port, 
      bus_sel_savedwin_data_94_port, bus_sel_savedwin_data_93_port, 
      bus_sel_savedwin_data_92_port, bus_sel_savedwin_data_91_port, 
      bus_sel_savedwin_data_90_port, bus_sel_savedwin_data_89_port, 
      bus_sel_savedwin_data_88_port, bus_sel_savedwin_data_87_port, 
      bus_sel_savedwin_data_86_port, bus_sel_savedwin_data_85_port, 
      bus_sel_savedwin_data_84_port, bus_sel_savedwin_data_83_port, 
      bus_sel_savedwin_data_82_port, bus_sel_savedwin_data_81_port, 
      bus_sel_savedwin_data_80_port, bus_sel_savedwin_data_79_port, 
      bus_sel_savedwin_data_78_port, bus_sel_savedwin_data_77_port, 
      bus_sel_savedwin_data_76_port, bus_sel_savedwin_data_75_port, 
      bus_sel_savedwin_data_74_port, bus_sel_savedwin_data_73_port, 
      bus_sel_savedwin_data_72_port, bus_sel_savedwin_data_71_port, 
      bus_sel_savedwin_data_70_port, bus_sel_savedwin_data_69_port, 
      bus_sel_savedwin_data_68_port, bus_sel_savedwin_data_67_port, 
      bus_sel_savedwin_data_66_port, bus_sel_savedwin_data_65_port, 
      bus_sel_savedwin_data_64_port, bus_sel_savedwin_data_63_port, 
      bus_sel_savedwin_data_62_port, bus_sel_savedwin_data_61_port, 
      bus_sel_savedwin_data_60_port, bus_sel_savedwin_data_59_port, 
      bus_sel_savedwin_data_58_port, bus_sel_savedwin_data_57_port, 
      bus_sel_savedwin_data_56_port, bus_sel_savedwin_data_55_port, 
      bus_sel_savedwin_data_54_port, bus_sel_savedwin_data_53_port, 
      bus_sel_savedwin_data_52_port, bus_sel_savedwin_data_51_port, 
      bus_sel_savedwin_data_50_port, bus_sel_savedwin_data_49_port, 
      bus_sel_savedwin_data_48_port, bus_sel_savedwin_data_47_port, 
      bus_sel_savedwin_data_46_port, bus_sel_savedwin_data_45_port, 
      bus_sel_savedwin_data_44_port, bus_sel_savedwin_data_43_port, 
      bus_sel_savedwin_data_42_port, bus_sel_savedwin_data_41_port, 
      bus_sel_savedwin_data_40_port, bus_sel_savedwin_data_39_port, 
      bus_sel_savedwin_data_38_port, bus_sel_savedwin_data_37_port, 
      bus_sel_savedwin_data_36_port, bus_sel_savedwin_data_35_port, 
      bus_sel_savedwin_data_34_port, bus_sel_savedwin_data_33_port, 
      bus_sel_savedwin_data_32_port, bus_sel_savedwin_data_31_port, 
      bus_sel_savedwin_data_30_port, bus_sel_savedwin_data_29_port, 
      bus_sel_savedwin_data_28_port, bus_sel_savedwin_data_27_port, 
      bus_sel_savedwin_data_26_port, bus_sel_savedwin_data_25_port, 
      bus_sel_savedwin_data_24_port, bus_sel_savedwin_data_23_port, 
      bus_sel_savedwin_data_22_port, bus_sel_savedwin_data_21_port, 
      bus_sel_savedwin_data_20_port, bus_sel_savedwin_data_19_port, 
      bus_sel_savedwin_data_18_port, bus_sel_savedwin_data_17_port, 
      bus_sel_savedwin_data_16_port, bus_sel_savedwin_data_15_port, 
      bus_sel_savedwin_data_14_port, bus_sel_savedwin_data_13_port, 
      bus_sel_savedwin_data_12_port, bus_sel_savedwin_data_11_port, 
      bus_sel_savedwin_data_10_port, bus_sel_savedwin_data_9_port, 
      bus_sel_savedwin_data_8_port, bus_sel_savedwin_data_7_port, 
      bus_sel_savedwin_data_6_port, bus_sel_savedwin_data_5_port, 
      bus_sel_savedwin_data_4_port, bus_sel_savedwin_data_3_port, 
      bus_sel_savedwin_data_2_port, bus_sel_savedwin_data_1_port, 
      bus_sel_savedwin_data_0_port, spill_address_ext_15_port, 
      spill_address_ext_14_port, spill_address_ext_13_port, 
      spill_address_ext_12_port, spill_address_ext_11_port, 
      spill_address_ext_10_port, spill_address_ext_9_port, 
      spill_address_ext_8_port, spill_address_ext_7_port, 
      spill_address_ext_6_port, spill_address_ext_5_port, 
      spill_address_ext_4_port, spill_address_ext_3_port, 
      spill_address_ext_2_port, spill_address_ext_1_port, 
      spill_address_ext_0_port, spill_address_3_port, spill_address_2_port, 
      spill_address_1_port, spill_address_0_port, working_POP, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, FILL_port, n340, 
      n341, SPILL_port, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
      n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
      n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
      n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
      n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
      n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
      n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
      n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
      n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
      n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
      n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
      n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
      n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
      n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
      n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
      n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
      n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
      n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
      n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
      n1620, n1621, n1622 : std_logic;

begin
   FILL <= FILL_port;
   SPILL <= SPILL_port;
   
   X_Logic1_port <= '1';
   CWP_NEXT_CALC : nwin_calc_F5_0 port map( c_win(4) => c_win_4_port, c_win(3) 
                           => c_win_3_port, c_win(2) => c_win_2_port, c_win(1) 
                           => c_win_1_port, c_win(0) => c_win_0_port, sel(1) =>
                           n340, sel(0) => n341, n_win(4) => next_cwp_4_port, 
                           n_win(3) => next_cwp_3_port, n_win(2) => 
                           next_cwp_2_port, n_win(1) => next_cwp_1_port, 
                           n_win(0) => next_cwp_0_port);
   CWP : reg_generic_N5_RSTVAL1_0 port map( D(4) => next_cwp_4_port, D(3) => 
                           next_cwp_3_port, D(2) => next_cwp_2_port, D(1) => 
                           next_cwp_1_port, D(0) => next_cwp_0_port, Q(4) => 
                           c_win_4_port, Q(3) => c_win_3_port, Q(2) => 
                           c_win_2_port, Q(1) => c_win_1_port, Q(0) => 
                           c_win_0_port, Clk => CLK, Rst => RESET, Enable => 
                           X_Logic1_port);
   SEL_BLK : select_block_NBIT_DATA32_N8_F5 port map( regs(2559) => 
                           bus_reg_dataout_2559_port, regs(2558) => 
                           bus_reg_dataout_2558_port, regs(2557) => 
                           bus_reg_dataout_2557_port, regs(2556) => 
                           bus_reg_dataout_2556_port, regs(2555) => 
                           bus_reg_dataout_2555_port, regs(2554) => 
                           bus_reg_dataout_2554_port, regs(2553) => 
                           bus_reg_dataout_2553_port, regs(2552) => 
                           bus_reg_dataout_2552_port, regs(2551) => 
                           bus_reg_dataout_2551_port, regs(2550) => 
                           bus_reg_dataout_2550_port, regs(2549) => 
                           bus_reg_dataout_2549_port, regs(2548) => 
                           bus_reg_dataout_2548_port, regs(2547) => 
                           bus_reg_dataout_2547_port, regs(2546) => 
                           bus_reg_dataout_2546_port, regs(2545) => 
                           bus_reg_dataout_2545_port, regs(2544) => 
                           bus_reg_dataout_2544_port, regs(2543) => 
                           bus_reg_dataout_2543_port, regs(2542) => 
                           bus_reg_dataout_2542_port, regs(2541) => 
                           bus_reg_dataout_2541_port, regs(2540) => 
                           bus_reg_dataout_2540_port, regs(2539) => 
                           bus_reg_dataout_2539_port, regs(2538) => 
                           bus_reg_dataout_2538_port, regs(2537) => 
                           bus_reg_dataout_2537_port, regs(2536) => 
                           bus_reg_dataout_2536_port, regs(2535) => 
                           bus_reg_dataout_2535_port, regs(2534) => 
                           bus_reg_dataout_2534_port, regs(2533) => 
                           bus_reg_dataout_2533_port, regs(2532) => 
                           bus_reg_dataout_2532_port, regs(2531) => 
                           bus_reg_dataout_2531_port, regs(2530) => 
                           bus_reg_dataout_2530_port, regs(2529) => 
                           bus_reg_dataout_2529_port, regs(2528) => 
                           bus_reg_dataout_2528_port, regs(2527) => 
                           bus_reg_dataout_2527_port, regs(2526) => 
                           bus_reg_dataout_2526_port, regs(2525) => 
                           bus_reg_dataout_2525_port, regs(2524) => 
                           bus_reg_dataout_2524_port, regs(2523) => 
                           bus_reg_dataout_2523_port, regs(2522) => 
                           bus_reg_dataout_2522_port, regs(2521) => 
                           bus_reg_dataout_2521_port, regs(2520) => 
                           bus_reg_dataout_2520_port, regs(2519) => 
                           bus_reg_dataout_2519_port, regs(2518) => 
                           bus_reg_dataout_2518_port, regs(2517) => 
                           bus_reg_dataout_2517_port, regs(2516) => 
                           bus_reg_dataout_2516_port, regs(2515) => 
                           bus_reg_dataout_2515_port, regs(2514) => 
                           bus_reg_dataout_2514_port, regs(2513) => 
                           bus_reg_dataout_2513_port, regs(2512) => 
                           bus_reg_dataout_2512_port, regs(2511) => 
                           bus_reg_dataout_2511_port, regs(2510) => 
                           bus_reg_dataout_2510_port, regs(2509) => 
                           bus_reg_dataout_2509_port, regs(2508) => 
                           bus_reg_dataout_2508_port, regs(2507) => 
                           bus_reg_dataout_2507_port, regs(2506) => 
                           bus_reg_dataout_2506_port, regs(2505) => 
                           bus_reg_dataout_2505_port, regs(2504) => 
                           bus_reg_dataout_2504_port, regs(2503) => 
                           bus_reg_dataout_2503_port, regs(2502) => 
                           bus_reg_dataout_2502_port, regs(2501) => 
                           bus_reg_dataout_2501_port, regs(2500) => 
                           bus_reg_dataout_2500_port, regs(2499) => 
                           bus_reg_dataout_2499_port, regs(2498) => 
                           bus_reg_dataout_2498_port, regs(2497) => 
                           bus_reg_dataout_2497_port, regs(2496) => 
                           bus_reg_dataout_2496_port, regs(2495) => 
                           bus_reg_dataout_2495_port, regs(2494) => 
                           bus_reg_dataout_2494_port, regs(2493) => 
                           bus_reg_dataout_2493_port, regs(2492) => 
                           bus_reg_dataout_2492_port, regs(2491) => 
                           bus_reg_dataout_2491_port, regs(2490) => 
                           bus_reg_dataout_2490_port, regs(2489) => 
                           bus_reg_dataout_2489_port, regs(2488) => 
                           bus_reg_dataout_2488_port, regs(2487) => 
                           bus_reg_dataout_2487_port, regs(2486) => 
                           bus_reg_dataout_2486_port, regs(2485) => 
                           bus_reg_dataout_2485_port, regs(2484) => 
                           bus_reg_dataout_2484_port, regs(2483) => 
                           bus_reg_dataout_2483_port, regs(2482) => 
                           bus_reg_dataout_2482_port, regs(2481) => 
                           bus_reg_dataout_2481_port, regs(2480) => 
                           bus_reg_dataout_2480_port, regs(2479) => 
                           bus_reg_dataout_2479_port, regs(2478) => 
                           bus_reg_dataout_2478_port, regs(2477) => 
                           bus_reg_dataout_2477_port, regs(2476) => 
                           bus_reg_dataout_2476_port, regs(2475) => 
                           bus_reg_dataout_2475_port, regs(2474) => 
                           bus_reg_dataout_2474_port, regs(2473) => 
                           bus_reg_dataout_2473_port, regs(2472) => 
                           bus_reg_dataout_2472_port, regs(2471) => 
                           bus_reg_dataout_2471_port, regs(2470) => 
                           bus_reg_dataout_2470_port, regs(2469) => 
                           bus_reg_dataout_2469_port, regs(2468) => 
                           bus_reg_dataout_2468_port, regs(2467) => 
                           bus_reg_dataout_2467_port, regs(2466) => 
                           bus_reg_dataout_2466_port, regs(2465) => 
                           bus_reg_dataout_2465_port, regs(2464) => 
                           bus_reg_dataout_2464_port, regs(2463) => 
                           bus_reg_dataout_2463_port, regs(2462) => 
                           bus_reg_dataout_2462_port, regs(2461) => 
                           bus_reg_dataout_2461_port, regs(2460) => 
                           bus_reg_dataout_2460_port, regs(2459) => 
                           bus_reg_dataout_2459_port, regs(2458) => 
                           bus_reg_dataout_2458_port, regs(2457) => 
                           bus_reg_dataout_2457_port, regs(2456) => 
                           bus_reg_dataout_2456_port, regs(2455) => 
                           bus_reg_dataout_2455_port, regs(2454) => 
                           bus_reg_dataout_2454_port, regs(2453) => 
                           bus_reg_dataout_2453_port, regs(2452) => 
                           bus_reg_dataout_2452_port, regs(2451) => 
                           bus_reg_dataout_2451_port, regs(2450) => 
                           bus_reg_dataout_2450_port, regs(2449) => 
                           bus_reg_dataout_2449_port, regs(2448) => 
                           bus_reg_dataout_2448_port, regs(2447) => 
                           bus_reg_dataout_2447_port, regs(2446) => 
                           bus_reg_dataout_2446_port, regs(2445) => 
                           bus_reg_dataout_2445_port, regs(2444) => 
                           bus_reg_dataout_2444_port, regs(2443) => 
                           bus_reg_dataout_2443_port, regs(2442) => 
                           bus_reg_dataout_2442_port, regs(2441) => 
                           bus_reg_dataout_2441_port, regs(2440) => 
                           bus_reg_dataout_2440_port, regs(2439) => 
                           bus_reg_dataout_2439_port, regs(2438) => 
                           bus_reg_dataout_2438_port, regs(2437) => 
                           bus_reg_dataout_2437_port, regs(2436) => 
                           bus_reg_dataout_2436_port, regs(2435) => 
                           bus_reg_dataout_2435_port, regs(2434) => 
                           bus_reg_dataout_2434_port, regs(2433) => 
                           bus_reg_dataout_2433_port, regs(2432) => 
                           bus_reg_dataout_2432_port, regs(2431) => 
                           bus_reg_dataout_2431_port, regs(2430) => 
                           bus_reg_dataout_2430_port, regs(2429) => 
                           bus_reg_dataout_2429_port, regs(2428) => 
                           bus_reg_dataout_2428_port, regs(2427) => 
                           bus_reg_dataout_2427_port, regs(2426) => 
                           bus_reg_dataout_2426_port, regs(2425) => 
                           bus_reg_dataout_2425_port, regs(2424) => 
                           bus_reg_dataout_2424_port, regs(2423) => 
                           bus_reg_dataout_2423_port, regs(2422) => 
                           bus_reg_dataout_2422_port, regs(2421) => 
                           bus_reg_dataout_2421_port, regs(2420) => 
                           bus_reg_dataout_2420_port, regs(2419) => 
                           bus_reg_dataout_2419_port, regs(2418) => 
                           bus_reg_dataout_2418_port, regs(2417) => 
                           bus_reg_dataout_2417_port, regs(2416) => 
                           bus_reg_dataout_2416_port, regs(2415) => 
                           bus_reg_dataout_2415_port, regs(2414) => 
                           bus_reg_dataout_2414_port, regs(2413) => 
                           bus_reg_dataout_2413_port, regs(2412) => 
                           bus_reg_dataout_2412_port, regs(2411) => 
                           bus_reg_dataout_2411_port, regs(2410) => 
                           bus_reg_dataout_2410_port, regs(2409) => 
                           bus_reg_dataout_2409_port, regs(2408) => 
                           bus_reg_dataout_2408_port, regs(2407) => 
                           bus_reg_dataout_2407_port, regs(2406) => 
                           bus_reg_dataout_2406_port, regs(2405) => 
                           bus_reg_dataout_2405_port, regs(2404) => 
                           bus_reg_dataout_2404_port, regs(2403) => 
                           bus_reg_dataout_2403_port, regs(2402) => 
                           bus_reg_dataout_2402_port, regs(2401) => 
                           bus_reg_dataout_2401_port, regs(2400) => 
                           bus_reg_dataout_2400_port, regs(2399) => 
                           bus_reg_dataout_2399_port, regs(2398) => 
                           bus_reg_dataout_2398_port, regs(2397) => 
                           bus_reg_dataout_2397_port, regs(2396) => 
                           bus_reg_dataout_2396_port, regs(2395) => 
                           bus_reg_dataout_2395_port, regs(2394) => 
                           bus_reg_dataout_2394_port, regs(2393) => 
                           bus_reg_dataout_2393_port, regs(2392) => 
                           bus_reg_dataout_2392_port, regs(2391) => 
                           bus_reg_dataout_2391_port, regs(2390) => 
                           bus_reg_dataout_2390_port, regs(2389) => 
                           bus_reg_dataout_2389_port, regs(2388) => 
                           bus_reg_dataout_2388_port, regs(2387) => 
                           bus_reg_dataout_2387_port, regs(2386) => 
                           bus_reg_dataout_2386_port, regs(2385) => 
                           bus_reg_dataout_2385_port, regs(2384) => 
                           bus_reg_dataout_2384_port, regs(2383) => 
                           bus_reg_dataout_2383_port, regs(2382) => 
                           bus_reg_dataout_2382_port, regs(2381) => 
                           bus_reg_dataout_2381_port, regs(2380) => 
                           bus_reg_dataout_2380_port, regs(2379) => 
                           bus_reg_dataout_2379_port, regs(2378) => 
                           bus_reg_dataout_2378_port, regs(2377) => 
                           bus_reg_dataout_2377_port, regs(2376) => 
                           bus_reg_dataout_2376_port, regs(2375) => 
                           bus_reg_dataout_2375_port, regs(2374) => 
                           bus_reg_dataout_2374_port, regs(2373) => 
                           bus_reg_dataout_2373_port, regs(2372) => 
                           bus_reg_dataout_2372_port, regs(2371) => 
                           bus_reg_dataout_2371_port, regs(2370) => 
                           bus_reg_dataout_2370_port, regs(2369) => 
                           bus_reg_dataout_2369_port, regs(2368) => 
                           bus_reg_dataout_2368_port, regs(2367) => 
                           bus_reg_dataout_2367_port, regs(2366) => 
                           bus_reg_dataout_2366_port, regs(2365) => 
                           bus_reg_dataout_2365_port, regs(2364) => 
                           bus_reg_dataout_2364_port, regs(2363) => 
                           bus_reg_dataout_2363_port, regs(2362) => 
                           bus_reg_dataout_2362_port, regs(2361) => 
                           bus_reg_dataout_2361_port, regs(2360) => 
                           bus_reg_dataout_2360_port, regs(2359) => 
                           bus_reg_dataout_2359_port, regs(2358) => 
                           bus_reg_dataout_2358_port, regs(2357) => 
                           bus_reg_dataout_2357_port, regs(2356) => 
                           bus_reg_dataout_2356_port, regs(2355) => 
                           bus_reg_dataout_2355_port, regs(2354) => 
                           bus_reg_dataout_2354_port, regs(2353) => 
                           bus_reg_dataout_2353_port, regs(2352) => 
                           bus_reg_dataout_2352_port, regs(2351) => 
                           bus_reg_dataout_2351_port, regs(2350) => 
                           bus_reg_dataout_2350_port, regs(2349) => 
                           bus_reg_dataout_2349_port, regs(2348) => 
                           bus_reg_dataout_2348_port, regs(2347) => 
                           bus_reg_dataout_2347_port, regs(2346) => 
                           bus_reg_dataout_2346_port, regs(2345) => 
                           bus_reg_dataout_2345_port, regs(2344) => 
                           bus_reg_dataout_2344_port, regs(2343) => 
                           bus_reg_dataout_2343_port, regs(2342) => 
                           bus_reg_dataout_2342_port, regs(2341) => 
                           bus_reg_dataout_2341_port, regs(2340) => 
                           bus_reg_dataout_2340_port, regs(2339) => 
                           bus_reg_dataout_2339_port, regs(2338) => 
                           bus_reg_dataout_2338_port, regs(2337) => 
                           bus_reg_dataout_2337_port, regs(2336) => 
                           bus_reg_dataout_2336_port, regs(2335) => 
                           bus_reg_dataout_2335_port, regs(2334) => 
                           bus_reg_dataout_2334_port, regs(2333) => 
                           bus_reg_dataout_2333_port, regs(2332) => 
                           bus_reg_dataout_2332_port, regs(2331) => 
                           bus_reg_dataout_2331_port, regs(2330) => 
                           bus_reg_dataout_2330_port, regs(2329) => 
                           bus_reg_dataout_2329_port, regs(2328) => 
                           bus_reg_dataout_2328_port, regs(2327) => 
                           bus_reg_dataout_2327_port, regs(2326) => 
                           bus_reg_dataout_2326_port, regs(2325) => 
                           bus_reg_dataout_2325_port, regs(2324) => 
                           bus_reg_dataout_2324_port, regs(2323) => 
                           bus_reg_dataout_2323_port, regs(2322) => 
                           bus_reg_dataout_2322_port, regs(2321) => 
                           bus_reg_dataout_2321_port, regs(2320) => 
                           bus_reg_dataout_2320_port, regs(2319) => 
                           bus_reg_dataout_2319_port, regs(2318) => 
                           bus_reg_dataout_2318_port, regs(2317) => 
                           bus_reg_dataout_2317_port, regs(2316) => 
                           bus_reg_dataout_2316_port, regs(2315) => 
                           bus_reg_dataout_2315_port, regs(2314) => 
                           bus_reg_dataout_2314_port, regs(2313) => 
                           bus_reg_dataout_2313_port, regs(2312) => 
                           bus_reg_dataout_2312_port, regs(2311) => 
                           bus_reg_dataout_2311_port, regs(2310) => 
                           bus_reg_dataout_2310_port, regs(2309) => 
                           bus_reg_dataout_2309_port, regs(2308) => 
                           bus_reg_dataout_2308_port, regs(2307) => 
                           bus_reg_dataout_2307_port, regs(2306) => 
                           bus_reg_dataout_2306_port, regs(2305) => 
                           bus_reg_dataout_2305_port, regs(2304) => 
                           bus_reg_dataout_2304_port, regs(2303) => 
                           bus_reg_dataout_2303_port, regs(2302) => 
                           bus_reg_dataout_2302_port, regs(2301) => 
                           bus_reg_dataout_2301_port, regs(2300) => 
                           bus_reg_dataout_2300_port, regs(2299) => 
                           bus_reg_dataout_2299_port, regs(2298) => 
                           bus_reg_dataout_2298_port, regs(2297) => 
                           bus_reg_dataout_2297_port, regs(2296) => 
                           bus_reg_dataout_2296_port, regs(2295) => 
                           bus_reg_dataout_2295_port, regs(2294) => 
                           bus_reg_dataout_2294_port, regs(2293) => 
                           bus_reg_dataout_2293_port, regs(2292) => 
                           bus_reg_dataout_2292_port, regs(2291) => 
                           bus_reg_dataout_2291_port, regs(2290) => 
                           bus_reg_dataout_2290_port, regs(2289) => 
                           bus_reg_dataout_2289_port, regs(2288) => 
                           bus_reg_dataout_2288_port, regs(2287) => 
                           bus_reg_dataout_2287_port, regs(2286) => 
                           bus_reg_dataout_2286_port, regs(2285) => 
                           bus_reg_dataout_2285_port, regs(2284) => 
                           bus_reg_dataout_2284_port, regs(2283) => 
                           bus_reg_dataout_2283_port, regs(2282) => 
                           bus_reg_dataout_2282_port, regs(2281) => 
                           bus_reg_dataout_2281_port, regs(2280) => 
                           bus_reg_dataout_2280_port, regs(2279) => 
                           bus_reg_dataout_2279_port, regs(2278) => 
                           bus_reg_dataout_2278_port, regs(2277) => 
                           bus_reg_dataout_2277_port, regs(2276) => 
                           bus_reg_dataout_2276_port, regs(2275) => 
                           bus_reg_dataout_2275_port, regs(2274) => 
                           bus_reg_dataout_2274_port, regs(2273) => 
                           bus_reg_dataout_2273_port, regs(2272) => 
                           bus_reg_dataout_2272_port, regs(2271) => 
                           bus_reg_dataout_2271_port, regs(2270) => 
                           bus_reg_dataout_2270_port, regs(2269) => 
                           bus_reg_dataout_2269_port, regs(2268) => 
                           bus_reg_dataout_2268_port, regs(2267) => 
                           bus_reg_dataout_2267_port, regs(2266) => 
                           bus_reg_dataout_2266_port, regs(2265) => 
                           bus_reg_dataout_2265_port, regs(2264) => 
                           bus_reg_dataout_2264_port, regs(2263) => 
                           bus_reg_dataout_2263_port, regs(2262) => 
                           bus_reg_dataout_2262_port, regs(2261) => 
                           bus_reg_dataout_2261_port, regs(2260) => 
                           bus_reg_dataout_2260_port, regs(2259) => 
                           bus_reg_dataout_2259_port, regs(2258) => 
                           bus_reg_dataout_2258_port, regs(2257) => 
                           bus_reg_dataout_2257_port, regs(2256) => 
                           bus_reg_dataout_2256_port, regs(2255) => 
                           bus_reg_dataout_2255_port, regs(2254) => 
                           bus_reg_dataout_2254_port, regs(2253) => 
                           bus_reg_dataout_2253_port, regs(2252) => 
                           bus_reg_dataout_2252_port, regs(2251) => 
                           bus_reg_dataout_2251_port, regs(2250) => 
                           bus_reg_dataout_2250_port, regs(2249) => 
                           bus_reg_dataout_2249_port, regs(2248) => 
                           bus_reg_dataout_2248_port, regs(2247) => 
                           bus_reg_dataout_2247_port, regs(2246) => 
                           bus_reg_dataout_2246_port, regs(2245) => 
                           bus_reg_dataout_2245_port, regs(2244) => 
                           bus_reg_dataout_2244_port, regs(2243) => 
                           bus_reg_dataout_2243_port, regs(2242) => 
                           bus_reg_dataout_2242_port, regs(2241) => 
                           bus_reg_dataout_2241_port, regs(2240) => 
                           bus_reg_dataout_2240_port, regs(2239) => 
                           bus_reg_dataout_2239_port, regs(2238) => 
                           bus_reg_dataout_2238_port, regs(2237) => 
                           bus_reg_dataout_2237_port, regs(2236) => 
                           bus_reg_dataout_2236_port, regs(2235) => 
                           bus_reg_dataout_2235_port, regs(2234) => 
                           bus_reg_dataout_2234_port, regs(2233) => 
                           bus_reg_dataout_2233_port, regs(2232) => 
                           bus_reg_dataout_2232_port, regs(2231) => 
                           bus_reg_dataout_2231_port, regs(2230) => 
                           bus_reg_dataout_2230_port, regs(2229) => 
                           bus_reg_dataout_2229_port, regs(2228) => 
                           bus_reg_dataout_2228_port, regs(2227) => 
                           bus_reg_dataout_2227_port, regs(2226) => 
                           bus_reg_dataout_2226_port, regs(2225) => 
                           bus_reg_dataout_2225_port, regs(2224) => 
                           bus_reg_dataout_2224_port, regs(2223) => 
                           bus_reg_dataout_2223_port, regs(2222) => 
                           bus_reg_dataout_2222_port, regs(2221) => 
                           bus_reg_dataout_2221_port, regs(2220) => 
                           bus_reg_dataout_2220_port, regs(2219) => 
                           bus_reg_dataout_2219_port, regs(2218) => 
                           bus_reg_dataout_2218_port, regs(2217) => 
                           bus_reg_dataout_2217_port, regs(2216) => 
                           bus_reg_dataout_2216_port, regs(2215) => 
                           bus_reg_dataout_2215_port, regs(2214) => 
                           bus_reg_dataout_2214_port, regs(2213) => 
                           bus_reg_dataout_2213_port, regs(2212) => 
                           bus_reg_dataout_2212_port, regs(2211) => 
                           bus_reg_dataout_2211_port, regs(2210) => 
                           bus_reg_dataout_2210_port, regs(2209) => 
                           bus_reg_dataout_2209_port, regs(2208) => 
                           bus_reg_dataout_2208_port, regs(2207) => 
                           bus_reg_dataout_2207_port, regs(2206) => 
                           bus_reg_dataout_2206_port, regs(2205) => 
                           bus_reg_dataout_2205_port, regs(2204) => 
                           bus_reg_dataout_2204_port, regs(2203) => 
                           bus_reg_dataout_2203_port, regs(2202) => 
                           bus_reg_dataout_2202_port, regs(2201) => 
                           bus_reg_dataout_2201_port, regs(2200) => 
                           bus_reg_dataout_2200_port, regs(2199) => 
                           bus_reg_dataout_2199_port, regs(2198) => 
                           bus_reg_dataout_2198_port, regs(2197) => 
                           bus_reg_dataout_2197_port, regs(2196) => 
                           bus_reg_dataout_2196_port, regs(2195) => 
                           bus_reg_dataout_2195_port, regs(2194) => 
                           bus_reg_dataout_2194_port, regs(2193) => 
                           bus_reg_dataout_2193_port, regs(2192) => 
                           bus_reg_dataout_2192_port, regs(2191) => 
                           bus_reg_dataout_2191_port, regs(2190) => 
                           bus_reg_dataout_2190_port, regs(2189) => 
                           bus_reg_dataout_2189_port, regs(2188) => 
                           bus_reg_dataout_2188_port, regs(2187) => 
                           bus_reg_dataout_2187_port, regs(2186) => 
                           bus_reg_dataout_2186_port, regs(2185) => 
                           bus_reg_dataout_2185_port, regs(2184) => 
                           bus_reg_dataout_2184_port, regs(2183) => 
                           bus_reg_dataout_2183_port, regs(2182) => 
                           bus_reg_dataout_2182_port, regs(2181) => 
                           bus_reg_dataout_2181_port, regs(2180) => 
                           bus_reg_dataout_2180_port, regs(2179) => 
                           bus_reg_dataout_2179_port, regs(2178) => 
                           bus_reg_dataout_2178_port, regs(2177) => 
                           bus_reg_dataout_2177_port, regs(2176) => 
                           bus_reg_dataout_2176_port, regs(2175) => 
                           bus_reg_dataout_2175_port, regs(2174) => 
                           bus_reg_dataout_2174_port, regs(2173) => 
                           bus_reg_dataout_2173_port, regs(2172) => 
                           bus_reg_dataout_2172_port, regs(2171) => 
                           bus_reg_dataout_2171_port, regs(2170) => 
                           bus_reg_dataout_2170_port, regs(2169) => 
                           bus_reg_dataout_2169_port, regs(2168) => 
                           bus_reg_dataout_2168_port, regs(2167) => 
                           bus_reg_dataout_2167_port, regs(2166) => 
                           bus_reg_dataout_2166_port, regs(2165) => 
                           bus_reg_dataout_2165_port, regs(2164) => 
                           bus_reg_dataout_2164_port, regs(2163) => 
                           bus_reg_dataout_2163_port, regs(2162) => 
                           bus_reg_dataout_2162_port, regs(2161) => 
                           bus_reg_dataout_2161_port, regs(2160) => 
                           bus_reg_dataout_2160_port, regs(2159) => 
                           bus_reg_dataout_2159_port, regs(2158) => 
                           bus_reg_dataout_2158_port, regs(2157) => 
                           bus_reg_dataout_2157_port, regs(2156) => 
                           bus_reg_dataout_2156_port, regs(2155) => 
                           bus_reg_dataout_2155_port, regs(2154) => 
                           bus_reg_dataout_2154_port, regs(2153) => 
                           bus_reg_dataout_2153_port, regs(2152) => 
                           bus_reg_dataout_2152_port, regs(2151) => 
                           bus_reg_dataout_2151_port, regs(2150) => 
                           bus_reg_dataout_2150_port, regs(2149) => 
                           bus_reg_dataout_2149_port, regs(2148) => 
                           bus_reg_dataout_2148_port, regs(2147) => 
                           bus_reg_dataout_2147_port, regs(2146) => 
                           bus_reg_dataout_2146_port, regs(2145) => 
                           bus_reg_dataout_2145_port, regs(2144) => 
                           bus_reg_dataout_2144_port, regs(2143) => 
                           bus_reg_dataout_2143_port, regs(2142) => 
                           bus_reg_dataout_2142_port, regs(2141) => 
                           bus_reg_dataout_2141_port, regs(2140) => 
                           bus_reg_dataout_2140_port, regs(2139) => 
                           bus_reg_dataout_2139_port, regs(2138) => 
                           bus_reg_dataout_2138_port, regs(2137) => 
                           bus_reg_dataout_2137_port, regs(2136) => 
                           bus_reg_dataout_2136_port, regs(2135) => 
                           bus_reg_dataout_2135_port, regs(2134) => 
                           bus_reg_dataout_2134_port, regs(2133) => 
                           bus_reg_dataout_2133_port, regs(2132) => 
                           bus_reg_dataout_2132_port, regs(2131) => 
                           bus_reg_dataout_2131_port, regs(2130) => 
                           bus_reg_dataout_2130_port, regs(2129) => 
                           bus_reg_dataout_2129_port, regs(2128) => 
                           bus_reg_dataout_2128_port, regs(2127) => 
                           bus_reg_dataout_2127_port, regs(2126) => 
                           bus_reg_dataout_2126_port, regs(2125) => 
                           bus_reg_dataout_2125_port, regs(2124) => 
                           bus_reg_dataout_2124_port, regs(2123) => 
                           bus_reg_dataout_2123_port, regs(2122) => 
                           bus_reg_dataout_2122_port, regs(2121) => 
                           bus_reg_dataout_2121_port, regs(2120) => 
                           bus_reg_dataout_2120_port, regs(2119) => 
                           bus_reg_dataout_2119_port, regs(2118) => 
                           bus_reg_dataout_2118_port, regs(2117) => 
                           bus_reg_dataout_2117_port, regs(2116) => 
                           bus_reg_dataout_2116_port, regs(2115) => 
                           bus_reg_dataout_2115_port, regs(2114) => 
                           bus_reg_dataout_2114_port, regs(2113) => 
                           bus_reg_dataout_2113_port, regs(2112) => 
                           bus_reg_dataout_2112_port, regs(2111) => 
                           bus_reg_dataout_2111_port, regs(2110) => 
                           bus_reg_dataout_2110_port, regs(2109) => 
                           bus_reg_dataout_2109_port, regs(2108) => 
                           bus_reg_dataout_2108_port, regs(2107) => 
                           bus_reg_dataout_2107_port, regs(2106) => 
                           bus_reg_dataout_2106_port, regs(2105) => 
                           bus_reg_dataout_2105_port, regs(2104) => 
                           bus_reg_dataout_2104_port, regs(2103) => 
                           bus_reg_dataout_2103_port, regs(2102) => 
                           bus_reg_dataout_2102_port, regs(2101) => 
                           bus_reg_dataout_2101_port, regs(2100) => 
                           bus_reg_dataout_2100_port, regs(2099) => 
                           bus_reg_dataout_2099_port, regs(2098) => 
                           bus_reg_dataout_2098_port, regs(2097) => 
                           bus_reg_dataout_2097_port, regs(2096) => 
                           bus_reg_dataout_2096_port, regs(2095) => 
                           bus_reg_dataout_2095_port, regs(2094) => 
                           bus_reg_dataout_2094_port, regs(2093) => 
                           bus_reg_dataout_2093_port, regs(2092) => 
                           bus_reg_dataout_2092_port, regs(2091) => 
                           bus_reg_dataout_2091_port, regs(2090) => 
                           bus_reg_dataout_2090_port, regs(2089) => 
                           bus_reg_dataout_2089_port, regs(2088) => 
                           bus_reg_dataout_2088_port, regs(2087) => 
                           bus_reg_dataout_2087_port, regs(2086) => 
                           bus_reg_dataout_2086_port, regs(2085) => 
                           bus_reg_dataout_2085_port, regs(2084) => 
                           bus_reg_dataout_2084_port, regs(2083) => 
                           bus_reg_dataout_2083_port, regs(2082) => 
                           bus_reg_dataout_2082_port, regs(2081) => 
                           bus_reg_dataout_2081_port, regs(2080) => 
                           bus_reg_dataout_2080_port, regs(2079) => 
                           bus_reg_dataout_2079_port, regs(2078) => 
                           bus_reg_dataout_2078_port, regs(2077) => 
                           bus_reg_dataout_2077_port, regs(2076) => 
                           bus_reg_dataout_2076_port, regs(2075) => 
                           bus_reg_dataout_2075_port, regs(2074) => 
                           bus_reg_dataout_2074_port, regs(2073) => 
                           bus_reg_dataout_2073_port, regs(2072) => 
                           bus_reg_dataout_2072_port, regs(2071) => 
                           bus_reg_dataout_2071_port, regs(2070) => 
                           bus_reg_dataout_2070_port, regs(2069) => 
                           bus_reg_dataout_2069_port, regs(2068) => 
                           bus_reg_dataout_2068_port, regs(2067) => 
                           bus_reg_dataout_2067_port, regs(2066) => 
                           bus_reg_dataout_2066_port, regs(2065) => 
                           bus_reg_dataout_2065_port, regs(2064) => 
                           bus_reg_dataout_2064_port, regs(2063) => 
                           bus_reg_dataout_2063_port, regs(2062) => 
                           bus_reg_dataout_2062_port, regs(2061) => 
                           bus_reg_dataout_2061_port, regs(2060) => 
                           bus_reg_dataout_2060_port, regs(2059) => 
                           bus_reg_dataout_2059_port, regs(2058) => 
                           bus_reg_dataout_2058_port, regs(2057) => 
                           bus_reg_dataout_2057_port, regs(2056) => 
                           bus_reg_dataout_2056_port, regs(2055) => 
                           bus_reg_dataout_2055_port, regs(2054) => 
                           bus_reg_dataout_2054_port, regs(2053) => 
                           bus_reg_dataout_2053_port, regs(2052) => 
                           bus_reg_dataout_2052_port, regs(2051) => 
                           bus_reg_dataout_2051_port, regs(2050) => 
                           bus_reg_dataout_2050_port, regs(2049) => 
                           bus_reg_dataout_2049_port, regs(2048) => 
                           bus_reg_dataout_2048_port, regs(2047) => 
                           bus_reg_dataout_2047_port, regs(2046) => 
                           bus_reg_dataout_2046_port, regs(2045) => 
                           bus_reg_dataout_2045_port, regs(2044) => 
                           bus_reg_dataout_2044_port, regs(2043) => 
                           bus_reg_dataout_2043_port, regs(2042) => 
                           bus_reg_dataout_2042_port, regs(2041) => 
                           bus_reg_dataout_2041_port, regs(2040) => 
                           bus_reg_dataout_2040_port, regs(2039) => 
                           bus_reg_dataout_2039_port, regs(2038) => 
                           bus_reg_dataout_2038_port, regs(2037) => 
                           bus_reg_dataout_2037_port, regs(2036) => 
                           bus_reg_dataout_2036_port, regs(2035) => 
                           bus_reg_dataout_2035_port, regs(2034) => 
                           bus_reg_dataout_2034_port, regs(2033) => 
                           bus_reg_dataout_2033_port, regs(2032) => 
                           bus_reg_dataout_2032_port, regs(2031) => 
                           bus_reg_dataout_2031_port, regs(2030) => 
                           bus_reg_dataout_2030_port, regs(2029) => 
                           bus_reg_dataout_2029_port, regs(2028) => 
                           bus_reg_dataout_2028_port, regs(2027) => 
                           bus_reg_dataout_2027_port, regs(2026) => 
                           bus_reg_dataout_2026_port, regs(2025) => 
                           bus_reg_dataout_2025_port, regs(2024) => 
                           bus_reg_dataout_2024_port, regs(2023) => 
                           bus_reg_dataout_2023_port, regs(2022) => 
                           bus_reg_dataout_2022_port, regs(2021) => 
                           bus_reg_dataout_2021_port, regs(2020) => 
                           bus_reg_dataout_2020_port, regs(2019) => 
                           bus_reg_dataout_2019_port, regs(2018) => 
                           bus_reg_dataout_2018_port, regs(2017) => 
                           bus_reg_dataout_2017_port, regs(2016) => 
                           bus_reg_dataout_2016_port, regs(2015) => 
                           bus_reg_dataout_2015_port, regs(2014) => 
                           bus_reg_dataout_2014_port, regs(2013) => 
                           bus_reg_dataout_2013_port, regs(2012) => 
                           bus_reg_dataout_2012_port, regs(2011) => 
                           bus_reg_dataout_2011_port, regs(2010) => 
                           bus_reg_dataout_2010_port, regs(2009) => 
                           bus_reg_dataout_2009_port, regs(2008) => 
                           bus_reg_dataout_2008_port, regs(2007) => 
                           bus_reg_dataout_2007_port, regs(2006) => 
                           bus_reg_dataout_2006_port, regs(2005) => 
                           bus_reg_dataout_2005_port, regs(2004) => 
                           bus_reg_dataout_2004_port, regs(2003) => 
                           bus_reg_dataout_2003_port, regs(2002) => 
                           bus_reg_dataout_2002_port, regs(2001) => 
                           bus_reg_dataout_2001_port, regs(2000) => 
                           bus_reg_dataout_2000_port, regs(1999) => 
                           bus_reg_dataout_1999_port, regs(1998) => 
                           bus_reg_dataout_1998_port, regs(1997) => 
                           bus_reg_dataout_1997_port, regs(1996) => 
                           bus_reg_dataout_1996_port, regs(1995) => 
                           bus_reg_dataout_1995_port, regs(1994) => 
                           bus_reg_dataout_1994_port, regs(1993) => 
                           bus_reg_dataout_1993_port, regs(1992) => 
                           bus_reg_dataout_1992_port, regs(1991) => 
                           bus_reg_dataout_1991_port, regs(1990) => 
                           bus_reg_dataout_1990_port, regs(1989) => 
                           bus_reg_dataout_1989_port, regs(1988) => 
                           bus_reg_dataout_1988_port, regs(1987) => 
                           bus_reg_dataout_1987_port, regs(1986) => 
                           bus_reg_dataout_1986_port, regs(1985) => 
                           bus_reg_dataout_1985_port, regs(1984) => 
                           bus_reg_dataout_1984_port, regs(1983) => 
                           bus_reg_dataout_1983_port, regs(1982) => 
                           bus_reg_dataout_1982_port, regs(1981) => 
                           bus_reg_dataout_1981_port, regs(1980) => 
                           bus_reg_dataout_1980_port, regs(1979) => 
                           bus_reg_dataout_1979_port, regs(1978) => 
                           bus_reg_dataout_1978_port, regs(1977) => 
                           bus_reg_dataout_1977_port, regs(1976) => 
                           bus_reg_dataout_1976_port, regs(1975) => 
                           bus_reg_dataout_1975_port, regs(1974) => 
                           bus_reg_dataout_1974_port, regs(1973) => 
                           bus_reg_dataout_1973_port, regs(1972) => 
                           bus_reg_dataout_1972_port, regs(1971) => 
                           bus_reg_dataout_1971_port, regs(1970) => 
                           bus_reg_dataout_1970_port, regs(1969) => 
                           bus_reg_dataout_1969_port, regs(1968) => 
                           bus_reg_dataout_1968_port, regs(1967) => 
                           bus_reg_dataout_1967_port, regs(1966) => 
                           bus_reg_dataout_1966_port, regs(1965) => 
                           bus_reg_dataout_1965_port, regs(1964) => 
                           bus_reg_dataout_1964_port, regs(1963) => 
                           bus_reg_dataout_1963_port, regs(1962) => 
                           bus_reg_dataout_1962_port, regs(1961) => 
                           bus_reg_dataout_1961_port, regs(1960) => 
                           bus_reg_dataout_1960_port, regs(1959) => 
                           bus_reg_dataout_1959_port, regs(1958) => 
                           bus_reg_dataout_1958_port, regs(1957) => 
                           bus_reg_dataout_1957_port, regs(1956) => 
                           bus_reg_dataout_1956_port, regs(1955) => 
                           bus_reg_dataout_1955_port, regs(1954) => 
                           bus_reg_dataout_1954_port, regs(1953) => 
                           bus_reg_dataout_1953_port, regs(1952) => 
                           bus_reg_dataout_1952_port, regs(1951) => 
                           bus_reg_dataout_1951_port, regs(1950) => 
                           bus_reg_dataout_1950_port, regs(1949) => 
                           bus_reg_dataout_1949_port, regs(1948) => 
                           bus_reg_dataout_1948_port, regs(1947) => 
                           bus_reg_dataout_1947_port, regs(1946) => 
                           bus_reg_dataout_1946_port, regs(1945) => 
                           bus_reg_dataout_1945_port, regs(1944) => 
                           bus_reg_dataout_1944_port, regs(1943) => 
                           bus_reg_dataout_1943_port, regs(1942) => 
                           bus_reg_dataout_1942_port, regs(1941) => 
                           bus_reg_dataout_1941_port, regs(1940) => 
                           bus_reg_dataout_1940_port, regs(1939) => 
                           bus_reg_dataout_1939_port, regs(1938) => 
                           bus_reg_dataout_1938_port, regs(1937) => 
                           bus_reg_dataout_1937_port, regs(1936) => 
                           bus_reg_dataout_1936_port, regs(1935) => 
                           bus_reg_dataout_1935_port, regs(1934) => 
                           bus_reg_dataout_1934_port, regs(1933) => 
                           bus_reg_dataout_1933_port, regs(1932) => 
                           bus_reg_dataout_1932_port, regs(1931) => 
                           bus_reg_dataout_1931_port, regs(1930) => 
                           bus_reg_dataout_1930_port, regs(1929) => 
                           bus_reg_dataout_1929_port, regs(1928) => 
                           bus_reg_dataout_1928_port, regs(1927) => 
                           bus_reg_dataout_1927_port, regs(1926) => 
                           bus_reg_dataout_1926_port, regs(1925) => 
                           bus_reg_dataout_1925_port, regs(1924) => 
                           bus_reg_dataout_1924_port, regs(1923) => 
                           bus_reg_dataout_1923_port, regs(1922) => 
                           bus_reg_dataout_1922_port, regs(1921) => 
                           bus_reg_dataout_1921_port, regs(1920) => 
                           bus_reg_dataout_1920_port, regs(1919) => 
                           bus_reg_dataout_1919_port, regs(1918) => 
                           bus_reg_dataout_1918_port, regs(1917) => 
                           bus_reg_dataout_1917_port, regs(1916) => 
                           bus_reg_dataout_1916_port, regs(1915) => 
                           bus_reg_dataout_1915_port, regs(1914) => 
                           bus_reg_dataout_1914_port, regs(1913) => 
                           bus_reg_dataout_1913_port, regs(1912) => 
                           bus_reg_dataout_1912_port, regs(1911) => 
                           bus_reg_dataout_1911_port, regs(1910) => 
                           bus_reg_dataout_1910_port, regs(1909) => 
                           bus_reg_dataout_1909_port, regs(1908) => 
                           bus_reg_dataout_1908_port, regs(1907) => 
                           bus_reg_dataout_1907_port, regs(1906) => 
                           bus_reg_dataout_1906_port, regs(1905) => 
                           bus_reg_dataout_1905_port, regs(1904) => 
                           bus_reg_dataout_1904_port, regs(1903) => 
                           bus_reg_dataout_1903_port, regs(1902) => 
                           bus_reg_dataout_1902_port, regs(1901) => 
                           bus_reg_dataout_1901_port, regs(1900) => 
                           bus_reg_dataout_1900_port, regs(1899) => 
                           bus_reg_dataout_1899_port, regs(1898) => 
                           bus_reg_dataout_1898_port, regs(1897) => 
                           bus_reg_dataout_1897_port, regs(1896) => 
                           bus_reg_dataout_1896_port, regs(1895) => 
                           bus_reg_dataout_1895_port, regs(1894) => 
                           bus_reg_dataout_1894_port, regs(1893) => 
                           bus_reg_dataout_1893_port, regs(1892) => 
                           bus_reg_dataout_1892_port, regs(1891) => 
                           bus_reg_dataout_1891_port, regs(1890) => 
                           bus_reg_dataout_1890_port, regs(1889) => 
                           bus_reg_dataout_1889_port, regs(1888) => 
                           bus_reg_dataout_1888_port, regs(1887) => 
                           bus_reg_dataout_1887_port, regs(1886) => 
                           bus_reg_dataout_1886_port, regs(1885) => 
                           bus_reg_dataout_1885_port, regs(1884) => 
                           bus_reg_dataout_1884_port, regs(1883) => 
                           bus_reg_dataout_1883_port, regs(1882) => 
                           bus_reg_dataout_1882_port, regs(1881) => 
                           bus_reg_dataout_1881_port, regs(1880) => 
                           bus_reg_dataout_1880_port, regs(1879) => 
                           bus_reg_dataout_1879_port, regs(1878) => 
                           bus_reg_dataout_1878_port, regs(1877) => 
                           bus_reg_dataout_1877_port, regs(1876) => 
                           bus_reg_dataout_1876_port, regs(1875) => 
                           bus_reg_dataout_1875_port, regs(1874) => 
                           bus_reg_dataout_1874_port, regs(1873) => 
                           bus_reg_dataout_1873_port, regs(1872) => 
                           bus_reg_dataout_1872_port, regs(1871) => 
                           bus_reg_dataout_1871_port, regs(1870) => 
                           bus_reg_dataout_1870_port, regs(1869) => 
                           bus_reg_dataout_1869_port, regs(1868) => 
                           bus_reg_dataout_1868_port, regs(1867) => 
                           bus_reg_dataout_1867_port, regs(1866) => 
                           bus_reg_dataout_1866_port, regs(1865) => 
                           bus_reg_dataout_1865_port, regs(1864) => 
                           bus_reg_dataout_1864_port, regs(1863) => 
                           bus_reg_dataout_1863_port, regs(1862) => 
                           bus_reg_dataout_1862_port, regs(1861) => 
                           bus_reg_dataout_1861_port, regs(1860) => 
                           bus_reg_dataout_1860_port, regs(1859) => 
                           bus_reg_dataout_1859_port, regs(1858) => 
                           bus_reg_dataout_1858_port, regs(1857) => 
                           bus_reg_dataout_1857_port, regs(1856) => 
                           bus_reg_dataout_1856_port, regs(1855) => 
                           bus_reg_dataout_1855_port, regs(1854) => 
                           bus_reg_dataout_1854_port, regs(1853) => 
                           bus_reg_dataout_1853_port, regs(1852) => 
                           bus_reg_dataout_1852_port, regs(1851) => 
                           bus_reg_dataout_1851_port, regs(1850) => 
                           bus_reg_dataout_1850_port, regs(1849) => 
                           bus_reg_dataout_1849_port, regs(1848) => 
                           bus_reg_dataout_1848_port, regs(1847) => 
                           bus_reg_dataout_1847_port, regs(1846) => 
                           bus_reg_dataout_1846_port, regs(1845) => 
                           bus_reg_dataout_1845_port, regs(1844) => 
                           bus_reg_dataout_1844_port, regs(1843) => 
                           bus_reg_dataout_1843_port, regs(1842) => 
                           bus_reg_dataout_1842_port, regs(1841) => 
                           bus_reg_dataout_1841_port, regs(1840) => 
                           bus_reg_dataout_1840_port, regs(1839) => 
                           bus_reg_dataout_1839_port, regs(1838) => 
                           bus_reg_dataout_1838_port, regs(1837) => 
                           bus_reg_dataout_1837_port, regs(1836) => 
                           bus_reg_dataout_1836_port, regs(1835) => 
                           bus_reg_dataout_1835_port, regs(1834) => 
                           bus_reg_dataout_1834_port, regs(1833) => 
                           bus_reg_dataout_1833_port, regs(1832) => 
                           bus_reg_dataout_1832_port, regs(1831) => 
                           bus_reg_dataout_1831_port, regs(1830) => 
                           bus_reg_dataout_1830_port, regs(1829) => 
                           bus_reg_dataout_1829_port, regs(1828) => 
                           bus_reg_dataout_1828_port, regs(1827) => 
                           bus_reg_dataout_1827_port, regs(1826) => 
                           bus_reg_dataout_1826_port, regs(1825) => 
                           bus_reg_dataout_1825_port, regs(1824) => 
                           bus_reg_dataout_1824_port, regs(1823) => 
                           bus_reg_dataout_1823_port, regs(1822) => 
                           bus_reg_dataout_1822_port, regs(1821) => 
                           bus_reg_dataout_1821_port, regs(1820) => 
                           bus_reg_dataout_1820_port, regs(1819) => 
                           bus_reg_dataout_1819_port, regs(1818) => 
                           bus_reg_dataout_1818_port, regs(1817) => 
                           bus_reg_dataout_1817_port, regs(1816) => 
                           bus_reg_dataout_1816_port, regs(1815) => 
                           bus_reg_dataout_1815_port, regs(1814) => 
                           bus_reg_dataout_1814_port, regs(1813) => 
                           bus_reg_dataout_1813_port, regs(1812) => 
                           bus_reg_dataout_1812_port, regs(1811) => 
                           bus_reg_dataout_1811_port, regs(1810) => 
                           bus_reg_dataout_1810_port, regs(1809) => 
                           bus_reg_dataout_1809_port, regs(1808) => 
                           bus_reg_dataout_1808_port, regs(1807) => 
                           bus_reg_dataout_1807_port, regs(1806) => 
                           bus_reg_dataout_1806_port, regs(1805) => 
                           bus_reg_dataout_1805_port, regs(1804) => 
                           bus_reg_dataout_1804_port, regs(1803) => 
                           bus_reg_dataout_1803_port, regs(1802) => 
                           bus_reg_dataout_1802_port, regs(1801) => 
                           bus_reg_dataout_1801_port, regs(1800) => 
                           bus_reg_dataout_1800_port, regs(1799) => 
                           bus_reg_dataout_1799_port, regs(1798) => 
                           bus_reg_dataout_1798_port, regs(1797) => 
                           bus_reg_dataout_1797_port, regs(1796) => 
                           bus_reg_dataout_1796_port, regs(1795) => 
                           bus_reg_dataout_1795_port, regs(1794) => 
                           bus_reg_dataout_1794_port, regs(1793) => 
                           bus_reg_dataout_1793_port, regs(1792) => 
                           bus_reg_dataout_1792_port, regs(1791) => 
                           bus_reg_dataout_1791_port, regs(1790) => 
                           bus_reg_dataout_1790_port, regs(1789) => 
                           bus_reg_dataout_1789_port, regs(1788) => 
                           bus_reg_dataout_1788_port, regs(1787) => 
                           bus_reg_dataout_1787_port, regs(1786) => 
                           bus_reg_dataout_1786_port, regs(1785) => 
                           bus_reg_dataout_1785_port, regs(1784) => 
                           bus_reg_dataout_1784_port, regs(1783) => 
                           bus_reg_dataout_1783_port, regs(1782) => 
                           bus_reg_dataout_1782_port, regs(1781) => 
                           bus_reg_dataout_1781_port, regs(1780) => 
                           bus_reg_dataout_1780_port, regs(1779) => 
                           bus_reg_dataout_1779_port, regs(1778) => 
                           bus_reg_dataout_1778_port, regs(1777) => 
                           bus_reg_dataout_1777_port, regs(1776) => 
                           bus_reg_dataout_1776_port, regs(1775) => 
                           bus_reg_dataout_1775_port, regs(1774) => 
                           bus_reg_dataout_1774_port, regs(1773) => 
                           bus_reg_dataout_1773_port, regs(1772) => 
                           bus_reg_dataout_1772_port, regs(1771) => 
                           bus_reg_dataout_1771_port, regs(1770) => 
                           bus_reg_dataout_1770_port, regs(1769) => 
                           bus_reg_dataout_1769_port, regs(1768) => 
                           bus_reg_dataout_1768_port, regs(1767) => 
                           bus_reg_dataout_1767_port, regs(1766) => 
                           bus_reg_dataout_1766_port, regs(1765) => 
                           bus_reg_dataout_1765_port, regs(1764) => 
                           bus_reg_dataout_1764_port, regs(1763) => 
                           bus_reg_dataout_1763_port, regs(1762) => 
                           bus_reg_dataout_1762_port, regs(1761) => 
                           bus_reg_dataout_1761_port, regs(1760) => 
                           bus_reg_dataout_1760_port, regs(1759) => 
                           bus_reg_dataout_1759_port, regs(1758) => 
                           bus_reg_dataout_1758_port, regs(1757) => 
                           bus_reg_dataout_1757_port, regs(1756) => 
                           bus_reg_dataout_1756_port, regs(1755) => 
                           bus_reg_dataout_1755_port, regs(1754) => 
                           bus_reg_dataout_1754_port, regs(1753) => 
                           bus_reg_dataout_1753_port, regs(1752) => 
                           bus_reg_dataout_1752_port, regs(1751) => 
                           bus_reg_dataout_1751_port, regs(1750) => 
                           bus_reg_dataout_1750_port, regs(1749) => 
                           bus_reg_dataout_1749_port, regs(1748) => 
                           bus_reg_dataout_1748_port, regs(1747) => 
                           bus_reg_dataout_1747_port, regs(1746) => 
                           bus_reg_dataout_1746_port, regs(1745) => 
                           bus_reg_dataout_1745_port, regs(1744) => 
                           bus_reg_dataout_1744_port, regs(1743) => 
                           bus_reg_dataout_1743_port, regs(1742) => 
                           bus_reg_dataout_1742_port, regs(1741) => 
                           bus_reg_dataout_1741_port, regs(1740) => 
                           bus_reg_dataout_1740_port, regs(1739) => 
                           bus_reg_dataout_1739_port, regs(1738) => 
                           bus_reg_dataout_1738_port, regs(1737) => 
                           bus_reg_dataout_1737_port, regs(1736) => 
                           bus_reg_dataout_1736_port, regs(1735) => 
                           bus_reg_dataout_1735_port, regs(1734) => 
                           bus_reg_dataout_1734_port, regs(1733) => 
                           bus_reg_dataout_1733_port, regs(1732) => 
                           bus_reg_dataout_1732_port, regs(1731) => 
                           bus_reg_dataout_1731_port, regs(1730) => 
                           bus_reg_dataout_1730_port, regs(1729) => 
                           bus_reg_dataout_1729_port, regs(1728) => 
                           bus_reg_dataout_1728_port, regs(1727) => 
                           bus_reg_dataout_1727_port, regs(1726) => 
                           bus_reg_dataout_1726_port, regs(1725) => 
                           bus_reg_dataout_1725_port, regs(1724) => 
                           bus_reg_dataout_1724_port, regs(1723) => 
                           bus_reg_dataout_1723_port, regs(1722) => 
                           bus_reg_dataout_1722_port, regs(1721) => 
                           bus_reg_dataout_1721_port, regs(1720) => 
                           bus_reg_dataout_1720_port, regs(1719) => 
                           bus_reg_dataout_1719_port, regs(1718) => 
                           bus_reg_dataout_1718_port, regs(1717) => 
                           bus_reg_dataout_1717_port, regs(1716) => 
                           bus_reg_dataout_1716_port, regs(1715) => 
                           bus_reg_dataout_1715_port, regs(1714) => 
                           bus_reg_dataout_1714_port, regs(1713) => 
                           bus_reg_dataout_1713_port, regs(1712) => 
                           bus_reg_dataout_1712_port, regs(1711) => 
                           bus_reg_dataout_1711_port, regs(1710) => 
                           bus_reg_dataout_1710_port, regs(1709) => 
                           bus_reg_dataout_1709_port, regs(1708) => 
                           bus_reg_dataout_1708_port, regs(1707) => 
                           bus_reg_dataout_1707_port, regs(1706) => 
                           bus_reg_dataout_1706_port, regs(1705) => 
                           bus_reg_dataout_1705_port, regs(1704) => 
                           bus_reg_dataout_1704_port, regs(1703) => 
                           bus_reg_dataout_1703_port, regs(1702) => 
                           bus_reg_dataout_1702_port, regs(1701) => 
                           bus_reg_dataout_1701_port, regs(1700) => 
                           bus_reg_dataout_1700_port, regs(1699) => 
                           bus_reg_dataout_1699_port, regs(1698) => 
                           bus_reg_dataout_1698_port, regs(1697) => 
                           bus_reg_dataout_1697_port, regs(1696) => 
                           bus_reg_dataout_1696_port, regs(1695) => 
                           bus_reg_dataout_1695_port, regs(1694) => 
                           bus_reg_dataout_1694_port, regs(1693) => 
                           bus_reg_dataout_1693_port, regs(1692) => 
                           bus_reg_dataout_1692_port, regs(1691) => 
                           bus_reg_dataout_1691_port, regs(1690) => 
                           bus_reg_dataout_1690_port, regs(1689) => 
                           bus_reg_dataout_1689_port, regs(1688) => 
                           bus_reg_dataout_1688_port, regs(1687) => 
                           bus_reg_dataout_1687_port, regs(1686) => 
                           bus_reg_dataout_1686_port, regs(1685) => 
                           bus_reg_dataout_1685_port, regs(1684) => 
                           bus_reg_dataout_1684_port, regs(1683) => 
                           bus_reg_dataout_1683_port, regs(1682) => 
                           bus_reg_dataout_1682_port, regs(1681) => 
                           bus_reg_dataout_1681_port, regs(1680) => 
                           bus_reg_dataout_1680_port, regs(1679) => 
                           bus_reg_dataout_1679_port, regs(1678) => 
                           bus_reg_dataout_1678_port, regs(1677) => 
                           bus_reg_dataout_1677_port, regs(1676) => 
                           bus_reg_dataout_1676_port, regs(1675) => 
                           bus_reg_dataout_1675_port, regs(1674) => 
                           bus_reg_dataout_1674_port, regs(1673) => 
                           bus_reg_dataout_1673_port, regs(1672) => 
                           bus_reg_dataout_1672_port, regs(1671) => 
                           bus_reg_dataout_1671_port, regs(1670) => 
                           bus_reg_dataout_1670_port, regs(1669) => 
                           bus_reg_dataout_1669_port, regs(1668) => 
                           bus_reg_dataout_1668_port, regs(1667) => 
                           bus_reg_dataout_1667_port, regs(1666) => 
                           bus_reg_dataout_1666_port, regs(1665) => 
                           bus_reg_dataout_1665_port, regs(1664) => 
                           bus_reg_dataout_1664_port, regs(1663) => 
                           bus_reg_dataout_1663_port, regs(1662) => 
                           bus_reg_dataout_1662_port, regs(1661) => 
                           bus_reg_dataout_1661_port, regs(1660) => 
                           bus_reg_dataout_1660_port, regs(1659) => 
                           bus_reg_dataout_1659_port, regs(1658) => 
                           bus_reg_dataout_1658_port, regs(1657) => 
                           bus_reg_dataout_1657_port, regs(1656) => 
                           bus_reg_dataout_1656_port, regs(1655) => 
                           bus_reg_dataout_1655_port, regs(1654) => 
                           bus_reg_dataout_1654_port, regs(1653) => 
                           bus_reg_dataout_1653_port, regs(1652) => 
                           bus_reg_dataout_1652_port, regs(1651) => 
                           bus_reg_dataout_1651_port, regs(1650) => 
                           bus_reg_dataout_1650_port, regs(1649) => 
                           bus_reg_dataout_1649_port, regs(1648) => 
                           bus_reg_dataout_1648_port, regs(1647) => 
                           bus_reg_dataout_1647_port, regs(1646) => 
                           bus_reg_dataout_1646_port, regs(1645) => 
                           bus_reg_dataout_1645_port, regs(1644) => 
                           bus_reg_dataout_1644_port, regs(1643) => 
                           bus_reg_dataout_1643_port, regs(1642) => 
                           bus_reg_dataout_1642_port, regs(1641) => 
                           bus_reg_dataout_1641_port, regs(1640) => 
                           bus_reg_dataout_1640_port, regs(1639) => 
                           bus_reg_dataout_1639_port, regs(1638) => 
                           bus_reg_dataout_1638_port, regs(1637) => 
                           bus_reg_dataout_1637_port, regs(1636) => 
                           bus_reg_dataout_1636_port, regs(1635) => 
                           bus_reg_dataout_1635_port, regs(1634) => 
                           bus_reg_dataout_1634_port, regs(1633) => 
                           bus_reg_dataout_1633_port, regs(1632) => 
                           bus_reg_dataout_1632_port, regs(1631) => 
                           bus_reg_dataout_1631_port, regs(1630) => 
                           bus_reg_dataout_1630_port, regs(1629) => 
                           bus_reg_dataout_1629_port, regs(1628) => 
                           bus_reg_dataout_1628_port, regs(1627) => 
                           bus_reg_dataout_1627_port, regs(1626) => 
                           bus_reg_dataout_1626_port, regs(1625) => 
                           bus_reg_dataout_1625_port, regs(1624) => 
                           bus_reg_dataout_1624_port, regs(1623) => 
                           bus_reg_dataout_1623_port, regs(1622) => 
                           bus_reg_dataout_1622_port, regs(1621) => 
                           bus_reg_dataout_1621_port, regs(1620) => 
                           bus_reg_dataout_1620_port, regs(1619) => 
                           bus_reg_dataout_1619_port, regs(1618) => 
                           bus_reg_dataout_1618_port, regs(1617) => 
                           bus_reg_dataout_1617_port, regs(1616) => 
                           bus_reg_dataout_1616_port, regs(1615) => 
                           bus_reg_dataout_1615_port, regs(1614) => 
                           bus_reg_dataout_1614_port, regs(1613) => 
                           bus_reg_dataout_1613_port, regs(1612) => 
                           bus_reg_dataout_1612_port, regs(1611) => 
                           bus_reg_dataout_1611_port, regs(1610) => 
                           bus_reg_dataout_1610_port, regs(1609) => 
                           bus_reg_dataout_1609_port, regs(1608) => 
                           bus_reg_dataout_1608_port, regs(1607) => 
                           bus_reg_dataout_1607_port, regs(1606) => 
                           bus_reg_dataout_1606_port, regs(1605) => 
                           bus_reg_dataout_1605_port, regs(1604) => 
                           bus_reg_dataout_1604_port, regs(1603) => 
                           bus_reg_dataout_1603_port, regs(1602) => 
                           bus_reg_dataout_1602_port, regs(1601) => 
                           bus_reg_dataout_1601_port, regs(1600) => 
                           bus_reg_dataout_1600_port, regs(1599) => 
                           bus_reg_dataout_1599_port, regs(1598) => 
                           bus_reg_dataout_1598_port, regs(1597) => 
                           bus_reg_dataout_1597_port, regs(1596) => 
                           bus_reg_dataout_1596_port, regs(1595) => 
                           bus_reg_dataout_1595_port, regs(1594) => 
                           bus_reg_dataout_1594_port, regs(1593) => 
                           bus_reg_dataout_1593_port, regs(1592) => 
                           bus_reg_dataout_1592_port, regs(1591) => 
                           bus_reg_dataout_1591_port, regs(1590) => 
                           bus_reg_dataout_1590_port, regs(1589) => 
                           bus_reg_dataout_1589_port, regs(1588) => 
                           bus_reg_dataout_1588_port, regs(1587) => 
                           bus_reg_dataout_1587_port, regs(1586) => 
                           bus_reg_dataout_1586_port, regs(1585) => 
                           bus_reg_dataout_1585_port, regs(1584) => 
                           bus_reg_dataout_1584_port, regs(1583) => 
                           bus_reg_dataout_1583_port, regs(1582) => 
                           bus_reg_dataout_1582_port, regs(1581) => 
                           bus_reg_dataout_1581_port, regs(1580) => 
                           bus_reg_dataout_1580_port, regs(1579) => 
                           bus_reg_dataout_1579_port, regs(1578) => 
                           bus_reg_dataout_1578_port, regs(1577) => 
                           bus_reg_dataout_1577_port, regs(1576) => 
                           bus_reg_dataout_1576_port, regs(1575) => 
                           bus_reg_dataout_1575_port, regs(1574) => 
                           bus_reg_dataout_1574_port, regs(1573) => 
                           bus_reg_dataout_1573_port, regs(1572) => 
                           bus_reg_dataout_1572_port, regs(1571) => 
                           bus_reg_dataout_1571_port, regs(1570) => 
                           bus_reg_dataout_1570_port, regs(1569) => 
                           bus_reg_dataout_1569_port, regs(1568) => 
                           bus_reg_dataout_1568_port, regs(1567) => 
                           bus_reg_dataout_1567_port, regs(1566) => 
                           bus_reg_dataout_1566_port, regs(1565) => 
                           bus_reg_dataout_1565_port, regs(1564) => 
                           bus_reg_dataout_1564_port, regs(1563) => 
                           bus_reg_dataout_1563_port, regs(1562) => 
                           bus_reg_dataout_1562_port, regs(1561) => 
                           bus_reg_dataout_1561_port, regs(1560) => 
                           bus_reg_dataout_1560_port, regs(1559) => 
                           bus_reg_dataout_1559_port, regs(1558) => 
                           bus_reg_dataout_1558_port, regs(1557) => 
                           bus_reg_dataout_1557_port, regs(1556) => 
                           bus_reg_dataout_1556_port, regs(1555) => 
                           bus_reg_dataout_1555_port, regs(1554) => 
                           bus_reg_dataout_1554_port, regs(1553) => 
                           bus_reg_dataout_1553_port, regs(1552) => 
                           bus_reg_dataout_1552_port, regs(1551) => 
                           bus_reg_dataout_1551_port, regs(1550) => 
                           bus_reg_dataout_1550_port, regs(1549) => 
                           bus_reg_dataout_1549_port, regs(1548) => 
                           bus_reg_dataout_1548_port, regs(1547) => 
                           bus_reg_dataout_1547_port, regs(1546) => 
                           bus_reg_dataout_1546_port, regs(1545) => 
                           bus_reg_dataout_1545_port, regs(1544) => 
                           bus_reg_dataout_1544_port, regs(1543) => 
                           bus_reg_dataout_1543_port, regs(1542) => 
                           bus_reg_dataout_1542_port, regs(1541) => 
                           bus_reg_dataout_1541_port, regs(1540) => 
                           bus_reg_dataout_1540_port, regs(1539) => 
                           bus_reg_dataout_1539_port, regs(1538) => 
                           bus_reg_dataout_1538_port, regs(1537) => 
                           bus_reg_dataout_1537_port, regs(1536) => 
                           bus_reg_dataout_1536_port, regs(1535) => 
                           bus_reg_dataout_1535_port, regs(1534) => 
                           bus_reg_dataout_1534_port, regs(1533) => 
                           bus_reg_dataout_1533_port, regs(1532) => 
                           bus_reg_dataout_1532_port, regs(1531) => 
                           bus_reg_dataout_1531_port, regs(1530) => 
                           bus_reg_dataout_1530_port, regs(1529) => 
                           bus_reg_dataout_1529_port, regs(1528) => 
                           bus_reg_dataout_1528_port, regs(1527) => 
                           bus_reg_dataout_1527_port, regs(1526) => 
                           bus_reg_dataout_1526_port, regs(1525) => 
                           bus_reg_dataout_1525_port, regs(1524) => 
                           bus_reg_dataout_1524_port, regs(1523) => 
                           bus_reg_dataout_1523_port, regs(1522) => 
                           bus_reg_dataout_1522_port, regs(1521) => 
                           bus_reg_dataout_1521_port, regs(1520) => 
                           bus_reg_dataout_1520_port, regs(1519) => 
                           bus_reg_dataout_1519_port, regs(1518) => 
                           bus_reg_dataout_1518_port, regs(1517) => 
                           bus_reg_dataout_1517_port, regs(1516) => 
                           bus_reg_dataout_1516_port, regs(1515) => 
                           bus_reg_dataout_1515_port, regs(1514) => 
                           bus_reg_dataout_1514_port, regs(1513) => 
                           bus_reg_dataout_1513_port, regs(1512) => 
                           bus_reg_dataout_1512_port, regs(1511) => 
                           bus_reg_dataout_1511_port, regs(1510) => 
                           bus_reg_dataout_1510_port, regs(1509) => 
                           bus_reg_dataout_1509_port, regs(1508) => 
                           bus_reg_dataout_1508_port, regs(1507) => 
                           bus_reg_dataout_1507_port, regs(1506) => 
                           bus_reg_dataout_1506_port, regs(1505) => 
                           bus_reg_dataout_1505_port, regs(1504) => 
                           bus_reg_dataout_1504_port, regs(1503) => 
                           bus_reg_dataout_1503_port, regs(1502) => 
                           bus_reg_dataout_1502_port, regs(1501) => 
                           bus_reg_dataout_1501_port, regs(1500) => 
                           bus_reg_dataout_1500_port, regs(1499) => 
                           bus_reg_dataout_1499_port, regs(1498) => 
                           bus_reg_dataout_1498_port, regs(1497) => 
                           bus_reg_dataout_1497_port, regs(1496) => 
                           bus_reg_dataout_1496_port, regs(1495) => 
                           bus_reg_dataout_1495_port, regs(1494) => 
                           bus_reg_dataout_1494_port, regs(1493) => 
                           bus_reg_dataout_1493_port, regs(1492) => 
                           bus_reg_dataout_1492_port, regs(1491) => 
                           bus_reg_dataout_1491_port, regs(1490) => 
                           bus_reg_dataout_1490_port, regs(1489) => 
                           bus_reg_dataout_1489_port, regs(1488) => 
                           bus_reg_dataout_1488_port, regs(1487) => 
                           bus_reg_dataout_1487_port, regs(1486) => 
                           bus_reg_dataout_1486_port, regs(1485) => 
                           bus_reg_dataout_1485_port, regs(1484) => 
                           bus_reg_dataout_1484_port, regs(1483) => 
                           bus_reg_dataout_1483_port, regs(1482) => 
                           bus_reg_dataout_1482_port, regs(1481) => 
                           bus_reg_dataout_1481_port, regs(1480) => 
                           bus_reg_dataout_1480_port, regs(1479) => 
                           bus_reg_dataout_1479_port, regs(1478) => 
                           bus_reg_dataout_1478_port, regs(1477) => 
                           bus_reg_dataout_1477_port, regs(1476) => 
                           bus_reg_dataout_1476_port, regs(1475) => 
                           bus_reg_dataout_1475_port, regs(1474) => 
                           bus_reg_dataout_1474_port, regs(1473) => 
                           bus_reg_dataout_1473_port, regs(1472) => 
                           bus_reg_dataout_1472_port, regs(1471) => 
                           bus_reg_dataout_1471_port, regs(1470) => 
                           bus_reg_dataout_1470_port, regs(1469) => 
                           bus_reg_dataout_1469_port, regs(1468) => 
                           bus_reg_dataout_1468_port, regs(1467) => 
                           bus_reg_dataout_1467_port, regs(1466) => 
                           bus_reg_dataout_1466_port, regs(1465) => 
                           bus_reg_dataout_1465_port, regs(1464) => 
                           bus_reg_dataout_1464_port, regs(1463) => 
                           bus_reg_dataout_1463_port, regs(1462) => 
                           bus_reg_dataout_1462_port, regs(1461) => 
                           bus_reg_dataout_1461_port, regs(1460) => 
                           bus_reg_dataout_1460_port, regs(1459) => 
                           bus_reg_dataout_1459_port, regs(1458) => 
                           bus_reg_dataout_1458_port, regs(1457) => 
                           bus_reg_dataout_1457_port, regs(1456) => 
                           bus_reg_dataout_1456_port, regs(1455) => 
                           bus_reg_dataout_1455_port, regs(1454) => 
                           bus_reg_dataout_1454_port, regs(1453) => 
                           bus_reg_dataout_1453_port, regs(1452) => 
                           bus_reg_dataout_1452_port, regs(1451) => 
                           bus_reg_dataout_1451_port, regs(1450) => 
                           bus_reg_dataout_1450_port, regs(1449) => 
                           bus_reg_dataout_1449_port, regs(1448) => 
                           bus_reg_dataout_1448_port, regs(1447) => 
                           bus_reg_dataout_1447_port, regs(1446) => 
                           bus_reg_dataout_1446_port, regs(1445) => 
                           bus_reg_dataout_1445_port, regs(1444) => 
                           bus_reg_dataout_1444_port, regs(1443) => 
                           bus_reg_dataout_1443_port, regs(1442) => 
                           bus_reg_dataout_1442_port, regs(1441) => 
                           bus_reg_dataout_1441_port, regs(1440) => 
                           bus_reg_dataout_1440_port, regs(1439) => 
                           bus_reg_dataout_1439_port, regs(1438) => 
                           bus_reg_dataout_1438_port, regs(1437) => 
                           bus_reg_dataout_1437_port, regs(1436) => 
                           bus_reg_dataout_1436_port, regs(1435) => 
                           bus_reg_dataout_1435_port, regs(1434) => 
                           bus_reg_dataout_1434_port, regs(1433) => 
                           bus_reg_dataout_1433_port, regs(1432) => 
                           bus_reg_dataout_1432_port, regs(1431) => 
                           bus_reg_dataout_1431_port, regs(1430) => 
                           bus_reg_dataout_1430_port, regs(1429) => 
                           bus_reg_dataout_1429_port, regs(1428) => 
                           bus_reg_dataout_1428_port, regs(1427) => 
                           bus_reg_dataout_1427_port, regs(1426) => 
                           bus_reg_dataout_1426_port, regs(1425) => 
                           bus_reg_dataout_1425_port, regs(1424) => 
                           bus_reg_dataout_1424_port, regs(1423) => 
                           bus_reg_dataout_1423_port, regs(1422) => 
                           bus_reg_dataout_1422_port, regs(1421) => 
                           bus_reg_dataout_1421_port, regs(1420) => 
                           bus_reg_dataout_1420_port, regs(1419) => 
                           bus_reg_dataout_1419_port, regs(1418) => 
                           bus_reg_dataout_1418_port, regs(1417) => 
                           bus_reg_dataout_1417_port, regs(1416) => 
                           bus_reg_dataout_1416_port, regs(1415) => 
                           bus_reg_dataout_1415_port, regs(1414) => 
                           bus_reg_dataout_1414_port, regs(1413) => 
                           bus_reg_dataout_1413_port, regs(1412) => 
                           bus_reg_dataout_1412_port, regs(1411) => 
                           bus_reg_dataout_1411_port, regs(1410) => 
                           bus_reg_dataout_1410_port, regs(1409) => 
                           bus_reg_dataout_1409_port, regs(1408) => 
                           bus_reg_dataout_1408_port, regs(1407) => 
                           bus_reg_dataout_1407_port, regs(1406) => 
                           bus_reg_dataout_1406_port, regs(1405) => 
                           bus_reg_dataout_1405_port, regs(1404) => 
                           bus_reg_dataout_1404_port, regs(1403) => 
                           bus_reg_dataout_1403_port, regs(1402) => 
                           bus_reg_dataout_1402_port, regs(1401) => 
                           bus_reg_dataout_1401_port, regs(1400) => 
                           bus_reg_dataout_1400_port, regs(1399) => 
                           bus_reg_dataout_1399_port, regs(1398) => 
                           bus_reg_dataout_1398_port, regs(1397) => 
                           bus_reg_dataout_1397_port, regs(1396) => 
                           bus_reg_dataout_1396_port, regs(1395) => 
                           bus_reg_dataout_1395_port, regs(1394) => 
                           bus_reg_dataout_1394_port, regs(1393) => 
                           bus_reg_dataout_1393_port, regs(1392) => 
                           bus_reg_dataout_1392_port, regs(1391) => 
                           bus_reg_dataout_1391_port, regs(1390) => 
                           bus_reg_dataout_1390_port, regs(1389) => 
                           bus_reg_dataout_1389_port, regs(1388) => 
                           bus_reg_dataout_1388_port, regs(1387) => 
                           bus_reg_dataout_1387_port, regs(1386) => 
                           bus_reg_dataout_1386_port, regs(1385) => 
                           bus_reg_dataout_1385_port, regs(1384) => 
                           bus_reg_dataout_1384_port, regs(1383) => 
                           bus_reg_dataout_1383_port, regs(1382) => 
                           bus_reg_dataout_1382_port, regs(1381) => 
                           bus_reg_dataout_1381_port, regs(1380) => 
                           bus_reg_dataout_1380_port, regs(1379) => 
                           bus_reg_dataout_1379_port, regs(1378) => 
                           bus_reg_dataout_1378_port, regs(1377) => 
                           bus_reg_dataout_1377_port, regs(1376) => 
                           bus_reg_dataout_1376_port, regs(1375) => 
                           bus_reg_dataout_1375_port, regs(1374) => 
                           bus_reg_dataout_1374_port, regs(1373) => 
                           bus_reg_dataout_1373_port, regs(1372) => 
                           bus_reg_dataout_1372_port, regs(1371) => 
                           bus_reg_dataout_1371_port, regs(1370) => 
                           bus_reg_dataout_1370_port, regs(1369) => 
                           bus_reg_dataout_1369_port, regs(1368) => 
                           bus_reg_dataout_1368_port, regs(1367) => 
                           bus_reg_dataout_1367_port, regs(1366) => 
                           bus_reg_dataout_1366_port, regs(1365) => 
                           bus_reg_dataout_1365_port, regs(1364) => 
                           bus_reg_dataout_1364_port, regs(1363) => 
                           bus_reg_dataout_1363_port, regs(1362) => 
                           bus_reg_dataout_1362_port, regs(1361) => 
                           bus_reg_dataout_1361_port, regs(1360) => 
                           bus_reg_dataout_1360_port, regs(1359) => 
                           bus_reg_dataout_1359_port, regs(1358) => 
                           bus_reg_dataout_1358_port, regs(1357) => 
                           bus_reg_dataout_1357_port, regs(1356) => 
                           bus_reg_dataout_1356_port, regs(1355) => 
                           bus_reg_dataout_1355_port, regs(1354) => 
                           bus_reg_dataout_1354_port, regs(1353) => 
                           bus_reg_dataout_1353_port, regs(1352) => 
                           bus_reg_dataout_1352_port, regs(1351) => 
                           bus_reg_dataout_1351_port, regs(1350) => 
                           bus_reg_dataout_1350_port, regs(1349) => 
                           bus_reg_dataout_1349_port, regs(1348) => 
                           bus_reg_dataout_1348_port, regs(1347) => 
                           bus_reg_dataout_1347_port, regs(1346) => 
                           bus_reg_dataout_1346_port, regs(1345) => 
                           bus_reg_dataout_1345_port, regs(1344) => 
                           bus_reg_dataout_1344_port, regs(1343) => 
                           bus_reg_dataout_1343_port, regs(1342) => 
                           bus_reg_dataout_1342_port, regs(1341) => 
                           bus_reg_dataout_1341_port, regs(1340) => 
                           bus_reg_dataout_1340_port, regs(1339) => 
                           bus_reg_dataout_1339_port, regs(1338) => 
                           bus_reg_dataout_1338_port, regs(1337) => 
                           bus_reg_dataout_1337_port, regs(1336) => 
                           bus_reg_dataout_1336_port, regs(1335) => 
                           bus_reg_dataout_1335_port, regs(1334) => 
                           bus_reg_dataout_1334_port, regs(1333) => 
                           bus_reg_dataout_1333_port, regs(1332) => 
                           bus_reg_dataout_1332_port, regs(1331) => 
                           bus_reg_dataout_1331_port, regs(1330) => 
                           bus_reg_dataout_1330_port, regs(1329) => 
                           bus_reg_dataout_1329_port, regs(1328) => 
                           bus_reg_dataout_1328_port, regs(1327) => 
                           bus_reg_dataout_1327_port, regs(1326) => 
                           bus_reg_dataout_1326_port, regs(1325) => 
                           bus_reg_dataout_1325_port, regs(1324) => 
                           bus_reg_dataout_1324_port, regs(1323) => 
                           bus_reg_dataout_1323_port, regs(1322) => 
                           bus_reg_dataout_1322_port, regs(1321) => 
                           bus_reg_dataout_1321_port, regs(1320) => 
                           bus_reg_dataout_1320_port, regs(1319) => 
                           bus_reg_dataout_1319_port, regs(1318) => 
                           bus_reg_dataout_1318_port, regs(1317) => 
                           bus_reg_dataout_1317_port, regs(1316) => 
                           bus_reg_dataout_1316_port, regs(1315) => 
                           bus_reg_dataout_1315_port, regs(1314) => 
                           bus_reg_dataout_1314_port, regs(1313) => 
                           bus_reg_dataout_1313_port, regs(1312) => 
                           bus_reg_dataout_1312_port, regs(1311) => 
                           bus_reg_dataout_1311_port, regs(1310) => 
                           bus_reg_dataout_1310_port, regs(1309) => 
                           bus_reg_dataout_1309_port, regs(1308) => 
                           bus_reg_dataout_1308_port, regs(1307) => 
                           bus_reg_dataout_1307_port, regs(1306) => 
                           bus_reg_dataout_1306_port, regs(1305) => 
                           bus_reg_dataout_1305_port, regs(1304) => 
                           bus_reg_dataout_1304_port, regs(1303) => 
                           bus_reg_dataout_1303_port, regs(1302) => 
                           bus_reg_dataout_1302_port, regs(1301) => 
                           bus_reg_dataout_1301_port, regs(1300) => 
                           bus_reg_dataout_1300_port, regs(1299) => 
                           bus_reg_dataout_1299_port, regs(1298) => 
                           bus_reg_dataout_1298_port, regs(1297) => 
                           bus_reg_dataout_1297_port, regs(1296) => 
                           bus_reg_dataout_1296_port, regs(1295) => 
                           bus_reg_dataout_1295_port, regs(1294) => 
                           bus_reg_dataout_1294_port, regs(1293) => 
                           bus_reg_dataout_1293_port, regs(1292) => 
                           bus_reg_dataout_1292_port, regs(1291) => 
                           bus_reg_dataout_1291_port, regs(1290) => 
                           bus_reg_dataout_1290_port, regs(1289) => 
                           bus_reg_dataout_1289_port, regs(1288) => 
                           bus_reg_dataout_1288_port, regs(1287) => 
                           bus_reg_dataout_1287_port, regs(1286) => 
                           bus_reg_dataout_1286_port, regs(1285) => 
                           bus_reg_dataout_1285_port, regs(1284) => 
                           bus_reg_dataout_1284_port, regs(1283) => 
                           bus_reg_dataout_1283_port, regs(1282) => 
                           bus_reg_dataout_1282_port, regs(1281) => 
                           bus_reg_dataout_1281_port, regs(1280) => 
                           bus_reg_dataout_1280_port, regs(1279) => 
                           bus_reg_dataout_1279_port, regs(1278) => 
                           bus_reg_dataout_1278_port, regs(1277) => 
                           bus_reg_dataout_1277_port, regs(1276) => 
                           bus_reg_dataout_1276_port, regs(1275) => 
                           bus_reg_dataout_1275_port, regs(1274) => 
                           bus_reg_dataout_1274_port, regs(1273) => 
                           bus_reg_dataout_1273_port, regs(1272) => 
                           bus_reg_dataout_1272_port, regs(1271) => 
                           bus_reg_dataout_1271_port, regs(1270) => 
                           bus_reg_dataout_1270_port, regs(1269) => 
                           bus_reg_dataout_1269_port, regs(1268) => 
                           bus_reg_dataout_1268_port, regs(1267) => 
                           bus_reg_dataout_1267_port, regs(1266) => 
                           bus_reg_dataout_1266_port, regs(1265) => 
                           bus_reg_dataout_1265_port, regs(1264) => 
                           bus_reg_dataout_1264_port, regs(1263) => 
                           bus_reg_dataout_1263_port, regs(1262) => 
                           bus_reg_dataout_1262_port, regs(1261) => 
                           bus_reg_dataout_1261_port, regs(1260) => 
                           bus_reg_dataout_1260_port, regs(1259) => 
                           bus_reg_dataout_1259_port, regs(1258) => 
                           bus_reg_dataout_1258_port, regs(1257) => 
                           bus_reg_dataout_1257_port, regs(1256) => 
                           bus_reg_dataout_1256_port, regs(1255) => 
                           bus_reg_dataout_1255_port, regs(1254) => 
                           bus_reg_dataout_1254_port, regs(1253) => 
                           bus_reg_dataout_1253_port, regs(1252) => 
                           bus_reg_dataout_1252_port, regs(1251) => 
                           bus_reg_dataout_1251_port, regs(1250) => 
                           bus_reg_dataout_1250_port, regs(1249) => 
                           bus_reg_dataout_1249_port, regs(1248) => 
                           bus_reg_dataout_1248_port, regs(1247) => 
                           bus_reg_dataout_1247_port, regs(1246) => 
                           bus_reg_dataout_1246_port, regs(1245) => 
                           bus_reg_dataout_1245_port, regs(1244) => 
                           bus_reg_dataout_1244_port, regs(1243) => 
                           bus_reg_dataout_1243_port, regs(1242) => 
                           bus_reg_dataout_1242_port, regs(1241) => 
                           bus_reg_dataout_1241_port, regs(1240) => 
                           bus_reg_dataout_1240_port, regs(1239) => 
                           bus_reg_dataout_1239_port, regs(1238) => 
                           bus_reg_dataout_1238_port, regs(1237) => 
                           bus_reg_dataout_1237_port, regs(1236) => 
                           bus_reg_dataout_1236_port, regs(1235) => 
                           bus_reg_dataout_1235_port, regs(1234) => 
                           bus_reg_dataout_1234_port, regs(1233) => 
                           bus_reg_dataout_1233_port, regs(1232) => 
                           bus_reg_dataout_1232_port, regs(1231) => 
                           bus_reg_dataout_1231_port, regs(1230) => 
                           bus_reg_dataout_1230_port, regs(1229) => 
                           bus_reg_dataout_1229_port, regs(1228) => 
                           bus_reg_dataout_1228_port, regs(1227) => 
                           bus_reg_dataout_1227_port, regs(1226) => 
                           bus_reg_dataout_1226_port, regs(1225) => 
                           bus_reg_dataout_1225_port, regs(1224) => 
                           bus_reg_dataout_1224_port, regs(1223) => 
                           bus_reg_dataout_1223_port, regs(1222) => 
                           bus_reg_dataout_1222_port, regs(1221) => 
                           bus_reg_dataout_1221_port, regs(1220) => 
                           bus_reg_dataout_1220_port, regs(1219) => 
                           bus_reg_dataout_1219_port, regs(1218) => 
                           bus_reg_dataout_1218_port, regs(1217) => 
                           bus_reg_dataout_1217_port, regs(1216) => 
                           bus_reg_dataout_1216_port, regs(1215) => 
                           bus_reg_dataout_1215_port, regs(1214) => 
                           bus_reg_dataout_1214_port, regs(1213) => 
                           bus_reg_dataout_1213_port, regs(1212) => 
                           bus_reg_dataout_1212_port, regs(1211) => 
                           bus_reg_dataout_1211_port, regs(1210) => 
                           bus_reg_dataout_1210_port, regs(1209) => 
                           bus_reg_dataout_1209_port, regs(1208) => 
                           bus_reg_dataout_1208_port, regs(1207) => 
                           bus_reg_dataout_1207_port, regs(1206) => 
                           bus_reg_dataout_1206_port, regs(1205) => 
                           bus_reg_dataout_1205_port, regs(1204) => 
                           bus_reg_dataout_1204_port, regs(1203) => 
                           bus_reg_dataout_1203_port, regs(1202) => 
                           bus_reg_dataout_1202_port, regs(1201) => 
                           bus_reg_dataout_1201_port, regs(1200) => 
                           bus_reg_dataout_1200_port, regs(1199) => 
                           bus_reg_dataout_1199_port, regs(1198) => 
                           bus_reg_dataout_1198_port, regs(1197) => 
                           bus_reg_dataout_1197_port, regs(1196) => 
                           bus_reg_dataout_1196_port, regs(1195) => 
                           bus_reg_dataout_1195_port, regs(1194) => 
                           bus_reg_dataout_1194_port, regs(1193) => 
                           bus_reg_dataout_1193_port, regs(1192) => 
                           bus_reg_dataout_1192_port, regs(1191) => 
                           bus_reg_dataout_1191_port, regs(1190) => 
                           bus_reg_dataout_1190_port, regs(1189) => 
                           bus_reg_dataout_1189_port, regs(1188) => 
                           bus_reg_dataout_1188_port, regs(1187) => 
                           bus_reg_dataout_1187_port, regs(1186) => 
                           bus_reg_dataout_1186_port, regs(1185) => 
                           bus_reg_dataout_1185_port, regs(1184) => 
                           bus_reg_dataout_1184_port, regs(1183) => 
                           bus_reg_dataout_1183_port, regs(1182) => 
                           bus_reg_dataout_1182_port, regs(1181) => 
                           bus_reg_dataout_1181_port, regs(1180) => 
                           bus_reg_dataout_1180_port, regs(1179) => 
                           bus_reg_dataout_1179_port, regs(1178) => 
                           bus_reg_dataout_1178_port, regs(1177) => 
                           bus_reg_dataout_1177_port, regs(1176) => 
                           bus_reg_dataout_1176_port, regs(1175) => 
                           bus_reg_dataout_1175_port, regs(1174) => 
                           bus_reg_dataout_1174_port, regs(1173) => 
                           bus_reg_dataout_1173_port, regs(1172) => 
                           bus_reg_dataout_1172_port, regs(1171) => 
                           bus_reg_dataout_1171_port, regs(1170) => 
                           bus_reg_dataout_1170_port, regs(1169) => 
                           bus_reg_dataout_1169_port, regs(1168) => 
                           bus_reg_dataout_1168_port, regs(1167) => 
                           bus_reg_dataout_1167_port, regs(1166) => 
                           bus_reg_dataout_1166_port, regs(1165) => 
                           bus_reg_dataout_1165_port, regs(1164) => 
                           bus_reg_dataout_1164_port, regs(1163) => 
                           bus_reg_dataout_1163_port, regs(1162) => 
                           bus_reg_dataout_1162_port, regs(1161) => 
                           bus_reg_dataout_1161_port, regs(1160) => 
                           bus_reg_dataout_1160_port, regs(1159) => 
                           bus_reg_dataout_1159_port, regs(1158) => 
                           bus_reg_dataout_1158_port, regs(1157) => 
                           bus_reg_dataout_1157_port, regs(1156) => 
                           bus_reg_dataout_1156_port, regs(1155) => 
                           bus_reg_dataout_1155_port, regs(1154) => 
                           bus_reg_dataout_1154_port, regs(1153) => 
                           bus_reg_dataout_1153_port, regs(1152) => 
                           bus_reg_dataout_1152_port, regs(1151) => 
                           bus_reg_dataout_1151_port, regs(1150) => 
                           bus_reg_dataout_1150_port, regs(1149) => 
                           bus_reg_dataout_1149_port, regs(1148) => 
                           bus_reg_dataout_1148_port, regs(1147) => 
                           bus_reg_dataout_1147_port, regs(1146) => 
                           bus_reg_dataout_1146_port, regs(1145) => 
                           bus_reg_dataout_1145_port, regs(1144) => 
                           bus_reg_dataout_1144_port, regs(1143) => 
                           bus_reg_dataout_1143_port, regs(1142) => 
                           bus_reg_dataout_1142_port, regs(1141) => 
                           bus_reg_dataout_1141_port, regs(1140) => 
                           bus_reg_dataout_1140_port, regs(1139) => 
                           bus_reg_dataout_1139_port, regs(1138) => 
                           bus_reg_dataout_1138_port, regs(1137) => 
                           bus_reg_dataout_1137_port, regs(1136) => 
                           bus_reg_dataout_1136_port, regs(1135) => 
                           bus_reg_dataout_1135_port, regs(1134) => 
                           bus_reg_dataout_1134_port, regs(1133) => 
                           bus_reg_dataout_1133_port, regs(1132) => 
                           bus_reg_dataout_1132_port, regs(1131) => 
                           bus_reg_dataout_1131_port, regs(1130) => 
                           bus_reg_dataout_1130_port, regs(1129) => 
                           bus_reg_dataout_1129_port, regs(1128) => 
                           bus_reg_dataout_1128_port, regs(1127) => 
                           bus_reg_dataout_1127_port, regs(1126) => 
                           bus_reg_dataout_1126_port, regs(1125) => 
                           bus_reg_dataout_1125_port, regs(1124) => 
                           bus_reg_dataout_1124_port, regs(1123) => 
                           bus_reg_dataout_1123_port, regs(1122) => 
                           bus_reg_dataout_1122_port, regs(1121) => 
                           bus_reg_dataout_1121_port, regs(1120) => 
                           bus_reg_dataout_1120_port, regs(1119) => 
                           bus_reg_dataout_1119_port, regs(1118) => 
                           bus_reg_dataout_1118_port, regs(1117) => 
                           bus_reg_dataout_1117_port, regs(1116) => 
                           bus_reg_dataout_1116_port, regs(1115) => 
                           bus_reg_dataout_1115_port, regs(1114) => 
                           bus_reg_dataout_1114_port, regs(1113) => 
                           bus_reg_dataout_1113_port, regs(1112) => 
                           bus_reg_dataout_1112_port, regs(1111) => 
                           bus_reg_dataout_1111_port, regs(1110) => 
                           bus_reg_dataout_1110_port, regs(1109) => 
                           bus_reg_dataout_1109_port, regs(1108) => 
                           bus_reg_dataout_1108_port, regs(1107) => 
                           bus_reg_dataout_1107_port, regs(1106) => 
                           bus_reg_dataout_1106_port, regs(1105) => 
                           bus_reg_dataout_1105_port, regs(1104) => 
                           bus_reg_dataout_1104_port, regs(1103) => 
                           bus_reg_dataout_1103_port, regs(1102) => 
                           bus_reg_dataout_1102_port, regs(1101) => 
                           bus_reg_dataout_1101_port, regs(1100) => 
                           bus_reg_dataout_1100_port, regs(1099) => 
                           bus_reg_dataout_1099_port, regs(1098) => 
                           bus_reg_dataout_1098_port, regs(1097) => 
                           bus_reg_dataout_1097_port, regs(1096) => 
                           bus_reg_dataout_1096_port, regs(1095) => 
                           bus_reg_dataout_1095_port, regs(1094) => 
                           bus_reg_dataout_1094_port, regs(1093) => 
                           bus_reg_dataout_1093_port, regs(1092) => 
                           bus_reg_dataout_1092_port, regs(1091) => 
                           bus_reg_dataout_1091_port, regs(1090) => 
                           bus_reg_dataout_1090_port, regs(1089) => 
                           bus_reg_dataout_1089_port, regs(1088) => 
                           bus_reg_dataout_1088_port, regs(1087) => 
                           bus_reg_dataout_1087_port, regs(1086) => 
                           bus_reg_dataout_1086_port, regs(1085) => 
                           bus_reg_dataout_1085_port, regs(1084) => 
                           bus_reg_dataout_1084_port, regs(1083) => 
                           bus_reg_dataout_1083_port, regs(1082) => 
                           bus_reg_dataout_1082_port, regs(1081) => 
                           bus_reg_dataout_1081_port, regs(1080) => 
                           bus_reg_dataout_1080_port, regs(1079) => 
                           bus_reg_dataout_1079_port, regs(1078) => 
                           bus_reg_dataout_1078_port, regs(1077) => 
                           bus_reg_dataout_1077_port, regs(1076) => 
                           bus_reg_dataout_1076_port, regs(1075) => 
                           bus_reg_dataout_1075_port, regs(1074) => 
                           bus_reg_dataout_1074_port, regs(1073) => 
                           bus_reg_dataout_1073_port, regs(1072) => 
                           bus_reg_dataout_1072_port, regs(1071) => 
                           bus_reg_dataout_1071_port, regs(1070) => 
                           bus_reg_dataout_1070_port, regs(1069) => 
                           bus_reg_dataout_1069_port, regs(1068) => 
                           bus_reg_dataout_1068_port, regs(1067) => 
                           bus_reg_dataout_1067_port, regs(1066) => 
                           bus_reg_dataout_1066_port, regs(1065) => 
                           bus_reg_dataout_1065_port, regs(1064) => 
                           bus_reg_dataout_1064_port, regs(1063) => 
                           bus_reg_dataout_1063_port, regs(1062) => 
                           bus_reg_dataout_1062_port, regs(1061) => 
                           bus_reg_dataout_1061_port, regs(1060) => 
                           bus_reg_dataout_1060_port, regs(1059) => 
                           bus_reg_dataout_1059_port, regs(1058) => 
                           bus_reg_dataout_1058_port, regs(1057) => 
                           bus_reg_dataout_1057_port, regs(1056) => 
                           bus_reg_dataout_1056_port, regs(1055) => 
                           bus_reg_dataout_1055_port, regs(1054) => 
                           bus_reg_dataout_1054_port, regs(1053) => 
                           bus_reg_dataout_1053_port, regs(1052) => 
                           bus_reg_dataout_1052_port, regs(1051) => 
                           bus_reg_dataout_1051_port, regs(1050) => 
                           bus_reg_dataout_1050_port, regs(1049) => 
                           bus_reg_dataout_1049_port, regs(1048) => 
                           bus_reg_dataout_1048_port, regs(1047) => 
                           bus_reg_dataout_1047_port, regs(1046) => 
                           bus_reg_dataout_1046_port, regs(1045) => 
                           bus_reg_dataout_1045_port, regs(1044) => 
                           bus_reg_dataout_1044_port, regs(1043) => 
                           bus_reg_dataout_1043_port, regs(1042) => 
                           bus_reg_dataout_1042_port, regs(1041) => 
                           bus_reg_dataout_1041_port, regs(1040) => 
                           bus_reg_dataout_1040_port, regs(1039) => 
                           bus_reg_dataout_1039_port, regs(1038) => 
                           bus_reg_dataout_1038_port, regs(1037) => 
                           bus_reg_dataout_1037_port, regs(1036) => 
                           bus_reg_dataout_1036_port, regs(1035) => 
                           bus_reg_dataout_1035_port, regs(1034) => 
                           bus_reg_dataout_1034_port, regs(1033) => 
                           bus_reg_dataout_1033_port, regs(1032) => 
                           bus_reg_dataout_1032_port, regs(1031) => 
                           bus_reg_dataout_1031_port, regs(1030) => 
                           bus_reg_dataout_1030_port, regs(1029) => 
                           bus_reg_dataout_1029_port, regs(1028) => 
                           bus_reg_dataout_1028_port, regs(1027) => 
                           bus_reg_dataout_1027_port, regs(1026) => 
                           bus_reg_dataout_1026_port, regs(1025) => 
                           bus_reg_dataout_1025_port, regs(1024) => 
                           bus_reg_dataout_1024_port, regs(1023) => 
                           bus_reg_dataout_1023_port, regs(1022) => 
                           bus_reg_dataout_1022_port, regs(1021) => 
                           bus_reg_dataout_1021_port, regs(1020) => 
                           bus_reg_dataout_1020_port, regs(1019) => 
                           bus_reg_dataout_1019_port, regs(1018) => 
                           bus_reg_dataout_1018_port, regs(1017) => 
                           bus_reg_dataout_1017_port, regs(1016) => 
                           bus_reg_dataout_1016_port, regs(1015) => 
                           bus_reg_dataout_1015_port, regs(1014) => 
                           bus_reg_dataout_1014_port, regs(1013) => 
                           bus_reg_dataout_1013_port, regs(1012) => 
                           bus_reg_dataout_1012_port, regs(1011) => 
                           bus_reg_dataout_1011_port, regs(1010) => 
                           bus_reg_dataout_1010_port, regs(1009) => 
                           bus_reg_dataout_1009_port, regs(1008) => 
                           bus_reg_dataout_1008_port, regs(1007) => 
                           bus_reg_dataout_1007_port, regs(1006) => 
                           bus_reg_dataout_1006_port, regs(1005) => 
                           bus_reg_dataout_1005_port, regs(1004) => 
                           bus_reg_dataout_1004_port, regs(1003) => 
                           bus_reg_dataout_1003_port, regs(1002) => 
                           bus_reg_dataout_1002_port, regs(1001) => 
                           bus_reg_dataout_1001_port, regs(1000) => 
                           bus_reg_dataout_1000_port, regs(999) => 
                           bus_reg_dataout_999_port, regs(998) => 
                           bus_reg_dataout_998_port, regs(997) => 
                           bus_reg_dataout_997_port, regs(996) => 
                           bus_reg_dataout_996_port, regs(995) => 
                           bus_reg_dataout_995_port, regs(994) => 
                           bus_reg_dataout_994_port, regs(993) => 
                           bus_reg_dataout_993_port, regs(992) => 
                           bus_reg_dataout_992_port, regs(991) => 
                           bus_reg_dataout_991_port, regs(990) => 
                           bus_reg_dataout_990_port, regs(989) => 
                           bus_reg_dataout_989_port, regs(988) => 
                           bus_reg_dataout_988_port, regs(987) => 
                           bus_reg_dataout_987_port, regs(986) => 
                           bus_reg_dataout_986_port, regs(985) => 
                           bus_reg_dataout_985_port, regs(984) => 
                           bus_reg_dataout_984_port, regs(983) => 
                           bus_reg_dataout_983_port, regs(982) => 
                           bus_reg_dataout_982_port, regs(981) => 
                           bus_reg_dataout_981_port, regs(980) => 
                           bus_reg_dataout_980_port, regs(979) => 
                           bus_reg_dataout_979_port, regs(978) => 
                           bus_reg_dataout_978_port, regs(977) => 
                           bus_reg_dataout_977_port, regs(976) => 
                           bus_reg_dataout_976_port, regs(975) => 
                           bus_reg_dataout_975_port, regs(974) => 
                           bus_reg_dataout_974_port, regs(973) => 
                           bus_reg_dataout_973_port, regs(972) => 
                           bus_reg_dataout_972_port, regs(971) => 
                           bus_reg_dataout_971_port, regs(970) => 
                           bus_reg_dataout_970_port, regs(969) => 
                           bus_reg_dataout_969_port, regs(968) => 
                           bus_reg_dataout_968_port, regs(967) => 
                           bus_reg_dataout_967_port, regs(966) => 
                           bus_reg_dataout_966_port, regs(965) => 
                           bus_reg_dataout_965_port, regs(964) => 
                           bus_reg_dataout_964_port, regs(963) => 
                           bus_reg_dataout_963_port, regs(962) => 
                           bus_reg_dataout_962_port, regs(961) => 
                           bus_reg_dataout_961_port, regs(960) => 
                           bus_reg_dataout_960_port, regs(959) => 
                           bus_reg_dataout_959_port, regs(958) => 
                           bus_reg_dataout_958_port, regs(957) => 
                           bus_reg_dataout_957_port, regs(956) => 
                           bus_reg_dataout_956_port, regs(955) => 
                           bus_reg_dataout_955_port, regs(954) => 
                           bus_reg_dataout_954_port, regs(953) => 
                           bus_reg_dataout_953_port, regs(952) => 
                           bus_reg_dataout_952_port, regs(951) => 
                           bus_reg_dataout_951_port, regs(950) => 
                           bus_reg_dataout_950_port, regs(949) => 
                           bus_reg_dataout_949_port, regs(948) => 
                           bus_reg_dataout_948_port, regs(947) => 
                           bus_reg_dataout_947_port, regs(946) => 
                           bus_reg_dataout_946_port, regs(945) => 
                           bus_reg_dataout_945_port, regs(944) => 
                           bus_reg_dataout_944_port, regs(943) => 
                           bus_reg_dataout_943_port, regs(942) => 
                           bus_reg_dataout_942_port, regs(941) => 
                           bus_reg_dataout_941_port, regs(940) => 
                           bus_reg_dataout_940_port, regs(939) => 
                           bus_reg_dataout_939_port, regs(938) => 
                           bus_reg_dataout_938_port, regs(937) => 
                           bus_reg_dataout_937_port, regs(936) => 
                           bus_reg_dataout_936_port, regs(935) => 
                           bus_reg_dataout_935_port, regs(934) => 
                           bus_reg_dataout_934_port, regs(933) => 
                           bus_reg_dataout_933_port, regs(932) => 
                           bus_reg_dataout_932_port, regs(931) => 
                           bus_reg_dataout_931_port, regs(930) => 
                           bus_reg_dataout_930_port, regs(929) => 
                           bus_reg_dataout_929_port, regs(928) => 
                           bus_reg_dataout_928_port, regs(927) => 
                           bus_reg_dataout_927_port, regs(926) => 
                           bus_reg_dataout_926_port, regs(925) => 
                           bus_reg_dataout_925_port, regs(924) => 
                           bus_reg_dataout_924_port, regs(923) => 
                           bus_reg_dataout_923_port, regs(922) => 
                           bus_reg_dataout_922_port, regs(921) => 
                           bus_reg_dataout_921_port, regs(920) => 
                           bus_reg_dataout_920_port, regs(919) => 
                           bus_reg_dataout_919_port, regs(918) => 
                           bus_reg_dataout_918_port, regs(917) => 
                           bus_reg_dataout_917_port, regs(916) => 
                           bus_reg_dataout_916_port, regs(915) => 
                           bus_reg_dataout_915_port, regs(914) => 
                           bus_reg_dataout_914_port, regs(913) => 
                           bus_reg_dataout_913_port, regs(912) => 
                           bus_reg_dataout_912_port, regs(911) => 
                           bus_reg_dataout_911_port, regs(910) => 
                           bus_reg_dataout_910_port, regs(909) => 
                           bus_reg_dataout_909_port, regs(908) => 
                           bus_reg_dataout_908_port, regs(907) => 
                           bus_reg_dataout_907_port, regs(906) => 
                           bus_reg_dataout_906_port, regs(905) => 
                           bus_reg_dataout_905_port, regs(904) => 
                           bus_reg_dataout_904_port, regs(903) => 
                           bus_reg_dataout_903_port, regs(902) => 
                           bus_reg_dataout_902_port, regs(901) => 
                           bus_reg_dataout_901_port, regs(900) => 
                           bus_reg_dataout_900_port, regs(899) => 
                           bus_reg_dataout_899_port, regs(898) => 
                           bus_reg_dataout_898_port, regs(897) => 
                           bus_reg_dataout_897_port, regs(896) => 
                           bus_reg_dataout_896_port, regs(895) => 
                           bus_reg_dataout_895_port, regs(894) => 
                           bus_reg_dataout_894_port, regs(893) => 
                           bus_reg_dataout_893_port, regs(892) => 
                           bus_reg_dataout_892_port, regs(891) => 
                           bus_reg_dataout_891_port, regs(890) => 
                           bus_reg_dataout_890_port, regs(889) => 
                           bus_reg_dataout_889_port, regs(888) => 
                           bus_reg_dataout_888_port, regs(887) => 
                           bus_reg_dataout_887_port, regs(886) => 
                           bus_reg_dataout_886_port, regs(885) => 
                           bus_reg_dataout_885_port, regs(884) => 
                           bus_reg_dataout_884_port, regs(883) => 
                           bus_reg_dataout_883_port, regs(882) => 
                           bus_reg_dataout_882_port, regs(881) => 
                           bus_reg_dataout_881_port, regs(880) => 
                           bus_reg_dataout_880_port, regs(879) => 
                           bus_reg_dataout_879_port, regs(878) => 
                           bus_reg_dataout_878_port, regs(877) => 
                           bus_reg_dataout_877_port, regs(876) => 
                           bus_reg_dataout_876_port, regs(875) => 
                           bus_reg_dataout_875_port, regs(874) => 
                           bus_reg_dataout_874_port, regs(873) => 
                           bus_reg_dataout_873_port, regs(872) => 
                           bus_reg_dataout_872_port, regs(871) => 
                           bus_reg_dataout_871_port, regs(870) => 
                           bus_reg_dataout_870_port, regs(869) => 
                           bus_reg_dataout_869_port, regs(868) => 
                           bus_reg_dataout_868_port, regs(867) => 
                           bus_reg_dataout_867_port, regs(866) => 
                           bus_reg_dataout_866_port, regs(865) => 
                           bus_reg_dataout_865_port, regs(864) => 
                           bus_reg_dataout_864_port, regs(863) => 
                           bus_reg_dataout_863_port, regs(862) => 
                           bus_reg_dataout_862_port, regs(861) => 
                           bus_reg_dataout_861_port, regs(860) => 
                           bus_reg_dataout_860_port, regs(859) => 
                           bus_reg_dataout_859_port, regs(858) => 
                           bus_reg_dataout_858_port, regs(857) => 
                           bus_reg_dataout_857_port, regs(856) => 
                           bus_reg_dataout_856_port, regs(855) => 
                           bus_reg_dataout_855_port, regs(854) => 
                           bus_reg_dataout_854_port, regs(853) => 
                           bus_reg_dataout_853_port, regs(852) => 
                           bus_reg_dataout_852_port, regs(851) => 
                           bus_reg_dataout_851_port, regs(850) => 
                           bus_reg_dataout_850_port, regs(849) => 
                           bus_reg_dataout_849_port, regs(848) => 
                           bus_reg_dataout_848_port, regs(847) => 
                           bus_reg_dataout_847_port, regs(846) => 
                           bus_reg_dataout_846_port, regs(845) => 
                           bus_reg_dataout_845_port, regs(844) => 
                           bus_reg_dataout_844_port, regs(843) => 
                           bus_reg_dataout_843_port, regs(842) => 
                           bus_reg_dataout_842_port, regs(841) => 
                           bus_reg_dataout_841_port, regs(840) => 
                           bus_reg_dataout_840_port, regs(839) => 
                           bus_reg_dataout_839_port, regs(838) => 
                           bus_reg_dataout_838_port, regs(837) => 
                           bus_reg_dataout_837_port, regs(836) => 
                           bus_reg_dataout_836_port, regs(835) => 
                           bus_reg_dataout_835_port, regs(834) => 
                           bus_reg_dataout_834_port, regs(833) => 
                           bus_reg_dataout_833_port, regs(832) => 
                           bus_reg_dataout_832_port, regs(831) => 
                           bus_reg_dataout_831_port, regs(830) => 
                           bus_reg_dataout_830_port, regs(829) => 
                           bus_reg_dataout_829_port, regs(828) => 
                           bus_reg_dataout_828_port, regs(827) => 
                           bus_reg_dataout_827_port, regs(826) => 
                           bus_reg_dataout_826_port, regs(825) => 
                           bus_reg_dataout_825_port, regs(824) => 
                           bus_reg_dataout_824_port, regs(823) => 
                           bus_reg_dataout_823_port, regs(822) => 
                           bus_reg_dataout_822_port, regs(821) => 
                           bus_reg_dataout_821_port, regs(820) => 
                           bus_reg_dataout_820_port, regs(819) => 
                           bus_reg_dataout_819_port, regs(818) => 
                           bus_reg_dataout_818_port, regs(817) => 
                           bus_reg_dataout_817_port, regs(816) => 
                           bus_reg_dataout_816_port, regs(815) => 
                           bus_reg_dataout_815_port, regs(814) => 
                           bus_reg_dataout_814_port, regs(813) => 
                           bus_reg_dataout_813_port, regs(812) => 
                           bus_reg_dataout_812_port, regs(811) => 
                           bus_reg_dataout_811_port, regs(810) => 
                           bus_reg_dataout_810_port, regs(809) => 
                           bus_reg_dataout_809_port, regs(808) => 
                           bus_reg_dataout_808_port, regs(807) => 
                           bus_reg_dataout_807_port, regs(806) => 
                           bus_reg_dataout_806_port, regs(805) => 
                           bus_reg_dataout_805_port, regs(804) => 
                           bus_reg_dataout_804_port, regs(803) => 
                           bus_reg_dataout_803_port, regs(802) => 
                           bus_reg_dataout_802_port, regs(801) => 
                           bus_reg_dataout_801_port, regs(800) => 
                           bus_reg_dataout_800_port, regs(799) => 
                           bus_reg_dataout_799_port, regs(798) => 
                           bus_reg_dataout_798_port, regs(797) => 
                           bus_reg_dataout_797_port, regs(796) => 
                           bus_reg_dataout_796_port, regs(795) => 
                           bus_reg_dataout_795_port, regs(794) => 
                           bus_reg_dataout_794_port, regs(793) => 
                           bus_reg_dataout_793_port, regs(792) => 
                           bus_reg_dataout_792_port, regs(791) => 
                           bus_reg_dataout_791_port, regs(790) => 
                           bus_reg_dataout_790_port, regs(789) => 
                           bus_reg_dataout_789_port, regs(788) => 
                           bus_reg_dataout_788_port, regs(787) => 
                           bus_reg_dataout_787_port, regs(786) => 
                           bus_reg_dataout_786_port, regs(785) => 
                           bus_reg_dataout_785_port, regs(784) => 
                           bus_reg_dataout_784_port, regs(783) => 
                           bus_reg_dataout_783_port, regs(782) => 
                           bus_reg_dataout_782_port, regs(781) => 
                           bus_reg_dataout_781_port, regs(780) => 
                           bus_reg_dataout_780_port, regs(779) => 
                           bus_reg_dataout_779_port, regs(778) => 
                           bus_reg_dataout_778_port, regs(777) => 
                           bus_reg_dataout_777_port, regs(776) => 
                           bus_reg_dataout_776_port, regs(775) => 
                           bus_reg_dataout_775_port, regs(774) => 
                           bus_reg_dataout_774_port, regs(773) => 
                           bus_reg_dataout_773_port, regs(772) => 
                           bus_reg_dataout_772_port, regs(771) => 
                           bus_reg_dataout_771_port, regs(770) => 
                           bus_reg_dataout_770_port, regs(769) => 
                           bus_reg_dataout_769_port, regs(768) => 
                           bus_reg_dataout_768_port, regs(767) => 
                           bus_reg_dataout_767_port, regs(766) => 
                           bus_reg_dataout_766_port, regs(765) => 
                           bus_reg_dataout_765_port, regs(764) => 
                           bus_reg_dataout_764_port, regs(763) => 
                           bus_reg_dataout_763_port, regs(762) => 
                           bus_reg_dataout_762_port, regs(761) => 
                           bus_reg_dataout_761_port, regs(760) => 
                           bus_reg_dataout_760_port, regs(759) => 
                           bus_reg_dataout_759_port, regs(758) => 
                           bus_reg_dataout_758_port, regs(757) => 
                           bus_reg_dataout_757_port, regs(756) => 
                           bus_reg_dataout_756_port, regs(755) => 
                           bus_reg_dataout_755_port, regs(754) => 
                           bus_reg_dataout_754_port, regs(753) => 
                           bus_reg_dataout_753_port, regs(752) => 
                           bus_reg_dataout_752_port, regs(751) => 
                           bus_reg_dataout_751_port, regs(750) => 
                           bus_reg_dataout_750_port, regs(749) => 
                           bus_reg_dataout_749_port, regs(748) => 
                           bus_reg_dataout_748_port, regs(747) => 
                           bus_reg_dataout_747_port, regs(746) => 
                           bus_reg_dataout_746_port, regs(745) => 
                           bus_reg_dataout_745_port, regs(744) => 
                           bus_reg_dataout_744_port, regs(743) => 
                           bus_reg_dataout_743_port, regs(742) => 
                           bus_reg_dataout_742_port, regs(741) => 
                           bus_reg_dataout_741_port, regs(740) => 
                           bus_reg_dataout_740_port, regs(739) => 
                           bus_reg_dataout_739_port, regs(738) => 
                           bus_reg_dataout_738_port, regs(737) => 
                           bus_reg_dataout_737_port, regs(736) => 
                           bus_reg_dataout_736_port, regs(735) => 
                           bus_reg_dataout_735_port, regs(734) => 
                           bus_reg_dataout_734_port, regs(733) => 
                           bus_reg_dataout_733_port, regs(732) => 
                           bus_reg_dataout_732_port, regs(731) => 
                           bus_reg_dataout_731_port, regs(730) => 
                           bus_reg_dataout_730_port, regs(729) => 
                           bus_reg_dataout_729_port, regs(728) => 
                           bus_reg_dataout_728_port, regs(727) => 
                           bus_reg_dataout_727_port, regs(726) => 
                           bus_reg_dataout_726_port, regs(725) => 
                           bus_reg_dataout_725_port, regs(724) => 
                           bus_reg_dataout_724_port, regs(723) => 
                           bus_reg_dataout_723_port, regs(722) => 
                           bus_reg_dataout_722_port, regs(721) => 
                           bus_reg_dataout_721_port, regs(720) => 
                           bus_reg_dataout_720_port, regs(719) => 
                           bus_reg_dataout_719_port, regs(718) => 
                           bus_reg_dataout_718_port, regs(717) => 
                           bus_reg_dataout_717_port, regs(716) => 
                           bus_reg_dataout_716_port, regs(715) => 
                           bus_reg_dataout_715_port, regs(714) => 
                           bus_reg_dataout_714_port, regs(713) => 
                           bus_reg_dataout_713_port, regs(712) => 
                           bus_reg_dataout_712_port, regs(711) => 
                           bus_reg_dataout_711_port, regs(710) => 
                           bus_reg_dataout_710_port, regs(709) => 
                           bus_reg_dataout_709_port, regs(708) => 
                           bus_reg_dataout_708_port, regs(707) => 
                           bus_reg_dataout_707_port, regs(706) => 
                           bus_reg_dataout_706_port, regs(705) => 
                           bus_reg_dataout_705_port, regs(704) => 
                           bus_reg_dataout_704_port, regs(703) => 
                           bus_reg_dataout_703_port, regs(702) => 
                           bus_reg_dataout_702_port, regs(701) => 
                           bus_reg_dataout_701_port, regs(700) => 
                           bus_reg_dataout_700_port, regs(699) => 
                           bus_reg_dataout_699_port, regs(698) => 
                           bus_reg_dataout_698_port, regs(697) => 
                           bus_reg_dataout_697_port, regs(696) => 
                           bus_reg_dataout_696_port, regs(695) => 
                           bus_reg_dataout_695_port, regs(694) => 
                           bus_reg_dataout_694_port, regs(693) => 
                           bus_reg_dataout_693_port, regs(692) => 
                           bus_reg_dataout_692_port, regs(691) => 
                           bus_reg_dataout_691_port, regs(690) => 
                           bus_reg_dataout_690_port, regs(689) => 
                           bus_reg_dataout_689_port, regs(688) => 
                           bus_reg_dataout_688_port, regs(687) => 
                           bus_reg_dataout_687_port, regs(686) => 
                           bus_reg_dataout_686_port, regs(685) => 
                           bus_reg_dataout_685_port, regs(684) => 
                           bus_reg_dataout_684_port, regs(683) => 
                           bus_reg_dataout_683_port, regs(682) => 
                           bus_reg_dataout_682_port, regs(681) => 
                           bus_reg_dataout_681_port, regs(680) => 
                           bus_reg_dataout_680_port, regs(679) => 
                           bus_reg_dataout_679_port, regs(678) => 
                           bus_reg_dataout_678_port, regs(677) => 
                           bus_reg_dataout_677_port, regs(676) => 
                           bus_reg_dataout_676_port, regs(675) => 
                           bus_reg_dataout_675_port, regs(674) => 
                           bus_reg_dataout_674_port, regs(673) => 
                           bus_reg_dataout_673_port, regs(672) => 
                           bus_reg_dataout_672_port, regs(671) => 
                           bus_reg_dataout_671_port, regs(670) => 
                           bus_reg_dataout_670_port, regs(669) => 
                           bus_reg_dataout_669_port, regs(668) => 
                           bus_reg_dataout_668_port, regs(667) => 
                           bus_reg_dataout_667_port, regs(666) => 
                           bus_reg_dataout_666_port, regs(665) => 
                           bus_reg_dataout_665_port, regs(664) => 
                           bus_reg_dataout_664_port, regs(663) => 
                           bus_reg_dataout_663_port, regs(662) => 
                           bus_reg_dataout_662_port, regs(661) => 
                           bus_reg_dataout_661_port, regs(660) => 
                           bus_reg_dataout_660_port, regs(659) => 
                           bus_reg_dataout_659_port, regs(658) => 
                           bus_reg_dataout_658_port, regs(657) => 
                           bus_reg_dataout_657_port, regs(656) => 
                           bus_reg_dataout_656_port, regs(655) => 
                           bus_reg_dataout_655_port, regs(654) => 
                           bus_reg_dataout_654_port, regs(653) => 
                           bus_reg_dataout_653_port, regs(652) => 
                           bus_reg_dataout_652_port, regs(651) => 
                           bus_reg_dataout_651_port, regs(650) => 
                           bus_reg_dataout_650_port, regs(649) => 
                           bus_reg_dataout_649_port, regs(648) => 
                           bus_reg_dataout_648_port, regs(647) => 
                           bus_reg_dataout_647_port, regs(646) => 
                           bus_reg_dataout_646_port, regs(645) => 
                           bus_reg_dataout_645_port, regs(644) => 
                           bus_reg_dataout_644_port, regs(643) => 
                           bus_reg_dataout_643_port, regs(642) => 
                           bus_reg_dataout_642_port, regs(641) => 
                           bus_reg_dataout_641_port, regs(640) => 
                           bus_reg_dataout_640_port, regs(639) => 
                           bus_reg_dataout_639_port, regs(638) => 
                           bus_reg_dataout_638_port, regs(637) => 
                           bus_reg_dataout_637_port, regs(636) => 
                           bus_reg_dataout_636_port, regs(635) => 
                           bus_reg_dataout_635_port, regs(634) => 
                           bus_reg_dataout_634_port, regs(633) => 
                           bus_reg_dataout_633_port, regs(632) => 
                           bus_reg_dataout_632_port, regs(631) => 
                           bus_reg_dataout_631_port, regs(630) => 
                           bus_reg_dataout_630_port, regs(629) => 
                           bus_reg_dataout_629_port, regs(628) => 
                           bus_reg_dataout_628_port, regs(627) => 
                           bus_reg_dataout_627_port, regs(626) => 
                           bus_reg_dataout_626_port, regs(625) => 
                           bus_reg_dataout_625_port, regs(624) => 
                           bus_reg_dataout_624_port, regs(623) => 
                           bus_reg_dataout_623_port, regs(622) => 
                           bus_reg_dataout_622_port, regs(621) => 
                           bus_reg_dataout_621_port, regs(620) => 
                           bus_reg_dataout_620_port, regs(619) => 
                           bus_reg_dataout_619_port, regs(618) => 
                           bus_reg_dataout_618_port, regs(617) => 
                           bus_reg_dataout_617_port, regs(616) => 
                           bus_reg_dataout_616_port, regs(615) => 
                           bus_reg_dataout_615_port, regs(614) => 
                           bus_reg_dataout_614_port, regs(613) => 
                           bus_reg_dataout_613_port, regs(612) => 
                           bus_reg_dataout_612_port, regs(611) => 
                           bus_reg_dataout_611_port, regs(610) => 
                           bus_reg_dataout_610_port, regs(609) => 
                           bus_reg_dataout_609_port, regs(608) => 
                           bus_reg_dataout_608_port, regs(607) => 
                           bus_reg_dataout_607_port, regs(606) => 
                           bus_reg_dataout_606_port, regs(605) => 
                           bus_reg_dataout_605_port, regs(604) => 
                           bus_reg_dataout_604_port, regs(603) => 
                           bus_reg_dataout_603_port, regs(602) => 
                           bus_reg_dataout_602_port, regs(601) => 
                           bus_reg_dataout_601_port, regs(600) => 
                           bus_reg_dataout_600_port, regs(599) => 
                           bus_reg_dataout_599_port, regs(598) => 
                           bus_reg_dataout_598_port, regs(597) => 
                           bus_reg_dataout_597_port, regs(596) => 
                           bus_reg_dataout_596_port, regs(595) => 
                           bus_reg_dataout_595_port, regs(594) => 
                           bus_reg_dataout_594_port, regs(593) => 
                           bus_reg_dataout_593_port, regs(592) => 
                           bus_reg_dataout_592_port, regs(591) => 
                           bus_reg_dataout_591_port, regs(590) => 
                           bus_reg_dataout_590_port, regs(589) => 
                           bus_reg_dataout_589_port, regs(588) => 
                           bus_reg_dataout_588_port, regs(587) => 
                           bus_reg_dataout_587_port, regs(586) => 
                           bus_reg_dataout_586_port, regs(585) => 
                           bus_reg_dataout_585_port, regs(584) => 
                           bus_reg_dataout_584_port, regs(583) => 
                           bus_reg_dataout_583_port, regs(582) => 
                           bus_reg_dataout_582_port, regs(581) => 
                           bus_reg_dataout_581_port, regs(580) => 
                           bus_reg_dataout_580_port, regs(579) => 
                           bus_reg_dataout_579_port, regs(578) => 
                           bus_reg_dataout_578_port, regs(577) => 
                           bus_reg_dataout_577_port, regs(576) => 
                           bus_reg_dataout_576_port, regs(575) => 
                           bus_reg_dataout_575_port, regs(574) => 
                           bus_reg_dataout_574_port, regs(573) => 
                           bus_reg_dataout_573_port, regs(572) => 
                           bus_reg_dataout_572_port, regs(571) => 
                           bus_reg_dataout_571_port, regs(570) => 
                           bus_reg_dataout_570_port, regs(569) => 
                           bus_reg_dataout_569_port, regs(568) => 
                           bus_reg_dataout_568_port, regs(567) => 
                           bus_reg_dataout_567_port, regs(566) => 
                           bus_reg_dataout_566_port, regs(565) => 
                           bus_reg_dataout_565_port, regs(564) => 
                           bus_reg_dataout_564_port, regs(563) => 
                           bus_reg_dataout_563_port, regs(562) => 
                           bus_reg_dataout_562_port, regs(561) => 
                           bus_reg_dataout_561_port, regs(560) => 
                           bus_reg_dataout_560_port, regs(559) => 
                           bus_reg_dataout_559_port, regs(558) => 
                           bus_reg_dataout_558_port, regs(557) => 
                           bus_reg_dataout_557_port, regs(556) => 
                           bus_reg_dataout_556_port, regs(555) => 
                           bus_reg_dataout_555_port, regs(554) => 
                           bus_reg_dataout_554_port, regs(553) => 
                           bus_reg_dataout_553_port, regs(552) => 
                           bus_reg_dataout_552_port, regs(551) => 
                           bus_reg_dataout_551_port, regs(550) => 
                           bus_reg_dataout_550_port, regs(549) => 
                           bus_reg_dataout_549_port, regs(548) => 
                           bus_reg_dataout_548_port, regs(547) => 
                           bus_reg_dataout_547_port, regs(546) => 
                           bus_reg_dataout_546_port, regs(545) => 
                           bus_reg_dataout_545_port, regs(544) => 
                           bus_reg_dataout_544_port, regs(543) => 
                           bus_reg_dataout_543_port, regs(542) => 
                           bus_reg_dataout_542_port, regs(541) => 
                           bus_reg_dataout_541_port, regs(540) => 
                           bus_reg_dataout_540_port, regs(539) => 
                           bus_reg_dataout_539_port, regs(538) => 
                           bus_reg_dataout_538_port, regs(537) => 
                           bus_reg_dataout_537_port, regs(536) => 
                           bus_reg_dataout_536_port, regs(535) => 
                           bus_reg_dataout_535_port, regs(534) => 
                           bus_reg_dataout_534_port, regs(533) => 
                           bus_reg_dataout_533_port, regs(532) => 
                           bus_reg_dataout_532_port, regs(531) => 
                           bus_reg_dataout_531_port, regs(530) => 
                           bus_reg_dataout_530_port, regs(529) => 
                           bus_reg_dataout_529_port, regs(528) => 
                           bus_reg_dataout_528_port, regs(527) => 
                           bus_reg_dataout_527_port, regs(526) => 
                           bus_reg_dataout_526_port, regs(525) => 
                           bus_reg_dataout_525_port, regs(524) => 
                           bus_reg_dataout_524_port, regs(523) => 
                           bus_reg_dataout_523_port, regs(522) => 
                           bus_reg_dataout_522_port, regs(521) => 
                           bus_reg_dataout_521_port, regs(520) => 
                           bus_reg_dataout_520_port, regs(519) => 
                           bus_reg_dataout_519_port, regs(518) => 
                           bus_reg_dataout_518_port, regs(517) => 
                           bus_reg_dataout_517_port, regs(516) => 
                           bus_reg_dataout_516_port, regs(515) => 
                           bus_reg_dataout_515_port, regs(514) => 
                           bus_reg_dataout_514_port, regs(513) => 
                           bus_reg_dataout_513_port, regs(512) => 
                           bus_reg_dataout_512_port, regs(511) => 
                           bus_reg_dataout_511_port, regs(510) => 
                           bus_reg_dataout_510_port, regs(509) => 
                           bus_reg_dataout_509_port, regs(508) => 
                           bus_reg_dataout_508_port, regs(507) => 
                           bus_reg_dataout_507_port, regs(506) => 
                           bus_reg_dataout_506_port, regs(505) => 
                           bus_reg_dataout_505_port, regs(504) => 
                           bus_reg_dataout_504_port, regs(503) => 
                           bus_reg_dataout_503_port, regs(502) => 
                           bus_reg_dataout_502_port, regs(501) => 
                           bus_reg_dataout_501_port, regs(500) => 
                           bus_reg_dataout_500_port, regs(499) => 
                           bus_reg_dataout_499_port, regs(498) => 
                           bus_reg_dataout_498_port, regs(497) => 
                           bus_reg_dataout_497_port, regs(496) => 
                           bus_reg_dataout_496_port, regs(495) => 
                           bus_reg_dataout_495_port, regs(494) => 
                           bus_reg_dataout_494_port, regs(493) => 
                           bus_reg_dataout_493_port, regs(492) => 
                           bus_reg_dataout_492_port, regs(491) => 
                           bus_reg_dataout_491_port, regs(490) => 
                           bus_reg_dataout_490_port, regs(489) => 
                           bus_reg_dataout_489_port, regs(488) => 
                           bus_reg_dataout_488_port, regs(487) => 
                           bus_reg_dataout_487_port, regs(486) => 
                           bus_reg_dataout_486_port, regs(485) => 
                           bus_reg_dataout_485_port, regs(484) => 
                           bus_reg_dataout_484_port, regs(483) => 
                           bus_reg_dataout_483_port, regs(482) => 
                           bus_reg_dataout_482_port, regs(481) => 
                           bus_reg_dataout_481_port, regs(480) => 
                           bus_reg_dataout_480_port, regs(479) => 
                           bus_reg_dataout_479_port, regs(478) => 
                           bus_reg_dataout_478_port, regs(477) => 
                           bus_reg_dataout_477_port, regs(476) => 
                           bus_reg_dataout_476_port, regs(475) => 
                           bus_reg_dataout_475_port, regs(474) => 
                           bus_reg_dataout_474_port, regs(473) => 
                           bus_reg_dataout_473_port, regs(472) => 
                           bus_reg_dataout_472_port, regs(471) => 
                           bus_reg_dataout_471_port, regs(470) => 
                           bus_reg_dataout_470_port, regs(469) => 
                           bus_reg_dataout_469_port, regs(468) => 
                           bus_reg_dataout_468_port, regs(467) => 
                           bus_reg_dataout_467_port, regs(466) => 
                           bus_reg_dataout_466_port, regs(465) => 
                           bus_reg_dataout_465_port, regs(464) => 
                           bus_reg_dataout_464_port, regs(463) => 
                           bus_reg_dataout_463_port, regs(462) => 
                           bus_reg_dataout_462_port, regs(461) => 
                           bus_reg_dataout_461_port, regs(460) => 
                           bus_reg_dataout_460_port, regs(459) => 
                           bus_reg_dataout_459_port, regs(458) => 
                           bus_reg_dataout_458_port, regs(457) => 
                           bus_reg_dataout_457_port, regs(456) => 
                           bus_reg_dataout_456_port, regs(455) => 
                           bus_reg_dataout_455_port, regs(454) => 
                           bus_reg_dataout_454_port, regs(453) => 
                           bus_reg_dataout_453_port, regs(452) => 
                           bus_reg_dataout_452_port, regs(451) => 
                           bus_reg_dataout_451_port, regs(450) => 
                           bus_reg_dataout_450_port, regs(449) => 
                           bus_reg_dataout_449_port, regs(448) => 
                           bus_reg_dataout_448_port, regs(447) => 
                           bus_reg_dataout_447_port, regs(446) => 
                           bus_reg_dataout_446_port, regs(445) => 
                           bus_reg_dataout_445_port, regs(444) => 
                           bus_reg_dataout_444_port, regs(443) => 
                           bus_reg_dataout_443_port, regs(442) => 
                           bus_reg_dataout_442_port, regs(441) => 
                           bus_reg_dataout_441_port, regs(440) => 
                           bus_reg_dataout_440_port, regs(439) => 
                           bus_reg_dataout_439_port, regs(438) => 
                           bus_reg_dataout_438_port, regs(437) => 
                           bus_reg_dataout_437_port, regs(436) => 
                           bus_reg_dataout_436_port, regs(435) => 
                           bus_reg_dataout_435_port, regs(434) => 
                           bus_reg_dataout_434_port, regs(433) => 
                           bus_reg_dataout_433_port, regs(432) => 
                           bus_reg_dataout_432_port, regs(431) => 
                           bus_reg_dataout_431_port, regs(430) => 
                           bus_reg_dataout_430_port, regs(429) => 
                           bus_reg_dataout_429_port, regs(428) => 
                           bus_reg_dataout_428_port, regs(427) => 
                           bus_reg_dataout_427_port, regs(426) => 
                           bus_reg_dataout_426_port, regs(425) => 
                           bus_reg_dataout_425_port, regs(424) => 
                           bus_reg_dataout_424_port, regs(423) => 
                           bus_reg_dataout_423_port, regs(422) => 
                           bus_reg_dataout_422_port, regs(421) => 
                           bus_reg_dataout_421_port, regs(420) => 
                           bus_reg_dataout_420_port, regs(419) => 
                           bus_reg_dataout_419_port, regs(418) => 
                           bus_reg_dataout_418_port, regs(417) => 
                           bus_reg_dataout_417_port, regs(416) => 
                           bus_reg_dataout_416_port, regs(415) => 
                           bus_reg_dataout_415_port, regs(414) => 
                           bus_reg_dataout_414_port, regs(413) => 
                           bus_reg_dataout_413_port, regs(412) => 
                           bus_reg_dataout_412_port, regs(411) => 
                           bus_reg_dataout_411_port, regs(410) => 
                           bus_reg_dataout_410_port, regs(409) => 
                           bus_reg_dataout_409_port, regs(408) => 
                           bus_reg_dataout_408_port, regs(407) => 
                           bus_reg_dataout_407_port, regs(406) => 
                           bus_reg_dataout_406_port, regs(405) => 
                           bus_reg_dataout_405_port, regs(404) => 
                           bus_reg_dataout_404_port, regs(403) => 
                           bus_reg_dataout_403_port, regs(402) => 
                           bus_reg_dataout_402_port, regs(401) => 
                           bus_reg_dataout_401_port, regs(400) => 
                           bus_reg_dataout_400_port, regs(399) => 
                           bus_reg_dataout_399_port, regs(398) => 
                           bus_reg_dataout_398_port, regs(397) => 
                           bus_reg_dataout_397_port, regs(396) => 
                           bus_reg_dataout_396_port, regs(395) => 
                           bus_reg_dataout_395_port, regs(394) => 
                           bus_reg_dataout_394_port, regs(393) => 
                           bus_reg_dataout_393_port, regs(392) => 
                           bus_reg_dataout_392_port, regs(391) => 
                           bus_reg_dataout_391_port, regs(390) => 
                           bus_reg_dataout_390_port, regs(389) => 
                           bus_reg_dataout_389_port, regs(388) => 
                           bus_reg_dataout_388_port, regs(387) => 
                           bus_reg_dataout_387_port, regs(386) => 
                           bus_reg_dataout_386_port, regs(385) => 
                           bus_reg_dataout_385_port, regs(384) => 
                           bus_reg_dataout_384_port, regs(383) => 
                           bus_reg_dataout_383_port, regs(382) => 
                           bus_reg_dataout_382_port, regs(381) => 
                           bus_reg_dataout_381_port, regs(380) => 
                           bus_reg_dataout_380_port, regs(379) => 
                           bus_reg_dataout_379_port, regs(378) => 
                           bus_reg_dataout_378_port, regs(377) => 
                           bus_reg_dataout_377_port, regs(376) => 
                           bus_reg_dataout_376_port, regs(375) => 
                           bus_reg_dataout_375_port, regs(374) => 
                           bus_reg_dataout_374_port, regs(373) => 
                           bus_reg_dataout_373_port, regs(372) => 
                           bus_reg_dataout_372_port, regs(371) => 
                           bus_reg_dataout_371_port, regs(370) => 
                           bus_reg_dataout_370_port, regs(369) => 
                           bus_reg_dataout_369_port, regs(368) => 
                           bus_reg_dataout_368_port, regs(367) => 
                           bus_reg_dataout_367_port, regs(366) => 
                           bus_reg_dataout_366_port, regs(365) => 
                           bus_reg_dataout_365_port, regs(364) => 
                           bus_reg_dataout_364_port, regs(363) => 
                           bus_reg_dataout_363_port, regs(362) => 
                           bus_reg_dataout_362_port, regs(361) => 
                           bus_reg_dataout_361_port, regs(360) => 
                           bus_reg_dataout_360_port, regs(359) => 
                           bus_reg_dataout_359_port, regs(358) => 
                           bus_reg_dataout_358_port, regs(357) => 
                           bus_reg_dataout_357_port, regs(356) => 
                           bus_reg_dataout_356_port, regs(355) => 
                           bus_reg_dataout_355_port, regs(354) => 
                           bus_reg_dataout_354_port, regs(353) => 
                           bus_reg_dataout_353_port, regs(352) => 
                           bus_reg_dataout_352_port, regs(351) => 
                           bus_reg_dataout_351_port, regs(350) => 
                           bus_reg_dataout_350_port, regs(349) => 
                           bus_reg_dataout_349_port, regs(348) => 
                           bus_reg_dataout_348_port, regs(347) => 
                           bus_reg_dataout_347_port, regs(346) => 
                           bus_reg_dataout_346_port, regs(345) => 
                           bus_reg_dataout_345_port, regs(344) => 
                           bus_reg_dataout_344_port, regs(343) => 
                           bus_reg_dataout_343_port, regs(342) => 
                           bus_reg_dataout_342_port, regs(341) => 
                           bus_reg_dataout_341_port, regs(340) => 
                           bus_reg_dataout_340_port, regs(339) => 
                           bus_reg_dataout_339_port, regs(338) => 
                           bus_reg_dataout_338_port, regs(337) => 
                           bus_reg_dataout_337_port, regs(336) => 
                           bus_reg_dataout_336_port, regs(335) => 
                           bus_reg_dataout_335_port, regs(334) => 
                           bus_reg_dataout_334_port, regs(333) => 
                           bus_reg_dataout_333_port, regs(332) => 
                           bus_reg_dataout_332_port, regs(331) => 
                           bus_reg_dataout_331_port, regs(330) => 
                           bus_reg_dataout_330_port, regs(329) => 
                           bus_reg_dataout_329_port, regs(328) => 
                           bus_reg_dataout_328_port, regs(327) => 
                           bus_reg_dataout_327_port, regs(326) => 
                           bus_reg_dataout_326_port, regs(325) => 
                           bus_reg_dataout_325_port, regs(324) => 
                           bus_reg_dataout_324_port, regs(323) => 
                           bus_reg_dataout_323_port, regs(322) => 
                           bus_reg_dataout_322_port, regs(321) => 
                           bus_reg_dataout_321_port, regs(320) => 
                           bus_reg_dataout_320_port, regs(319) => 
                           bus_reg_dataout_319_port, regs(318) => 
                           bus_reg_dataout_318_port, regs(317) => 
                           bus_reg_dataout_317_port, regs(316) => 
                           bus_reg_dataout_316_port, regs(315) => 
                           bus_reg_dataout_315_port, regs(314) => 
                           bus_reg_dataout_314_port, regs(313) => 
                           bus_reg_dataout_313_port, regs(312) => 
                           bus_reg_dataout_312_port, regs(311) => 
                           bus_reg_dataout_311_port, regs(310) => 
                           bus_reg_dataout_310_port, regs(309) => 
                           bus_reg_dataout_309_port, regs(308) => 
                           bus_reg_dataout_308_port, regs(307) => 
                           bus_reg_dataout_307_port, regs(306) => 
                           bus_reg_dataout_306_port, regs(305) => 
                           bus_reg_dataout_305_port, regs(304) => 
                           bus_reg_dataout_304_port, regs(303) => 
                           bus_reg_dataout_303_port, regs(302) => 
                           bus_reg_dataout_302_port, regs(301) => 
                           bus_reg_dataout_301_port, regs(300) => 
                           bus_reg_dataout_300_port, regs(299) => 
                           bus_reg_dataout_299_port, regs(298) => 
                           bus_reg_dataout_298_port, regs(297) => 
                           bus_reg_dataout_297_port, regs(296) => 
                           bus_reg_dataout_296_port, regs(295) => 
                           bus_reg_dataout_295_port, regs(294) => 
                           bus_reg_dataout_294_port, regs(293) => 
                           bus_reg_dataout_293_port, regs(292) => 
                           bus_reg_dataout_292_port, regs(291) => 
                           bus_reg_dataout_291_port, regs(290) => 
                           bus_reg_dataout_290_port, regs(289) => 
                           bus_reg_dataout_289_port, regs(288) => 
                           bus_reg_dataout_288_port, regs(287) => 
                           bus_reg_dataout_287_port, regs(286) => 
                           bus_reg_dataout_286_port, regs(285) => 
                           bus_reg_dataout_285_port, regs(284) => 
                           bus_reg_dataout_284_port, regs(283) => 
                           bus_reg_dataout_283_port, regs(282) => 
                           bus_reg_dataout_282_port, regs(281) => 
                           bus_reg_dataout_281_port, regs(280) => 
                           bus_reg_dataout_280_port, regs(279) => 
                           bus_reg_dataout_279_port, regs(278) => 
                           bus_reg_dataout_278_port, regs(277) => 
                           bus_reg_dataout_277_port, regs(276) => 
                           bus_reg_dataout_276_port, regs(275) => 
                           bus_reg_dataout_275_port, regs(274) => 
                           bus_reg_dataout_274_port, regs(273) => 
                           bus_reg_dataout_273_port, regs(272) => 
                           bus_reg_dataout_272_port, regs(271) => 
                           bus_reg_dataout_271_port, regs(270) => 
                           bus_reg_dataout_270_port, regs(269) => 
                           bus_reg_dataout_269_port, regs(268) => 
                           bus_reg_dataout_268_port, regs(267) => 
                           bus_reg_dataout_267_port, regs(266) => 
                           bus_reg_dataout_266_port, regs(265) => 
                           bus_reg_dataout_265_port, regs(264) => 
                           bus_reg_dataout_264_port, regs(263) => 
                           bus_reg_dataout_263_port, regs(262) => 
                           bus_reg_dataout_262_port, regs(261) => 
                           bus_reg_dataout_261_port, regs(260) => 
                           bus_reg_dataout_260_port, regs(259) => 
                           bus_reg_dataout_259_port, regs(258) => 
                           bus_reg_dataout_258_port, regs(257) => 
                           bus_reg_dataout_257_port, regs(256) => 
                           bus_reg_dataout_256_port, regs(255) => 
                           bus_reg_dataout_255_port, regs(254) => 
                           bus_reg_dataout_254_port, regs(253) => 
                           bus_reg_dataout_253_port, regs(252) => 
                           bus_reg_dataout_252_port, regs(251) => 
                           bus_reg_dataout_251_port, regs(250) => 
                           bus_reg_dataout_250_port, regs(249) => 
                           bus_reg_dataout_249_port, regs(248) => 
                           bus_reg_dataout_248_port, regs(247) => 
                           bus_reg_dataout_247_port, regs(246) => 
                           bus_reg_dataout_246_port, regs(245) => 
                           bus_reg_dataout_245_port, regs(244) => 
                           bus_reg_dataout_244_port, regs(243) => 
                           bus_reg_dataout_243_port, regs(242) => 
                           bus_reg_dataout_242_port, regs(241) => 
                           bus_reg_dataout_241_port, regs(240) => 
                           bus_reg_dataout_240_port, regs(239) => 
                           bus_reg_dataout_239_port, regs(238) => 
                           bus_reg_dataout_238_port, regs(237) => 
                           bus_reg_dataout_237_port, regs(236) => 
                           bus_reg_dataout_236_port, regs(235) => 
                           bus_reg_dataout_235_port, regs(234) => 
                           bus_reg_dataout_234_port, regs(233) => 
                           bus_reg_dataout_233_port, regs(232) => 
                           bus_reg_dataout_232_port, regs(231) => 
                           bus_reg_dataout_231_port, regs(230) => 
                           bus_reg_dataout_230_port, regs(229) => 
                           bus_reg_dataout_229_port, regs(228) => 
                           bus_reg_dataout_228_port, regs(227) => 
                           bus_reg_dataout_227_port, regs(226) => 
                           bus_reg_dataout_226_port, regs(225) => 
                           bus_reg_dataout_225_port, regs(224) => 
                           bus_reg_dataout_224_port, regs(223) => 
                           bus_reg_dataout_223_port, regs(222) => 
                           bus_reg_dataout_222_port, regs(221) => 
                           bus_reg_dataout_221_port, regs(220) => 
                           bus_reg_dataout_220_port, regs(219) => 
                           bus_reg_dataout_219_port, regs(218) => 
                           bus_reg_dataout_218_port, regs(217) => 
                           bus_reg_dataout_217_port, regs(216) => 
                           bus_reg_dataout_216_port, regs(215) => 
                           bus_reg_dataout_215_port, regs(214) => 
                           bus_reg_dataout_214_port, regs(213) => 
                           bus_reg_dataout_213_port, regs(212) => 
                           bus_reg_dataout_212_port, regs(211) => 
                           bus_reg_dataout_211_port, regs(210) => 
                           bus_reg_dataout_210_port, regs(209) => 
                           bus_reg_dataout_209_port, regs(208) => 
                           bus_reg_dataout_208_port, regs(207) => 
                           bus_reg_dataout_207_port, regs(206) => 
                           bus_reg_dataout_206_port, regs(205) => 
                           bus_reg_dataout_205_port, regs(204) => 
                           bus_reg_dataout_204_port, regs(203) => 
                           bus_reg_dataout_203_port, regs(202) => 
                           bus_reg_dataout_202_port, regs(201) => 
                           bus_reg_dataout_201_port, regs(200) => 
                           bus_reg_dataout_200_port, regs(199) => 
                           bus_reg_dataout_199_port, regs(198) => 
                           bus_reg_dataout_198_port, regs(197) => 
                           bus_reg_dataout_197_port, regs(196) => 
                           bus_reg_dataout_196_port, regs(195) => 
                           bus_reg_dataout_195_port, regs(194) => 
                           bus_reg_dataout_194_port, regs(193) => 
                           bus_reg_dataout_193_port, regs(192) => 
                           bus_reg_dataout_192_port, regs(191) => 
                           bus_reg_dataout_191_port, regs(190) => 
                           bus_reg_dataout_190_port, regs(189) => 
                           bus_reg_dataout_189_port, regs(188) => 
                           bus_reg_dataout_188_port, regs(187) => 
                           bus_reg_dataout_187_port, regs(186) => 
                           bus_reg_dataout_186_port, regs(185) => 
                           bus_reg_dataout_185_port, regs(184) => 
                           bus_reg_dataout_184_port, regs(183) => 
                           bus_reg_dataout_183_port, regs(182) => 
                           bus_reg_dataout_182_port, regs(181) => 
                           bus_reg_dataout_181_port, regs(180) => 
                           bus_reg_dataout_180_port, regs(179) => 
                           bus_reg_dataout_179_port, regs(178) => 
                           bus_reg_dataout_178_port, regs(177) => 
                           bus_reg_dataout_177_port, regs(176) => 
                           bus_reg_dataout_176_port, regs(175) => 
                           bus_reg_dataout_175_port, regs(174) => 
                           bus_reg_dataout_174_port, regs(173) => 
                           bus_reg_dataout_173_port, regs(172) => 
                           bus_reg_dataout_172_port, regs(171) => 
                           bus_reg_dataout_171_port, regs(170) => 
                           bus_reg_dataout_170_port, regs(169) => 
                           bus_reg_dataout_169_port, regs(168) => 
                           bus_reg_dataout_168_port, regs(167) => 
                           bus_reg_dataout_167_port, regs(166) => 
                           bus_reg_dataout_166_port, regs(165) => 
                           bus_reg_dataout_165_port, regs(164) => 
                           bus_reg_dataout_164_port, regs(163) => 
                           bus_reg_dataout_163_port, regs(162) => 
                           bus_reg_dataout_162_port, regs(161) => 
                           bus_reg_dataout_161_port, regs(160) => 
                           bus_reg_dataout_160_port, regs(159) => 
                           bus_reg_dataout_159_port, regs(158) => 
                           bus_reg_dataout_158_port, regs(157) => 
                           bus_reg_dataout_157_port, regs(156) => 
                           bus_reg_dataout_156_port, regs(155) => 
                           bus_reg_dataout_155_port, regs(154) => 
                           bus_reg_dataout_154_port, regs(153) => 
                           bus_reg_dataout_153_port, regs(152) => 
                           bus_reg_dataout_152_port, regs(151) => 
                           bus_reg_dataout_151_port, regs(150) => 
                           bus_reg_dataout_150_port, regs(149) => 
                           bus_reg_dataout_149_port, regs(148) => 
                           bus_reg_dataout_148_port, regs(147) => 
                           bus_reg_dataout_147_port, regs(146) => 
                           bus_reg_dataout_146_port, regs(145) => 
                           bus_reg_dataout_145_port, regs(144) => 
                           bus_reg_dataout_144_port, regs(143) => 
                           bus_reg_dataout_143_port, regs(142) => 
                           bus_reg_dataout_142_port, regs(141) => 
                           bus_reg_dataout_141_port, regs(140) => 
                           bus_reg_dataout_140_port, regs(139) => 
                           bus_reg_dataout_139_port, regs(138) => 
                           bus_reg_dataout_138_port, regs(137) => 
                           bus_reg_dataout_137_port, regs(136) => 
                           bus_reg_dataout_136_port, regs(135) => 
                           bus_reg_dataout_135_port, regs(134) => 
                           bus_reg_dataout_134_port, regs(133) => 
                           bus_reg_dataout_133_port, regs(132) => 
                           bus_reg_dataout_132_port, regs(131) => 
                           bus_reg_dataout_131_port, regs(130) => 
                           bus_reg_dataout_130_port, regs(129) => 
                           bus_reg_dataout_129_port, regs(128) => 
                           bus_reg_dataout_128_port, regs(127) => 
                           bus_reg_dataout_127_port, regs(126) => 
                           bus_reg_dataout_126_port, regs(125) => 
                           bus_reg_dataout_125_port, regs(124) => 
                           bus_reg_dataout_124_port, regs(123) => 
                           bus_reg_dataout_123_port, regs(122) => 
                           bus_reg_dataout_122_port, regs(121) => 
                           bus_reg_dataout_121_port, regs(120) => 
                           bus_reg_dataout_120_port, regs(119) => 
                           bus_reg_dataout_119_port, regs(118) => 
                           bus_reg_dataout_118_port, regs(117) => 
                           bus_reg_dataout_117_port, regs(116) => 
                           bus_reg_dataout_116_port, regs(115) => 
                           bus_reg_dataout_115_port, regs(114) => 
                           bus_reg_dataout_114_port, regs(113) => 
                           bus_reg_dataout_113_port, regs(112) => 
                           bus_reg_dataout_112_port, regs(111) => 
                           bus_reg_dataout_111_port, regs(110) => 
                           bus_reg_dataout_110_port, regs(109) => 
                           bus_reg_dataout_109_port, regs(108) => 
                           bus_reg_dataout_108_port, regs(107) => 
                           bus_reg_dataout_107_port, regs(106) => 
                           bus_reg_dataout_106_port, regs(105) => 
                           bus_reg_dataout_105_port, regs(104) => 
                           bus_reg_dataout_104_port, regs(103) => 
                           bus_reg_dataout_103_port, regs(102) => 
                           bus_reg_dataout_102_port, regs(101) => 
                           bus_reg_dataout_101_port, regs(100) => 
                           bus_reg_dataout_100_port, regs(99) => 
                           bus_reg_dataout_99_port, regs(98) => 
                           bus_reg_dataout_98_port, regs(97) => 
                           bus_reg_dataout_97_port, regs(96) => 
                           bus_reg_dataout_96_port, regs(95) => 
                           bus_reg_dataout_95_port, regs(94) => 
                           bus_reg_dataout_94_port, regs(93) => 
                           bus_reg_dataout_93_port, regs(92) => 
                           bus_reg_dataout_92_port, regs(91) => 
                           bus_reg_dataout_91_port, regs(90) => 
                           bus_reg_dataout_90_port, regs(89) => 
                           bus_reg_dataout_89_port, regs(88) => 
                           bus_reg_dataout_88_port, regs(87) => 
                           bus_reg_dataout_87_port, regs(86) => 
                           bus_reg_dataout_86_port, regs(85) => 
                           bus_reg_dataout_85_port, regs(84) => 
                           bus_reg_dataout_84_port, regs(83) => 
                           bus_reg_dataout_83_port, regs(82) => 
                           bus_reg_dataout_82_port, regs(81) => 
                           bus_reg_dataout_81_port, regs(80) => 
                           bus_reg_dataout_80_port, regs(79) => 
                           bus_reg_dataout_79_port, regs(78) => 
                           bus_reg_dataout_78_port, regs(77) => 
                           bus_reg_dataout_77_port, regs(76) => 
                           bus_reg_dataout_76_port, regs(75) => 
                           bus_reg_dataout_75_port, regs(74) => 
                           bus_reg_dataout_74_port, regs(73) => 
                           bus_reg_dataout_73_port, regs(72) => 
                           bus_reg_dataout_72_port, regs(71) => 
                           bus_reg_dataout_71_port, regs(70) => 
                           bus_reg_dataout_70_port, regs(69) => 
                           bus_reg_dataout_69_port, regs(68) => 
                           bus_reg_dataout_68_port, regs(67) => 
                           bus_reg_dataout_67_port, regs(66) => 
                           bus_reg_dataout_66_port, regs(65) => 
                           bus_reg_dataout_65_port, regs(64) => 
                           bus_reg_dataout_64_port, regs(63) => 
                           bus_reg_dataout_63_port, regs(62) => 
                           bus_reg_dataout_62_port, regs(61) => 
                           bus_reg_dataout_61_port, regs(60) => 
                           bus_reg_dataout_60_port, regs(59) => 
                           bus_reg_dataout_59_port, regs(58) => 
                           bus_reg_dataout_58_port, regs(57) => 
                           bus_reg_dataout_57_port, regs(56) => 
                           bus_reg_dataout_56_port, regs(55) => 
                           bus_reg_dataout_55_port, regs(54) => 
                           bus_reg_dataout_54_port, regs(53) => 
                           bus_reg_dataout_53_port, regs(52) => 
                           bus_reg_dataout_52_port, regs(51) => 
                           bus_reg_dataout_51_port, regs(50) => 
                           bus_reg_dataout_50_port, regs(49) => 
                           bus_reg_dataout_49_port, regs(48) => 
                           bus_reg_dataout_48_port, regs(47) => 
                           bus_reg_dataout_47_port, regs(46) => 
                           bus_reg_dataout_46_port, regs(45) => 
                           bus_reg_dataout_45_port, regs(44) => 
                           bus_reg_dataout_44_port, regs(43) => 
                           bus_reg_dataout_43_port, regs(42) => 
                           bus_reg_dataout_42_port, regs(41) => 
                           bus_reg_dataout_41_port, regs(40) => 
                           bus_reg_dataout_40_port, regs(39) => 
                           bus_reg_dataout_39_port, regs(38) => 
                           bus_reg_dataout_38_port, regs(37) => 
                           bus_reg_dataout_37_port, regs(36) => 
                           bus_reg_dataout_36_port, regs(35) => 
                           bus_reg_dataout_35_port, regs(34) => 
                           bus_reg_dataout_34_port, regs(33) => 
                           bus_reg_dataout_33_port, regs(32) => 
                           bus_reg_dataout_32_port, regs(31) => 
                           bus_reg_dataout_31_port, regs(30) => 
                           bus_reg_dataout_30_port, regs(29) => 
                           bus_reg_dataout_29_port, regs(28) => 
                           bus_reg_dataout_28_port, regs(27) => 
                           bus_reg_dataout_27_port, regs(26) => 
                           bus_reg_dataout_26_port, regs(25) => 
                           bus_reg_dataout_25_port, regs(24) => 
                           bus_reg_dataout_24_port, regs(23) => 
                           bus_reg_dataout_23_port, regs(22) => 
                           bus_reg_dataout_22_port, regs(21) => 
                           bus_reg_dataout_21_port, regs(20) => 
                           bus_reg_dataout_20_port, regs(19) => 
                           bus_reg_dataout_19_port, regs(18) => 
                           bus_reg_dataout_18_port, regs(17) => 
                           bus_reg_dataout_17_port, regs(16) => 
                           bus_reg_dataout_16_port, regs(15) => 
                           bus_reg_dataout_15_port, regs(14) => 
                           bus_reg_dataout_14_port, regs(13) => 
                           bus_reg_dataout_13_port, regs(12) => 
                           bus_reg_dataout_12_port, regs(11) => 
                           bus_reg_dataout_11_port, regs(10) => 
                           bus_reg_dataout_10_port, regs(9) => 
                           bus_reg_dataout_9_port, regs(8) => 
                           bus_reg_dataout_8_port, regs(7) => 
                           bus_reg_dataout_7_port, regs(6) => 
                           bus_reg_dataout_6_port, regs(5) => 
                           bus_reg_dataout_5_port, regs(4) => 
                           bus_reg_dataout_4_port, regs(3) => 
                           bus_reg_dataout_3_port, regs(2) => 
                           bus_reg_dataout_2_port, regs(1) => 
                           bus_reg_dataout_1_port, regs(0) => 
                           bus_reg_dataout_0_port, win(4) => c_win_4_port, 
                           win(3) => c_win_3_port, win(2) => c_win_2_port, 
                           win(1) => c_win_1_port, win(0) => c_win_0_port, 
                           curr_proc_regs(767) => 
                           bus_selected_win_data_767_port, curr_proc_regs(766) 
                           => bus_selected_win_data_766_port, 
                           curr_proc_regs(765) => 
                           bus_selected_win_data_765_port, curr_proc_regs(764) 
                           => bus_selected_win_data_764_port, 
                           curr_proc_regs(763) => 
                           bus_selected_win_data_763_port, curr_proc_regs(762) 
                           => bus_selected_win_data_762_port, 
                           curr_proc_regs(761) => 
                           bus_selected_win_data_761_port, curr_proc_regs(760) 
                           => bus_selected_win_data_760_port, 
                           curr_proc_regs(759) => 
                           bus_selected_win_data_759_port, curr_proc_regs(758) 
                           => bus_selected_win_data_758_port, 
                           curr_proc_regs(757) => 
                           bus_selected_win_data_757_port, curr_proc_regs(756) 
                           => bus_selected_win_data_756_port, 
                           curr_proc_regs(755) => 
                           bus_selected_win_data_755_port, curr_proc_regs(754) 
                           => bus_selected_win_data_754_port, 
                           curr_proc_regs(753) => 
                           bus_selected_win_data_753_port, curr_proc_regs(752) 
                           => bus_selected_win_data_752_port, 
                           curr_proc_regs(751) => 
                           bus_selected_win_data_751_port, curr_proc_regs(750) 
                           => bus_selected_win_data_750_port, 
                           curr_proc_regs(749) => 
                           bus_selected_win_data_749_port, curr_proc_regs(748) 
                           => bus_selected_win_data_748_port, 
                           curr_proc_regs(747) => 
                           bus_selected_win_data_747_port, curr_proc_regs(746) 
                           => bus_selected_win_data_746_port, 
                           curr_proc_regs(745) => 
                           bus_selected_win_data_745_port, curr_proc_regs(744) 
                           => bus_selected_win_data_744_port, 
                           curr_proc_regs(743) => 
                           bus_selected_win_data_743_port, curr_proc_regs(742) 
                           => bus_selected_win_data_742_port, 
                           curr_proc_regs(741) => 
                           bus_selected_win_data_741_port, curr_proc_regs(740) 
                           => bus_selected_win_data_740_port, 
                           curr_proc_regs(739) => 
                           bus_selected_win_data_739_port, curr_proc_regs(738) 
                           => bus_selected_win_data_738_port, 
                           curr_proc_regs(737) => 
                           bus_selected_win_data_737_port, curr_proc_regs(736) 
                           => bus_selected_win_data_736_port, 
                           curr_proc_regs(735) => 
                           bus_selected_win_data_735_port, curr_proc_regs(734) 
                           => bus_selected_win_data_734_port, 
                           curr_proc_regs(733) => 
                           bus_selected_win_data_733_port, curr_proc_regs(732) 
                           => bus_selected_win_data_732_port, 
                           curr_proc_regs(731) => 
                           bus_selected_win_data_731_port, curr_proc_regs(730) 
                           => bus_selected_win_data_730_port, 
                           curr_proc_regs(729) => 
                           bus_selected_win_data_729_port, curr_proc_regs(728) 
                           => bus_selected_win_data_728_port, 
                           curr_proc_regs(727) => 
                           bus_selected_win_data_727_port, curr_proc_regs(726) 
                           => bus_selected_win_data_726_port, 
                           curr_proc_regs(725) => 
                           bus_selected_win_data_725_port, curr_proc_regs(724) 
                           => bus_selected_win_data_724_port, 
                           curr_proc_regs(723) => 
                           bus_selected_win_data_723_port, curr_proc_regs(722) 
                           => bus_selected_win_data_722_port, 
                           curr_proc_regs(721) => 
                           bus_selected_win_data_721_port, curr_proc_regs(720) 
                           => bus_selected_win_data_720_port, 
                           curr_proc_regs(719) => 
                           bus_selected_win_data_719_port, curr_proc_regs(718) 
                           => bus_selected_win_data_718_port, 
                           curr_proc_regs(717) => 
                           bus_selected_win_data_717_port, curr_proc_regs(716) 
                           => bus_selected_win_data_716_port, 
                           curr_proc_regs(715) => 
                           bus_selected_win_data_715_port, curr_proc_regs(714) 
                           => bus_selected_win_data_714_port, 
                           curr_proc_regs(713) => 
                           bus_selected_win_data_713_port, curr_proc_regs(712) 
                           => bus_selected_win_data_712_port, 
                           curr_proc_regs(711) => 
                           bus_selected_win_data_711_port, curr_proc_regs(710) 
                           => bus_selected_win_data_710_port, 
                           curr_proc_regs(709) => 
                           bus_selected_win_data_709_port, curr_proc_regs(708) 
                           => bus_selected_win_data_708_port, 
                           curr_proc_regs(707) => 
                           bus_selected_win_data_707_port, curr_proc_regs(706) 
                           => bus_selected_win_data_706_port, 
                           curr_proc_regs(705) => 
                           bus_selected_win_data_705_port, curr_proc_regs(704) 
                           => bus_selected_win_data_704_port, 
                           curr_proc_regs(703) => 
                           bus_selected_win_data_703_port, curr_proc_regs(702) 
                           => bus_selected_win_data_702_port, 
                           curr_proc_regs(701) => 
                           bus_selected_win_data_701_port, curr_proc_regs(700) 
                           => bus_selected_win_data_700_port, 
                           curr_proc_regs(699) => 
                           bus_selected_win_data_699_port, curr_proc_regs(698) 
                           => bus_selected_win_data_698_port, 
                           curr_proc_regs(697) => 
                           bus_selected_win_data_697_port, curr_proc_regs(696) 
                           => bus_selected_win_data_696_port, 
                           curr_proc_regs(695) => 
                           bus_selected_win_data_695_port, curr_proc_regs(694) 
                           => bus_selected_win_data_694_port, 
                           curr_proc_regs(693) => 
                           bus_selected_win_data_693_port, curr_proc_regs(692) 
                           => bus_selected_win_data_692_port, 
                           curr_proc_regs(691) => 
                           bus_selected_win_data_691_port, curr_proc_regs(690) 
                           => bus_selected_win_data_690_port, 
                           curr_proc_regs(689) => 
                           bus_selected_win_data_689_port, curr_proc_regs(688) 
                           => bus_selected_win_data_688_port, 
                           curr_proc_regs(687) => 
                           bus_selected_win_data_687_port, curr_proc_regs(686) 
                           => bus_selected_win_data_686_port, 
                           curr_proc_regs(685) => 
                           bus_selected_win_data_685_port, curr_proc_regs(684) 
                           => bus_selected_win_data_684_port, 
                           curr_proc_regs(683) => 
                           bus_selected_win_data_683_port, curr_proc_regs(682) 
                           => bus_selected_win_data_682_port, 
                           curr_proc_regs(681) => 
                           bus_selected_win_data_681_port, curr_proc_regs(680) 
                           => bus_selected_win_data_680_port, 
                           curr_proc_regs(679) => 
                           bus_selected_win_data_679_port, curr_proc_regs(678) 
                           => bus_selected_win_data_678_port, 
                           curr_proc_regs(677) => 
                           bus_selected_win_data_677_port, curr_proc_regs(676) 
                           => bus_selected_win_data_676_port, 
                           curr_proc_regs(675) => 
                           bus_selected_win_data_675_port, curr_proc_regs(674) 
                           => bus_selected_win_data_674_port, 
                           curr_proc_regs(673) => 
                           bus_selected_win_data_673_port, curr_proc_regs(672) 
                           => bus_selected_win_data_672_port, 
                           curr_proc_regs(671) => 
                           bus_selected_win_data_671_port, curr_proc_regs(670) 
                           => bus_selected_win_data_670_port, 
                           curr_proc_regs(669) => 
                           bus_selected_win_data_669_port, curr_proc_regs(668) 
                           => bus_selected_win_data_668_port, 
                           curr_proc_regs(667) => 
                           bus_selected_win_data_667_port, curr_proc_regs(666) 
                           => bus_selected_win_data_666_port, 
                           curr_proc_regs(665) => 
                           bus_selected_win_data_665_port, curr_proc_regs(664) 
                           => bus_selected_win_data_664_port, 
                           curr_proc_regs(663) => 
                           bus_selected_win_data_663_port, curr_proc_regs(662) 
                           => bus_selected_win_data_662_port, 
                           curr_proc_regs(661) => 
                           bus_selected_win_data_661_port, curr_proc_regs(660) 
                           => bus_selected_win_data_660_port, 
                           curr_proc_regs(659) => 
                           bus_selected_win_data_659_port, curr_proc_regs(658) 
                           => bus_selected_win_data_658_port, 
                           curr_proc_regs(657) => 
                           bus_selected_win_data_657_port, curr_proc_regs(656) 
                           => bus_selected_win_data_656_port, 
                           curr_proc_regs(655) => 
                           bus_selected_win_data_655_port, curr_proc_regs(654) 
                           => bus_selected_win_data_654_port, 
                           curr_proc_regs(653) => 
                           bus_selected_win_data_653_port, curr_proc_regs(652) 
                           => bus_selected_win_data_652_port, 
                           curr_proc_regs(651) => 
                           bus_selected_win_data_651_port, curr_proc_regs(650) 
                           => bus_selected_win_data_650_port, 
                           curr_proc_regs(649) => 
                           bus_selected_win_data_649_port, curr_proc_regs(648) 
                           => bus_selected_win_data_648_port, 
                           curr_proc_regs(647) => 
                           bus_selected_win_data_647_port, curr_proc_regs(646) 
                           => bus_selected_win_data_646_port, 
                           curr_proc_regs(645) => 
                           bus_selected_win_data_645_port, curr_proc_regs(644) 
                           => bus_selected_win_data_644_port, 
                           curr_proc_regs(643) => 
                           bus_selected_win_data_643_port, curr_proc_regs(642) 
                           => bus_selected_win_data_642_port, 
                           curr_proc_regs(641) => 
                           bus_selected_win_data_641_port, curr_proc_regs(640) 
                           => bus_selected_win_data_640_port, 
                           curr_proc_regs(639) => 
                           bus_selected_win_data_639_port, curr_proc_regs(638) 
                           => bus_selected_win_data_638_port, 
                           curr_proc_regs(637) => 
                           bus_selected_win_data_637_port, curr_proc_regs(636) 
                           => bus_selected_win_data_636_port, 
                           curr_proc_regs(635) => 
                           bus_selected_win_data_635_port, curr_proc_regs(634) 
                           => bus_selected_win_data_634_port, 
                           curr_proc_regs(633) => 
                           bus_selected_win_data_633_port, curr_proc_regs(632) 
                           => bus_selected_win_data_632_port, 
                           curr_proc_regs(631) => 
                           bus_selected_win_data_631_port, curr_proc_regs(630) 
                           => bus_selected_win_data_630_port, 
                           curr_proc_regs(629) => 
                           bus_selected_win_data_629_port, curr_proc_regs(628) 
                           => bus_selected_win_data_628_port, 
                           curr_proc_regs(627) => 
                           bus_selected_win_data_627_port, curr_proc_regs(626) 
                           => bus_selected_win_data_626_port, 
                           curr_proc_regs(625) => 
                           bus_selected_win_data_625_port, curr_proc_regs(624) 
                           => bus_selected_win_data_624_port, 
                           curr_proc_regs(623) => 
                           bus_selected_win_data_623_port, curr_proc_regs(622) 
                           => bus_selected_win_data_622_port, 
                           curr_proc_regs(621) => 
                           bus_selected_win_data_621_port, curr_proc_regs(620) 
                           => bus_selected_win_data_620_port, 
                           curr_proc_regs(619) => 
                           bus_selected_win_data_619_port, curr_proc_regs(618) 
                           => bus_selected_win_data_618_port, 
                           curr_proc_regs(617) => 
                           bus_selected_win_data_617_port, curr_proc_regs(616) 
                           => bus_selected_win_data_616_port, 
                           curr_proc_regs(615) => 
                           bus_selected_win_data_615_port, curr_proc_regs(614) 
                           => bus_selected_win_data_614_port, 
                           curr_proc_regs(613) => 
                           bus_selected_win_data_613_port, curr_proc_regs(612) 
                           => bus_selected_win_data_612_port, 
                           curr_proc_regs(611) => 
                           bus_selected_win_data_611_port, curr_proc_regs(610) 
                           => bus_selected_win_data_610_port, 
                           curr_proc_regs(609) => 
                           bus_selected_win_data_609_port, curr_proc_regs(608) 
                           => bus_selected_win_data_608_port, 
                           curr_proc_regs(607) => 
                           bus_selected_win_data_607_port, curr_proc_regs(606) 
                           => bus_selected_win_data_606_port, 
                           curr_proc_regs(605) => 
                           bus_selected_win_data_605_port, curr_proc_regs(604) 
                           => bus_selected_win_data_604_port, 
                           curr_proc_regs(603) => 
                           bus_selected_win_data_603_port, curr_proc_regs(602) 
                           => bus_selected_win_data_602_port, 
                           curr_proc_regs(601) => 
                           bus_selected_win_data_601_port, curr_proc_regs(600) 
                           => bus_selected_win_data_600_port, 
                           curr_proc_regs(599) => 
                           bus_selected_win_data_599_port, curr_proc_regs(598) 
                           => bus_selected_win_data_598_port, 
                           curr_proc_regs(597) => 
                           bus_selected_win_data_597_port, curr_proc_regs(596) 
                           => bus_selected_win_data_596_port, 
                           curr_proc_regs(595) => 
                           bus_selected_win_data_595_port, curr_proc_regs(594) 
                           => bus_selected_win_data_594_port, 
                           curr_proc_regs(593) => 
                           bus_selected_win_data_593_port, curr_proc_regs(592) 
                           => bus_selected_win_data_592_port, 
                           curr_proc_regs(591) => 
                           bus_selected_win_data_591_port, curr_proc_regs(590) 
                           => bus_selected_win_data_590_port, 
                           curr_proc_regs(589) => 
                           bus_selected_win_data_589_port, curr_proc_regs(588) 
                           => bus_selected_win_data_588_port, 
                           curr_proc_regs(587) => 
                           bus_selected_win_data_587_port, curr_proc_regs(586) 
                           => bus_selected_win_data_586_port, 
                           curr_proc_regs(585) => 
                           bus_selected_win_data_585_port, curr_proc_regs(584) 
                           => bus_selected_win_data_584_port, 
                           curr_proc_regs(583) => 
                           bus_selected_win_data_583_port, curr_proc_regs(582) 
                           => bus_selected_win_data_582_port, 
                           curr_proc_regs(581) => 
                           bus_selected_win_data_581_port, curr_proc_regs(580) 
                           => bus_selected_win_data_580_port, 
                           curr_proc_regs(579) => 
                           bus_selected_win_data_579_port, curr_proc_regs(578) 
                           => bus_selected_win_data_578_port, 
                           curr_proc_regs(577) => 
                           bus_selected_win_data_577_port, curr_proc_regs(576) 
                           => bus_selected_win_data_576_port, 
                           curr_proc_regs(575) => 
                           bus_selected_win_data_575_port, curr_proc_regs(574) 
                           => bus_selected_win_data_574_port, 
                           curr_proc_regs(573) => 
                           bus_selected_win_data_573_port, curr_proc_regs(572) 
                           => bus_selected_win_data_572_port, 
                           curr_proc_regs(571) => 
                           bus_selected_win_data_571_port, curr_proc_regs(570) 
                           => bus_selected_win_data_570_port, 
                           curr_proc_regs(569) => 
                           bus_selected_win_data_569_port, curr_proc_regs(568) 
                           => bus_selected_win_data_568_port, 
                           curr_proc_regs(567) => 
                           bus_selected_win_data_567_port, curr_proc_regs(566) 
                           => bus_selected_win_data_566_port, 
                           curr_proc_regs(565) => 
                           bus_selected_win_data_565_port, curr_proc_regs(564) 
                           => bus_selected_win_data_564_port, 
                           curr_proc_regs(563) => 
                           bus_selected_win_data_563_port, curr_proc_regs(562) 
                           => bus_selected_win_data_562_port, 
                           curr_proc_regs(561) => 
                           bus_selected_win_data_561_port, curr_proc_regs(560) 
                           => bus_selected_win_data_560_port, 
                           curr_proc_regs(559) => 
                           bus_selected_win_data_559_port, curr_proc_regs(558) 
                           => bus_selected_win_data_558_port, 
                           curr_proc_regs(557) => 
                           bus_selected_win_data_557_port, curr_proc_regs(556) 
                           => bus_selected_win_data_556_port, 
                           curr_proc_regs(555) => 
                           bus_selected_win_data_555_port, curr_proc_regs(554) 
                           => bus_selected_win_data_554_port, 
                           curr_proc_regs(553) => 
                           bus_selected_win_data_553_port, curr_proc_regs(552) 
                           => bus_selected_win_data_552_port, 
                           curr_proc_regs(551) => 
                           bus_selected_win_data_551_port, curr_proc_regs(550) 
                           => bus_selected_win_data_550_port, 
                           curr_proc_regs(549) => 
                           bus_selected_win_data_549_port, curr_proc_regs(548) 
                           => bus_selected_win_data_548_port, 
                           curr_proc_regs(547) => 
                           bus_selected_win_data_547_port, curr_proc_regs(546) 
                           => bus_selected_win_data_546_port, 
                           curr_proc_regs(545) => 
                           bus_selected_win_data_545_port, curr_proc_regs(544) 
                           => bus_selected_win_data_544_port, 
                           curr_proc_regs(543) => 
                           bus_selected_win_data_543_port, curr_proc_regs(542) 
                           => bus_selected_win_data_542_port, 
                           curr_proc_regs(541) => 
                           bus_selected_win_data_541_port, curr_proc_regs(540) 
                           => bus_selected_win_data_540_port, 
                           curr_proc_regs(539) => 
                           bus_selected_win_data_539_port, curr_proc_regs(538) 
                           => bus_selected_win_data_538_port, 
                           curr_proc_regs(537) => 
                           bus_selected_win_data_537_port, curr_proc_regs(536) 
                           => bus_selected_win_data_536_port, 
                           curr_proc_regs(535) => 
                           bus_selected_win_data_535_port, curr_proc_regs(534) 
                           => bus_selected_win_data_534_port, 
                           curr_proc_regs(533) => 
                           bus_selected_win_data_533_port, curr_proc_regs(532) 
                           => bus_selected_win_data_532_port, 
                           curr_proc_regs(531) => 
                           bus_selected_win_data_531_port, curr_proc_regs(530) 
                           => bus_selected_win_data_530_port, 
                           curr_proc_regs(529) => 
                           bus_selected_win_data_529_port, curr_proc_regs(528) 
                           => bus_selected_win_data_528_port, 
                           curr_proc_regs(527) => 
                           bus_selected_win_data_527_port, curr_proc_regs(526) 
                           => bus_selected_win_data_526_port, 
                           curr_proc_regs(525) => 
                           bus_selected_win_data_525_port, curr_proc_regs(524) 
                           => bus_selected_win_data_524_port, 
                           curr_proc_regs(523) => 
                           bus_selected_win_data_523_port, curr_proc_regs(522) 
                           => bus_selected_win_data_522_port, 
                           curr_proc_regs(521) => 
                           bus_selected_win_data_521_port, curr_proc_regs(520) 
                           => bus_selected_win_data_520_port, 
                           curr_proc_regs(519) => 
                           bus_selected_win_data_519_port, curr_proc_regs(518) 
                           => bus_selected_win_data_518_port, 
                           curr_proc_regs(517) => 
                           bus_selected_win_data_517_port, curr_proc_regs(516) 
                           => bus_selected_win_data_516_port, 
                           curr_proc_regs(515) => 
                           bus_selected_win_data_515_port, curr_proc_regs(514) 
                           => bus_selected_win_data_514_port, 
                           curr_proc_regs(513) => 
                           bus_selected_win_data_513_port, curr_proc_regs(512) 
                           => bus_selected_win_data_512_port, 
                           curr_proc_regs(511) => 
                           bus_selected_win_data_511_port, curr_proc_regs(510) 
                           => bus_selected_win_data_510_port, 
                           curr_proc_regs(509) => 
                           bus_selected_win_data_509_port, curr_proc_regs(508) 
                           => bus_selected_win_data_508_port, 
                           curr_proc_regs(507) => 
                           bus_selected_win_data_507_port, curr_proc_regs(506) 
                           => bus_selected_win_data_506_port, 
                           curr_proc_regs(505) => 
                           bus_selected_win_data_505_port, curr_proc_regs(504) 
                           => bus_selected_win_data_504_port, 
                           curr_proc_regs(503) => 
                           bus_selected_win_data_503_port, curr_proc_regs(502) 
                           => bus_selected_win_data_502_port, 
                           curr_proc_regs(501) => 
                           bus_selected_win_data_501_port, curr_proc_regs(500) 
                           => bus_selected_win_data_500_port, 
                           curr_proc_regs(499) => 
                           bus_selected_win_data_499_port, curr_proc_regs(498) 
                           => bus_selected_win_data_498_port, 
                           curr_proc_regs(497) => 
                           bus_selected_win_data_497_port, curr_proc_regs(496) 
                           => bus_selected_win_data_496_port, 
                           curr_proc_regs(495) => 
                           bus_selected_win_data_495_port, curr_proc_regs(494) 
                           => bus_selected_win_data_494_port, 
                           curr_proc_regs(493) => 
                           bus_selected_win_data_493_port, curr_proc_regs(492) 
                           => bus_selected_win_data_492_port, 
                           curr_proc_regs(491) => 
                           bus_selected_win_data_491_port, curr_proc_regs(490) 
                           => bus_selected_win_data_490_port, 
                           curr_proc_regs(489) => 
                           bus_selected_win_data_489_port, curr_proc_regs(488) 
                           => bus_selected_win_data_488_port, 
                           curr_proc_regs(487) => 
                           bus_selected_win_data_487_port, curr_proc_regs(486) 
                           => bus_selected_win_data_486_port, 
                           curr_proc_regs(485) => 
                           bus_selected_win_data_485_port, curr_proc_regs(484) 
                           => bus_selected_win_data_484_port, 
                           curr_proc_regs(483) => 
                           bus_selected_win_data_483_port, curr_proc_regs(482) 
                           => bus_selected_win_data_482_port, 
                           curr_proc_regs(481) => 
                           bus_selected_win_data_481_port, curr_proc_regs(480) 
                           => bus_selected_win_data_480_port, 
                           curr_proc_regs(479) => 
                           bus_selected_win_data_479_port, curr_proc_regs(478) 
                           => bus_selected_win_data_478_port, 
                           curr_proc_regs(477) => 
                           bus_selected_win_data_477_port, curr_proc_regs(476) 
                           => bus_selected_win_data_476_port, 
                           curr_proc_regs(475) => 
                           bus_selected_win_data_475_port, curr_proc_regs(474) 
                           => bus_selected_win_data_474_port, 
                           curr_proc_regs(473) => 
                           bus_selected_win_data_473_port, curr_proc_regs(472) 
                           => bus_selected_win_data_472_port, 
                           curr_proc_regs(471) => 
                           bus_selected_win_data_471_port, curr_proc_regs(470) 
                           => bus_selected_win_data_470_port, 
                           curr_proc_regs(469) => 
                           bus_selected_win_data_469_port, curr_proc_regs(468) 
                           => bus_selected_win_data_468_port, 
                           curr_proc_regs(467) => 
                           bus_selected_win_data_467_port, curr_proc_regs(466) 
                           => bus_selected_win_data_466_port, 
                           curr_proc_regs(465) => 
                           bus_selected_win_data_465_port, curr_proc_regs(464) 
                           => bus_selected_win_data_464_port, 
                           curr_proc_regs(463) => 
                           bus_selected_win_data_463_port, curr_proc_regs(462) 
                           => bus_selected_win_data_462_port, 
                           curr_proc_regs(461) => 
                           bus_selected_win_data_461_port, curr_proc_regs(460) 
                           => bus_selected_win_data_460_port, 
                           curr_proc_regs(459) => 
                           bus_selected_win_data_459_port, curr_proc_regs(458) 
                           => bus_selected_win_data_458_port, 
                           curr_proc_regs(457) => 
                           bus_selected_win_data_457_port, curr_proc_regs(456) 
                           => bus_selected_win_data_456_port, 
                           curr_proc_regs(455) => 
                           bus_selected_win_data_455_port, curr_proc_regs(454) 
                           => bus_selected_win_data_454_port, 
                           curr_proc_regs(453) => 
                           bus_selected_win_data_453_port, curr_proc_regs(452) 
                           => bus_selected_win_data_452_port, 
                           curr_proc_regs(451) => 
                           bus_selected_win_data_451_port, curr_proc_regs(450) 
                           => bus_selected_win_data_450_port, 
                           curr_proc_regs(449) => 
                           bus_selected_win_data_449_port, curr_proc_regs(448) 
                           => bus_selected_win_data_448_port, 
                           curr_proc_regs(447) => 
                           bus_selected_win_data_447_port, curr_proc_regs(446) 
                           => bus_selected_win_data_446_port, 
                           curr_proc_regs(445) => 
                           bus_selected_win_data_445_port, curr_proc_regs(444) 
                           => bus_selected_win_data_444_port, 
                           curr_proc_regs(443) => 
                           bus_selected_win_data_443_port, curr_proc_regs(442) 
                           => bus_selected_win_data_442_port, 
                           curr_proc_regs(441) => 
                           bus_selected_win_data_441_port, curr_proc_regs(440) 
                           => bus_selected_win_data_440_port, 
                           curr_proc_regs(439) => 
                           bus_selected_win_data_439_port, curr_proc_regs(438) 
                           => bus_selected_win_data_438_port, 
                           curr_proc_regs(437) => 
                           bus_selected_win_data_437_port, curr_proc_regs(436) 
                           => bus_selected_win_data_436_port, 
                           curr_proc_regs(435) => 
                           bus_selected_win_data_435_port, curr_proc_regs(434) 
                           => bus_selected_win_data_434_port, 
                           curr_proc_regs(433) => 
                           bus_selected_win_data_433_port, curr_proc_regs(432) 
                           => bus_selected_win_data_432_port, 
                           curr_proc_regs(431) => 
                           bus_selected_win_data_431_port, curr_proc_regs(430) 
                           => bus_selected_win_data_430_port, 
                           curr_proc_regs(429) => 
                           bus_selected_win_data_429_port, curr_proc_regs(428) 
                           => bus_selected_win_data_428_port, 
                           curr_proc_regs(427) => 
                           bus_selected_win_data_427_port, curr_proc_regs(426) 
                           => bus_selected_win_data_426_port, 
                           curr_proc_regs(425) => 
                           bus_selected_win_data_425_port, curr_proc_regs(424) 
                           => bus_selected_win_data_424_port, 
                           curr_proc_regs(423) => 
                           bus_selected_win_data_423_port, curr_proc_regs(422) 
                           => bus_selected_win_data_422_port, 
                           curr_proc_regs(421) => 
                           bus_selected_win_data_421_port, curr_proc_regs(420) 
                           => bus_selected_win_data_420_port, 
                           curr_proc_regs(419) => 
                           bus_selected_win_data_419_port, curr_proc_regs(418) 
                           => bus_selected_win_data_418_port, 
                           curr_proc_regs(417) => 
                           bus_selected_win_data_417_port, curr_proc_regs(416) 
                           => bus_selected_win_data_416_port, 
                           curr_proc_regs(415) => 
                           bus_selected_win_data_415_port, curr_proc_regs(414) 
                           => bus_selected_win_data_414_port, 
                           curr_proc_regs(413) => 
                           bus_selected_win_data_413_port, curr_proc_regs(412) 
                           => bus_selected_win_data_412_port, 
                           curr_proc_regs(411) => 
                           bus_selected_win_data_411_port, curr_proc_regs(410) 
                           => bus_selected_win_data_410_port, 
                           curr_proc_regs(409) => 
                           bus_selected_win_data_409_port, curr_proc_regs(408) 
                           => bus_selected_win_data_408_port, 
                           curr_proc_regs(407) => 
                           bus_selected_win_data_407_port, curr_proc_regs(406) 
                           => bus_selected_win_data_406_port, 
                           curr_proc_regs(405) => 
                           bus_selected_win_data_405_port, curr_proc_regs(404) 
                           => bus_selected_win_data_404_port, 
                           curr_proc_regs(403) => 
                           bus_selected_win_data_403_port, curr_proc_regs(402) 
                           => bus_selected_win_data_402_port, 
                           curr_proc_regs(401) => 
                           bus_selected_win_data_401_port, curr_proc_regs(400) 
                           => bus_selected_win_data_400_port, 
                           curr_proc_regs(399) => 
                           bus_selected_win_data_399_port, curr_proc_regs(398) 
                           => bus_selected_win_data_398_port, 
                           curr_proc_regs(397) => 
                           bus_selected_win_data_397_port, curr_proc_regs(396) 
                           => bus_selected_win_data_396_port, 
                           curr_proc_regs(395) => 
                           bus_selected_win_data_395_port, curr_proc_regs(394) 
                           => bus_selected_win_data_394_port, 
                           curr_proc_regs(393) => 
                           bus_selected_win_data_393_port, curr_proc_regs(392) 
                           => bus_selected_win_data_392_port, 
                           curr_proc_regs(391) => 
                           bus_selected_win_data_391_port, curr_proc_regs(390) 
                           => bus_selected_win_data_390_port, 
                           curr_proc_regs(389) => 
                           bus_selected_win_data_389_port, curr_proc_regs(388) 
                           => bus_selected_win_data_388_port, 
                           curr_proc_regs(387) => 
                           bus_selected_win_data_387_port, curr_proc_regs(386) 
                           => bus_selected_win_data_386_port, 
                           curr_proc_regs(385) => 
                           bus_selected_win_data_385_port, curr_proc_regs(384) 
                           => bus_selected_win_data_384_port, 
                           curr_proc_regs(383) => 
                           bus_selected_win_data_383_port, curr_proc_regs(382) 
                           => bus_selected_win_data_382_port, 
                           curr_proc_regs(381) => 
                           bus_selected_win_data_381_port, curr_proc_regs(380) 
                           => bus_selected_win_data_380_port, 
                           curr_proc_regs(379) => 
                           bus_selected_win_data_379_port, curr_proc_regs(378) 
                           => bus_selected_win_data_378_port, 
                           curr_proc_regs(377) => 
                           bus_selected_win_data_377_port, curr_proc_regs(376) 
                           => bus_selected_win_data_376_port, 
                           curr_proc_regs(375) => 
                           bus_selected_win_data_375_port, curr_proc_regs(374) 
                           => bus_selected_win_data_374_port, 
                           curr_proc_regs(373) => 
                           bus_selected_win_data_373_port, curr_proc_regs(372) 
                           => bus_selected_win_data_372_port, 
                           curr_proc_regs(371) => 
                           bus_selected_win_data_371_port, curr_proc_regs(370) 
                           => bus_selected_win_data_370_port, 
                           curr_proc_regs(369) => 
                           bus_selected_win_data_369_port, curr_proc_regs(368) 
                           => bus_selected_win_data_368_port, 
                           curr_proc_regs(367) => 
                           bus_selected_win_data_367_port, curr_proc_regs(366) 
                           => bus_selected_win_data_366_port, 
                           curr_proc_regs(365) => 
                           bus_selected_win_data_365_port, curr_proc_regs(364) 
                           => bus_selected_win_data_364_port, 
                           curr_proc_regs(363) => 
                           bus_selected_win_data_363_port, curr_proc_regs(362) 
                           => bus_selected_win_data_362_port, 
                           curr_proc_regs(361) => 
                           bus_selected_win_data_361_port, curr_proc_regs(360) 
                           => bus_selected_win_data_360_port, 
                           curr_proc_regs(359) => 
                           bus_selected_win_data_359_port, curr_proc_regs(358) 
                           => bus_selected_win_data_358_port, 
                           curr_proc_regs(357) => 
                           bus_selected_win_data_357_port, curr_proc_regs(356) 
                           => bus_selected_win_data_356_port, 
                           curr_proc_regs(355) => 
                           bus_selected_win_data_355_port, curr_proc_regs(354) 
                           => bus_selected_win_data_354_port, 
                           curr_proc_regs(353) => 
                           bus_selected_win_data_353_port, curr_proc_regs(352) 
                           => bus_selected_win_data_352_port, 
                           curr_proc_regs(351) => 
                           bus_selected_win_data_351_port, curr_proc_regs(350) 
                           => bus_selected_win_data_350_port, 
                           curr_proc_regs(349) => 
                           bus_selected_win_data_349_port, curr_proc_regs(348) 
                           => bus_selected_win_data_348_port, 
                           curr_proc_regs(347) => 
                           bus_selected_win_data_347_port, curr_proc_regs(346) 
                           => bus_selected_win_data_346_port, 
                           curr_proc_regs(345) => 
                           bus_selected_win_data_345_port, curr_proc_regs(344) 
                           => bus_selected_win_data_344_port, 
                           curr_proc_regs(343) => 
                           bus_selected_win_data_343_port, curr_proc_regs(342) 
                           => bus_selected_win_data_342_port, 
                           curr_proc_regs(341) => 
                           bus_selected_win_data_341_port, curr_proc_regs(340) 
                           => bus_selected_win_data_340_port, 
                           curr_proc_regs(339) => 
                           bus_selected_win_data_339_port, curr_proc_regs(338) 
                           => bus_selected_win_data_338_port, 
                           curr_proc_regs(337) => 
                           bus_selected_win_data_337_port, curr_proc_regs(336) 
                           => bus_selected_win_data_336_port, 
                           curr_proc_regs(335) => 
                           bus_selected_win_data_335_port, curr_proc_regs(334) 
                           => bus_selected_win_data_334_port, 
                           curr_proc_regs(333) => 
                           bus_selected_win_data_333_port, curr_proc_regs(332) 
                           => bus_selected_win_data_332_port, 
                           curr_proc_regs(331) => 
                           bus_selected_win_data_331_port, curr_proc_regs(330) 
                           => bus_selected_win_data_330_port, 
                           curr_proc_regs(329) => 
                           bus_selected_win_data_329_port, curr_proc_regs(328) 
                           => bus_selected_win_data_328_port, 
                           curr_proc_regs(327) => 
                           bus_selected_win_data_327_port, curr_proc_regs(326) 
                           => bus_selected_win_data_326_port, 
                           curr_proc_regs(325) => 
                           bus_selected_win_data_325_port, curr_proc_regs(324) 
                           => bus_selected_win_data_324_port, 
                           curr_proc_regs(323) => 
                           bus_selected_win_data_323_port, curr_proc_regs(322) 
                           => bus_selected_win_data_322_port, 
                           curr_proc_regs(321) => 
                           bus_selected_win_data_321_port, curr_proc_regs(320) 
                           => bus_selected_win_data_320_port, 
                           curr_proc_regs(319) => 
                           bus_selected_win_data_319_port, curr_proc_regs(318) 
                           => bus_selected_win_data_318_port, 
                           curr_proc_regs(317) => 
                           bus_selected_win_data_317_port, curr_proc_regs(316) 
                           => bus_selected_win_data_316_port, 
                           curr_proc_regs(315) => 
                           bus_selected_win_data_315_port, curr_proc_regs(314) 
                           => bus_selected_win_data_314_port, 
                           curr_proc_regs(313) => 
                           bus_selected_win_data_313_port, curr_proc_regs(312) 
                           => bus_selected_win_data_312_port, 
                           curr_proc_regs(311) => 
                           bus_selected_win_data_311_port, curr_proc_regs(310) 
                           => bus_selected_win_data_310_port, 
                           curr_proc_regs(309) => 
                           bus_selected_win_data_309_port, curr_proc_regs(308) 
                           => bus_selected_win_data_308_port, 
                           curr_proc_regs(307) => 
                           bus_selected_win_data_307_port, curr_proc_regs(306) 
                           => bus_selected_win_data_306_port, 
                           curr_proc_regs(305) => 
                           bus_selected_win_data_305_port, curr_proc_regs(304) 
                           => bus_selected_win_data_304_port, 
                           curr_proc_regs(303) => 
                           bus_selected_win_data_303_port, curr_proc_regs(302) 
                           => bus_selected_win_data_302_port, 
                           curr_proc_regs(301) => 
                           bus_selected_win_data_301_port, curr_proc_regs(300) 
                           => bus_selected_win_data_300_port, 
                           curr_proc_regs(299) => 
                           bus_selected_win_data_299_port, curr_proc_regs(298) 
                           => bus_selected_win_data_298_port, 
                           curr_proc_regs(297) => 
                           bus_selected_win_data_297_port, curr_proc_regs(296) 
                           => bus_selected_win_data_296_port, 
                           curr_proc_regs(295) => 
                           bus_selected_win_data_295_port, curr_proc_regs(294) 
                           => bus_selected_win_data_294_port, 
                           curr_proc_regs(293) => 
                           bus_selected_win_data_293_port, curr_proc_regs(292) 
                           => bus_selected_win_data_292_port, 
                           curr_proc_regs(291) => 
                           bus_selected_win_data_291_port, curr_proc_regs(290) 
                           => bus_selected_win_data_290_port, 
                           curr_proc_regs(289) => 
                           bus_selected_win_data_289_port, curr_proc_regs(288) 
                           => bus_selected_win_data_288_port, 
                           curr_proc_regs(287) => 
                           bus_selected_win_data_287_port, curr_proc_regs(286) 
                           => bus_selected_win_data_286_port, 
                           curr_proc_regs(285) => 
                           bus_selected_win_data_285_port, curr_proc_regs(284) 
                           => bus_selected_win_data_284_port, 
                           curr_proc_regs(283) => 
                           bus_selected_win_data_283_port, curr_proc_regs(282) 
                           => bus_selected_win_data_282_port, 
                           curr_proc_regs(281) => 
                           bus_selected_win_data_281_port, curr_proc_regs(280) 
                           => bus_selected_win_data_280_port, 
                           curr_proc_regs(279) => 
                           bus_selected_win_data_279_port, curr_proc_regs(278) 
                           => bus_selected_win_data_278_port, 
                           curr_proc_regs(277) => 
                           bus_selected_win_data_277_port, curr_proc_regs(276) 
                           => bus_selected_win_data_276_port, 
                           curr_proc_regs(275) => 
                           bus_selected_win_data_275_port, curr_proc_regs(274) 
                           => bus_selected_win_data_274_port, 
                           curr_proc_regs(273) => 
                           bus_selected_win_data_273_port, curr_proc_regs(272) 
                           => bus_selected_win_data_272_port, 
                           curr_proc_regs(271) => 
                           bus_selected_win_data_271_port, curr_proc_regs(270) 
                           => bus_selected_win_data_270_port, 
                           curr_proc_regs(269) => 
                           bus_selected_win_data_269_port, curr_proc_regs(268) 
                           => bus_selected_win_data_268_port, 
                           curr_proc_regs(267) => 
                           bus_selected_win_data_267_port, curr_proc_regs(266) 
                           => bus_selected_win_data_266_port, 
                           curr_proc_regs(265) => 
                           bus_selected_win_data_265_port, curr_proc_regs(264) 
                           => bus_selected_win_data_264_port, 
                           curr_proc_regs(263) => 
                           bus_selected_win_data_263_port, curr_proc_regs(262) 
                           => bus_selected_win_data_262_port, 
                           curr_proc_regs(261) => 
                           bus_selected_win_data_261_port, curr_proc_regs(260) 
                           => bus_selected_win_data_260_port, 
                           curr_proc_regs(259) => 
                           bus_selected_win_data_259_port, curr_proc_regs(258) 
                           => bus_selected_win_data_258_port, 
                           curr_proc_regs(257) => 
                           bus_selected_win_data_257_port, curr_proc_regs(256) 
                           => bus_selected_win_data_256_port, 
                           curr_proc_regs(255) => 
                           bus_selected_win_data_255_port, curr_proc_regs(254) 
                           => bus_selected_win_data_254_port, 
                           curr_proc_regs(253) => 
                           bus_selected_win_data_253_port, curr_proc_regs(252) 
                           => bus_selected_win_data_252_port, 
                           curr_proc_regs(251) => 
                           bus_selected_win_data_251_port, curr_proc_regs(250) 
                           => bus_selected_win_data_250_port, 
                           curr_proc_regs(249) => 
                           bus_selected_win_data_249_port, curr_proc_regs(248) 
                           => bus_selected_win_data_248_port, 
                           curr_proc_regs(247) => 
                           bus_selected_win_data_247_port, curr_proc_regs(246) 
                           => bus_selected_win_data_246_port, 
                           curr_proc_regs(245) => 
                           bus_selected_win_data_245_port, curr_proc_regs(244) 
                           => bus_selected_win_data_244_port, 
                           curr_proc_regs(243) => 
                           bus_selected_win_data_243_port, curr_proc_regs(242) 
                           => bus_selected_win_data_242_port, 
                           curr_proc_regs(241) => 
                           bus_selected_win_data_241_port, curr_proc_regs(240) 
                           => bus_selected_win_data_240_port, 
                           curr_proc_regs(239) => 
                           bus_selected_win_data_239_port, curr_proc_regs(238) 
                           => bus_selected_win_data_238_port, 
                           curr_proc_regs(237) => 
                           bus_selected_win_data_237_port, curr_proc_regs(236) 
                           => bus_selected_win_data_236_port, 
                           curr_proc_regs(235) => 
                           bus_selected_win_data_235_port, curr_proc_regs(234) 
                           => bus_selected_win_data_234_port, 
                           curr_proc_regs(233) => 
                           bus_selected_win_data_233_port, curr_proc_regs(232) 
                           => bus_selected_win_data_232_port, 
                           curr_proc_regs(231) => 
                           bus_selected_win_data_231_port, curr_proc_regs(230) 
                           => bus_selected_win_data_230_port, 
                           curr_proc_regs(229) => 
                           bus_selected_win_data_229_port, curr_proc_regs(228) 
                           => bus_selected_win_data_228_port, 
                           curr_proc_regs(227) => 
                           bus_selected_win_data_227_port, curr_proc_regs(226) 
                           => bus_selected_win_data_226_port, 
                           curr_proc_regs(225) => 
                           bus_selected_win_data_225_port, curr_proc_regs(224) 
                           => bus_selected_win_data_224_port, 
                           curr_proc_regs(223) => 
                           bus_selected_win_data_223_port, curr_proc_regs(222) 
                           => bus_selected_win_data_222_port, 
                           curr_proc_regs(221) => 
                           bus_selected_win_data_221_port, curr_proc_regs(220) 
                           => bus_selected_win_data_220_port, 
                           curr_proc_regs(219) => 
                           bus_selected_win_data_219_port, curr_proc_regs(218) 
                           => bus_selected_win_data_218_port, 
                           curr_proc_regs(217) => 
                           bus_selected_win_data_217_port, curr_proc_regs(216) 
                           => bus_selected_win_data_216_port, 
                           curr_proc_regs(215) => 
                           bus_selected_win_data_215_port, curr_proc_regs(214) 
                           => bus_selected_win_data_214_port, 
                           curr_proc_regs(213) => 
                           bus_selected_win_data_213_port, curr_proc_regs(212) 
                           => bus_selected_win_data_212_port, 
                           curr_proc_regs(211) => 
                           bus_selected_win_data_211_port, curr_proc_regs(210) 
                           => bus_selected_win_data_210_port, 
                           curr_proc_regs(209) => 
                           bus_selected_win_data_209_port, curr_proc_regs(208) 
                           => bus_selected_win_data_208_port, 
                           curr_proc_regs(207) => 
                           bus_selected_win_data_207_port, curr_proc_regs(206) 
                           => bus_selected_win_data_206_port, 
                           curr_proc_regs(205) => 
                           bus_selected_win_data_205_port, curr_proc_regs(204) 
                           => bus_selected_win_data_204_port, 
                           curr_proc_regs(203) => 
                           bus_selected_win_data_203_port, curr_proc_regs(202) 
                           => bus_selected_win_data_202_port, 
                           curr_proc_regs(201) => 
                           bus_selected_win_data_201_port, curr_proc_regs(200) 
                           => bus_selected_win_data_200_port, 
                           curr_proc_regs(199) => 
                           bus_selected_win_data_199_port, curr_proc_regs(198) 
                           => bus_selected_win_data_198_port, 
                           curr_proc_regs(197) => 
                           bus_selected_win_data_197_port, curr_proc_regs(196) 
                           => bus_selected_win_data_196_port, 
                           curr_proc_regs(195) => 
                           bus_selected_win_data_195_port, curr_proc_regs(194) 
                           => bus_selected_win_data_194_port, 
                           curr_proc_regs(193) => 
                           bus_selected_win_data_193_port, curr_proc_regs(192) 
                           => bus_selected_win_data_192_port, 
                           curr_proc_regs(191) => 
                           bus_selected_win_data_191_port, curr_proc_regs(190) 
                           => bus_selected_win_data_190_port, 
                           curr_proc_regs(189) => 
                           bus_selected_win_data_189_port, curr_proc_regs(188) 
                           => bus_selected_win_data_188_port, 
                           curr_proc_regs(187) => 
                           bus_selected_win_data_187_port, curr_proc_regs(186) 
                           => bus_selected_win_data_186_port, 
                           curr_proc_regs(185) => 
                           bus_selected_win_data_185_port, curr_proc_regs(184) 
                           => bus_selected_win_data_184_port, 
                           curr_proc_regs(183) => 
                           bus_selected_win_data_183_port, curr_proc_regs(182) 
                           => bus_selected_win_data_182_port, 
                           curr_proc_regs(181) => 
                           bus_selected_win_data_181_port, curr_proc_regs(180) 
                           => bus_selected_win_data_180_port, 
                           curr_proc_regs(179) => 
                           bus_selected_win_data_179_port, curr_proc_regs(178) 
                           => bus_selected_win_data_178_port, 
                           curr_proc_regs(177) => 
                           bus_selected_win_data_177_port, curr_proc_regs(176) 
                           => bus_selected_win_data_176_port, 
                           curr_proc_regs(175) => 
                           bus_selected_win_data_175_port, curr_proc_regs(174) 
                           => bus_selected_win_data_174_port, 
                           curr_proc_regs(173) => 
                           bus_selected_win_data_173_port, curr_proc_regs(172) 
                           => bus_selected_win_data_172_port, 
                           curr_proc_regs(171) => 
                           bus_selected_win_data_171_port, curr_proc_regs(170) 
                           => bus_selected_win_data_170_port, 
                           curr_proc_regs(169) => 
                           bus_selected_win_data_169_port, curr_proc_regs(168) 
                           => bus_selected_win_data_168_port, 
                           curr_proc_regs(167) => 
                           bus_selected_win_data_167_port, curr_proc_regs(166) 
                           => bus_selected_win_data_166_port, 
                           curr_proc_regs(165) => 
                           bus_selected_win_data_165_port, curr_proc_regs(164) 
                           => bus_selected_win_data_164_port, 
                           curr_proc_regs(163) => 
                           bus_selected_win_data_163_port, curr_proc_regs(162) 
                           => bus_selected_win_data_162_port, 
                           curr_proc_regs(161) => 
                           bus_selected_win_data_161_port, curr_proc_regs(160) 
                           => bus_selected_win_data_160_port, 
                           curr_proc_regs(159) => 
                           bus_selected_win_data_159_port, curr_proc_regs(158) 
                           => bus_selected_win_data_158_port, 
                           curr_proc_regs(157) => 
                           bus_selected_win_data_157_port, curr_proc_regs(156) 
                           => bus_selected_win_data_156_port, 
                           curr_proc_regs(155) => 
                           bus_selected_win_data_155_port, curr_proc_regs(154) 
                           => bus_selected_win_data_154_port, 
                           curr_proc_regs(153) => 
                           bus_selected_win_data_153_port, curr_proc_regs(152) 
                           => bus_selected_win_data_152_port, 
                           curr_proc_regs(151) => 
                           bus_selected_win_data_151_port, curr_proc_regs(150) 
                           => bus_selected_win_data_150_port, 
                           curr_proc_regs(149) => 
                           bus_selected_win_data_149_port, curr_proc_regs(148) 
                           => bus_selected_win_data_148_port, 
                           curr_proc_regs(147) => 
                           bus_selected_win_data_147_port, curr_proc_regs(146) 
                           => bus_selected_win_data_146_port, 
                           curr_proc_regs(145) => 
                           bus_selected_win_data_145_port, curr_proc_regs(144) 
                           => bus_selected_win_data_144_port, 
                           curr_proc_regs(143) => 
                           bus_selected_win_data_143_port, curr_proc_regs(142) 
                           => bus_selected_win_data_142_port, 
                           curr_proc_regs(141) => 
                           bus_selected_win_data_141_port, curr_proc_regs(140) 
                           => bus_selected_win_data_140_port, 
                           curr_proc_regs(139) => 
                           bus_selected_win_data_139_port, curr_proc_regs(138) 
                           => bus_selected_win_data_138_port, 
                           curr_proc_regs(137) => 
                           bus_selected_win_data_137_port, curr_proc_regs(136) 
                           => bus_selected_win_data_136_port, 
                           curr_proc_regs(135) => 
                           bus_selected_win_data_135_port, curr_proc_regs(134) 
                           => bus_selected_win_data_134_port, 
                           curr_proc_regs(133) => 
                           bus_selected_win_data_133_port, curr_proc_regs(132) 
                           => bus_selected_win_data_132_port, 
                           curr_proc_regs(131) => 
                           bus_selected_win_data_131_port, curr_proc_regs(130) 
                           => bus_selected_win_data_130_port, 
                           curr_proc_regs(129) => 
                           bus_selected_win_data_129_port, curr_proc_regs(128) 
                           => bus_selected_win_data_128_port, 
                           curr_proc_regs(127) => 
                           bus_selected_win_data_127_port, curr_proc_regs(126) 
                           => bus_selected_win_data_126_port, 
                           curr_proc_regs(125) => 
                           bus_selected_win_data_125_port, curr_proc_regs(124) 
                           => bus_selected_win_data_124_port, 
                           curr_proc_regs(123) => 
                           bus_selected_win_data_123_port, curr_proc_regs(122) 
                           => bus_selected_win_data_122_port, 
                           curr_proc_regs(121) => 
                           bus_selected_win_data_121_port, curr_proc_regs(120) 
                           => bus_selected_win_data_120_port, 
                           curr_proc_regs(119) => 
                           bus_selected_win_data_119_port, curr_proc_regs(118) 
                           => bus_selected_win_data_118_port, 
                           curr_proc_regs(117) => 
                           bus_selected_win_data_117_port, curr_proc_regs(116) 
                           => bus_selected_win_data_116_port, 
                           curr_proc_regs(115) => 
                           bus_selected_win_data_115_port, curr_proc_regs(114) 
                           => bus_selected_win_data_114_port, 
                           curr_proc_regs(113) => 
                           bus_selected_win_data_113_port, curr_proc_regs(112) 
                           => bus_selected_win_data_112_port, 
                           curr_proc_regs(111) => 
                           bus_selected_win_data_111_port, curr_proc_regs(110) 
                           => bus_selected_win_data_110_port, 
                           curr_proc_regs(109) => 
                           bus_selected_win_data_109_port, curr_proc_regs(108) 
                           => bus_selected_win_data_108_port, 
                           curr_proc_regs(107) => 
                           bus_selected_win_data_107_port, curr_proc_regs(106) 
                           => bus_selected_win_data_106_port, 
                           curr_proc_regs(105) => 
                           bus_selected_win_data_105_port, curr_proc_regs(104) 
                           => bus_selected_win_data_104_port, 
                           curr_proc_regs(103) => 
                           bus_selected_win_data_103_port, curr_proc_regs(102) 
                           => bus_selected_win_data_102_port, 
                           curr_proc_regs(101) => 
                           bus_selected_win_data_101_port, curr_proc_regs(100) 
                           => bus_selected_win_data_100_port, 
                           curr_proc_regs(99) => bus_selected_win_data_99_port,
                           curr_proc_regs(98) => bus_selected_win_data_98_port,
                           curr_proc_regs(97) => bus_selected_win_data_97_port,
                           curr_proc_regs(96) => bus_selected_win_data_96_port,
                           curr_proc_regs(95) => bus_selected_win_data_95_port,
                           curr_proc_regs(94) => bus_selected_win_data_94_port,
                           curr_proc_regs(93) => bus_selected_win_data_93_port,
                           curr_proc_regs(92) => bus_selected_win_data_92_port,
                           curr_proc_regs(91) => bus_selected_win_data_91_port,
                           curr_proc_regs(90) => bus_selected_win_data_90_port,
                           curr_proc_regs(89) => bus_selected_win_data_89_port,
                           curr_proc_regs(88) => bus_selected_win_data_88_port,
                           curr_proc_regs(87) => bus_selected_win_data_87_port,
                           curr_proc_regs(86) => bus_selected_win_data_86_port,
                           curr_proc_regs(85) => bus_selected_win_data_85_port,
                           curr_proc_regs(84) => bus_selected_win_data_84_port,
                           curr_proc_regs(83) => bus_selected_win_data_83_port,
                           curr_proc_regs(82) => bus_selected_win_data_82_port,
                           curr_proc_regs(81) => bus_selected_win_data_81_port,
                           curr_proc_regs(80) => bus_selected_win_data_80_port,
                           curr_proc_regs(79) => bus_selected_win_data_79_port,
                           curr_proc_regs(78) => bus_selected_win_data_78_port,
                           curr_proc_regs(77) => bus_selected_win_data_77_port,
                           curr_proc_regs(76) => bus_selected_win_data_76_port,
                           curr_proc_regs(75) => bus_selected_win_data_75_port,
                           curr_proc_regs(74) => bus_selected_win_data_74_port,
                           curr_proc_regs(73) => bus_selected_win_data_73_port,
                           curr_proc_regs(72) => bus_selected_win_data_72_port,
                           curr_proc_regs(71) => bus_selected_win_data_71_port,
                           curr_proc_regs(70) => bus_selected_win_data_70_port,
                           curr_proc_regs(69) => bus_selected_win_data_69_port,
                           curr_proc_regs(68) => bus_selected_win_data_68_port,
                           curr_proc_regs(67) => bus_selected_win_data_67_port,
                           curr_proc_regs(66) => bus_selected_win_data_66_port,
                           curr_proc_regs(65) => bus_selected_win_data_65_port,
                           curr_proc_regs(64) => bus_selected_win_data_64_port,
                           curr_proc_regs(63) => bus_selected_win_data_63_port,
                           curr_proc_regs(62) => bus_selected_win_data_62_port,
                           curr_proc_regs(61) => bus_selected_win_data_61_port,
                           curr_proc_regs(60) => bus_selected_win_data_60_port,
                           curr_proc_regs(59) => bus_selected_win_data_59_port,
                           curr_proc_regs(58) => bus_selected_win_data_58_port,
                           curr_proc_regs(57) => bus_selected_win_data_57_port,
                           curr_proc_regs(56) => bus_selected_win_data_56_port,
                           curr_proc_regs(55) => bus_selected_win_data_55_port,
                           curr_proc_regs(54) => bus_selected_win_data_54_port,
                           curr_proc_regs(53) => bus_selected_win_data_53_port,
                           curr_proc_regs(52) => bus_selected_win_data_52_port,
                           curr_proc_regs(51) => bus_selected_win_data_51_port,
                           curr_proc_regs(50) => bus_selected_win_data_50_port,
                           curr_proc_regs(49) => bus_selected_win_data_49_port,
                           curr_proc_regs(48) => bus_selected_win_data_48_port,
                           curr_proc_regs(47) => bus_selected_win_data_47_port,
                           curr_proc_regs(46) => bus_selected_win_data_46_port,
                           curr_proc_regs(45) => bus_selected_win_data_45_port,
                           curr_proc_regs(44) => bus_selected_win_data_44_port,
                           curr_proc_regs(43) => bus_selected_win_data_43_port,
                           curr_proc_regs(42) => bus_selected_win_data_42_port,
                           curr_proc_regs(41) => bus_selected_win_data_41_port,
                           curr_proc_regs(40) => bus_selected_win_data_40_port,
                           curr_proc_regs(39) => bus_selected_win_data_39_port,
                           curr_proc_regs(38) => bus_selected_win_data_38_port,
                           curr_proc_regs(37) => bus_selected_win_data_37_port,
                           curr_proc_regs(36) => bus_selected_win_data_36_port,
                           curr_proc_regs(35) => bus_selected_win_data_35_port,
                           curr_proc_regs(34) => bus_selected_win_data_34_port,
                           curr_proc_regs(33) => bus_selected_win_data_33_port,
                           curr_proc_regs(32) => bus_selected_win_data_32_port,
                           curr_proc_regs(31) => bus_selected_win_data_31_port,
                           curr_proc_regs(30) => bus_selected_win_data_30_port,
                           curr_proc_regs(29) => bus_selected_win_data_29_port,
                           curr_proc_regs(28) => bus_selected_win_data_28_port,
                           curr_proc_regs(27) => bus_selected_win_data_27_port,
                           curr_proc_regs(26) => bus_selected_win_data_26_port,
                           curr_proc_regs(25) => bus_selected_win_data_25_port,
                           curr_proc_regs(24) => bus_selected_win_data_24_port,
                           curr_proc_regs(23) => bus_selected_win_data_23_port,
                           curr_proc_regs(22) => bus_selected_win_data_22_port,
                           curr_proc_regs(21) => bus_selected_win_data_21_port,
                           curr_proc_regs(20) => bus_selected_win_data_20_port,
                           curr_proc_regs(19) => bus_selected_win_data_19_port,
                           curr_proc_regs(18) => bus_selected_win_data_18_port,
                           curr_proc_regs(17) => bus_selected_win_data_17_port,
                           curr_proc_regs(16) => bus_selected_win_data_16_port,
                           curr_proc_regs(15) => bus_selected_win_data_15_port,
                           curr_proc_regs(14) => bus_selected_win_data_14_port,
                           curr_proc_regs(13) => bus_selected_win_data_13_port,
                           curr_proc_regs(12) => bus_selected_win_data_12_port,
                           curr_proc_regs(11) => bus_selected_win_data_11_port,
                           curr_proc_regs(10) => bus_selected_win_data_10_port,
                           curr_proc_regs(9) => bus_selected_win_data_9_port, 
                           curr_proc_regs(8) => bus_selected_win_data_8_port, 
                           curr_proc_regs(7) => bus_selected_win_data_7_port, 
                           curr_proc_regs(6) => bus_selected_win_data_6_port, 
                           curr_proc_regs(5) => bus_selected_win_data_5_port, 
                           curr_proc_regs(4) => bus_selected_win_data_4_port, 
                           curr_proc_regs(3) => bus_selected_win_data_3_port, 
                           curr_proc_regs(2) => bus_selected_win_data_2_port, 
                           curr_proc_regs(1) => bus_selected_win_data_1_port, 
                           curr_proc_regs(0) => bus_selected_win_data_0_port);
   RDPORT0 : mux_N32_M5_0 port map( S(4) => ADD_RD1(4), S(3) => ADD_RD1(3), 
                           S(2) => ADD_RD1(2), S(1) => ADD_RD1(1), S(0) => 
                           ADD_RD1(0), Q(1023) => 
                           bus_selected_win_data_767_port, Q(1022) => 
                           bus_selected_win_data_766_port, Q(1021) => 
                           bus_selected_win_data_765_port, Q(1020) => 
                           bus_selected_win_data_764_port, Q(1019) => 
                           bus_selected_win_data_763_port, Q(1018) => 
                           bus_selected_win_data_762_port, Q(1017) => 
                           bus_selected_win_data_761_port, Q(1016) => 
                           bus_selected_win_data_760_port, Q(1015) => 
                           bus_selected_win_data_759_port, Q(1014) => 
                           bus_selected_win_data_758_port, Q(1013) => 
                           bus_selected_win_data_757_port, Q(1012) => 
                           bus_selected_win_data_756_port, Q(1011) => 
                           bus_selected_win_data_755_port, Q(1010) => 
                           bus_selected_win_data_754_port, Q(1009) => 
                           bus_selected_win_data_753_port, Q(1008) => 
                           bus_selected_win_data_752_port, Q(1007) => 
                           bus_selected_win_data_751_port, Q(1006) => 
                           bus_selected_win_data_750_port, Q(1005) => 
                           bus_selected_win_data_749_port, Q(1004) => 
                           bus_selected_win_data_748_port, Q(1003) => 
                           bus_selected_win_data_747_port, Q(1002) => 
                           bus_selected_win_data_746_port, Q(1001) => 
                           bus_selected_win_data_745_port, Q(1000) => 
                           bus_selected_win_data_744_port, Q(999) => 
                           bus_selected_win_data_743_port, Q(998) => 
                           bus_selected_win_data_742_port, Q(997) => 
                           bus_selected_win_data_741_port, Q(996) => 
                           bus_selected_win_data_740_port, Q(995) => 
                           bus_selected_win_data_739_port, Q(994) => 
                           bus_selected_win_data_738_port, Q(993) => 
                           bus_selected_win_data_737_port, Q(992) => 
                           bus_selected_win_data_736_port, Q(991) => 
                           bus_selected_win_data_735_port, Q(990) => 
                           bus_selected_win_data_734_port, Q(989) => 
                           bus_selected_win_data_733_port, Q(988) => 
                           bus_selected_win_data_732_port, Q(987) => 
                           bus_selected_win_data_731_port, Q(986) => 
                           bus_selected_win_data_730_port, Q(985) => 
                           bus_selected_win_data_729_port, Q(984) => 
                           bus_selected_win_data_728_port, Q(983) => 
                           bus_selected_win_data_727_port, Q(982) => 
                           bus_selected_win_data_726_port, Q(981) => 
                           bus_selected_win_data_725_port, Q(980) => 
                           bus_selected_win_data_724_port, Q(979) => 
                           bus_selected_win_data_723_port, Q(978) => 
                           bus_selected_win_data_722_port, Q(977) => 
                           bus_selected_win_data_721_port, Q(976) => 
                           bus_selected_win_data_720_port, Q(975) => 
                           bus_selected_win_data_719_port, Q(974) => 
                           bus_selected_win_data_718_port, Q(973) => 
                           bus_selected_win_data_717_port, Q(972) => 
                           bus_selected_win_data_716_port, Q(971) => 
                           bus_selected_win_data_715_port, Q(970) => 
                           bus_selected_win_data_714_port, Q(969) => 
                           bus_selected_win_data_713_port, Q(968) => 
                           bus_selected_win_data_712_port, Q(967) => 
                           bus_selected_win_data_711_port, Q(966) => 
                           bus_selected_win_data_710_port, Q(965) => 
                           bus_selected_win_data_709_port, Q(964) => 
                           bus_selected_win_data_708_port, Q(963) => 
                           bus_selected_win_data_707_port, Q(962) => 
                           bus_selected_win_data_706_port, Q(961) => 
                           bus_selected_win_data_705_port, Q(960) => 
                           bus_selected_win_data_704_port, Q(959) => 
                           bus_selected_win_data_703_port, Q(958) => 
                           bus_selected_win_data_702_port, Q(957) => 
                           bus_selected_win_data_701_port, Q(956) => 
                           bus_selected_win_data_700_port, Q(955) => 
                           bus_selected_win_data_699_port, Q(954) => 
                           bus_selected_win_data_698_port, Q(953) => 
                           bus_selected_win_data_697_port, Q(952) => 
                           bus_selected_win_data_696_port, Q(951) => 
                           bus_selected_win_data_695_port, Q(950) => 
                           bus_selected_win_data_694_port, Q(949) => 
                           bus_selected_win_data_693_port, Q(948) => 
                           bus_selected_win_data_692_port, Q(947) => 
                           bus_selected_win_data_691_port, Q(946) => 
                           bus_selected_win_data_690_port, Q(945) => 
                           bus_selected_win_data_689_port, Q(944) => 
                           bus_selected_win_data_688_port, Q(943) => 
                           bus_selected_win_data_687_port, Q(942) => 
                           bus_selected_win_data_686_port, Q(941) => 
                           bus_selected_win_data_685_port, Q(940) => 
                           bus_selected_win_data_684_port, Q(939) => 
                           bus_selected_win_data_683_port, Q(938) => 
                           bus_selected_win_data_682_port, Q(937) => 
                           bus_selected_win_data_681_port, Q(936) => 
                           bus_selected_win_data_680_port, Q(935) => 
                           bus_selected_win_data_679_port, Q(934) => 
                           bus_selected_win_data_678_port, Q(933) => 
                           bus_selected_win_data_677_port, Q(932) => 
                           bus_selected_win_data_676_port, Q(931) => 
                           bus_selected_win_data_675_port, Q(930) => 
                           bus_selected_win_data_674_port, Q(929) => 
                           bus_selected_win_data_673_port, Q(928) => 
                           bus_selected_win_data_672_port, Q(927) => 
                           bus_selected_win_data_671_port, Q(926) => 
                           bus_selected_win_data_670_port, Q(925) => 
                           bus_selected_win_data_669_port, Q(924) => 
                           bus_selected_win_data_668_port, Q(923) => 
                           bus_selected_win_data_667_port, Q(922) => 
                           bus_selected_win_data_666_port, Q(921) => 
                           bus_selected_win_data_665_port, Q(920) => 
                           bus_selected_win_data_664_port, Q(919) => 
                           bus_selected_win_data_663_port, Q(918) => 
                           bus_selected_win_data_662_port, Q(917) => 
                           bus_selected_win_data_661_port, Q(916) => 
                           bus_selected_win_data_660_port, Q(915) => 
                           bus_selected_win_data_659_port, Q(914) => 
                           bus_selected_win_data_658_port, Q(913) => 
                           bus_selected_win_data_657_port, Q(912) => 
                           bus_selected_win_data_656_port, Q(911) => 
                           bus_selected_win_data_655_port, Q(910) => 
                           bus_selected_win_data_654_port, Q(909) => 
                           bus_selected_win_data_653_port, Q(908) => 
                           bus_selected_win_data_652_port, Q(907) => 
                           bus_selected_win_data_651_port, Q(906) => 
                           bus_selected_win_data_650_port, Q(905) => 
                           bus_selected_win_data_649_port, Q(904) => 
                           bus_selected_win_data_648_port, Q(903) => 
                           bus_selected_win_data_647_port, Q(902) => 
                           bus_selected_win_data_646_port, Q(901) => 
                           bus_selected_win_data_645_port, Q(900) => 
                           bus_selected_win_data_644_port, Q(899) => 
                           bus_selected_win_data_643_port, Q(898) => 
                           bus_selected_win_data_642_port, Q(897) => 
                           bus_selected_win_data_641_port, Q(896) => 
                           bus_selected_win_data_640_port, Q(895) => 
                           bus_selected_win_data_639_port, Q(894) => 
                           bus_selected_win_data_638_port, Q(893) => 
                           bus_selected_win_data_637_port, Q(892) => 
                           bus_selected_win_data_636_port, Q(891) => 
                           bus_selected_win_data_635_port, Q(890) => 
                           bus_selected_win_data_634_port, Q(889) => 
                           bus_selected_win_data_633_port, Q(888) => 
                           bus_selected_win_data_632_port, Q(887) => 
                           bus_selected_win_data_631_port, Q(886) => 
                           bus_selected_win_data_630_port, Q(885) => 
                           bus_selected_win_data_629_port, Q(884) => 
                           bus_selected_win_data_628_port, Q(883) => 
                           bus_selected_win_data_627_port, Q(882) => 
                           bus_selected_win_data_626_port, Q(881) => 
                           bus_selected_win_data_625_port, Q(880) => 
                           bus_selected_win_data_624_port, Q(879) => 
                           bus_selected_win_data_623_port, Q(878) => 
                           bus_selected_win_data_622_port, Q(877) => 
                           bus_selected_win_data_621_port, Q(876) => 
                           bus_selected_win_data_620_port, Q(875) => 
                           bus_selected_win_data_619_port, Q(874) => 
                           bus_selected_win_data_618_port, Q(873) => 
                           bus_selected_win_data_617_port, Q(872) => 
                           bus_selected_win_data_616_port, Q(871) => 
                           bus_selected_win_data_615_port, Q(870) => 
                           bus_selected_win_data_614_port, Q(869) => 
                           bus_selected_win_data_613_port, Q(868) => 
                           bus_selected_win_data_612_port, Q(867) => 
                           bus_selected_win_data_611_port, Q(866) => 
                           bus_selected_win_data_610_port, Q(865) => 
                           bus_selected_win_data_609_port, Q(864) => 
                           bus_selected_win_data_608_port, Q(863) => 
                           bus_selected_win_data_607_port, Q(862) => 
                           bus_selected_win_data_606_port, Q(861) => 
                           bus_selected_win_data_605_port, Q(860) => 
                           bus_selected_win_data_604_port, Q(859) => 
                           bus_selected_win_data_603_port, Q(858) => 
                           bus_selected_win_data_602_port, Q(857) => 
                           bus_selected_win_data_601_port, Q(856) => 
                           bus_selected_win_data_600_port, Q(855) => 
                           bus_selected_win_data_599_port, Q(854) => 
                           bus_selected_win_data_598_port, Q(853) => 
                           bus_selected_win_data_597_port, Q(852) => 
                           bus_selected_win_data_596_port, Q(851) => 
                           bus_selected_win_data_595_port, Q(850) => 
                           bus_selected_win_data_594_port, Q(849) => 
                           bus_selected_win_data_593_port, Q(848) => 
                           bus_selected_win_data_592_port, Q(847) => 
                           bus_selected_win_data_591_port, Q(846) => 
                           bus_selected_win_data_590_port, Q(845) => 
                           bus_selected_win_data_589_port, Q(844) => 
                           bus_selected_win_data_588_port, Q(843) => 
                           bus_selected_win_data_587_port, Q(842) => 
                           bus_selected_win_data_586_port, Q(841) => 
                           bus_selected_win_data_585_port, Q(840) => 
                           bus_selected_win_data_584_port, Q(839) => 
                           bus_selected_win_data_583_port, Q(838) => 
                           bus_selected_win_data_582_port, Q(837) => 
                           bus_selected_win_data_581_port, Q(836) => 
                           bus_selected_win_data_580_port, Q(835) => 
                           bus_selected_win_data_579_port, Q(834) => 
                           bus_selected_win_data_578_port, Q(833) => 
                           bus_selected_win_data_577_port, Q(832) => 
                           bus_selected_win_data_576_port, Q(831) => 
                           bus_selected_win_data_575_port, Q(830) => 
                           bus_selected_win_data_574_port, Q(829) => 
                           bus_selected_win_data_573_port, Q(828) => 
                           bus_selected_win_data_572_port, Q(827) => 
                           bus_selected_win_data_571_port, Q(826) => 
                           bus_selected_win_data_570_port, Q(825) => 
                           bus_selected_win_data_569_port, Q(824) => 
                           bus_selected_win_data_568_port, Q(823) => 
                           bus_selected_win_data_567_port, Q(822) => 
                           bus_selected_win_data_566_port, Q(821) => 
                           bus_selected_win_data_565_port, Q(820) => 
                           bus_selected_win_data_564_port, Q(819) => 
                           bus_selected_win_data_563_port, Q(818) => 
                           bus_selected_win_data_562_port, Q(817) => 
                           bus_selected_win_data_561_port, Q(816) => 
                           bus_selected_win_data_560_port, Q(815) => 
                           bus_selected_win_data_559_port, Q(814) => 
                           bus_selected_win_data_558_port, Q(813) => 
                           bus_selected_win_data_557_port, Q(812) => 
                           bus_selected_win_data_556_port, Q(811) => 
                           bus_selected_win_data_555_port, Q(810) => 
                           bus_selected_win_data_554_port, Q(809) => 
                           bus_selected_win_data_553_port, Q(808) => 
                           bus_selected_win_data_552_port, Q(807) => 
                           bus_selected_win_data_551_port, Q(806) => 
                           bus_selected_win_data_550_port, Q(805) => 
                           bus_selected_win_data_549_port, Q(804) => 
                           bus_selected_win_data_548_port, Q(803) => 
                           bus_selected_win_data_547_port, Q(802) => 
                           bus_selected_win_data_546_port, Q(801) => 
                           bus_selected_win_data_545_port, Q(800) => 
                           bus_selected_win_data_544_port, Q(799) => 
                           bus_selected_win_data_543_port, Q(798) => 
                           bus_selected_win_data_542_port, Q(797) => 
                           bus_selected_win_data_541_port, Q(796) => 
                           bus_selected_win_data_540_port, Q(795) => 
                           bus_selected_win_data_539_port, Q(794) => 
                           bus_selected_win_data_538_port, Q(793) => 
                           bus_selected_win_data_537_port, Q(792) => 
                           bus_selected_win_data_536_port, Q(791) => 
                           bus_selected_win_data_535_port, Q(790) => 
                           bus_selected_win_data_534_port, Q(789) => 
                           bus_selected_win_data_533_port, Q(788) => 
                           bus_selected_win_data_532_port, Q(787) => 
                           bus_selected_win_data_531_port, Q(786) => 
                           bus_selected_win_data_530_port, Q(785) => 
                           bus_selected_win_data_529_port, Q(784) => 
                           bus_selected_win_data_528_port, Q(783) => 
                           bus_selected_win_data_527_port, Q(782) => 
                           bus_selected_win_data_526_port, Q(781) => 
                           bus_selected_win_data_525_port, Q(780) => 
                           bus_selected_win_data_524_port, Q(779) => 
                           bus_selected_win_data_523_port, Q(778) => 
                           bus_selected_win_data_522_port, Q(777) => 
                           bus_selected_win_data_521_port, Q(776) => 
                           bus_selected_win_data_520_port, Q(775) => 
                           bus_selected_win_data_519_port, Q(774) => 
                           bus_selected_win_data_518_port, Q(773) => 
                           bus_selected_win_data_517_port, Q(772) => 
                           bus_selected_win_data_516_port, Q(771) => 
                           bus_selected_win_data_515_port, Q(770) => 
                           bus_selected_win_data_514_port, Q(769) => 
                           bus_selected_win_data_513_port, Q(768) => 
                           bus_selected_win_data_512_port, Q(767) => 
                           bus_selected_win_data_511_port, Q(766) => 
                           bus_selected_win_data_510_port, Q(765) => 
                           bus_selected_win_data_509_port, Q(764) => 
                           bus_selected_win_data_508_port, Q(763) => 
                           bus_selected_win_data_507_port, Q(762) => 
                           bus_selected_win_data_506_port, Q(761) => 
                           bus_selected_win_data_505_port, Q(760) => 
                           bus_selected_win_data_504_port, Q(759) => 
                           bus_selected_win_data_503_port, Q(758) => 
                           bus_selected_win_data_502_port, Q(757) => 
                           bus_selected_win_data_501_port, Q(756) => 
                           bus_selected_win_data_500_port, Q(755) => 
                           bus_selected_win_data_499_port, Q(754) => 
                           bus_selected_win_data_498_port, Q(753) => 
                           bus_selected_win_data_497_port, Q(752) => 
                           bus_selected_win_data_496_port, Q(751) => 
                           bus_selected_win_data_495_port, Q(750) => 
                           bus_selected_win_data_494_port, Q(749) => 
                           bus_selected_win_data_493_port, Q(748) => 
                           bus_selected_win_data_492_port, Q(747) => 
                           bus_selected_win_data_491_port, Q(746) => 
                           bus_selected_win_data_490_port, Q(745) => 
                           bus_selected_win_data_489_port, Q(744) => 
                           bus_selected_win_data_488_port, Q(743) => 
                           bus_selected_win_data_487_port, Q(742) => 
                           bus_selected_win_data_486_port, Q(741) => 
                           bus_selected_win_data_485_port, Q(740) => 
                           bus_selected_win_data_484_port, Q(739) => 
                           bus_selected_win_data_483_port, Q(738) => 
                           bus_selected_win_data_482_port, Q(737) => 
                           bus_selected_win_data_481_port, Q(736) => 
                           bus_selected_win_data_480_port, Q(735) => 
                           bus_selected_win_data_479_port, Q(734) => 
                           bus_selected_win_data_478_port, Q(733) => 
                           bus_selected_win_data_477_port, Q(732) => 
                           bus_selected_win_data_476_port, Q(731) => 
                           bus_selected_win_data_475_port, Q(730) => 
                           bus_selected_win_data_474_port, Q(729) => 
                           bus_selected_win_data_473_port, Q(728) => 
                           bus_selected_win_data_472_port, Q(727) => 
                           bus_selected_win_data_471_port, Q(726) => 
                           bus_selected_win_data_470_port, Q(725) => 
                           bus_selected_win_data_469_port, Q(724) => 
                           bus_selected_win_data_468_port, Q(723) => 
                           bus_selected_win_data_467_port, Q(722) => 
                           bus_selected_win_data_466_port, Q(721) => 
                           bus_selected_win_data_465_port, Q(720) => 
                           bus_selected_win_data_464_port, Q(719) => 
                           bus_selected_win_data_463_port, Q(718) => 
                           bus_selected_win_data_462_port, Q(717) => 
                           bus_selected_win_data_461_port, Q(716) => 
                           bus_selected_win_data_460_port, Q(715) => 
                           bus_selected_win_data_459_port, Q(714) => 
                           bus_selected_win_data_458_port, Q(713) => 
                           bus_selected_win_data_457_port, Q(712) => 
                           bus_selected_win_data_456_port, Q(711) => 
                           bus_selected_win_data_455_port, Q(710) => 
                           bus_selected_win_data_454_port, Q(709) => 
                           bus_selected_win_data_453_port, Q(708) => 
                           bus_selected_win_data_452_port, Q(707) => 
                           bus_selected_win_data_451_port, Q(706) => 
                           bus_selected_win_data_450_port, Q(705) => 
                           bus_selected_win_data_449_port, Q(704) => 
                           bus_selected_win_data_448_port, Q(703) => 
                           bus_selected_win_data_447_port, Q(702) => 
                           bus_selected_win_data_446_port, Q(701) => 
                           bus_selected_win_data_445_port, Q(700) => 
                           bus_selected_win_data_444_port, Q(699) => 
                           bus_selected_win_data_443_port, Q(698) => 
                           bus_selected_win_data_442_port, Q(697) => 
                           bus_selected_win_data_441_port, Q(696) => 
                           bus_selected_win_data_440_port, Q(695) => 
                           bus_selected_win_data_439_port, Q(694) => 
                           bus_selected_win_data_438_port, Q(693) => 
                           bus_selected_win_data_437_port, Q(692) => 
                           bus_selected_win_data_436_port, Q(691) => 
                           bus_selected_win_data_435_port, Q(690) => 
                           bus_selected_win_data_434_port, Q(689) => 
                           bus_selected_win_data_433_port, Q(688) => 
                           bus_selected_win_data_432_port, Q(687) => 
                           bus_selected_win_data_431_port, Q(686) => 
                           bus_selected_win_data_430_port, Q(685) => 
                           bus_selected_win_data_429_port, Q(684) => 
                           bus_selected_win_data_428_port, Q(683) => 
                           bus_selected_win_data_427_port, Q(682) => 
                           bus_selected_win_data_426_port, Q(681) => 
                           bus_selected_win_data_425_port, Q(680) => 
                           bus_selected_win_data_424_port, Q(679) => 
                           bus_selected_win_data_423_port, Q(678) => 
                           bus_selected_win_data_422_port, Q(677) => 
                           bus_selected_win_data_421_port, Q(676) => 
                           bus_selected_win_data_420_port, Q(675) => 
                           bus_selected_win_data_419_port, Q(674) => 
                           bus_selected_win_data_418_port, Q(673) => 
                           bus_selected_win_data_417_port, Q(672) => 
                           bus_selected_win_data_416_port, Q(671) => 
                           bus_selected_win_data_415_port, Q(670) => 
                           bus_selected_win_data_414_port, Q(669) => 
                           bus_selected_win_data_413_port, Q(668) => 
                           bus_selected_win_data_412_port, Q(667) => 
                           bus_selected_win_data_411_port, Q(666) => 
                           bus_selected_win_data_410_port, Q(665) => 
                           bus_selected_win_data_409_port, Q(664) => 
                           bus_selected_win_data_408_port, Q(663) => 
                           bus_selected_win_data_407_port, Q(662) => 
                           bus_selected_win_data_406_port, Q(661) => 
                           bus_selected_win_data_405_port, Q(660) => 
                           bus_selected_win_data_404_port, Q(659) => 
                           bus_selected_win_data_403_port, Q(658) => 
                           bus_selected_win_data_402_port, Q(657) => 
                           bus_selected_win_data_401_port, Q(656) => 
                           bus_selected_win_data_400_port, Q(655) => 
                           bus_selected_win_data_399_port, Q(654) => 
                           bus_selected_win_data_398_port, Q(653) => 
                           bus_selected_win_data_397_port, Q(652) => 
                           bus_selected_win_data_396_port, Q(651) => 
                           bus_selected_win_data_395_port, Q(650) => 
                           bus_selected_win_data_394_port, Q(649) => 
                           bus_selected_win_data_393_port, Q(648) => 
                           bus_selected_win_data_392_port, Q(647) => 
                           bus_selected_win_data_391_port, Q(646) => 
                           bus_selected_win_data_390_port, Q(645) => 
                           bus_selected_win_data_389_port, Q(644) => 
                           bus_selected_win_data_388_port, Q(643) => 
                           bus_selected_win_data_387_port, Q(642) => 
                           bus_selected_win_data_386_port, Q(641) => 
                           bus_selected_win_data_385_port, Q(640) => 
                           bus_selected_win_data_384_port, Q(639) => 
                           bus_selected_win_data_383_port, Q(638) => 
                           bus_selected_win_data_382_port, Q(637) => 
                           bus_selected_win_data_381_port, Q(636) => 
                           bus_selected_win_data_380_port, Q(635) => 
                           bus_selected_win_data_379_port, Q(634) => 
                           bus_selected_win_data_378_port, Q(633) => 
                           bus_selected_win_data_377_port, Q(632) => 
                           bus_selected_win_data_376_port, Q(631) => 
                           bus_selected_win_data_375_port, Q(630) => 
                           bus_selected_win_data_374_port, Q(629) => 
                           bus_selected_win_data_373_port, Q(628) => 
                           bus_selected_win_data_372_port, Q(627) => 
                           bus_selected_win_data_371_port, Q(626) => 
                           bus_selected_win_data_370_port, Q(625) => 
                           bus_selected_win_data_369_port, Q(624) => 
                           bus_selected_win_data_368_port, Q(623) => 
                           bus_selected_win_data_367_port, Q(622) => 
                           bus_selected_win_data_366_port, Q(621) => 
                           bus_selected_win_data_365_port, Q(620) => 
                           bus_selected_win_data_364_port, Q(619) => 
                           bus_selected_win_data_363_port, Q(618) => 
                           bus_selected_win_data_362_port, Q(617) => 
                           bus_selected_win_data_361_port, Q(616) => 
                           bus_selected_win_data_360_port, Q(615) => 
                           bus_selected_win_data_359_port, Q(614) => 
                           bus_selected_win_data_358_port, Q(613) => 
                           bus_selected_win_data_357_port, Q(612) => 
                           bus_selected_win_data_356_port, Q(611) => 
                           bus_selected_win_data_355_port, Q(610) => 
                           bus_selected_win_data_354_port, Q(609) => 
                           bus_selected_win_data_353_port, Q(608) => 
                           bus_selected_win_data_352_port, Q(607) => 
                           bus_selected_win_data_351_port, Q(606) => 
                           bus_selected_win_data_350_port, Q(605) => 
                           bus_selected_win_data_349_port, Q(604) => 
                           bus_selected_win_data_348_port, Q(603) => 
                           bus_selected_win_data_347_port, Q(602) => 
                           bus_selected_win_data_346_port, Q(601) => 
                           bus_selected_win_data_345_port, Q(600) => 
                           bus_selected_win_data_344_port, Q(599) => 
                           bus_selected_win_data_343_port, Q(598) => 
                           bus_selected_win_data_342_port, Q(597) => 
                           bus_selected_win_data_341_port, Q(596) => 
                           bus_selected_win_data_340_port, Q(595) => 
                           bus_selected_win_data_339_port, Q(594) => 
                           bus_selected_win_data_338_port, Q(593) => 
                           bus_selected_win_data_337_port, Q(592) => 
                           bus_selected_win_data_336_port, Q(591) => 
                           bus_selected_win_data_335_port, Q(590) => 
                           bus_selected_win_data_334_port, Q(589) => 
                           bus_selected_win_data_333_port, Q(588) => 
                           bus_selected_win_data_332_port, Q(587) => 
                           bus_selected_win_data_331_port, Q(586) => 
                           bus_selected_win_data_330_port, Q(585) => 
                           bus_selected_win_data_329_port, Q(584) => 
                           bus_selected_win_data_328_port, Q(583) => 
                           bus_selected_win_data_327_port, Q(582) => 
                           bus_selected_win_data_326_port, Q(581) => 
                           bus_selected_win_data_325_port, Q(580) => 
                           bus_selected_win_data_324_port, Q(579) => 
                           bus_selected_win_data_323_port, Q(578) => 
                           bus_selected_win_data_322_port, Q(577) => 
                           bus_selected_win_data_321_port, Q(576) => 
                           bus_selected_win_data_320_port, Q(575) => 
                           bus_selected_win_data_319_port, Q(574) => 
                           bus_selected_win_data_318_port, Q(573) => 
                           bus_selected_win_data_317_port, Q(572) => 
                           bus_selected_win_data_316_port, Q(571) => 
                           bus_selected_win_data_315_port, Q(570) => 
                           bus_selected_win_data_314_port, Q(569) => 
                           bus_selected_win_data_313_port, Q(568) => 
                           bus_selected_win_data_312_port, Q(567) => 
                           bus_selected_win_data_311_port, Q(566) => 
                           bus_selected_win_data_310_port, Q(565) => 
                           bus_selected_win_data_309_port, Q(564) => 
                           bus_selected_win_data_308_port, Q(563) => 
                           bus_selected_win_data_307_port, Q(562) => 
                           bus_selected_win_data_306_port, Q(561) => 
                           bus_selected_win_data_305_port, Q(560) => 
                           bus_selected_win_data_304_port, Q(559) => 
                           bus_selected_win_data_303_port, Q(558) => 
                           bus_selected_win_data_302_port, Q(557) => 
                           bus_selected_win_data_301_port, Q(556) => 
                           bus_selected_win_data_300_port, Q(555) => 
                           bus_selected_win_data_299_port, Q(554) => 
                           bus_selected_win_data_298_port, Q(553) => 
                           bus_selected_win_data_297_port, Q(552) => 
                           bus_selected_win_data_296_port, Q(551) => 
                           bus_selected_win_data_295_port, Q(550) => 
                           bus_selected_win_data_294_port, Q(549) => 
                           bus_selected_win_data_293_port, Q(548) => 
                           bus_selected_win_data_292_port, Q(547) => 
                           bus_selected_win_data_291_port, Q(546) => 
                           bus_selected_win_data_290_port, Q(545) => 
                           bus_selected_win_data_289_port, Q(544) => 
                           bus_selected_win_data_288_port, Q(543) => 
                           bus_selected_win_data_287_port, Q(542) => 
                           bus_selected_win_data_286_port, Q(541) => 
                           bus_selected_win_data_285_port, Q(540) => 
                           bus_selected_win_data_284_port, Q(539) => 
                           bus_selected_win_data_283_port, Q(538) => 
                           bus_selected_win_data_282_port, Q(537) => 
                           bus_selected_win_data_281_port, Q(536) => 
                           bus_selected_win_data_280_port, Q(535) => 
                           bus_selected_win_data_279_port, Q(534) => 
                           bus_selected_win_data_278_port, Q(533) => 
                           bus_selected_win_data_277_port, Q(532) => 
                           bus_selected_win_data_276_port, Q(531) => 
                           bus_selected_win_data_275_port, Q(530) => 
                           bus_selected_win_data_274_port, Q(529) => 
                           bus_selected_win_data_273_port, Q(528) => 
                           bus_selected_win_data_272_port, Q(527) => 
                           bus_selected_win_data_271_port, Q(526) => 
                           bus_selected_win_data_270_port, Q(525) => 
                           bus_selected_win_data_269_port, Q(524) => 
                           bus_selected_win_data_268_port, Q(523) => 
                           bus_selected_win_data_267_port, Q(522) => 
                           bus_selected_win_data_266_port, Q(521) => 
                           bus_selected_win_data_265_port, Q(520) => 
                           bus_selected_win_data_264_port, Q(519) => 
                           bus_selected_win_data_263_port, Q(518) => 
                           bus_selected_win_data_262_port, Q(517) => 
                           bus_selected_win_data_261_port, Q(516) => 
                           bus_selected_win_data_260_port, Q(515) => 
                           bus_selected_win_data_259_port, Q(514) => 
                           bus_selected_win_data_258_port, Q(513) => 
                           bus_selected_win_data_257_port, Q(512) => 
                           bus_selected_win_data_256_port, Q(511) => 
                           bus_selected_win_data_255_port, Q(510) => 
                           bus_selected_win_data_254_port, Q(509) => 
                           bus_selected_win_data_253_port, Q(508) => 
                           bus_selected_win_data_252_port, Q(507) => 
                           bus_selected_win_data_251_port, Q(506) => 
                           bus_selected_win_data_250_port, Q(505) => 
                           bus_selected_win_data_249_port, Q(504) => 
                           bus_selected_win_data_248_port, Q(503) => 
                           bus_selected_win_data_247_port, Q(502) => 
                           bus_selected_win_data_246_port, Q(501) => 
                           bus_selected_win_data_245_port, Q(500) => 
                           bus_selected_win_data_244_port, Q(499) => 
                           bus_selected_win_data_243_port, Q(498) => 
                           bus_selected_win_data_242_port, Q(497) => 
                           bus_selected_win_data_241_port, Q(496) => 
                           bus_selected_win_data_240_port, Q(495) => 
                           bus_selected_win_data_239_port, Q(494) => 
                           bus_selected_win_data_238_port, Q(493) => 
                           bus_selected_win_data_237_port, Q(492) => 
                           bus_selected_win_data_236_port, Q(491) => 
                           bus_selected_win_data_235_port, Q(490) => 
                           bus_selected_win_data_234_port, Q(489) => 
                           bus_selected_win_data_233_port, Q(488) => 
                           bus_selected_win_data_232_port, Q(487) => 
                           bus_selected_win_data_231_port, Q(486) => 
                           bus_selected_win_data_230_port, Q(485) => 
                           bus_selected_win_data_229_port, Q(484) => 
                           bus_selected_win_data_228_port, Q(483) => 
                           bus_selected_win_data_227_port, Q(482) => 
                           bus_selected_win_data_226_port, Q(481) => 
                           bus_selected_win_data_225_port, Q(480) => 
                           bus_selected_win_data_224_port, Q(479) => 
                           bus_selected_win_data_223_port, Q(478) => 
                           bus_selected_win_data_222_port, Q(477) => 
                           bus_selected_win_data_221_port, Q(476) => 
                           bus_selected_win_data_220_port, Q(475) => 
                           bus_selected_win_data_219_port, Q(474) => 
                           bus_selected_win_data_218_port, Q(473) => 
                           bus_selected_win_data_217_port, Q(472) => 
                           bus_selected_win_data_216_port, Q(471) => 
                           bus_selected_win_data_215_port, Q(470) => 
                           bus_selected_win_data_214_port, Q(469) => 
                           bus_selected_win_data_213_port, Q(468) => 
                           bus_selected_win_data_212_port, Q(467) => 
                           bus_selected_win_data_211_port, Q(466) => 
                           bus_selected_win_data_210_port, Q(465) => 
                           bus_selected_win_data_209_port, Q(464) => 
                           bus_selected_win_data_208_port, Q(463) => 
                           bus_selected_win_data_207_port, Q(462) => 
                           bus_selected_win_data_206_port, Q(461) => 
                           bus_selected_win_data_205_port, Q(460) => 
                           bus_selected_win_data_204_port, Q(459) => 
                           bus_selected_win_data_203_port, Q(458) => 
                           bus_selected_win_data_202_port, Q(457) => 
                           bus_selected_win_data_201_port, Q(456) => 
                           bus_selected_win_data_200_port, Q(455) => 
                           bus_selected_win_data_199_port, Q(454) => 
                           bus_selected_win_data_198_port, Q(453) => 
                           bus_selected_win_data_197_port, Q(452) => 
                           bus_selected_win_data_196_port, Q(451) => 
                           bus_selected_win_data_195_port, Q(450) => 
                           bus_selected_win_data_194_port, Q(449) => 
                           bus_selected_win_data_193_port, Q(448) => 
                           bus_selected_win_data_192_port, Q(447) => 
                           bus_selected_win_data_191_port, Q(446) => 
                           bus_selected_win_data_190_port, Q(445) => 
                           bus_selected_win_data_189_port, Q(444) => 
                           bus_selected_win_data_188_port, Q(443) => 
                           bus_selected_win_data_187_port, Q(442) => 
                           bus_selected_win_data_186_port, Q(441) => 
                           bus_selected_win_data_185_port, Q(440) => 
                           bus_selected_win_data_184_port, Q(439) => 
                           bus_selected_win_data_183_port, Q(438) => 
                           bus_selected_win_data_182_port, Q(437) => 
                           bus_selected_win_data_181_port, Q(436) => 
                           bus_selected_win_data_180_port, Q(435) => 
                           bus_selected_win_data_179_port, Q(434) => 
                           bus_selected_win_data_178_port, Q(433) => 
                           bus_selected_win_data_177_port, Q(432) => 
                           bus_selected_win_data_176_port, Q(431) => 
                           bus_selected_win_data_175_port, Q(430) => 
                           bus_selected_win_data_174_port, Q(429) => 
                           bus_selected_win_data_173_port, Q(428) => 
                           bus_selected_win_data_172_port, Q(427) => 
                           bus_selected_win_data_171_port, Q(426) => 
                           bus_selected_win_data_170_port, Q(425) => 
                           bus_selected_win_data_169_port, Q(424) => 
                           bus_selected_win_data_168_port, Q(423) => 
                           bus_selected_win_data_167_port, Q(422) => 
                           bus_selected_win_data_166_port, Q(421) => 
                           bus_selected_win_data_165_port, Q(420) => 
                           bus_selected_win_data_164_port, Q(419) => 
                           bus_selected_win_data_163_port, Q(418) => 
                           bus_selected_win_data_162_port, Q(417) => 
                           bus_selected_win_data_161_port, Q(416) => 
                           bus_selected_win_data_160_port, Q(415) => 
                           bus_selected_win_data_159_port, Q(414) => 
                           bus_selected_win_data_158_port, Q(413) => 
                           bus_selected_win_data_157_port, Q(412) => 
                           bus_selected_win_data_156_port, Q(411) => 
                           bus_selected_win_data_155_port, Q(410) => 
                           bus_selected_win_data_154_port, Q(409) => 
                           bus_selected_win_data_153_port, Q(408) => 
                           bus_selected_win_data_152_port, Q(407) => 
                           bus_selected_win_data_151_port, Q(406) => 
                           bus_selected_win_data_150_port, Q(405) => 
                           bus_selected_win_data_149_port, Q(404) => 
                           bus_selected_win_data_148_port, Q(403) => 
                           bus_selected_win_data_147_port, Q(402) => 
                           bus_selected_win_data_146_port, Q(401) => 
                           bus_selected_win_data_145_port, Q(400) => 
                           bus_selected_win_data_144_port, Q(399) => 
                           bus_selected_win_data_143_port, Q(398) => 
                           bus_selected_win_data_142_port, Q(397) => 
                           bus_selected_win_data_141_port, Q(396) => 
                           bus_selected_win_data_140_port, Q(395) => 
                           bus_selected_win_data_139_port, Q(394) => 
                           bus_selected_win_data_138_port, Q(393) => 
                           bus_selected_win_data_137_port, Q(392) => 
                           bus_selected_win_data_136_port, Q(391) => 
                           bus_selected_win_data_135_port, Q(390) => 
                           bus_selected_win_data_134_port, Q(389) => 
                           bus_selected_win_data_133_port, Q(388) => 
                           bus_selected_win_data_132_port, Q(387) => 
                           bus_selected_win_data_131_port, Q(386) => 
                           bus_selected_win_data_130_port, Q(385) => 
                           bus_selected_win_data_129_port, Q(384) => 
                           bus_selected_win_data_128_port, Q(383) => 
                           bus_selected_win_data_127_port, Q(382) => 
                           bus_selected_win_data_126_port, Q(381) => 
                           bus_selected_win_data_125_port, Q(380) => 
                           bus_selected_win_data_124_port, Q(379) => 
                           bus_selected_win_data_123_port, Q(378) => 
                           bus_selected_win_data_122_port, Q(377) => 
                           bus_selected_win_data_121_port, Q(376) => 
                           bus_selected_win_data_120_port, Q(375) => 
                           bus_selected_win_data_119_port, Q(374) => 
                           bus_selected_win_data_118_port, Q(373) => 
                           bus_selected_win_data_117_port, Q(372) => 
                           bus_selected_win_data_116_port, Q(371) => 
                           bus_selected_win_data_115_port, Q(370) => 
                           bus_selected_win_data_114_port, Q(369) => 
                           bus_selected_win_data_113_port, Q(368) => 
                           bus_selected_win_data_112_port, Q(367) => 
                           bus_selected_win_data_111_port, Q(366) => 
                           bus_selected_win_data_110_port, Q(365) => 
                           bus_selected_win_data_109_port, Q(364) => 
                           bus_selected_win_data_108_port, Q(363) => 
                           bus_selected_win_data_107_port, Q(362) => 
                           bus_selected_win_data_106_port, Q(361) => 
                           bus_selected_win_data_105_port, Q(360) => 
                           bus_selected_win_data_104_port, Q(359) => 
                           bus_selected_win_data_103_port, Q(358) => 
                           bus_selected_win_data_102_port, Q(357) => 
                           bus_selected_win_data_101_port, Q(356) => 
                           bus_selected_win_data_100_port, Q(355) => 
                           bus_selected_win_data_99_port, Q(354) => 
                           bus_selected_win_data_98_port, Q(353) => 
                           bus_selected_win_data_97_port, Q(352) => 
                           bus_selected_win_data_96_port, Q(351) => 
                           bus_selected_win_data_95_port, Q(350) => 
                           bus_selected_win_data_94_port, Q(349) => 
                           bus_selected_win_data_93_port, Q(348) => 
                           bus_selected_win_data_92_port, Q(347) => 
                           bus_selected_win_data_91_port, Q(346) => 
                           bus_selected_win_data_90_port, Q(345) => 
                           bus_selected_win_data_89_port, Q(344) => 
                           bus_selected_win_data_88_port, Q(343) => 
                           bus_selected_win_data_87_port, Q(342) => 
                           bus_selected_win_data_86_port, Q(341) => 
                           bus_selected_win_data_85_port, Q(340) => 
                           bus_selected_win_data_84_port, Q(339) => 
                           bus_selected_win_data_83_port, Q(338) => 
                           bus_selected_win_data_82_port, Q(337) => 
                           bus_selected_win_data_81_port, Q(336) => 
                           bus_selected_win_data_80_port, Q(335) => 
                           bus_selected_win_data_79_port, Q(334) => 
                           bus_selected_win_data_78_port, Q(333) => 
                           bus_selected_win_data_77_port, Q(332) => 
                           bus_selected_win_data_76_port, Q(331) => 
                           bus_selected_win_data_75_port, Q(330) => 
                           bus_selected_win_data_74_port, Q(329) => 
                           bus_selected_win_data_73_port, Q(328) => 
                           bus_selected_win_data_72_port, Q(327) => 
                           bus_selected_win_data_71_port, Q(326) => 
                           bus_selected_win_data_70_port, Q(325) => 
                           bus_selected_win_data_69_port, Q(324) => 
                           bus_selected_win_data_68_port, Q(323) => 
                           bus_selected_win_data_67_port, Q(322) => 
                           bus_selected_win_data_66_port, Q(321) => 
                           bus_selected_win_data_65_port, Q(320) => 
                           bus_selected_win_data_64_port, Q(319) => 
                           bus_selected_win_data_63_port, Q(318) => 
                           bus_selected_win_data_62_port, Q(317) => 
                           bus_selected_win_data_61_port, Q(316) => 
                           bus_selected_win_data_60_port, Q(315) => 
                           bus_selected_win_data_59_port, Q(314) => 
                           bus_selected_win_data_58_port, Q(313) => 
                           bus_selected_win_data_57_port, Q(312) => 
                           bus_selected_win_data_56_port, Q(311) => 
                           bus_selected_win_data_55_port, Q(310) => 
                           bus_selected_win_data_54_port, Q(309) => 
                           bus_selected_win_data_53_port, Q(308) => 
                           bus_selected_win_data_52_port, Q(307) => 
                           bus_selected_win_data_51_port, Q(306) => 
                           bus_selected_win_data_50_port, Q(305) => 
                           bus_selected_win_data_49_port, Q(304) => 
                           bus_selected_win_data_48_port, Q(303) => 
                           bus_selected_win_data_47_port, Q(302) => 
                           bus_selected_win_data_46_port, Q(301) => 
                           bus_selected_win_data_45_port, Q(300) => 
                           bus_selected_win_data_44_port, Q(299) => 
                           bus_selected_win_data_43_port, Q(298) => 
                           bus_selected_win_data_42_port, Q(297) => 
                           bus_selected_win_data_41_port, Q(296) => 
                           bus_selected_win_data_40_port, Q(295) => 
                           bus_selected_win_data_39_port, Q(294) => 
                           bus_selected_win_data_38_port, Q(293) => 
                           bus_selected_win_data_37_port, Q(292) => 
                           bus_selected_win_data_36_port, Q(291) => 
                           bus_selected_win_data_35_port, Q(290) => 
                           bus_selected_win_data_34_port, Q(289) => 
                           bus_selected_win_data_33_port, Q(288) => 
                           bus_selected_win_data_32_port, Q(287) => 
                           bus_selected_win_data_31_port, Q(286) => 
                           bus_selected_win_data_30_port, Q(285) => 
                           bus_selected_win_data_29_port, Q(284) => 
                           bus_selected_win_data_28_port, Q(283) => 
                           bus_selected_win_data_27_port, Q(282) => 
                           bus_selected_win_data_26_port, Q(281) => 
                           bus_selected_win_data_25_port, Q(280) => 
                           bus_selected_win_data_24_port, Q(279) => 
                           bus_selected_win_data_23_port, Q(278) => 
                           bus_selected_win_data_22_port, Q(277) => 
                           bus_selected_win_data_21_port, Q(276) => 
                           bus_selected_win_data_20_port, Q(275) => 
                           bus_selected_win_data_19_port, Q(274) => 
                           bus_selected_win_data_18_port, Q(273) => 
                           bus_selected_win_data_17_port, Q(272) => 
                           bus_selected_win_data_16_port, Q(271) => 
                           bus_selected_win_data_15_port, Q(270) => 
                           bus_selected_win_data_14_port, Q(269) => 
                           bus_selected_win_data_13_port, Q(268) => 
                           bus_selected_win_data_12_port, Q(267) => 
                           bus_selected_win_data_11_port, Q(266) => 
                           bus_selected_win_data_10_port, Q(265) => 
                           bus_selected_win_data_9_port, Q(264) => 
                           bus_selected_win_data_8_port, Q(263) => 
                           bus_selected_win_data_7_port, Q(262) => 
                           bus_selected_win_data_6_port, Q(261) => 
                           bus_selected_win_data_5_port, Q(260) => 
                           bus_selected_win_data_4_port, Q(259) => 
                           bus_selected_win_data_3_port, Q(258) => 
                           bus_selected_win_data_2_port, Q(257) => 
                           bus_selected_win_data_1_port, Q(256) => 
                           bus_selected_win_data_0_port, Q(255) => 
                           bus_complete_win_data_255_port, Q(254) => 
                           bus_complete_win_data_254_port, Q(253) => 
                           bus_complete_win_data_253_port, Q(252) => 
                           bus_complete_win_data_252_port, Q(251) => 
                           bus_complete_win_data_251_port, Q(250) => 
                           bus_complete_win_data_250_port, Q(249) => 
                           bus_complete_win_data_249_port, Q(248) => 
                           bus_complete_win_data_248_port, Q(247) => 
                           bus_complete_win_data_247_port, Q(246) => 
                           bus_complete_win_data_246_port, Q(245) => 
                           bus_complete_win_data_245_port, Q(244) => 
                           bus_complete_win_data_244_port, Q(243) => 
                           bus_complete_win_data_243_port, Q(242) => 
                           bus_complete_win_data_242_port, Q(241) => 
                           bus_complete_win_data_241_port, Q(240) => 
                           bus_complete_win_data_240_port, Q(239) => 
                           bus_complete_win_data_239_port, Q(238) => 
                           bus_complete_win_data_238_port, Q(237) => 
                           bus_complete_win_data_237_port, Q(236) => 
                           bus_complete_win_data_236_port, Q(235) => 
                           bus_complete_win_data_235_port, Q(234) => 
                           bus_complete_win_data_234_port, Q(233) => 
                           bus_complete_win_data_233_port, Q(232) => 
                           bus_complete_win_data_232_port, Q(231) => 
                           bus_complete_win_data_231_port, Q(230) => 
                           bus_complete_win_data_230_port, Q(229) => 
                           bus_complete_win_data_229_port, Q(228) => 
                           bus_complete_win_data_228_port, Q(227) => 
                           bus_complete_win_data_227_port, Q(226) => 
                           bus_complete_win_data_226_port, Q(225) => 
                           bus_complete_win_data_225_port, Q(224) => 
                           bus_complete_win_data_224_port, Q(223) => 
                           bus_complete_win_data_223_port, Q(222) => 
                           bus_complete_win_data_222_port, Q(221) => 
                           bus_complete_win_data_221_port, Q(220) => 
                           bus_complete_win_data_220_port, Q(219) => 
                           bus_complete_win_data_219_port, Q(218) => 
                           bus_complete_win_data_218_port, Q(217) => 
                           bus_complete_win_data_217_port, Q(216) => 
                           bus_complete_win_data_216_port, Q(215) => 
                           bus_complete_win_data_215_port, Q(214) => 
                           bus_complete_win_data_214_port, Q(213) => 
                           bus_complete_win_data_213_port, Q(212) => 
                           bus_complete_win_data_212_port, Q(211) => 
                           bus_complete_win_data_211_port, Q(210) => 
                           bus_complete_win_data_210_port, Q(209) => 
                           bus_complete_win_data_209_port, Q(208) => 
                           bus_complete_win_data_208_port, Q(207) => 
                           bus_complete_win_data_207_port, Q(206) => 
                           bus_complete_win_data_206_port, Q(205) => 
                           bus_complete_win_data_205_port, Q(204) => 
                           bus_complete_win_data_204_port, Q(203) => 
                           bus_complete_win_data_203_port, Q(202) => 
                           bus_complete_win_data_202_port, Q(201) => 
                           bus_complete_win_data_201_port, Q(200) => 
                           bus_complete_win_data_200_port, Q(199) => 
                           bus_complete_win_data_199_port, Q(198) => 
                           bus_complete_win_data_198_port, Q(197) => 
                           bus_complete_win_data_197_port, Q(196) => 
                           bus_complete_win_data_196_port, Q(195) => 
                           bus_complete_win_data_195_port, Q(194) => 
                           bus_complete_win_data_194_port, Q(193) => 
                           bus_complete_win_data_193_port, Q(192) => 
                           bus_complete_win_data_192_port, Q(191) => 
                           bus_complete_win_data_191_port, Q(190) => 
                           bus_complete_win_data_190_port, Q(189) => 
                           bus_complete_win_data_189_port, Q(188) => 
                           bus_complete_win_data_188_port, Q(187) => 
                           bus_complete_win_data_187_port, Q(186) => 
                           bus_complete_win_data_186_port, Q(185) => 
                           bus_complete_win_data_185_port, Q(184) => 
                           bus_complete_win_data_184_port, Q(183) => 
                           bus_complete_win_data_183_port, Q(182) => 
                           bus_complete_win_data_182_port, Q(181) => 
                           bus_complete_win_data_181_port, Q(180) => 
                           bus_complete_win_data_180_port, Q(179) => 
                           bus_complete_win_data_179_port, Q(178) => 
                           bus_complete_win_data_178_port, Q(177) => 
                           bus_complete_win_data_177_port, Q(176) => 
                           bus_complete_win_data_176_port, Q(175) => 
                           bus_complete_win_data_175_port, Q(174) => 
                           bus_complete_win_data_174_port, Q(173) => 
                           bus_complete_win_data_173_port, Q(172) => 
                           bus_complete_win_data_172_port, Q(171) => 
                           bus_complete_win_data_171_port, Q(170) => 
                           bus_complete_win_data_170_port, Q(169) => 
                           bus_complete_win_data_169_port, Q(168) => 
                           bus_complete_win_data_168_port, Q(167) => 
                           bus_complete_win_data_167_port, Q(166) => 
                           bus_complete_win_data_166_port, Q(165) => 
                           bus_complete_win_data_165_port, Q(164) => 
                           bus_complete_win_data_164_port, Q(163) => 
                           bus_complete_win_data_163_port, Q(162) => 
                           bus_complete_win_data_162_port, Q(161) => 
                           bus_complete_win_data_161_port, Q(160) => 
                           bus_complete_win_data_160_port, Q(159) => 
                           bus_complete_win_data_159_port, Q(158) => 
                           bus_complete_win_data_158_port, Q(157) => 
                           bus_complete_win_data_157_port, Q(156) => 
                           bus_complete_win_data_156_port, Q(155) => 
                           bus_complete_win_data_155_port, Q(154) => 
                           bus_complete_win_data_154_port, Q(153) => 
                           bus_complete_win_data_153_port, Q(152) => 
                           bus_complete_win_data_152_port, Q(151) => 
                           bus_complete_win_data_151_port, Q(150) => 
                           bus_complete_win_data_150_port, Q(149) => 
                           bus_complete_win_data_149_port, Q(148) => 
                           bus_complete_win_data_148_port, Q(147) => 
                           bus_complete_win_data_147_port, Q(146) => 
                           bus_complete_win_data_146_port, Q(145) => 
                           bus_complete_win_data_145_port, Q(144) => 
                           bus_complete_win_data_144_port, Q(143) => 
                           bus_complete_win_data_143_port, Q(142) => 
                           bus_complete_win_data_142_port, Q(141) => 
                           bus_complete_win_data_141_port, Q(140) => 
                           bus_complete_win_data_140_port, Q(139) => 
                           bus_complete_win_data_139_port, Q(138) => 
                           bus_complete_win_data_138_port, Q(137) => 
                           bus_complete_win_data_137_port, Q(136) => 
                           bus_complete_win_data_136_port, Q(135) => 
                           bus_complete_win_data_135_port, Q(134) => 
                           bus_complete_win_data_134_port, Q(133) => 
                           bus_complete_win_data_133_port, Q(132) => 
                           bus_complete_win_data_132_port, Q(131) => 
                           bus_complete_win_data_131_port, Q(130) => 
                           bus_complete_win_data_130_port, Q(129) => 
                           bus_complete_win_data_129_port, Q(128) => 
                           bus_complete_win_data_128_port, Q(127) => 
                           bus_complete_win_data_127_port, Q(126) => 
                           bus_complete_win_data_126_port, Q(125) => 
                           bus_complete_win_data_125_port, Q(124) => 
                           bus_complete_win_data_124_port, Q(123) => 
                           bus_complete_win_data_123_port, Q(122) => 
                           bus_complete_win_data_122_port, Q(121) => 
                           bus_complete_win_data_121_port, Q(120) => 
                           bus_complete_win_data_120_port, Q(119) => 
                           bus_complete_win_data_119_port, Q(118) => 
                           bus_complete_win_data_118_port, Q(117) => 
                           bus_complete_win_data_117_port, Q(116) => 
                           bus_complete_win_data_116_port, Q(115) => 
                           bus_complete_win_data_115_port, Q(114) => 
                           bus_complete_win_data_114_port, Q(113) => 
                           bus_complete_win_data_113_port, Q(112) => 
                           bus_complete_win_data_112_port, Q(111) => 
                           bus_complete_win_data_111_port, Q(110) => 
                           bus_complete_win_data_110_port, Q(109) => 
                           bus_complete_win_data_109_port, Q(108) => 
                           bus_complete_win_data_108_port, Q(107) => 
                           bus_complete_win_data_107_port, Q(106) => 
                           bus_complete_win_data_106_port, Q(105) => 
                           bus_complete_win_data_105_port, Q(104) => 
                           bus_complete_win_data_104_port, Q(103) => 
                           bus_complete_win_data_103_port, Q(102) => 
                           bus_complete_win_data_102_port, Q(101) => 
                           bus_complete_win_data_101_port, Q(100) => 
                           bus_complete_win_data_100_port, Q(99) => 
                           bus_complete_win_data_99_port, Q(98) => 
                           bus_complete_win_data_98_port, Q(97) => 
                           bus_complete_win_data_97_port, Q(96) => 
                           bus_complete_win_data_96_port, Q(95) => 
                           bus_complete_win_data_95_port, Q(94) => 
                           bus_complete_win_data_94_port, Q(93) => 
                           bus_complete_win_data_93_port, Q(92) => 
                           bus_complete_win_data_92_port, Q(91) => 
                           bus_complete_win_data_91_port, Q(90) => 
                           bus_complete_win_data_90_port, Q(89) => 
                           bus_complete_win_data_89_port, Q(88) => 
                           bus_complete_win_data_88_port, Q(87) => 
                           bus_complete_win_data_87_port, Q(86) => 
                           bus_complete_win_data_86_port, Q(85) => 
                           bus_complete_win_data_85_port, Q(84) => 
                           bus_complete_win_data_84_port, Q(83) => 
                           bus_complete_win_data_83_port, Q(82) => 
                           bus_complete_win_data_82_port, Q(81) => 
                           bus_complete_win_data_81_port, Q(80) => 
                           bus_complete_win_data_80_port, Q(79) => 
                           bus_complete_win_data_79_port, Q(78) => 
                           bus_complete_win_data_78_port, Q(77) => 
                           bus_complete_win_data_77_port, Q(76) => 
                           bus_complete_win_data_76_port, Q(75) => 
                           bus_complete_win_data_75_port, Q(74) => 
                           bus_complete_win_data_74_port, Q(73) => 
                           bus_complete_win_data_73_port, Q(72) => 
                           bus_complete_win_data_72_port, Q(71) => 
                           bus_complete_win_data_71_port, Q(70) => 
                           bus_complete_win_data_70_port, Q(69) => 
                           bus_complete_win_data_69_port, Q(68) => 
                           bus_complete_win_data_68_port, Q(67) => 
                           bus_complete_win_data_67_port, Q(66) => 
                           bus_complete_win_data_66_port, Q(65) => 
                           bus_complete_win_data_65_port, Q(64) => 
                           bus_complete_win_data_64_port, Q(63) => 
                           bus_complete_win_data_63_port, Q(62) => 
                           bus_complete_win_data_62_port, Q(61) => 
                           bus_complete_win_data_61_port, Q(60) => 
                           bus_complete_win_data_60_port, Q(59) => 
                           bus_complete_win_data_59_port, Q(58) => 
                           bus_complete_win_data_58_port, Q(57) => 
                           bus_complete_win_data_57_port, Q(56) => 
                           bus_complete_win_data_56_port, Q(55) => 
                           bus_complete_win_data_55_port, Q(54) => 
                           bus_complete_win_data_54_port, Q(53) => 
                           bus_complete_win_data_53_port, Q(52) => 
                           bus_complete_win_data_52_port, Q(51) => 
                           bus_complete_win_data_51_port, Q(50) => 
                           bus_complete_win_data_50_port, Q(49) => 
                           bus_complete_win_data_49_port, Q(48) => 
                           bus_complete_win_data_48_port, Q(47) => 
                           bus_complete_win_data_47_port, Q(46) => 
                           bus_complete_win_data_46_port, Q(45) => 
                           bus_complete_win_data_45_port, Q(44) => 
                           bus_complete_win_data_44_port, Q(43) => 
                           bus_complete_win_data_43_port, Q(42) => 
                           bus_complete_win_data_42_port, Q(41) => 
                           bus_complete_win_data_41_port, Q(40) => 
                           bus_complete_win_data_40_port, Q(39) => 
                           bus_complete_win_data_39_port, Q(38) => 
                           bus_complete_win_data_38_port, Q(37) => 
                           bus_complete_win_data_37_port, Q(36) => 
                           bus_complete_win_data_36_port, Q(35) => 
                           bus_complete_win_data_35_port, Q(34) => 
                           bus_complete_win_data_34_port, Q(33) => 
                           bus_complete_win_data_33_port, Q(32) => 
                           bus_complete_win_data_32_port, Q(31) => 
                           bus_complete_win_data_31_port, Q(30) => 
                           bus_complete_win_data_30_port, Q(29) => 
                           bus_complete_win_data_29_port, Q(28) => 
                           bus_complete_win_data_28_port, Q(27) => 
                           bus_complete_win_data_27_port, Q(26) => 
                           bus_complete_win_data_26_port, Q(25) => 
                           bus_complete_win_data_25_port, Q(24) => 
                           bus_complete_win_data_24_port, Q(23) => 
                           bus_complete_win_data_23_port, Q(22) => 
                           bus_complete_win_data_22_port, Q(21) => 
                           bus_complete_win_data_21_port, Q(20) => 
                           bus_complete_win_data_20_port, Q(19) => 
                           bus_complete_win_data_19_port, Q(18) => 
                           bus_complete_win_data_18_port, Q(17) => 
                           bus_complete_win_data_17_port, Q(16) => 
                           bus_complete_win_data_16_port, Q(15) => 
                           bus_complete_win_data_15_port, Q(14) => 
                           bus_complete_win_data_14_port, Q(13) => 
                           bus_complete_win_data_13_port, Q(12) => 
                           bus_complete_win_data_12_port, Q(11) => 
                           bus_complete_win_data_11_port, Q(10) => 
                           bus_complete_win_data_10_port, Q(9) => 
                           bus_complete_win_data_9_port, Q(8) => 
                           bus_complete_win_data_8_port, Q(7) => 
                           bus_complete_win_data_7_port, Q(6) => 
                           bus_complete_win_data_6_port, Q(5) => 
                           bus_complete_win_data_5_port, Q(4) => 
                           bus_complete_win_data_4_port, Q(3) => 
                           bus_complete_win_data_3_port, Q(2) => 
                           bus_complete_win_data_2_port, Q(1) => 
                           bus_complete_win_data_1_port, Q(0) => 
                           bus_complete_win_data_0_port, Y(31) => 
                           internal_out1_31_port, Y(30) => 
                           internal_out1_30_port, Y(29) => 
                           internal_out1_29_port, Y(28) => 
                           internal_out1_28_port, Y(27) => 
                           internal_out1_27_port, Y(26) => 
                           internal_out1_26_port, Y(25) => 
                           internal_out1_25_port, Y(24) => 
                           internal_out1_24_port, Y(23) => 
                           internal_out1_23_port, Y(22) => 
                           internal_out1_22_port, Y(21) => 
                           internal_out1_21_port, Y(20) => 
                           internal_out1_20_port, Y(19) => 
                           internal_out1_19_port, Y(18) => 
                           internal_out1_18_port, Y(17) => 
                           internal_out1_17_port, Y(16) => 
                           internal_out1_16_port, Y(15) => 
                           internal_out1_15_port, Y(14) => 
                           internal_out1_14_port, Y(13) => 
                           internal_out1_13_port, Y(12) => 
                           internal_out1_12_port, Y(11) => 
                           internal_out1_11_port, Y(10) => 
                           internal_out1_10_port, Y(9) => internal_out1_9_port,
                           Y(8) => internal_out1_8_port, Y(7) => 
                           internal_out1_7_port, Y(6) => internal_out1_6_port, 
                           Y(5) => internal_out1_5_port, Y(4) => 
                           internal_out1_4_port, Y(3) => internal_out1_3_port, 
                           Y(2) => internal_out1_2_port, Y(1) => 
                           internal_out1_1_port, Y(0) => internal_out1_0_port);
   RDPORT0_OUTREG : reg_generic_N32_RSTVAL0_0 port map( D(31) => 
                           internal_out1_31_port, D(30) => 
                           internal_out1_30_port, D(29) => 
                           internal_out1_29_port, D(28) => 
                           internal_out1_28_port, D(27) => 
                           internal_out1_27_port, D(26) => 
                           internal_out1_26_port, D(25) => 
                           internal_out1_25_port, D(24) => 
                           internal_out1_24_port, D(23) => 
                           internal_out1_23_port, D(22) => 
                           internal_out1_22_port, D(21) => 
                           internal_out1_21_port, D(20) => 
                           internal_out1_20_port, D(19) => 
                           internal_out1_19_port, D(18) => 
                           internal_out1_18_port, D(17) => 
                           internal_out1_17_port, D(16) => 
                           internal_out1_16_port, D(15) => 
                           internal_out1_15_port, D(14) => 
                           internal_out1_14_port, D(13) => 
                           internal_out1_13_port, D(12) => 
                           internal_out1_12_port, D(11) => 
                           internal_out1_11_port, D(10) => 
                           internal_out1_10_port, D(9) => internal_out1_9_port,
                           D(8) => internal_out1_8_port, D(7) => 
                           internal_out1_7_port, D(6) => internal_out1_6_port, 
                           D(5) => internal_out1_5_port, D(4) => 
                           internal_out1_4_port, D(3) => internal_out1_3_port, 
                           D(2) => internal_out1_2_port, D(1) => 
                           internal_out1_1_port, D(0) => internal_out1_0_port, 
                           Q(31) => OUT1(31), Q(30) => OUT1(30), Q(29) => 
                           OUT1(29), Q(28) => OUT1(28), Q(27) => OUT1(27), 
                           Q(26) => OUT1(26), Q(25) => OUT1(25), Q(24) => 
                           OUT1(24), Q(23) => OUT1(23), Q(22) => OUT1(22), 
                           Q(21) => OUT1(21), Q(20) => OUT1(20), Q(19) => 
                           OUT1(19), Q(18) => OUT1(18), Q(17) => OUT1(17), 
                           Q(16) => OUT1(16), Q(15) => OUT1(15), Q(14) => 
                           OUT1(14), Q(13) => OUT1(13), Q(12) => OUT1(12), 
                           Q(11) => OUT1(11), Q(10) => OUT1(10), Q(9) => 
                           OUT1(9), Q(8) => OUT1(8), Q(7) => OUT1(7), Q(6) => 
                           OUT1(6), Q(5) => OUT1(5), Q(4) => OUT1(4), Q(3) => 
                           OUT1(3), Q(2) => OUT1(2), Q(1) => OUT1(1), Q(0) => 
                           OUT1(0), Clk => CLK, Rst => RESET, Enable => int_RD1
                           );
   RDPORT1 : mux_N32_M5_1 port map( S(4) => ADD_RD2(4), S(3) => ADD_RD2(3), 
                           S(2) => ADD_RD2(2), S(1) => ADD_RD2(1), S(0) => 
                           ADD_RD2(0), Q(1023) => 
                           bus_selected_win_data_767_port, Q(1022) => 
                           bus_selected_win_data_766_port, Q(1021) => 
                           bus_selected_win_data_765_port, Q(1020) => 
                           bus_selected_win_data_764_port, Q(1019) => 
                           bus_selected_win_data_763_port, Q(1018) => 
                           bus_selected_win_data_762_port, Q(1017) => 
                           bus_selected_win_data_761_port, Q(1016) => 
                           bus_selected_win_data_760_port, Q(1015) => 
                           bus_selected_win_data_759_port, Q(1014) => 
                           bus_selected_win_data_758_port, Q(1013) => 
                           bus_selected_win_data_757_port, Q(1012) => 
                           bus_selected_win_data_756_port, Q(1011) => 
                           bus_selected_win_data_755_port, Q(1010) => 
                           bus_selected_win_data_754_port, Q(1009) => 
                           bus_selected_win_data_753_port, Q(1008) => 
                           bus_selected_win_data_752_port, Q(1007) => 
                           bus_selected_win_data_751_port, Q(1006) => 
                           bus_selected_win_data_750_port, Q(1005) => 
                           bus_selected_win_data_749_port, Q(1004) => 
                           bus_selected_win_data_748_port, Q(1003) => 
                           bus_selected_win_data_747_port, Q(1002) => 
                           bus_selected_win_data_746_port, Q(1001) => 
                           bus_selected_win_data_745_port, Q(1000) => 
                           bus_selected_win_data_744_port, Q(999) => 
                           bus_selected_win_data_743_port, Q(998) => 
                           bus_selected_win_data_742_port, Q(997) => 
                           bus_selected_win_data_741_port, Q(996) => 
                           bus_selected_win_data_740_port, Q(995) => 
                           bus_selected_win_data_739_port, Q(994) => 
                           bus_selected_win_data_738_port, Q(993) => 
                           bus_selected_win_data_737_port, Q(992) => 
                           bus_selected_win_data_736_port, Q(991) => 
                           bus_selected_win_data_735_port, Q(990) => 
                           bus_selected_win_data_734_port, Q(989) => 
                           bus_selected_win_data_733_port, Q(988) => 
                           bus_selected_win_data_732_port, Q(987) => 
                           bus_selected_win_data_731_port, Q(986) => 
                           bus_selected_win_data_730_port, Q(985) => 
                           bus_selected_win_data_729_port, Q(984) => 
                           bus_selected_win_data_728_port, Q(983) => 
                           bus_selected_win_data_727_port, Q(982) => 
                           bus_selected_win_data_726_port, Q(981) => 
                           bus_selected_win_data_725_port, Q(980) => 
                           bus_selected_win_data_724_port, Q(979) => 
                           bus_selected_win_data_723_port, Q(978) => 
                           bus_selected_win_data_722_port, Q(977) => 
                           bus_selected_win_data_721_port, Q(976) => 
                           bus_selected_win_data_720_port, Q(975) => 
                           bus_selected_win_data_719_port, Q(974) => 
                           bus_selected_win_data_718_port, Q(973) => 
                           bus_selected_win_data_717_port, Q(972) => 
                           bus_selected_win_data_716_port, Q(971) => 
                           bus_selected_win_data_715_port, Q(970) => 
                           bus_selected_win_data_714_port, Q(969) => 
                           bus_selected_win_data_713_port, Q(968) => 
                           bus_selected_win_data_712_port, Q(967) => 
                           bus_selected_win_data_711_port, Q(966) => 
                           bus_selected_win_data_710_port, Q(965) => 
                           bus_selected_win_data_709_port, Q(964) => 
                           bus_selected_win_data_708_port, Q(963) => 
                           bus_selected_win_data_707_port, Q(962) => 
                           bus_selected_win_data_706_port, Q(961) => 
                           bus_selected_win_data_705_port, Q(960) => 
                           bus_selected_win_data_704_port, Q(959) => 
                           bus_selected_win_data_703_port, Q(958) => 
                           bus_selected_win_data_702_port, Q(957) => 
                           bus_selected_win_data_701_port, Q(956) => 
                           bus_selected_win_data_700_port, Q(955) => 
                           bus_selected_win_data_699_port, Q(954) => 
                           bus_selected_win_data_698_port, Q(953) => 
                           bus_selected_win_data_697_port, Q(952) => 
                           bus_selected_win_data_696_port, Q(951) => 
                           bus_selected_win_data_695_port, Q(950) => 
                           bus_selected_win_data_694_port, Q(949) => 
                           bus_selected_win_data_693_port, Q(948) => 
                           bus_selected_win_data_692_port, Q(947) => 
                           bus_selected_win_data_691_port, Q(946) => 
                           bus_selected_win_data_690_port, Q(945) => 
                           bus_selected_win_data_689_port, Q(944) => 
                           bus_selected_win_data_688_port, Q(943) => 
                           bus_selected_win_data_687_port, Q(942) => 
                           bus_selected_win_data_686_port, Q(941) => 
                           bus_selected_win_data_685_port, Q(940) => 
                           bus_selected_win_data_684_port, Q(939) => 
                           bus_selected_win_data_683_port, Q(938) => 
                           bus_selected_win_data_682_port, Q(937) => 
                           bus_selected_win_data_681_port, Q(936) => 
                           bus_selected_win_data_680_port, Q(935) => 
                           bus_selected_win_data_679_port, Q(934) => 
                           bus_selected_win_data_678_port, Q(933) => 
                           bus_selected_win_data_677_port, Q(932) => 
                           bus_selected_win_data_676_port, Q(931) => 
                           bus_selected_win_data_675_port, Q(930) => 
                           bus_selected_win_data_674_port, Q(929) => 
                           bus_selected_win_data_673_port, Q(928) => 
                           bus_selected_win_data_672_port, Q(927) => 
                           bus_selected_win_data_671_port, Q(926) => 
                           bus_selected_win_data_670_port, Q(925) => 
                           bus_selected_win_data_669_port, Q(924) => 
                           bus_selected_win_data_668_port, Q(923) => 
                           bus_selected_win_data_667_port, Q(922) => 
                           bus_selected_win_data_666_port, Q(921) => 
                           bus_selected_win_data_665_port, Q(920) => 
                           bus_selected_win_data_664_port, Q(919) => 
                           bus_selected_win_data_663_port, Q(918) => 
                           bus_selected_win_data_662_port, Q(917) => 
                           bus_selected_win_data_661_port, Q(916) => 
                           bus_selected_win_data_660_port, Q(915) => 
                           bus_selected_win_data_659_port, Q(914) => 
                           bus_selected_win_data_658_port, Q(913) => 
                           bus_selected_win_data_657_port, Q(912) => 
                           bus_selected_win_data_656_port, Q(911) => 
                           bus_selected_win_data_655_port, Q(910) => 
                           bus_selected_win_data_654_port, Q(909) => 
                           bus_selected_win_data_653_port, Q(908) => 
                           bus_selected_win_data_652_port, Q(907) => 
                           bus_selected_win_data_651_port, Q(906) => 
                           bus_selected_win_data_650_port, Q(905) => 
                           bus_selected_win_data_649_port, Q(904) => 
                           bus_selected_win_data_648_port, Q(903) => 
                           bus_selected_win_data_647_port, Q(902) => 
                           bus_selected_win_data_646_port, Q(901) => 
                           bus_selected_win_data_645_port, Q(900) => 
                           bus_selected_win_data_644_port, Q(899) => 
                           bus_selected_win_data_643_port, Q(898) => 
                           bus_selected_win_data_642_port, Q(897) => 
                           bus_selected_win_data_641_port, Q(896) => 
                           bus_selected_win_data_640_port, Q(895) => 
                           bus_selected_win_data_639_port, Q(894) => 
                           bus_selected_win_data_638_port, Q(893) => 
                           bus_selected_win_data_637_port, Q(892) => 
                           bus_selected_win_data_636_port, Q(891) => 
                           bus_selected_win_data_635_port, Q(890) => 
                           bus_selected_win_data_634_port, Q(889) => 
                           bus_selected_win_data_633_port, Q(888) => 
                           bus_selected_win_data_632_port, Q(887) => 
                           bus_selected_win_data_631_port, Q(886) => 
                           bus_selected_win_data_630_port, Q(885) => 
                           bus_selected_win_data_629_port, Q(884) => 
                           bus_selected_win_data_628_port, Q(883) => 
                           bus_selected_win_data_627_port, Q(882) => 
                           bus_selected_win_data_626_port, Q(881) => 
                           bus_selected_win_data_625_port, Q(880) => 
                           bus_selected_win_data_624_port, Q(879) => 
                           bus_selected_win_data_623_port, Q(878) => 
                           bus_selected_win_data_622_port, Q(877) => 
                           bus_selected_win_data_621_port, Q(876) => 
                           bus_selected_win_data_620_port, Q(875) => 
                           bus_selected_win_data_619_port, Q(874) => 
                           bus_selected_win_data_618_port, Q(873) => 
                           bus_selected_win_data_617_port, Q(872) => 
                           bus_selected_win_data_616_port, Q(871) => 
                           bus_selected_win_data_615_port, Q(870) => 
                           bus_selected_win_data_614_port, Q(869) => 
                           bus_selected_win_data_613_port, Q(868) => 
                           bus_selected_win_data_612_port, Q(867) => 
                           bus_selected_win_data_611_port, Q(866) => 
                           bus_selected_win_data_610_port, Q(865) => 
                           bus_selected_win_data_609_port, Q(864) => 
                           bus_selected_win_data_608_port, Q(863) => 
                           bus_selected_win_data_607_port, Q(862) => 
                           bus_selected_win_data_606_port, Q(861) => 
                           bus_selected_win_data_605_port, Q(860) => 
                           bus_selected_win_data_604_port, Q(859) => 
                           bus_selected_win_data_603_port, Q(858) => 
                           bus_selected_win_data_602_port, Q(857) => 
                           bus_selected_win_data_601_port, Q(856) => 
                           bus_selected_win_data_600_port, Q(855) => 
                           bus_selected_win_data_599_port, Q(854) => 
                           bus_selected_win_data_598_port, Q(853) => 
                           bus_selected_win_data_597_port, Q(852) => 
                           bus_selected_win_data_596_port, Q(851) => 
                           bus_selected_win_data_595_port, Q(850) => 
                           bus_selected_win_data_594_port, Q(849) => 
                           bus_selected_win_data_593_port, Q(848) => 
                           bus_selected_win_data_592_port, Q(847) => 
                           bus_selected_win_data_591_port, Q(846) => 
                           bus_selected_win_data_590_port, Q(845) => 
                           bus_selected_win_data_589_port, Q(844) => 
                           bus_selected_win_data_588_port, Q(843) => 
                           bus_selected_win_data_587_port, Q(842) => 
                           bus_selected_win_data_586_port, Q(841) => 
                           bus_selected_win_data_585_port, Q(840) => 
                           bus_selected_win_data_584_port, Q(839) => 
                           bus_selected_win_data_583_port, Q(838) => 
                           bus_selected_win_data_582_port, Q(837) => 
                           bus_selected_win_data_581_port, Q(836) => 
                           bus_selected_win_data_580_port, Q(835) => 
                           bus_selected_win_data_579_port, Q(834) => 
                           bus_selected_win_data_578_port, Q(833) => 
                           bus_selected_win_data_577_port, Q(832) => 
                           bus_selected_win_data_576_port, Q(831) => 
                           bus_selected_win_data_575_port, Q(830) => 
                           bus_selected_win_data_574_port, Q(829) => 
                           bus_selected_win_data_573_port, Q(828) => 
                           bus_selected_win_data_572_port, Q(827) => 
                           bus_selected_win_data_571_port, Q(826) => 
                           bus_selected_win_data_570_port, Q(825) => 
                           bus_selected_win_data_569_port, Q(824) => 
                           bus_selected_win_data_568_port, Q(823) => 
                           bus_selected_win_data_567_port, Q(822) => 
                           bus_selected_win_data_566_port, Q(821) => 
                           bus_selected_win_data_565_port, Q(820) => 
                           bus_selected_win_data_564_port, Q(819) => 
                           bus_selected_win_data_563_port, Q(818) => 
                           bus_selected_win_data_562_port, Q(817) => 
                           bus_selected_win_data_561_port, Q(816) => 
                           bus_selected_win_data_560_port, Q(815) => 
                           bus_selected_win_data_559_port, Q(814) => 
                           bus_selected_win_data_558_port, Q(813) => 
                           bus_selected_win_data_557_port, Q(812) => 
                           bus_selected_win_data_556_port, Q(811) => 
                           bus_selected_win_data_555_port, Q(810) => 
                           bus_selected_win_data_554_port, Q(809) => 
                           bus_selected_win_data_553_port, Q(808) => 
                           bus_selected_win_data_552_port, Q(807) => 
                           bus_selected_win_data_551_port, Q(806) => 
                           bus_selected_win_data_550_port, Q(805) => 
                           bus_selected_win_data_549_port, Q(804) => 
                           bus_selected_win_data_548_port, Q(803) => 
                           bus_selected_win_data_547_port, Q(802) => 
                           bus_selected_win_data_546_port, Q(801) => 
                           bus_selected_win_data_545_port, Q(800) => 
                           bus_selected_win_data_544_port, Q(799) => 
                           bus_selected_win_data_543_port, Q(798) => 
                           bus_selected_win_data_542_port, Q(797) => 
                           bus_selected_win_data_541_port, Q(796) => 
                           bus_selected_win_data_540_port, Q(795) => 
                           bus_selected_win_data_539_port, Q(794) => 
                           bus_selected_win_data_538_port, Q(793) => 
                           bus_selected_win_data_537_port, Q(792) => 
                           bus_selected_win_data_536_port, Q(791) => 
                           bus_selected_win_data_535_port, Q(790) => 
                           bus_selected_win_data_534_port, Q(789) => 
                           bus_selected_win_data_533_port, Q(788) => 
                           bus_selected_win_data_532_port, Q(787) => 
                           bus_selected_win_data_531_port, Q(786) => 
                           bus_selected_win_data_530_port, Q(785) => 
                           bus_selected_win_data_529_port, Q(784) => 
                           bus_selected_win_data_528_port, Q(783) => 
                           bus_selected_win_data_527_port, Q(782) => 
                           bus_selected_win_data_526_port, Q(781) => 
                           bus_selected_win_data_525_port, Q(780) => 
                           bus_selected_win_data_524_port, Q(779) => 
                           bus_selected_win_data_523_port, Q(778) => 
                           bus_selected_win_data_522_port, Q(777) => 
                           bus_selected_win_data_521_port, Q(776) => 
                           bus_selected_win_data_520_port, Q(775) => 
                           bus_selected_win_data_519_port, Q(774) => 
                           bus_selected_win_data_518_port, Q(773) => 
                           bus_selected_win_data_517_port, Q(772) => 
                           bus_selected_win_data_516_port, Q(771) => 
                           bus_selected_win_data_515_port, Q(770) => 
                           bus_selected_win_data_514_port, Q(769) => 
                           bus_selected_win_data_513_port, Q(768) => 
                           bus_selected_win_data_512_port, Q(767) => 
                           bus_selected_win_data_511_port, Q(766) => 
                           bus_selected_win_data_510_port, Q(765) => 
                           bus_selected_win_data_509_port, Q(764) => 
                           bus_selected_win_data_508_port, Q(763) => 
                           bus_selected_win_data_507_port, Q(762) => 
                           bus_selected_win_data_506_port, Q(761) => 
                           bus_selected_win_data_505_port, Q(760) => 
                           bus_selected_win_data_504_port, Q(759) => 
                           bus_selected_win_data_503_port, Q(758) => 
                           bus_selected_win_data_502_port, Q(757) => 
                           bus_selected_win_data_501_port, Q(756) => 
                           bus_selected_win_data_500_port, Q(755) => 
                           bus_selected_win_data_499_port, Q(754) => 
                           bus_selected_win_data_498_port, Q(753) => 
                           bus_selected_win_data_497_port, Q(752) => 
                           bus_selected_win_data_496_port, Q(751) => 
                           bus_selected_win_data_495_port, Q(750) => 
                           bus_selected_win_data_494_port, Q(749) => 
                           bus_selected_win_data_493_port, Q(748) => 
                           bus_selected_win_data_492_port, Q(747) => 
                           bus_selected_win_data_491_port, Q(746) => 
                           bus_selected_win_data_490_port, Q(745) => 
                           bus_selected_win_data_489_port, Q(744) => 
                           bus_selected_win_data_488_port, Q(743) => 
                           bus_selected_win_data_487_port, Q(742) => 
                           bus_selected_win_data_486_port, Q(741) => 
                           bus_selected_win_data_485_port, Q(740) => 
                           bus_selected_win_data_484_port, Q(739) => 
                           bus_selected_win_data_483_port, Q(738) => 
                           bus_selected_win_data_482_port, Q(737) => 
                           bus_selected_win_data_481_port, Q(736) => 
                           bus_selected_win_data_480_port, Q(735) => 
                           bus_selected_win_data_479_port, Q(734) => 
                           bus_selected_win_data_478_port, Q(733) => 
                           bus_selected_win_data_477_port, Q(732) => 
                           bus_selected_win_data_476_port, Q(731) => 
                           bus_selected_win_data_475_port, Q(730) => 
                           bus_selected_win_data_474_port, Q(729) => 
                           bus_selected_win_data_473_port, Q(728) => 
                           bus_selected_win_data_472_port, Q(727) => 
                           bus_selected_win_data_471_port, Q(726) => 
                           bus_selected_win_data_470_port, Q(725) => 
                           bus_selected_win_data_469_port, Q(724) => 
                           bus_selected_win_data_468_port, Q(723) => 
                           bus_selected_win_data_467_port, Q(722) => 
                           bus_selected_win_data_466_port, Q(721) => 
                           bus_selected_win_data_465_port, Q(720) => 
                           bus_selected_win_data_464_port, Q(719) => 
                           bus_selected_win_data_463_port, Q(718) => 
                           bus_selected_win_data_462_port, Q(717) => 
                           bus_selected_win_data_461_port, Q(716) => 
                           bus_selected_win_data_460_port, Q(715) => 
                           bus_selected_win_data_459_port, Q(714) => 
                           bus_selected_win_data_458_port, Q(713) => 
                           bus_selected_win_data_457_port, Q(712) => 
                           bus_selected_win_data_456_port, Q(711) => 
                           bus_selected_win_data_455_port, Q(710) => 
                           bus_selected_win_data_454_port, Q(709) => 
                           bus_selected_win_data_453_port, Q(708) => 
                           bus_selected_win_data_452_port, Q(707) => 
                           bus_selected_win_data_451_port, Q(706) => 
                           bus_selected_win_data_450_port, Q(705) => 
                           bus_selected_win_data_449_port, Q(704) => 
                           bus_selected_win_data_448_port, Q(703) => 
                           bus_selected_win_data_447_port, Q(702) => 
                           bus_selected_win_data_446_port, Q(701) => 
                           bus_selected_win_data_445_port, Q(700) => 
                           bus_selected_win_data_444_port, Q(699) => 
                           bus_selected_win_data_443_port, Q(698) => 
                           bus_selected_win_data_442_port, Q(697) => 
                           bus_selected_win_data_441_port, Q(696) => 
                           bus_selected_win_data_440_port, Q(695) => 
                           bus_selected_win_data_439_port, Q(694) => 
                           bus_selected_win_data_438_port, Q(693) => 
                           bus_selected_win_data_437_port, Q(692) => 
                           bus_selected_win_data_436_port, Q(691) => 
                           bus_selected_win_data_435_port, Q(690) => 
                           bus_selected_win_data_434_port, Q(689) => 
                           bus_selected_win_data_433_port, Q(688) => 
                           bus_selected_win_data_432_port, Q(687) => 
                           bus_selected_win_data_431_port, Q(686) => 
                           bus_selected_win_data_430_port, Q(685) => 
                           bus_selected_win_data_429_port, Q(684) => 
                           bus_selected_win_data_428_port, Q(683) => 
                           bus_selected_win_data_427_port, Q(682) => 
                           bus_selected_win_data_426_port, Q(681) => 
                           bus_selected_win_data_425_port, Q(680) => 
                           bus_selected_win_data_424_port, Q(679) => 
                           bus_selected_win_data_423_port, Q(678) => 
                           bus_selected_win_data_422_port, Q(677) => 
                           bus_selected_win_data_421_port, Q(676) => 
                           bus_selected_win_data_420_port, Q(675) => 
                           bus_selected_win_data_419_port, Q(674) => 
                           bus_selected_win_data_418_port, Q(673) => 
                           bus_selected_win_data_417_port, Q(672) => 
                           bus_selected_win_data_416_port, Q(671) => 
                           bus_selected_win_data_415_port, Q(670) => 
                           bus_selected_win_data_414_port, Q(669) => 
                           bus_selected_win_data_413_port, Q(668) => 
                           bus_selected_win_data_412_port, Q(667) => 
                           bus_selected_win_data_411_port, Q(666) => 
                           bus_selected_win_data_410_port, Q(665) => 
                           bus_selected_win_data_409_port, Q(664) => 
                           bus_selected_win_data_408_port, Q(663) => 
                           bus_selected_win_data_407_port, Q(662) => 
                           bus_selected_win_data_406_port, Q(661) => 
                           bus_selected_win_data_405_port, Q(660) => 
                           bus_selected_win_data_404_port, Q(659) => 
                           bus_selected_win_data_403_port, Q(658) => 
                           bus_selected_win_data_402_port, Q(657) => 
                           bus_selected_win_data_401_port, Q(656) => 
                           bus_selected_win_data_400_port, Q(655) => 
                           bus_selected_win_data_399_port, Q(654) => 
                           bus_selected_win_data_398_port, Q(653) => 
                           bus_selected_win_data_397_port, Q(652) => 
                           bus_selected_win_data_396_port, Q(651) => 
                           bus_selected_win_data_395_port, Q(650) => 
                           bus_selected_win_data_394_port, Q(649) => 
                           bus_selected_win_data_393_port, Q(648) => 
                           bus_selected_win_data_392_port, Q(647) => 
                           bus_selected_win_data_391_port, Q(646) => 
                           bus_selected_win_data_390_port, Q(645) => 
                           bus_selected_win_data_389_port, Q(644) => 
                           bus_selected_win_data_388_port, Q(643) => 
                           bus_selected_win_data_387_port, Q(642) => 
                           bus_selected_win_data_386_port, Q(641) => 
                           bus_selected_win_data_385_port, Q(640) => 
                           bus_selected_win_data_384_port, Q(639) => 
                           bus_selected_win_data_383_port, Q(638) => 
                           bus_selected_win_data_382_port, Q(637) => 
                           bus_selected_win_data_381_port, Q(636) => 
                           bus_selected_win_data_380_port, Q(635) => 
                           bus_selected_win_data_379_port, Q(634) => 
                           bus_selected_win_data_378_port, Q(633) => 
                           bus_selected_win_data_377_port, Q(632) => 
                           bus_selected_win_data_376_port, Q(631) => 
                           bus_selected_win_data_375_port, Q(630) => 
                           bus_selected_win_data_374_port, Q(629) => 
                           bus_selected_win_data_373_port, Q(628) => 
                           bus_selected_win_data_372_port, Q(627) => 
                           bus_selected_win_data_371_port, Q(626) => 
                           bus_selected_win_data_370_port, Q(625) => 
                           bus_selected_win_data_369_port, Q(624) => 
                           bus_selected_win_data_368_port, Q(623) => 
                           bus_selected_win_data_367_port, Q(622) => 
                           bus_selected_win_data_366_port, Q(621) => 
                           bus_selected_win_data_365_port, Q(620) => 
                           bus_selected_win_data_364_port, Q(619) => 
                           bus_selected_win_data_363_port, Q(618) => 
                           bus_selected_win_data_362_port, Q(617) => 
                           bus_selected_win_data_361_port, Q(616) => 
                           bus_selected_win_data_360_port, Q(615) => 
                           bus_selected_win_data_359_port, Q(614) => 
                           bus_selected_win_data_358_port, Q(613) => 
                           bus_selected_win_data_357_port, Q(612) => 
                           bus_selected_win_data_356_port, Q(611) => 
                           bus_selected_win_data_355_port, Q(610) => 
                           bus_selected_win_data_354_port, Q(609) => 
                           bus_selected_win_data_353_port, Q(608) => 
                           bus_selected_win_data_352_port, Q(607) => 
                           bus_selected_win_data_351_port, Q(606) => 
                           bus_selected_win_data_350_port, Q(605) => 
                           bus_selected_win_data_349_port, Q(604) => 
                           bus_selected_win_data_348_port, Q(603) => 
                           bus_selected_win_data_347_port, Q(602) => 
                           bus_selected_win_data_346_port, Q(601) => 
                           bus_selected_win_data_345_port, Q(600) => 
                           bus_selected_win_data_344_port, Q(599) => 
                           bus_selected_win_data_343_port, Q(598) => 
                           bus_selected_win_data_342_port, Q(597) => 
                           bus_selected_win_data_341_port, Q(596) => 
                           bus_selected_win_data_340_port, Q(595) => 
                           bus_selected_win_data_339_port, Q(594) => 
                           bus_selected_win_data_338_port, Q(593) => 
                           bus_selected_win_data_337_port, Q(592) => 
                           bus_selected_win_data_336_port, Q(591) => 
                           bus_selected_win_data_335_port, Q(590) => 
                           bus_selected_win_data_334_port, Q(589) => 
                           bus_selected_win_data_333_port, Q(588) => 
                           bus_selected_win_data_332_port, Q(587) => 
                           bus_selected_win_data_331_port, Q(586) => 
                           bus_selected_win_data_330_port, Q(585) => 
                           bus_selected_win_data_329_port, Q(584) => 
                           bus_selected_win_data_328_port, Q(583) => 
                           bus_selected_win_data_327_port, Q(582) => 
                           bus_selected_win_data_326_port, Q(581) => 
                           bus_selected_win_data_325_port, Q(580) => 
                           bus_selected_win_data_324_port, Q(579) => 
                           bus_selected_win_data_323_port, Q(578) => 
                           bus_selected_win_data_322_port, Q(577) => 
                           bus_selected_win_data_321_port, Q(576) => 
                           bus_selected_win_data_320_port, Q(575) => 
                           bus_selected_win_data_319_port, Q(574) => 
                           bus_selected_win_data_318_port, Q(573) => 
                           bus_selected_win_data_317_port, Q(572) => 
                           bus_selected_win_data_316_port, Q(571) => 
                           bus_selected_win_data_315_port, Q(570) => 
                           bus_selected_win_data_314_port, Q(569) => 
                           bus_selected_win_data_313_port, Q(568) => 
                           bus_selected_win_data_312_port, Q(567) => 
                           bus_selected_win_data_311_port, Q(566) => 
                           bus_selected_win_data_310_port, Q(565) => 
                           bus_selected_win_data_309_port, Q(564) => 
                           bus_selected_win_data_308_port, Q(563) => 
                           bus_selected_win_data_307_port, Q(562) => 
                           bus_selected_win_data_306_port, Q(561) => 
                           bus_selected_win_data_305_port, Q(560) => 
                           bus_selected_win_data_304_port, Q(559) => 
                           bus_selected_win_data_303_port, Q(558) => 
                           bus_selected_win_data_302_port, Q(557) => 
                           bus_selected_win_data_301_port, Q(556) => 
                           bus_selected_win_data_300_port, Q(555) => 
                           bus_selected_win_data_299_port, Q(554) => 
                           bus_selected_win_data_298_port, Q(553) => 
                           bus_selected_win_data_297_port, Q(552) => 
                           bus_selected_win_data_296_port, Q(551) => 
                           bus_selected_win_data_295_port, Q(550) => 
                           bus_selected_win_data_294_port, Q(549) => 
                           bus_selected_win_data_293_port, Q(548) => 
                           bus_selected_win_data_292_port, Q(547) => 
                           bus_selected_win_data_291_port, Q(546) => 
                           bus_selected_win_data_290_port, Q(545) => 
                           bus_selected_win_data_289_port, Q(544) => 
                           bus_selected_win_data_288_port, Q(543) => 
                           bus_selected_win_data_287_port, Q(542) => 
                           bus_selected_win_data_286_port, Q(541) => 
                           bus_selected_win_data_285_port, Q(540) => 
                           bus_selected_win_data_284_port, Q(539) => 
                           bus_selected_win_data_283_port, Q(538) => 
                           bus_selected_win_data_282_port, Q(537) => 
                           bus_selected_win_data_281_port, Q(536) => 
                           bus_selected_win_data_280_port, Q(535) => 
                           bus_selected_win_data_279_port, Q(534) => 
                           bus_selected_win_data_278_port, Q(533) => 
                           bus_selected_win_data_277_port, Q(532) => 
                           bus_selected_win_data_276_port, Q(531) => 
                           bus_selected_win_data_275_port, Q(530) => 
                           bus_selected_win_data_274_port, Q(529) => 
                           bus_selected_win_data_273_port, Q(528) => 
                           bus_selected_win_data_272_port, Q(527) => 
                           bus_selected_win_data_271_port, Q(526) => 
                           bus_selected_win_data_270_port, Q(525) => 
                           bus_selected_win_data_269_port, Q(524) => 
                           bus_selected_win_data_268_port, Q(523) => 
                           bus_selected_win_data_267_port, Q(522) => 
                           bus_selected_win_data_266_port, Q(521) => 
                           bus_selected_win_data_265_port, Q(520) => 
                           bus_selected_win_data_264_port, Q(519) => 
                           bus_selected_win_data_263_port, Q(518) => 
                           bus_selected_win_data_262_port, Q(517) => 
                           bus_selected_win_data_261_port, Q(516) => 
                           bus_selected_win_data_260_port, Q(515) => 
                           bus_selected_win_data_259_port, Q(514) => 
                           bus_selected_win_data_258_port, Q(513) => 
                           bus_selected_win_data_257_port, Q(512) => 
                           bus_selected_win_data_256_port, Q(511) => 
                           bus_selected_win_data_255_port, Q(510) => 
                           bus_selected_win_data_254_port, Q(509) => 
                           bus_selected_win_data_253_port, Q(508) => 
                           bus_selected_win_data_252_port, Q(507) => 
                           bus_selected_win_data_251_port, Q(506) => 
                           bus_selected_win_data_250_port, Q(505) => 
                           bus_selected_win_data_249_port, Q(504) => 
                           bus_selected_win_data_248_port, Q(503) => 
                           bus_selected_win_data_247_port, Q(502) => 
                           bus_selected_win_data_246_port, Q(501) => 
                           bus_selected_win_data_245_port, Q(500) => 
                           bus_selected_win_data_244_port, Q(499) => 
                           bus_selected_win_data_243_port, Q(498) => 
                           bus_selected_win_data_242_port, Q(497) => 
                           bus_selected_win_data_241_port, Q(496) => 
                           bus_selected_win_data_240_port, Q(495) => 
                           bus_selected_win_data_239_port, Q(494) => 
                           bus_selected_win_data_238_port, Q(493) => 
                           bus_selected_win_data_237_port, Q(492) => 
                           bus_selected_win_data_236_port, Q(491) => 
                           bus_selected_win_data_235_port, Q(490) => 
                           bus_selected_win_data_234_port, Q(489) => 
                           bus_selected_win_data_233_port, Q(488) => 
                           bus_selected_win_data_232_port, Q(487) => 
                           bus_selected_win_data_231_port, Q(486) => 
                           bus_selected_win_data_230_port, Q(485) => 
                           bus_selected_win_data_229_port, Q(484) => 
                           bus_selected_win_data_228_port, Q(483) => 
                           bus_selected_win_data_227_port, Q(482) => 
                           bus_selected_win_data_226_port, Q(481) => 
                           bus_selected_win_data_225_port, Q(480) => 
                           bus_selected_win_data_224_port, Q(479) => 
                           bus_selected_win_data_223_port, Q(478) => 
                           bus_selected_win_data_222_port, Q(477) => 
                           bus_selected_win_data_221_port, Q(476) => 
                           bus_selected_win_data_220_port, Q(475) => 
                           bus_selected_win_data_219_port, Q(474) => 
                           bus_selected_win_data_218_port, Q(473) => 
                           bus_selected_win_data_217_port, Q(472) => 
                           bus_selected_win_data_216_port, Q(471) => 
                           bus_selected_win_data_215_port, Q(470) => 
                           bus_selected_win_data_214_port, Q(469) => 
                           bus_selected_win_data_213_port, Q(468) => 
                           bus_selected_win_data_212_port, Q(467) => 
                           bus_selected_win_data_211_port, Q(466) => 
                           bus_selected_win_data_210_port, Q(465) => 
                           bus_selected_win_data_209_port, Q(464) => 
                           bus_selected_win_data_208_port, Q(463) => 
                           bus_selected_win_data_207_port, Q(462) => 
                           bus_selected_win_data_206_port, Q(461) => 
                           bus_selected_win_data_205_port, Q(460) => 
                           bus_selected_win_data_204_port, Q(459) => 
                           bus_selected_win_data_203_port, Q(458) => 
                           bus_selected_win_data_202_port, Q(457) => 
                           bus_selected_win_data_201_port, Q(456) => 
                           bus_selected_win_data_200_port, Q(455) => 
                           bus_selected_win_data_199_port, Q(454) => 
                           bus_selected_win_data_198_port, Q(453) => 
                           bus_selected_win_data_197_port, Q(452) => 
                           bus_selected_win_data_196_port, Q(451) => 
                           bus_selected_win_data_195_port, Q(450) => 
                           bus_selected_win_data_194_port, Q(449) => 
                           bus_selected_win_data_193_port, Q(448) => 
                           bus_selected_win_data_192_port, Q(447) => 
                           bus_selected_win_data_191_port, Q(446) => 
                           bus_selected_win_data_190_port, Q(445) => 
                           bus_selected_win_data_189_port, Q(444) => 
                           bus_selected_win_data_188_port, Q(443) => 
                           bus_selected_win_data_187_port, Q(442) => 
                           bus_selected_win_data_186_port, Q(441) => 
                           bus_selected_win_data_185_port, Q(440) => 
                           bus_selected_win_data_184_port, Q(439) => 
                           bus_selected_win_data_183_port, Q(438) => 
                           bus_selected_win_data_182_port, Q(437) => 
                           bus_selected_win_data_181_port, Q(436) => 
                           bus_selected_win_data_180_port, Q(435) => 
                           bus_selected_win_data_179_port, Q(434) => 
                           bus_selected_win_data_178_port, Q(433) => 
                           bus_selected_win_data_177_port, Q(432) => 
                           bus_selected_win_data_176_port, Q(431) => 
                           bus_selected_win_data_175_port, Q(430) => 
                           bus_selected_win_data_174_port, Q(429) => 
                           bus_selected_win_data_173_port, Q(428) => 
                           bus_selected_win_data_172_port, Q(427) => 
                           bus_selected_win_data_171_port, Q(426) => 
                           bus_selected_win_data_170_port, Q(425) => 
                           bus_selected_win_data_169_port, Q(424) => 
                           bus_selected_win_data_168_port, Q(423) => 
                           bus_selected_win_data_167_port, Q(422) => 
                           bus_selected_win_data_166_port, Q(421) => 
                           bus_selected_win_data_165_port, Q(420) => 
                           bus_selected_win_data_164_port, Q(419) => 
                           bus_selected_win_data_163_port, Q(418) => 
                           bus_selected_win_data_162_port, Q(417) => 
                           bus_selected_win_data_161_port, Q(416) => 
                           bus_selected_win_data_160_port, Q(415) => 
                           bus_selected_win_data_159_port, Q(414) => 
                           bus_selected_win_data_158_port, Q(413) => 
                           bus_selected_win_data_157_port, Q(412) => 
                           bus_selected_win_data_156_port, Q(411) => 
                           bus_selected_win_data_155_port, Q(410) => 
                           bus_selected_win_data_154_port, Q(409) => 
                           bus_selected_win_data_153_port, Q(408) => 
                           bus_selected_win_data_152_port, Q(407) => 
                           bus_selected_win_data_151_port, Q(406) => 
                           bus_selected_win_data_150_port, Q(405) => 
                           bus_selected_win_data_149_port, Q(404) => 
                           bus_selected_win_data_148_port, Q(403) => 
                           bus_selected_win_data_147_port, Q(402) => 
                           bus_selected_win_data_146_port, Q(401) => 
                           bus_selected_win_data_145_port, Q(400) => 
                           bus_selected_win_data_144_port, Q(399) => 
                           bus_selected_win_data_143_port, Q(398) => 
                           bus_selected_win_data_142_port, Q(397) => 
                           bus_selected_win_data_141_port, Q(396) => 
                           bus_selected_win_data_140_port, Q(395) => 
                           bus_selected_win_data_139_port, Q(394) => 
                           bus_selected_win_data_138_port, Q(393) => 
                           bus_selected_win_data_137_port, Q(392) => 
                           bus_selected_win_data_136_port, Q(391) => 
                           bus_selected_win_data_135_port, Q(390) => 
                           bus_selected_win_data_134_port, Q(389) => 
                           bus_selected_win_data_133_port, Q(388) => 
                           bus_selected_win_data_132_port, Q(387) => 
                           bus_selected_win_data_131_port, Q(386) => 
                           bus_selected_win_data_130_port, Q(385) => 
                           bus_selected_win_data_129_port, Q(384) => 
                           bus_selected_win_data_128_port, Q(383) => 
                           bus_selected_win_data_127_port, Q(382) => 
                           bus_selected_win_data_126_port, Q(381) => 
                           bus_selected_win_data_125_port, Q(380) => 
                           bus_selected_win_data_124_port, Q(379) => 
                           bus_selected_win_data_123_port, Q(378) => 
                           bus_selected_win_data_122_port, Q(377) => 
                           bus_selected_win_data_121_port, Q(376) => 
                           bus_selected_win_data_120_port, Q(375) => 
                           bus_selected_win_data_119_port, Q(374) => 
                           bus_selected_win_data_118_port, Q(373) => 
                           bus_selected_win_data_117_port, Q(372) => 
                           bus_selected_win_data_116_port, Q(371) => 
                           bus_selected_win_data_115_port, Q(370) => 
                           bus_selected_win_data_114_port, Q(369) => 
                           bus_selected_win_data_113_port, Q(368) => 
                           bus_selected_win_data_112_port, Q(367) => 
                           bus_selected_win_data_111_port, Q(366) => 
                           bus_selected_win_data_110_port, Q(365) => 
                           bus_selected_win_data_109_port, Q(364) => 
                           bus_selected_win_data_108_port, Q(363) => 
                           bus_selected_win_data_107_port, Q(362) => 
                           bus_selected_win_data_106_port, Q(361) => 
                           bus_selected_win_data_105_port, Q(360) => 
                           bus_selected_win_data_104_port, Q(359) => 
                           bus_selected_win_data_103_port, Q(358) => 
                           bus_selected_win_data_102_port, Q(357) => 
                           bus_selected_win_data_101_port, Q(356) => 
                           bus_selected_win_data_100_port, Q(355) => 
                           bus_selected_win_data_99_port, Q(354) => 
                           bus_selected_win_data_98_port, Q(353) => 
                           bus_selected_win_data_97_port, Q(352) => 
                           bus_selected_win_data_96_port, Q(351) => 
                           bus_selected_win_data_95_port, Q(350) => 
                           bus_selected_win_data_94_port, Q(349) => 
                           bus_selected_win_data_93_port, Q(348) => 
                           bus_selected_win_data_92_port, Q(347) => 
                           bus_selected_win_data_91_port, Q(346) => 
                           bus_selected_win_data_90_port, Q(345) => 
                           bus_selected_win_data_89_port, Q(344) => 
                           bus_selected_win_data_88_port, Q(343) => 
                           bus_selected_win_data_87_port, Q(342) => 
                           bus_selected_win_data_86_port, Q(341) => 
                           bus_selected_win_data_85_port, Q(340) => 
                           bus_selected_win_data_84_port, Q(339) => 
                           bus_selected_win_data_83_port, Q(338) => 
                           bus_selected_win_data_82_port, Q(337) => 
                           bus_selected_win_data_81_port, Q(336) => 
                           bus_selected_win_data_80_port, Q(335) => 
                           bus_selected_win_data_79_port, Q(334) => 
                           bus_selected_win_data_78_port, Q(333) => 
                           bus_selected_win_data_77_port, Q(332) => 
                           bus_selected_win_data_76_port, Q(331) => 
                           bus_selected_win_data_75_port, Q(330) => 
                           bus_selected_win_data_74_port, Q(329) => 
                           bus_selected_win_data_73_port, Q(328) => 
                           bus_selected_win_data_72_port, Q(327) => 
                           bus_selected_win_data_71_port, Q(326) => 
                           bus_selected_win_data_70_port, Q(325) => 
                           bus_selected_win_data_69_port, Q(324) => 
                           bus_selected_win_data_68_port, Q(323) => 
                           bus_selected_win_data_67_port, Q(322) => 
                           bus_selected_win_data_66_port, Q(321) => 
                           bus_selected_win_data_65_port, Q(320) => 
                           bus_selected_win_data_64_port, Q(319) => 
                           bus_selected_win_data_63_port, Q(318) => 
                           bus_selected_win_data_62_port, Q(317) => 
                           bus_selected_win_data_61_port, Q(316) => 
                           bus_selected_win_data_60_port, Q(315) => 
                           bus_selected_win_data_59_port, Q(314) => 
                           bus_selected_win_data_58_port, Q(313) => 
                           bus_selected_win_data_57_port, Q(312) => 
                           bus_selected_win_data_56_port, Q(311) => 
                           bus_selected_win_data_55_port, Q(310) => 
                           bus_selected_win_data_54_port, Q(309) => 
                           bus_selected_win_data_53_port, Q(308) => 
                           bus_selected_win_data_52_port, Q(307) => 
                           bus_selected_win_data_51_port, Q(306) => 
                           bus_selected_win_data_50_port, Q(305) => 
                           bus_selected_win_data_49_port, Q(304) => 
                           bus_selected_win_data_48_port, Q(303) => 
                           bus_selected_win_data_47_port, Q(302) => 
                           bus_selected_win_data_46_port, Q(301) => 
                           bus_selected_win_data_45_port, Q(300) => 
                           bus_selected_win_data_44_port, Q(299) => 
                           bus_selected_win_data_43_port, Q(298) => 
                           bus_selected_win_data_42_port, Q(297) => 
                           bus_selected_win_data_41_port, Q(296) => 
                           bus_selected_win_data_40_port, Q(295) => 
                           bus_selected_win_data_39_port, Q(294) => 
                           bus_selected_win_data_38_port, Q(293) => 
                           bus_selected_win_data_37_port, Q(292) => 
                           bus_selected_win_data_36_port, Q(291) => 
                           bus_selected_win_data_35_port, Q(290) => 
                           bus_selected_win_data_34_port, Q(289) => 
                           bus_selected_win_data_33_port, Q(288) => 
                           bus_selected_win_data_32_port, Q(287) => 
                           bus_selected_win_data_31_port, Q(286) => 
                           bus_selected_win_data_30_port, Q(285) => 
                           bus_selected_win_data_29_port, Q(284) => 
                           bus_selected_win_data_28_port, Q(283) => 
                           bus_selected_win_data_27_port, Q(282) => 
                           bus_selected_win_data_26_port, Q(281) => 
                           bus_selected_win_data_25_port, Q(280) => 
                           bus_selected_win_data_24_port, Q(279) => 
                           bus_selected_win_data_23_port, Q(278) => 
                           bus_selected_win_data_22_port, Q(277) => 
                           bus_selected_win_data_21_port, Q(276) => 
                           bus_selected_win_data_20_port, Q(275) => 
                           bus_selected_win_data_19_port, Q(274) => 
                           bus_selected_win_data_18_port, Q(273) => 
                           bus_selected_win_data_17_port, Q(272) => 
                           bus_selected_win_data_16_port, Q(271) => 
                           bus_selected_win_data_15_port, Q(270) => 
                           bus_selected_win_data_14_port, Q(269) => 
                           bus_selected_win_data_13_port, Q(268) => 
                           bus_selected_win_data_12_port, Q(267) => 
                           bus_selected_win_data_11_port, Q(266) => 
                           bus_selected_win_data_10_port, Q(265) => 
                           bus_selected_win_data_9_port, Q(264) => 
                           bus_selected_win_data_8_port, Q(263) => 
                           bus_selected_win_data_7_port, Q(262) => 
                           bus_selected_win_data_6_port, Q(261) => 
                           bus_selected_win_data_5_port, Q(260) => 
                           bus_selected_win_data_4_port, Q(259) => 
                           bus_selected_win_data_3_port, Q(258) => 
                           bus_selected_win_data_2_port, Q(257) => 
                           bus_selected_win_data_1_port, Q(256) => 
                           bus_selected_win_data_0_port, Q(255) => 
                           bus_complete_win_data_255_port, Q(254) => 
                           bus_complete_win_data_254_port, Q(253) => 
                           bus_complete_win_data_253_port, Q(252) => 
                           bus_complete_win_data_252_port, Q(251) => 
                           bus_complete_win_data_251_port, Q(250) => 
                           bus_complete_win_data_250_port, Q(249) => 
                           bus_complete_win_data_249_port, Q(248) => 
                           bus_complete_win_data_248_port, Q(247) => 
                           bus_complete_win_data_247_port, Q(246) => 
                           bus_complete_win_data_246_port, Q(245) => 
                           bus_complete_win_data_245_port, Q(244) => 
                           bus_complete_win_data_244_port, Q(243) => 
                           bus_complete_win_data_243_port, Q(242) => 
                           bus_complete_win_data_242_port, Q(241) => 
                           bus_complete_win_data_241_port, Q(240) => 
                           bus_complete_win_data_240_port, Q(239) => 
                           bus_complete_win_data_239_port, Q(238) => 
                           bus_complete_win_data_238_port, Q(237) => 
                           bus_complete_win_data_237_port, Q(236) => 
                           bus_complete_win_data_236_port, Q(235) => 
                           bus_complete_win_data_235_port, Q(234) => 
                           bus_complete_win_data_234_port, Q(233) => 
                           bus_complete_win_data_233_port, Q(232) => 
                           bus_complete_win_data_232_port, Q(231) => 
                           bus_complete_win_data_231_port, Q(230) => 
                           bus_complete_win_data_230_port, Q(229) => 
                           bus_complete_win_data_229_port, Q(228) => 
                           bus_complete_win_data_228_port, Q(227) => 
                           bus_complete_win_data_227_port, Q(226) => 
                           bus_complete_win_data_226_port, Q(225) => 
                           bus_complete_win_data_225_port, Q(224) => 
                           bus_complete_win_data_224_port, Q(223) => 
                           bus_complete_win_data_223_port, Q(222) => 
                           bus_complete_win_data_222_port, Q(221) => 
                           bus_complete_win_data_221_port, Q(220) => 
                           bus_complete_win_data_220_port, Q(219) => 
                           bus_complete_win_data_219_port, Q(218) => 
                           bus_complete_win_data_218_port, Q(217) => 
                           bus_complete_win_data_217_port, Q(216) => 
                           bus_complete_win_data_216_port, Q(215) => 
                           bus_complete_win_data_215_port, Q(214) => 
                           bus_complete_win_data_214_port, Q(213) => 
                           bus_complete_win_data_213_port, Q(212) => 
                           bus_complete_win_data_212_port, Q(211) => 
                           bus_complete_win_data_211_port, Q(210) => 
                           bus_complete_win_data_210_port, Q(209) => 
                           bus_complete_win_data_209_port, Q(208) => 
                           bus_complete_win_data_208_port, Q(207) => 
                           bus_complete_win_data_207_port, Q(206) => 
                           bus_complete_win_data_206_port, Q(205) => 
                           bus_complete_win_data_205_port, Q(204) => 
                           bus_complete_win_data_204_port, Q(203) => 
                           bus_complete_win_data_203_port, Q(202) => 
                           bus_complete_win_data_202_port, Q(201) => 
                           bus_complete_win_data_201_port, Q(200) => 
                           bus_complete_win_data_200_port, Q(199) => 
                           bus_complete_win_data_199_port, Q(198) => 
                           bus_complete_win_data_198_port, Q(197) => 
                           bus_complete_win_data_197_port, Q(196) => 
                           bus_complete_win_data_196_port, Q(195) => 
                           bus_complete_win_data_195_port, Q(194) => 
                           bus_complete_win_data_194_port, Q(193) => 
                           bus_complete_win_data_193_port, Q(192) => 
                           bus_complete_win_data_192_port, Q(191) => 
                           bus_complete_win_data_191_port, Q(190) => 
                           bus_complete_win_data_190_port, Q(189) => 
                           bus_complete_win_data_189_port, Q(188) => 
                           bus_complete_win_data_188_port, Q(187) => 
                           bus_complete_win_data_187_port, Q(186) => 
                           bus_complete_win_data_186_port, Q(185) => 
                           bus_complete_win_data_185_port, Q(184) => 
                           bus_complete_win_data_184_port, Q(183) => 
                           bus_complete_win_data_183_port, Q(182) => 
                           bus_complete_win_data_182_port, Q(181) => 
                           bus_complete_win_data_181_port, Q(180) => 
                           bus_complete_win_data_180_port, Q(179) => 
                           bus_complete_win_data_179_port, Q(178) => 
                           bus_complete_win_data_178_port, Q(177) => 
                           bus_complete_win_data_177_port, Q(176) => 
                           bus_complete_win_data_176_port, Q(175) => 
                           bus_complete_win_data_175_port, Q(174) => 
                           bus_complete_win_data_174_port, Q(173) => 
                           bus_complete_win_data_173_port, Q(172) => 
                           bus_complete_win_data_172_port, Q(171) => 
                           bus_complete_win_data_171_port, Q(170) => 
                           bus_complete_win_data_170_port, Q(169) => 
                           bus_complete_win_data_169_port, Q(168) => 
                           bus_complete_win_data_168_port, Q(167) => 
                           bus_complete_win_data_167_port, Q(166) => 
                           bus_complete_win_data_166_port, Q(165) => 
                           bus_complete_win_data_165_port, Q(164) => 
                           bus_complete_win_data_164_port, Q(163) => 
                           bus_complete_win_data_163_port, Q(162) => 
                           bus_complete_win_data_162_port, Q(161) => 
                           bus_complete_win_data_161_port, Q(160) => 
                           bus_complete_win_data_160_port, Q(159) => 
                           bus_complete_win_data_159_port, Q(158) => 
                           bus_complete_win_data_158_port, Q(157) => 
                           bus_complete_win_data_157_port, Q(156) => 
                           bus_complete_win_data_156_port, Q(155) => 
                           bus_complete_win_data_155_port, Q(154) => 
                           bus_complete_win_data_154_port, Q(153) => 
                           bus_complete_win_data_153_port, Q(152) => 
                           bus_complete_win_data_152_port, Q(151) => 
                           bus_complete_win_data_151_port, Q(150) => 
                           bus_complete_win_data_150_port, Q(149) => 
                           bus_complete_win_data_149_port, Q(148) => 
                           bus_complete_win_data_148_port, Q(147) => 
                           bus_complete_win_data_147_port, Q(146) => 
                           bus_complete_win_data_146_port, Q(145) => 
                           bus_complete_win_data_145_port, Q(144) => 
                           bus_complete_win_data_144_port, Q(143) => 
                           bus_complete_win_data_143_port, Q(142) => 
                           bus_complete_win_data_142_port, Q(141) => 
                           bus_complete_win_data_141_port, Q(140) => 
                           bus_complete_win_data_140_port, Q(139) => 
                           bus_complete_win_data_139_port, Q(138) => 
                           bus_complete_win_data_138_port, Q(137) => 
                           bus_complete_win_data_137_port, Q(136) => 
                           bus_complete_win_data_136_port, Q(135) => 
                           bus_complete_win_data_135_port, Q(134) => 
                           bus_complete_win_data_134_port, Q(133) => 
                           bus_complete_win_data_133_port, Q(132) => 
                           bus_complete_win_data_132_port, Q(131) => 
                           bus_complete_win_data_131_port, Q(130) => 
                           bus_complete_win_data_130_port, Q(129) => 
                           bus_complete_win_data_129_port, Q(128) => 
                           bus_complete_win_data_128_port, Q(127) => 
                           bus_complete_win_data_127_port, Q(126) => 
                           bus_complete_win_data_126_port, Q(125) => 
                           bus_complete_win_data_125_port, Q(124) => 
                           bus_complete_win_data_124_port, Q(123) => 
                           bus_complete_win_data_123_port, Q(122) => 
                           bus_complete_win_data_122_port, Q(121) => 
                           bus_complete_win_data_121_port, Q(120) => 
                           bus_complete_win_data_120_port, Q(119) => 
                           bus_complete_win_data_119_port, Q(118) => 
                           bus_complete_win_data_118_port, Q(117) => 
                           bus_complete_win_data_117_port, Q(116) => 
                           bus_complete_win_data_116_port, Q(115) => 
                           bus_complete_win_data_115_port, Q(114) => 
                           bus_complete_win_data_114_port, Q(113) => 
                           bus_complete_win_data_113_port, Q(112) => 
                           bus_complete_win_data_112_port, Q(111) => 
                           bus_complete_win_data_111_port, Q(110) => 
                           bus_complete_win_data_110_port, Q(109) => 
                           bus_complete_win_data_109_port, Q(108) => 
                           bus_complete_win_data_108_port, Q(107) => 
                           bus_complete_win_data_107_port, Q(106) => 
                           bus_complete_win_data_106_port, Q(105) => 
                           bus_complete_win_data_105_port, Q(104) => 
                           bus_complete_win_data_104_port, Q(103) => 
                           bus_complete_win_data_103_port, Q(102) => 
                           bus_complete_win_data_102_port, Q(101) => 
                           bus_complete_win_data_101_port, Q(100) => 
                           bus_complete_win_data_100_port, Q(99) => 
                           bus_complete_win_data_99_port, Q(98) => 
                           bus_complete_win_data_98_port, Q(97) => 
                           bus_complete_win_data_97_port, Q(96) => 
                           bus_complete_win_data_96_port, Q(95) => 
                           bus_complete_win_data_95_port, Q(94) => 
                           bus_complete_win_data_94_port, Q(93) => 
                           bus_complete_win_data_93_port, Q(92) => 
                           bus_complete_win_data_92_port, Q(91) => 
                           bus_complete_win_data_91_port, Q(90) => 
                           bus_complete_win_data_90_port, Q(89) => 
                           bus_complete_win_data_89_port, Q(88) => 
                           bus_complete_win_data_88_port, Q(87) => 
                           bus_complete_win_data_87_port, Q(86) => 
                           bus_complete_win_data_86_port, Q(85) => 
                           bus_complete_win_data_85_port, Q(84) => 
                           bus_complete_win_data_84_port, Q(83) => 
                           bus_complete_win_data_83_port, Q(82) => 
                           bus_complete_win_data_82_port, Q(81) => 
                           bus_complete_win_data_81_port, Q(80) => 
                           bus_complete_win_data_80_port, Q(79) => 
                           bus_complete_win_data_79_port, Q(78) => 
                           bus_complete_win_data_78_port, Q(77) => 
                           bus_complete_win_data_77_port, Q(76) => 
                           bus_complete_win_data_76_port, Q(75) => 
                           bus_complete_win_data_75_port, Q(74) => 
                           bus_complete_win_data_74_port, Q(73) => 
                           bus_complete_win_data_73_port, Q(72) => 
                           bus_complete_win_data_72_port, Q(71) => 
                           bus_complete_win_data_71_port, Q(70) => 
                           bus_complete_win_data_70_port, Q(69) => 
                           bus_complete_win_data_69_port, Q(68) => 
                           bus_complete_win_data_68_port, Q(67) => 
                           bus_complete_win_data_67_port, Q(66) => 
                           bus_complete_win_data_66_port, Q(65) => 
                           bus_complete_win_data_65_port, Q(64) => 
                           bus_complete_win_data_64_port, Q(63) => 
                           bus_complete_win_data_63_port, Q(62) => 
                           bus_complete_win_data_62_port, Q(61) => 
                           bus_complete_win_data_61_port, Q(60) => 
                           bus_complete_win_data_60_port, Q(59) => 
                           bus_complete_win_data_59_port, Q(58) => 
                           bus_complete_win_data_58_port, Q(57) => 
                           bus_complete_win_data_57_port, Q(56) => 
                           bus_complete_win_data_56_port, Q(55) => 
                           bus_complete_win_data_55_port, Q(54) => 
                           bus_complete_win_data_54_port, Q(53) => 
                           bus_complete_win_data_53_port, Q(52) => 
                           bus_complete_win_data_52_port, Q(51) => 
                           bus_complete_win_data_51_port, Q(50) => 
                           bus_complete_win_data_50_port, Q(49) => 
                           bus_complete_win_data_49_port, Q(48) => 
                           bus_complete_win_data_48_port, Q(47) => 
                           bus_complete_win_data_47_port, Q(46) => 
                           bus_complete_win_data_46_port, Q(45) => 
                           bus_complete_win_data_45_port, Q(44) => 
                           bus_complete_win_data_44_port, Q(43) => 
                           bus_complete_win_data_43_port, Q(42) => 
                           bus_complete_win_data_42_port, Q(41) => 
                           bus_complete_win_data_41_port, Q(40) => 
                           bus_complete_win_data_40_port, Q(39) => 
                           bus_complete_win_data_39_port, Q(38) => 
                           bus_complete_win_data_38_port, Q(37) => 
                           bus_complete_win_data_37_port, Q(36) => 
                           bus_complete_win_data_36_port, Q(35) => 
                           bus_complete_win_data_35_port, Q(34) => 
                           bus_complete_win_data_34_port, Q(33) => 
                           bus_complete_win_data_33_port, Q(32) => 
                           bus_complete_win_data_32_port, Q(31) => 
                           bus_complete_win_data_31_port, Q(30) => 
                           bus_complete_win_data_30_port, Q(29) => 
                           bus_complete_win_data_29_port, Q(28) => 
                           bus_complete_win_data_28_port, Q(27) => 
                           bus_complete_win_data_27_port, Q(26) => 
                           bus_complete_win_data_26_port, Q(25) => 
                           bus_complete_win_data_25_port, Q(24) => 
                           bus_complete_win_data_24_port, Q(23) => 
                           bus_complete_win_data_23_port, Q(22) => 
                           bus_complete_win_data_22_port, Q(21) => 
                           bus_complete_win_data_21_port, Q(20) => 
                           bus_complete_win_data_20_port, Q(19) => 
                           bus_complete_win_data_19_port, Q(18) => 
                           bus_complete_win_data_18_port, Q(17) => 
                           bus_complete_win_data_17_port, Q(16) => 
                           bus_complete_win_data_16_port, Q(15) => 
                           bus_complete_win_data_15_port, Q(14) => 
                           bus_complete_win_data_14_port, Q(13) => 
                           bus_complete_win_data_13_port, Q(12) => 
                           bus_complete_win_data_12_port, Q(11) => 
                           bus_complete_win_data_11_port, Q(10) => 
                           bus_complete_win_data_10_port, Q(9) => 
                           bus_complete_win_data_9_port, Q(8) => 
                           bus_complete_win_data_8_port, Q(7) => 
                           bus_complete_win_data_7_port, Q(6) => 
                           bus_complete_win_data_6_port, Q(5) => 
                           bus_complete_win_data_5_port, Q(4) => 
                           bus_complete_win_data_4_port, Q(3) => 
                           bus_complete_win_data_3_port, Q(2) => 
                           bus_complete_win_data_2_port, Q(1) => 
                           bus_complete_win_data_1_port, Q(0) => 
                           bus_complete_win_data_0_port, Y(31) => 
                           internal_out2_31_port, Y(30) => 
                           internal_out2_30_port, Y(29) => 
                           internal_out2_29_port, Y(28) => 
                           internal_out2_28_port, Y(27) => 
                           internal_out2_27_port, Y(26) => 
                           internal_out2_26_port, Y(25) => 
                           internal_out2_25_port, Y(24) => 
                           internal_out2_24_port, Y(23) => 
                           internal_out2_23_port, Y(22) => 
                           internal_out2_22_port, Y(21) => 
                           internal_out2_21_port, Y(20) => 
                           internal_out2_20_port, Y(19) => 
                           internal_out2_19_port, Y(18) => 
                           internal_out2_18_port, Y(17) => 
                           internal_out2_17_port, Y(16) => 
                           internal_out2_16_port, Y(15) => 
                           internal_out2_15_port, Y(14) => 
                           internal_out2_14_port, Y(13) => 
                           internal_out2_13_port, Y(12) => 
                           internal_out2_12_port, Y(11) => 
                           internal_out2_11_port, Y(10) => 
                           internal_out2_10_port, Y(9) => internal_out2_9_port,
                           Y(8) => internal_out2_8_port, Y(7) => 
                           internal_out2_7_port, Y(6) => internal_out2_6_port, 
                           Y(5) => internal_out2_5_port, Y(4) => 
                           internal_out2_4_port, Y(3) => internal_out2_3_port, 
                           Y(2) => internal_out2_2_port, Y(1) => 
                           internal_out2_1_port, Y(0) => internal_out2_0_port);
   RDPORT1_OUTREG : reg_generic_N32_RSTVAL0_89 port map( D(31) => 
                           internal_out2_31_port, D(30) => 
                           internal_out2_30_port, D(29) => 
                           internal_out2_29_port, D(28) => 
                           internal_out2_28_port, D(27) => 
                           internal_out2_27_port, D(26) => 
                           internal_out2_26_port, D(25) => 
                           internal_out2_25_port, D(24) => 
                           internal_out2_24_port, D(23) => 
                           internal_out2_23_port, D(22) => 
                           internal_out2_22_port, D(21) => 
                           internal_out2_21_port, D(20) => 
                           internal_out2_20_port, D(19) => 
                           internal_out2_19_port, D(18) => 
                           internal_out2_18_port, D(17) => 
                           internal_out2_17_port, D(16) => 
                           internal_out2_16_port, D(15) => 
                           internal_out2_15_port, D(14) => 
                           internal_out2_14_port, D(13) => 
                           internal_out2_13_port, D(12) => 
                           internal_out2_12_port, D(11) => 
                           internal_out2_11_port, D(10) => 
                           internal_out2_10_port, D(9) => internal_out2_9_port,
                           D(8) => internal_out2_8_port, D(7) => 
                           internal_out2_7_port, D(6) => internal_out2_6_port, 
                           D(5) => internal_out2_5_port, D(4) => 
                           internal_out2_4_port, D(3) => internal_out2_3_port, 
                           D(2) => internal_out2_2_port, D(1) => 
                           internal_out2_1_port, D(0) => internal_out2_0_port, 
                           Q(31) => OUT2(31), Q(30) => OUT2(30), Q(29) => 
                           OUT2(29), Q(28) => OUT2(28), Q(27) => OUT2(27), 
                           Q(26) => OUT2(26), Q(25) => OUT2(25), Q(24) => 
                           OUT2(24), Q(23) => OUT2(23), Q(22) => OUT2(22), 
                           Q(21) => OUT2(21), Q(20) => OUT2(20), Q(19) => 
                           OUT2(19), Q(18) => OUT2(18), Q(17) => OUT2(17), 
                           Q(16) => OUT2(16), Q(15) => OUT2(15), Q(14) => 
                           OUT2(14), Q(13) => OUT2(13), Q(12) => OUT2(12), 
                           Q(11) => OUT2(11), Q(10) => OUT2(10), Q(9) => 
                           OUT2(9), Q(8) => OUT2(8), Q(7) => OUT2(7), Q(6) => 
                           OUT2(6), Q(5) => OUT2(5), Q(4) => OUT2(4), Q(3) => 
                           OUT2(3), Q(2) => OUT2(2), Q(1) => OUT2(1), Q(0) => 
                           OUT2(0), Clk => CLK, Rst => RESET, Enable => int_RD2
                           );
   BLOCK_GLOB_0 : reg_generic_N32_RSTVAL0_88 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_31_port, Q(30) => 
                           bus_complete_win_data_30_port, Q(29) => 
                           bus_complete_win_data_29_port, Q(28) => 
                           bus_complete_win_data_28_port, Q(27) => 
                           bus_complete_win_data_27_port, Q(26) => 
                           bus_complete_win_data_26_port, Q(25) => 
                           bus_complete_win_data_25_port, Q(24) => 
                           bus_complete_win_data_24_port, Q(23) => 
                           bus_complete_win_data_23_port, Q(22) => 
                           bus_complete_win_data_22_port, Q(21) => 
                           bus_complete_win_data_21_port, Q(20) => 
                           bus_complete_win_data_20_port, Q(19) => 
                           bus_complete_win_data_19_port, Q(18) => 
                           bus_complete_win_data_18_port, Q(17) => 
                           bus_complete_win_data_17_port, Q(16) => 
                           bus_complete_win_data_16_port, Q(15) => 
                           bus_complete_win_data_15_port, Q(14) => 
                           bus_complete_win_data_14_port, Q(13) => 
                           bus_complete_win_data_13_port, Q(12) => 
                           bus_complete_win_data_12_port, Q(11) => 
                           bus_complete_win_data_11_port, Q(10) => 
                           bus_complete_win_data_10_port, Q(9) => 
                           bus_complete_win_data_9_port, Q(8) => 
                           bus_complete_win_data_8_port, Q(7) => 
                           bus_complete_win_data_7_port, Q(6) => 
                           bus_complete_win_data_6_port, Q(5) => 
                           bus_complete_win_data_5_port, Q(4) => 
                           bus_complete_win_data_4_port, Q(3) => 
                           bus_complete_win_data_3_port, Q(2) => 
                           bus_complete_win_data_2_port, Q(1) => 
                           bus_complete_win_data_1_port, Q(0) => 
                           bus_complete_win_data_0_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_0_port);
   BLOCK_GLOB_1 : reg_generic_N32_RSTVAL0_87 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_63_port, Q(30) => 
                           bus_complete_win_data_62_port, Q(29) => 
                           bus_complete_win_data_61_port, Q(28) => 
                           bus_complete_win_data_60_port, Q(27) => 
                           bus_complete_win_data_59_port, Q(26) => 
                           bus_complete_win_data_58_port, Q(25) => 
                           bus_complete_win_data_57_port, Q(24) => 
                           bus_complete_win_data_56_port, Q(23) => 
                           bus_complete_win_data_55_port, Q(22) => 
                           bus_complete_win_data_54_port, Q(21) => 
                           bus_complete_win_data_53_port, Q(20) => 
                           bus_complete_win_data_52_port, Q(19) => 
                           bus_complete_win_data_51_port, Q(18) => 
                           bus_complete_win_data_50_port, Q(17) => 
                           bus_complete_win_data_49_port, Q(16) => 
                           bus_complete_win_data_48_port, Q(15) => 
                           bus_complete_win_data_47_port, Q(14) => 
                           bus_complete_win_data_46_port, Q(13) => 
                           bus_complete_win_data_45_port, Q(12) => 
                           bus_complete_win_data_44_port, Q(11) => 
                           bus_complete_win_data_43_port, Q(10) => 
                           bus_complete_win_data_42_port, Q(9) => 
                           bus_complete_win_data_41_port, Q(8) => 
                           bus_complete_win_data_40_port, Q(7) => 
                           bus_complete_win_data_39_port, Q(6) => 
                           bus_complete_win_data_38_port, Q(5) => 
                           bus_complete_win_data_37_port, Q(4) => 
                           bus_complete_win_data_36_port, Q(3) => 
                           bus_complete_win_data_35_port, Q(2) => 
                           bus_complete_win_data_34_port, Q(1) => 
                           bus_complete_win_data_33_port, Q(0) => 
                           bus_complete_win_data_32_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_1_port);
   BLOCK_GLOB_2 : reg_generic_N32_RSTVAL0_86 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_95_port, Q(30) => 
                           bus_complete_win_data_94_port, Q(29) => 
                           bus_complete_win_data_93_port, Q(28) => 
                           bus_complete_win_data_92_port, Q(27) => 
                           bus_complete_win_data_91_port, Q(26) => 
                           bus_complete_win_data_90_port, Q(25) => 
                           bus_complete_win_data_89_port, Q(24) => 
                           bus_complete_win_data_88_port, Q(23) => 
                           bus_complete_win_data_87_port, Q(22) => 
                           bus_complete_win_data_86_port, Q(21) => 
                           bus_complete_win_data_85_port, Q(20) => 
                           bus_complete_win_data_84_port, Q(19) => 
                           bus_complete_win_data_83_port, Q(18) => 
                           bus_complete_win_data_82_port, Q(17) => 
                           bus_complete_win_data_81_port, Q(16) => 
                           bus_complete_win_data_80_port, Q(15) => 
                           bus_complete_win_data_79_port, Q(14) => 
                           bus_complete_win_data_78_port, Q(13) => 
                           bus_complete_win_data_77_port, Q(12) => 
                           bus_complete_win_data_76_port, Q(11) => 
                           bus_complete_win_data_75_port, Q(10) => 
                           bus_complete_win_data_74_port, Q(9) => 
                           bus_complete_win_data_73_port, Q(8) => 
                           bus_complete_win_data_72_port, Q(7) => 
                           bus_complete_win_data_71_port, Q(6) => 
                           bus_complete_win_data_70_port, Q(5) => 
                           bus_complete_win_data_69_port, Q(4) => 
                           bus_complete_win_data_68_port, Q(3) => 
                           bus_complete_win_data_67_port, Q(2) => 
                           bus_complete_win_data_66_port, Q(1) => 
                           bus_complete_win_data_65_port, Q(0) => 
                           bus_complete_win_data_64_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_2_port);
   BLOCK_GLOB_3 : reg_generic_N32_RSTVAL0_85 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_127_port, Q(30) => 
                           bus_complete_win_data_126_port, Q(29) => 
                           bus_complete_win_data_125_port, Q(28) => 
                           bus_complete_win_data_124_port, Q(27) => 
                           bus_complete_win_data_123_port, Q(26) => 
                           bus_complete_win_data_122_port, Q(25) => 
                           bus_complete_win_data_121_port, Q(24) => 
                           bus_complete_win_data_120_port, Q(23) => 
                           bus_complete_win_data_119_port, Q(22) => 
                           bus_complete_win_data_118_port, Q(21) => 
                           bus_complete_win_data_117_port, Q(20) => 
                           bus_complete_win_data_116_port, Q(19) => 
                           bus_complete_win_data_115_port, Q(18) => 
                           bus_complete_win_data_114_port, Q(17) => 
                           bus_complete_win_data_113_port, Q(16) => 
                           bus_complete_win_data_112_port, Q(15) => 
                           bus_complete_win_data_111_port, Q(14) => 
                           bus_complete_win_data_110_port, Q(13) => 
                           bus_complete_win_data_109_port, Q(12) => 
                           bus_complete_win_data_108_port, Q(11) => 
                           bus_complete_win_data_107_port, Q(10) => 
                           bus_complete_win_data_106_port, Q(9) => 
                           bus_complete_win_data_105_port, Q(8) => 
                           bus_complete_win_data_104_port, Q(7) => 
                           bus_complete_win_data_103_port, Q(6) => 
                           bus_complete_win_data_102_port, Q(5) => 
                           bus_complete_win_data_101_port, Q(4) => 
                           bus_complete_win_data_100_port, Q(3) => 
                           bus_complete_win_data_99_port, Q(2) => 
                           bus_complete_win_data_98_port, Q(1) => 
                           bus_complete_win_data_97_port, Q(0) => 
                           bus_complete_win_data_96_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_3_port);
   BLOCK_GLOB_4 : reg_generic_N32_RSTVAL0_84 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_159_port, Q(30) => 
                           bus_complete_win_data_158_port, Q(29) => 
                           bus_complete_win_data_157_port, Q(28) => 
                           bus_complete_win_data_156_port, Q(27) => 
                           bus_complete_win_data_155_port, Q(26) => 
                           bus_complete_win_data_154_port, Q(25) => 
                           bus_complete_win_data_153_port, Q(24) => 
                           bus_complete_win_data_152_port, Q(23) => 
                           bus_complete_win_data_151_port, Q(22) => 
                           bus_complete_win_data_150_port, Q(21) => 
                           bus_complete_win_data_149_port, Q(20) => 
                           bus_complete_win_data_148_port, Q(19) => 
                           bus_complete_win_data_147_port, Q(18) => 
                           bus_complete_win_data_146_port, Q(17) => 
                           bus_complete_win_data_145_port, Q(16) => 
                           bus_complete_win_data_144_port, Q(15) => 
                           bus_complete_win_data_143_port, Q(14) => 
                           bus_complete_win_data_142_port, Q(13) => 
                           bus_complete_win_data_141_port, Q(12) => 
                           bus_complete_win_data_140_port, Q(11) => 
                           bus_complete_win_data_139_port, Q(10) => 
                           bus_complete_win_data_138_port, Q(9) => 
                           bus_complete_win_data_137_port, Q(8) => 
                           bus_complete_win_data_136_port, Q(7) => 
                           bus_complete_win_data_135_port, Q(6) => 
                           bus_complete_win_data_134_port, Q(5) => 
                           bus_complete_win_data_133_port, Q(4) => 
                           bus_complete_win_data_132_port, Q(3) => 
                           bus_complete_win_data_131_port, Q(2) => 
                           bus_complete_win_data_130_port, Q(1) => 
                           bus_complete_win_data_129_port, Q(0) => 
                           bus_complete_win_data_128_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_4_port);
   BLOCK_GLOB_5 : reg_generic_N32_RSTVAL0_83 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_191_port, Q(30) => 
                           bus_complete_win_data_190_port, Q(29) => 
                           bus_complete_win_data_189_port, Q(28) => 
                           bus_complete_win_data_188_port, Q(27) => 
                           bus_complete_win_data_187_port, Q(26) => 
                           bus_complete_win_data_186_port, Q(25) => 
                           bus_complete_win_data_185_port, Q(24) => 
                           bus_complete_win_data_184_port, Q(23) => 
                           bus_complete_win_data_183_port, Q(22) => 
                           bus_complete_win_data_182_port, Q(21) => 
                           bus_complete_win_data_181_port, Q(20) => 
                           bus_complete_win_data_180_port, Q(19) => 
                           bus_complete_win_data_179_port, Q(18) => 
                           bus_complete_win_data_178_port, Q(17) => 
                           bus_complete_win_data_177_port, Q(16) => 
                           bus_complete_win_data_176_port, Q(15) => 
                           bus_complete_win_data_175_port, Q(14) => 
                           bus_complete_win_data_174_port, Q(13) => 
                           bus_complete_win_data_173_port, Q(12) => 
                           bus_complete_win_data_172_port, Q(11) => 
                           bus_complete_win_data_171_port, Q(10) => 
                           bus_complete_win_data_170_port, Q(9) => 
                           bus_complete_win_data_169_port, Q(8) => 
                           bus_complete_win_data_168_port, Q(7) => 
                           bus_complete_win_data_167_port, Q(6) => 
                           bus_complete_win_data_166_port, Q(5) => 
                           bus_complete_win_data_165_port, Q(4) => 
                           bus_complete_win_data_164_port, Q(3) => 
                           bus_complete_win_data_163_port, Q(2) => 
                           bus_complete_win_data_162_port, Q(1) => 
                           bus_complete_win_data_161_port, Q(0) => 
                           bus_complete_win_data_160_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_5_port);
   BLOCK_GLOB_6 : reg_generic_N32_RSTVAL0_82 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_223_port, Q(30) => 
                           bus_complete_win_data_222_port, Q(29) => 
                           bus_complete_win_data_221_port, Q(28) => 
                           bus_complete_win_data_220_port, Q(27) => 
                           bus_complete_win_data_219_port, Q(26) => 
                           bus_complete_win_data_218_port, Q(25) => 
                           bus_complete_win_data_217_port, Q(24) => 
                           bus_complete_win_data_216_port, Q(23) => 
                           bus_complete_win_data_215_port, Q(22) => 
                           bus_complete_win_data_214_port, Q(21) => 
                           bus_complete_win_data_213_port, Q(20) => 
                           bus_complete_win_data_212_port, Q(19) => 
                           bus_complete_win_data_211_port, Q(18) => 
                           bus_complete_win_data_210_port, Q(17) => 
                           bus_complete_win_data_209_port, Q(16) => 
                           bus_complete_win_data_208_port, Q(15) => 
                           bus_complete_win_data_207_port, Q(14) => 
                           bus_complete_win_data_206_port, Q(13) => 
                           bus_complete_win_data_205_port, Q(12) => 
                           bus_complete_win_data_204_port, Q(11) => 
                           bus_complete_win_data_203_port, Q(10) => 
                           bus_complete_win_data_202_port, Q(9) => 
                           bus_complete_win_data_201_port, Q(8) => 
                           bus_complete_win_data_200_port, Q(7) => 
                           bus_complete_win_data_199_port, Q(6) => 
                           bus_complete_win_data_198_port, Q(5) => 
                           bus_complete_win_data_197_port, Q(4) => 
                           bus_complete_win_data_196_port, Q(3) => 
                           bus_complete_win_data_195_port, Q(2) => 
                           bus_complete_win_data_194_port, Q(1) => 
                           bus_complete_win_data_193_port, Q(0) => 
                           bus_complete_win_data_192_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_6_port);
   BLOCK_GLOB_7 : reg_generic_N32_RSTVAL0_81 port map( D(31) => DATAIN(31), 
                           D(30) => DATAIN(30), D(29) => DATAIN(29), D(28) => 
                           DATAIN(28), D(27) => DATAIN(27), D(26) => DATAIN(26)
                           , D(25) => DATAIN(25), D(24) => DATAIN(24), D(23) =>
                           DATAIN(23), D(22) => DATAIN(22), D(21) => DATAIN(21)
                           , D(20) => DATAIN(20), D(19) => DATAIN(19), D(18) =>
                           DATAIN(18), D(17) => DATAIN(17), D(16) => DATAIN(16)
                           , D(15) => DATAIN(15), D(14) => DATAIN(14), D(13) =>
                           DATAIN(13), D(12) => DATAIN(12), D(11) => DATAIN(11)
                           , D(10) => DATAIN(10), D(9) => DATAIN(9), D(8) => 
                           DATAIN(8), D(7) => DATAIN(7), D(6) => DATAIN(6), 
                           D(5) => DATAIN(5), D(4) => DATAIN(4), D(3) => 
                           DATAIN(3), D(2) => DATAIN(2), D(1) => DATAIN(1), 
                           D(0) => DATAIN(0), Q(31) => 
                           bus_complete_win_data_255_port, Q(30) => 
                           bus_complete_win_data_254_port, Q(29) => 
                           bus_complete_win_data_253_port, Q(28) => 
                           bus_complete_win_data_252_port, Q(27) => 
                           bus_complete_win_data_251_port, Q(26) => 
                           bus_complete_win_data_250_port, Q(25) => 
                           bus_complete_win_data_249_port, Q(24) => 
                           bus_complete_win_data_248_port, Q(23) => 
                           bus_complete_win_data_247_port, Q(22) => 
                           bus_complete_win_data_246_port, Q(21) => 
                           bus_complete_win_data_245_port, Q(20) => 
                           bus_complete_win_data_244_port, Q(19) => 
                           bus_complete_win_data_243_port, Q(18) => 
                           bus_complete_win_data_242_port, Q(17) => 
                           bus_complete_win_data_241_port, Q(16) => 
                           bus_complete_win_data_240_port, Q(15) => 
                           bus_complete_win_data_239_port, Q(14) => 
                           bus_complete_win_data_238_port, Q(13) => 
                           bus_complete_win_data_237_port, Q(12) => 
                           bus_complete_win_data_236_port, Q(11) => 
                           bus_complete_win_data_235_port, Q(10) => 
                           bus_complete_win_data_234_port, Q(9) => 
                           bus_complete_win_data_233_port, Q(8) => 
                           bus_complete_win_data_232_port, Q(7) => 
                           bus_complete_win_data_231_port, Q(6) => 
                           bus_complete_win_data_230_port, Q(5) => 
                           bus_complete_win_data_229_port, Q(4) => 
                           bus_complete_win_data_228_port, Q(3) => 
                           bus_complete_win_data_227_port, Q(2) => 
                           bus_complete_win_data_226_port, Q(1) => 
                           bus_complete_win_data_225_port, Q(0) => 
                           bus_complete_win_data_224_port, Clk => CLK, Rst => 
                           RESET, Enable => en_regi_7_port);
   MUX_SELINPUT_8 : mux_N32_M1_0 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1615
                           , Y(30) => n1607, Y(29) => n1599, Y(28) => n1591, 
                           Y(27) => n1583, Y(26) => n1575, Y(25) => n1567, 
                           Y(24) => n1559, Y(23) => n1551, Y(22) => n1543, 
                           Y(21) => n1535, Y(20) => n1527, Y(19) => n1519, 
                           Y(18) => n1511, Y(17) => n1503, Y(16) => n1495, 
                           Y(15) => n1487, Y(14) => n1479, Y(13) => n1471, 
                           Y(12) => n1463, Y(11) => n1455, Y(10) => n1447, Y(9)
                           => n1439, Y(8) => n1431, Y(7) => n1423, Y(6) => 
                           n1415, Y(5) => n1407, Y(4) => n1399, Y(3) => n1391, 
                           Y(2) => n1383, Y(1) => n1375, Y(0) => n1367);
   BLOCKi_8 : reg_generic_N32_RSTVAL0_80 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_31_port, Q(30) => 
                           bus_reg_dataout_30_port, Q(29) => 
                           bus_reg_dataout_29_port, Q(28) => 
                           bus_reg_dataout_28_port, Q(27) => 
                           bus_reg_dataout_27_port, Q(26) => 
                           bus_reg_dataout_26_port, Q(25) => 
                           bus_reg_dataout_25_port, Q(24) => 
                           bus_reg_dataout_24_port, Q(23) => 
                           bus_reg_dataout_23_port, Q(22) => 
                           bus_reg_dataout_22_port, Q(21) => 
                           bus_reg_dataout_21_port, Q(20) => 
                           bus_reg_dataout_20_port, Q(19) => 
                           bus_reg_dataout_19_port, Q(18) => 
                           bus_reg_dataout_18_port, Q(17) => 
                           bus_reg_dataout_17_port, Q(16) => 
                           bus_reg_dataout_16_port, Q(15) => 
                           bus_reg_dataout_15_port, Q(14) => 
                           bus_reg_dataout_14_port, Q(13) => 
                           bus_reg_dataout_13_port, Q(12) => 
                           bus_reg_dataout_12_port, Q(11) => 
                           bus_reg_dataout_11_port, Q(10) => 
                           bus_reg_dataout_10_port, Q(9) => 
                           bus_reg_dataout_9_port, Q(8) => 
                           bus_reg_dataout_8_port, Q(7) => 
                           bus_reg_dataout_7_port, Q(6) => 
                           bus_reg_dataout_6_port, Q(5) => 
                           bus_reg_dataout_5_port, Q(4) => 
                           bus_reg_dataout_4_port, Q(3) => 
                           bus_reg_dataout_3_port, Q(2) => 
                           bus_reg_dataout_2_port, Q(1) => 
                           bus_reg_dataout_1_port, Q(0) => 
                           bus_reg_dataout_0_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_8_port);
   BLOCKi_9 : reg_generic_N32_RSTVAL0_79 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_63_port, Q(30) => 
                           bus_reg_dataout_62_port, Q(29) => 
                           bus_reg_dataout_61_port, Q(28) => 
                           bus_reg_dataout_60_port, Q(27) => 
                           bus_reg_dataout_59_port, Q(26) => 
                           bus_reg_dataout_58_port, Q(25) => 
                           bus_reg_dataout_57_port, Q(24) => 
                           bus_reg_dataout_56_port, Q(23) => 
                           bus_reg_dataout_55_port, Q(22) => 
                           bus_reg_dataout_54_port, Q(21) => 
                           bus_reg_dataout_53_port, Q(20) => 
                           bus_reg_dataout_52_port, Q(19) => 
                           bus_reg_dataout_51_port, Q(18) => 
                           bus_reg_dataout_50_port, Q(17) => 
                           bus_reg_dataout_49_port, Q(16) => 
                           bus_reg_dataout_48_port, Q(15) => 
                           bus_reg_dataout_47_port, Q(14) => 
                           bus_reg_dataout_46_port, Q(13) => 
                           bus_reg_dataout_45_port, Q(12) => 
                           bus_reg_dataout_44_port, Q(11) => 
                           bus_reg_dataout_43_port, Q(10) => 
                           bus_reg_dataout_42_port, Q(9) => 
                           bus_reg_dataout_41_port, Q(8) => 
                           bus_reg_dataout_40_port, Q(7) => 
                           bus_reg_dataout_39_port, Q(6) => 
                           bus_reg_dataout_38_port, Q(5) => 
                           bus_reg_dataout_37_port, Q(4) => 
                           bus_reg_dataout_36_port, Q(3) => 
                           bus_reg_dataout_35_port, Q(2) => 
                           bus_reg_dataout_34_port, Q(1) => 
                           bus_reg_dataout_33_port, Q(0) => 
                           bus_reg_dataout_32_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_9_port);
   MUX_SELINPUT_10 : mux_N32_M1_39 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1622
                           , Y(30) => n1614, Y(29) => n1606, Y(28) => n1598, 
                           Y(27) => n1590, Y(26) => n1582, Y(25) => n1574, 
                           Y(24) => n1566, Y(23) => n1558, Y(22) => n1550, 
                           Y(21) => n1542, Y(20) => n1534, Y(19) => n1526, 
                           Y(18) => n1518, Y(17) => n1510, Y(16) => n1502, 
                           Y(15) => n1494, Y(14) => n1486, Y(13) => n1478, 
                           Y(12) => n1470, Y(11) => n1462, Y(10) => n1454, Y(9)
                           => n1446, Y(8) => n1438, Y(7) => n1430, Y(6) => 
                           n1422, Y(5) => n1414, Y(4) => n1406, Y(3) => n1398, 
                           Y(2) => n1390, Y(1) => n1382, Y(0) => n1374);
   BLOCKi_10 : reg_generic_N32_RSTVAL0_78 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_95_port, Q(30) => 
                           bus_reg_dataout_94_port, Q(29) => 
                           bus_reg_dataout_93_port, Q(28) => 
                           bus_reg_dataout_92_port, Q(27) => 
                           bus_reg_dataout_91_port, Q(26) => 
                           bus_reg_dataout_90_port, Q(25) => 
                           bus_reg_dataout_89_port, Q(24) => 
                           bus_reg_dataout_88_port, Q(23) => 
                           bus_reg_dataout_87_port, Q(22) => 
                           bus_reg_dataout_86_port, Q(21) => 
                           bus_reg_dataout_85_port, Q(20) => 
                           bus_reg_dataout_84_port, Q(19) => 
                           bus_reg_dataout_83_port, Q(18) => 
                           bus_reg_dataout_82_port, Q(17) => 
                           bus_reg_dataout_81_port, Q(16) => 
                           bus_reg_dataout_80_port, Q(15) => 
                           bus_reg_dataout_79_port, Q(14) => 
                           bus_reg_dataout_78_port, Q(13) => 
                           bus_reg_dataout_77_port, Q(12) => 
                           bus_reg_dataout_76_port, Q(11) => 
                           bus_reg_dataout_75_port, Q(10) => 
                           bus_reg_dataout_74_port, Q(9) => 
                           bus_reg_dataout_73_port, Q(8) => 
                           bus_reg_dataout_72_port, Q(7) => 
                           bus_reg_dataout_71_port, Q(6) => 
                           bus_reg_dataout_70_port, Q(5) => 
                           bus_reg_dataout_69_port, Q(4) => 
                           bus_reg_dataout_68_port, Q(3) => 
                           bus_reg_dataout_67_port, Q(2) => 
                           bus_reg_dataout_66_port, Q(1) => 
                           bus_reg_dataout_65_port, Q(0) => 
                           bus_reg_dataout_64_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_10_port);
   BLOCKi_11 : reg_generic_N32_RSTVAL0_77 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_127_port, Q(30) => 
                           bus_reg_dataout_126_port, Q(29) => 
                           bus_reg_dataout_125_port, Q(28) => 
                           bus_reg_dataout_124_port, Q(27) => 
                           bus_reg_dataout_123_port, Q(26) => 
                           bus_reg_dataout_122_port, Q(25) => 
                           bus_reg_dataout_121_port, Q(24) => 
                           bus_reg_dataout_120_port, Q(23) => 
                           bus_reg_dataout_119_port, Q(22) => 
                           bus_reg_dataout_118_port, Q(21) => 
                           bus_reg_dataout_117_port, Q(20) => 
                           bus_reg_dataout_116_port, Q(19) => 
                           bus_reg_dataout_115_port, Q(18) => 
                           bus_reg_dataout_114_port, Q(17) => 
                           bus_reg_dataout_113_port, Q(16) => 
                           bus_reg_dataout_112_port, Q(15) => 
                           bus_reg_dataout_111_port, Q(14) => 
                           bus_reg_dataout_110_port, Q(13) => 
                           bus_reg_dataout_109_port, Q(12) => 
                           bus_reg_dataout_108_port, Q(11) => 
                           bus_reg_dataout_107_port, Q(10) => 
                           bus_reg_dataout_106_port, Q(9) => 
                           bus_reg_dataout_105_port, Q(8) => 
                           bus_reg_dataout_104_port, Q(7) => 
                           bus_reg_dataout_103_port, Q(6) => 
                           bus_reg_dataout_102_port, Q(5) => 
                           bus_reg_dataout_101_port, Q(4) => 
                           bus_reg_dataout_100_port, Q(3) => 
                           bus_reg_dataout_99_port, Q(2) => 
                           bus_reg_dataout_98_port, Q(1) => 
                           bus_reg_dataout_97_port, Q(0) => 
                           bus_reg_dataout_96_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_11_port);
   MUX_SELINPUT_12 : mux_N32_M1_38 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1621
                           , Y(30) => n1613, Y(29) => n1605, Y(28) => n1597, 
                           Y(27) => n1589, Y(26) => n1581, Y(25) => n1573, 
                           Y(24) => n1565, Y(23) => n1557, Y(22) => n1549, 
                           Y(21) => n1541, Y(20) => n1533, Y(19) => n1525, 
                           Y(18) => n1517, Y(17) => n1509, Y(16) => n1501, 
                           Y(15) => n1493, Y(14) => n1485, Y(13) => n1477, 
                           Y(12) => n1469, Y(11) => n1461, Y(10) => n1453, Y(9)
                           => n1445, Y(8) => n1437, Y(7) => n1429, Y(6) => 
                           n1421, Y(5) => n1413, Y(4) => n1405, Y(3) => n1397, 
                           Y(2) => n1389, Y(1) => n1381, Y(0) => n1373);
   BLOCKi_12 : reg_generic_N32_RSTVAL0_76 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_159_port, Q(30) => 
                           bus_reg_dataout_158_port, Q(29) => 
                           bus_reg_dataout_157_port, Q(28) => 
                           bus_reg_dataout_156_port, Q(27) => 
                           bus_reg_dataout_155_port, Q(26) => 
                           bus_reg_dataout_154_port, Q(25) => 
                           bus_reg_dataout_153_port, Q(24) => 
                           bus_reg_dataout_152_port, Q(23) => 
                           bus_reg_dataout_151_port, Q(22) => 
                           bus_reg_dataout_150_port, Q(21) => 
                           bus_reg_dataout_149_port, Q(20) => 
                           bus_reg_dataout_148_port, Q(19) => 
                           bus_reg_dataout_147_port, Q(18) => 
                           bus_reg_dataout_146_port, Q(17) => 
                           bus_reg_dataout_145_port, Q(16) => 
                           bus_reg_dataout_144_port, Q(15) => 
                           bus_reg_dataout_143_port, Q(14) => 
                           bus_reg_dataout_142_port, Q(13) => 
                           bus_reg_dataout_141_port, Q(12) => 
                           bus_reg_dataout_140_port, Q(11) => 
                           bus_reg_dataout_139_port, Q(10) => 
                           bus_reg_dataout_138_port, Q(9) => 
                           bus_reg_dataout_137_port, Q(8) => 
                           bus_reg_dataout_136_port, Q(7) => 
                           bus_reg_dataout_135_port, Q(6) => 
                           bus_reg_dataout_134_port, Q(5) => 
                           bus_reg_dataout_133_port, Q(4) => 
                           bus_reg_dataout_132_port, Q(3) => 
                           bus_reg_dataout_131_port, Q(2) => 
                           bus_reg_dataout_130_port, Q(1) => 
                           bus_reg_dataout_129_port, Q(0) => 
                           bus_reg_dataout_128_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_12_port);
   BLOCKi_13 : reg_generic_N32_RSTVAL0_75 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_191_port, Q(30) => 
                           bus_reg_dataout_190_port, Q(29) => 
                           bus_reg_dataout_189_port, Q(28) => 
                           bus_reg_dataout_188_port, Q(27) => 
                           bus_reg_dataout_187_port, Q(26) => 
                           bus_reg_dataout_186_port, Q(25) => 
                           bus_reg_dataout_185_port, Q(24) => 
                           bus_reg_dataout_184_port, Q(23) => 
                           bus_reg_dataout_183_port, Q(22) => 
                           bus_reg_dataout_182_port, Q(21) => 
                           bus_reg_dataout_181_port, Q(20) => 
                           bus_reg_dataout_180_port, Q(19) => 
                           bus_reg_dataout_179_port, Q(18) => 
                           bus_reg_dataout_178_port, Q(17) => 
                           bus_reg_dataout_177_port, Q(16) => 
                           bus_reg_dataout_176_port, Q(15) => 
                           bus_reg_dataout_175_port, Q(14) => 
                           bus_reg_dataout_174_port, Q(13) => 
                           bus_reg_dataout_173_port, Q(12) => 
                           bus_reg_dataout_172_port, Q(11) => 
                           bus_reg_dataout_171_port, Q(10) => 
                           bus_reg_dataout_170_port, Q(9) => 
                           bus_reg_dataout_169_port, Q(8) => 
                           bus_reg_dataout_168_port, Q(7) => 
                           bus_reg_dataout_167_port, Q(6) => 
                           bus_reg_dataout_166_port, Q(5) => 
                           bus_reg_dataout_165_port, Q(4) => 
                           bus_reg_dataout_164_port, Q(3) => 
                           bus_reg_dataout_163_port, Q(2) => 
                           bus_reg_dataout_162_port, Q(1) => 
                           bus_reg_dataout_161_port, Q(0) => 
                           bus_reg_dataout_160_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_13_port);
   MUX_SELINPUT_14 : mux_N32_M1_37 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1620
                           , Y(30) => n1612, Y(29) => n1604, Y(28) => n1596, 
                           Y(27) => n1588, Y(26) => n1580, Y(25) => n1572, 
                           Y(24) => n1564, Y(23) => n1556, Y(22) => n1548, 
                           Y(21) => n1540, Y(20) => n1532, Y(19) => n1524, 
                           Y(18) => n1516, Y(17) => n1508, Y(16) => n1500, 
                           Y(15) => n1492, Y(14) => n1484, Y(13) => n1476, 
                           Y(12) => n1468, Y(11) => n1460, Y(10) => n1452, Y(9)
                           => n1444, Y(8) => n1436, Y(7) => n1428, Y(6) => 
                           n1420, Y(5) => n1412, Y(4) => n1404, Y(3) => n1396, 
                           Y(2) => n1388, Y(1) => n1380, Y(0) => n1372);
   BLOCKi_14 : reg_generic_N32_RSTVAL0_74 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_223_port, Q(30) => 
                           bus_reg_dataout_222_port, Q(29) => 
                           bus_reg_dataout_221_port, Q(28) => 
                           bus_reg_dataout_220_port, Q(27) => 
                           bus_reg_dataout_219_port, Q(26) => 
                           bus_reg_dataout_218_port, Q(25) => 
                           bus_reg_dataout_217_port, Q(24) => 
                           bus_reg_dataout_216_port, Q(23) => 
                           bus_reg_dataout_215_port, Q(22) => 
                           bus_reg_dataout_214_port, Q(21) => 
                           bus_reg_dataout_213_port, Q(20) => 
                           bus_reg_dataout_212_port, Q(19) => 
                           bus_reg_dataout_211_port, Q(18) => 
                           bus_reg_dataout_210_port, Q(17) => 
                           bus_reg_dataout_209_port, Q(16) => 
                           bus_reg_dataout_208_port, Q(15) => 
                           bus_reg_dataout_207_port, Q(14) => 
                           bus_reg_dataout_206_port, Q(13) => 
                           bus_reg_dataout_205_port, Q(12) => 
                           bus_reg_dataout_204_port, Q(11) => 
                           bus_reg_dataout_203_port, Q(10) => 
                           bus_reg_dataout_202_port, Q(9) => 
                           bus_reg_dataout_201_port, Q(8) => 
                           bus_reg_dataout_200_port, Q(7) => 
                           bus_reg_dataout_199_port, Q(6) => 
                           bus_reg_dataout_198_port, Q(5) => 
                           bus_reg_dataout_197_port, Q(4) => 
                           bus_reg_dataout_196_port, Q(3) => 
                           bus_reg_dataout_195_port, Q(2) => 
                           bus_reg_dataout_194_port, Q(1) => 
                           bus_reg_dataout_193_port, Q(0) => 
                           bus_reg_dataout_192_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_14_port);
   BLOCKi_15 : reg_generic_N32_RSTVAL0_73 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_255_port, Q(30) => 
                           bus_reg_dataout_254_port, Q(29) => 
                           bus_reg_dataout_253_port, Q(28) => 
                           bus_reg_dataout_252_port, Q(27) => 
                           bus_reg_dataout_251_port, Q(26) => 
                           bus_reg_dataout_250_port, Q(25) => 
                           bus_reg_dataout_249_port, Q(24) => 
                           bus_reg_dataout_248_port, Q(23) => 
                           bus_reg_dataout_247_port, Q(22) => 
                           bus_reg_dataout_246_port, Q(21) => 
                           bus_reg_dataout_245_port, Q(20) => 
                           bus_reg_dataout_244_port, Q(19) => 
                           bus_reg_dataout_243_port, Q(18) => 
                           bus_reg_dataout_242_port, Q(17) => 
                           bus_reg_dataout_241_port, Q(16) => 
                           bus_reg_dataout_240_port, Q(15) => 
                           bus_reg_dataout_239_port, Q(14) => 
                           bus_reg_dataout_238_port, Q(13) => 
                           bus_reg_dataout_237_port, Q(12) => 
                           bus_reg_dataout_236_port, Q(11) => 
                           bus_reg_dataout_235_port, Q(10) => 
                           bus_reg_dataout_234_port, Q(9) => 
                           bus_reg_dataout_233_port, Q(8) => 
                           bus_reg_dataout_232_port, Q(7) => 
                           bus_reg_dataout_231_port, Q(6) => 
                           bus_reg_dataout_230_port, Q(5) => 
                           bus_reg_dataout_229_port, Q(4) => 
                           bus_reg_dataout_228_port, Q(3) => 
                           bus_reg_dataout_227_port, Q(2) => 
                           bus_reg_dataout_226_port, Q(1) => 
                           bus_reg_dataout_225_port, Q(0) => 
                           bus_reg_dataout_224_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_15_port);
   MUX_SELINPUT_16 : mux_N32_M1_36 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1619
                           , Y(30) => n1611, Y(29) => n1603, Y(28) => n1595, 
                           Y(27) => n1587, Y(26) => n1579, Y(25) => n1571, 
                           Y(24) => n1563, Y(23) => n1555, Y(22) => n1547, 
                           Y(21) => n1539, Y(20) => n1531, Y(19) => n1523, 
                           Y(18) => n1515, Y(17) => n1507, Y(16) => n1499, 
                           Y(15) => n1491, Y(14) => n1483, Y(13) => n1475, 
                           Y(12) => n1467, Y(11) => n1459, Y(10) => n1451, Y(9)
                           => n1443, Y(8) => n1435, Y(7) => n1427, Y(6) => 
                           n1419, Y(5) => n1411, Y(4) => n1403, Y(3) => n1395, 
                           Y(2) => n1387, Y(1) => n1379, Y(0) => n1371);
   BLOCKi_16 : reg_generic_N32_RSTVAL0_72 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_287_port, Q(30) => 
                           bus_reg_dataout_286_port, Q(29) => 
                           bus_reg_dataout_285_port, Q(28) => 
                           bus_reg_dataout_284_port, Q(27) => 
                           bus_reg_dataout_283_port, Q(26) => 
                           bus_reg_dataout_282_port, Q(25) => 
                           bus_reg_dataout_281_port, Q(24) => 
                           bus_reg_dataout_280_port, Q(23) => 
                           bus_reg_dataout_279_port, Q(22) => 
                           bus_reg_dataout_278_port, Q(21) => 
                           bus_reg_dataout_277_port, Q(20) => 
                           bus_reg_dataout_276_port, Q(19) => 
                           bus_reg_dataout_275_port, Q(18) => 
                           bus_reg_dataout_274_port, Q(17) => 
                           bus_reg_dataout_273_port, Q(16) => 
                           bus_reg_dataout_272_port, Q(15) => 
                           bus_reg_dataout_271_port, Q(14) => 
                           bus_reg_dataout_270_port, Q(13) => 
                           bus_reg_dataout_269_port, Q(12) => 
                           bus_reg_dataout_268_port, Q(11) => 
                           bus_reg_dataout_267_port, Q(10) => 
                           bus_reg_dataout_266_port, Q(9) => 
                           bus_reg_dataout_265_port, Q(8) => 
                           bus_reg_dataout_264_port, Q(7) => 
                           bus_reg_dataout_263_port, Q(6) => 
                           bus_reg_dataout_262_port, Q(5) => 
                           bus_reg_dataout_261_port, Q(4) => 
                           bus_reg_dataout_260_port, Q(3) => 
                           bus_reg_dataout_259_port, Q(2) => 
                           bus_reg_dataout_258_port, Q(1) => 
                           bus_reg_dataout_257_port, Q(0) => 
                           bus_reg_dataout_256_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_16_port);
   BLOCKi_17 : reg_generic_N32_RSTVAL0_71 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_319_port, Q(30) => 
                           bus_reg_dataout_318_port, Q(29) => 
                           bus_reg_dataout_317_port, Q(28) => 
                           bus_reg_dataout_316_port, Q(27) => 
                           bus_reg_dataout_315_port, Q(26) => 
                           bus_reg_dataout_314_port, Q(25) => 
                           bus_reg_dataout_313_port, Q(24) => 
                           bus_reg_dataout_312_port, Q(23) => 
                           bus_reg_dataout_311_port, Q(22) => 
                           bus_reg_dataout_310_port, Q(21) => 
                           bus_reg_dataout_309_port, Q(20) => 
                           bus_reg_dataout_308_port, Q(19) => 
                           bus_reg_dataout_307_port, Q(18) => 
                           bus_reg_dataout_306_port, Q(17) => 
                           bus_reg_dataout_305_port, Q(16) => 
                           bus_reg_dataout_304_port, Q(15) => 
                           bus_reg_dataout_303_port, Q(14) => 
                           bus_reg_dataout_302_port, Q(13) => 
                           bus_reg_dataout_301_port, Q(12) => 
                           bus_reg_dataout_300_port, Q(11) => 
                           bus_reg_dataout_299_port, Q(10) => 
                           bus_reg_dataout_298_port, Q(9) => 
                           bus_reg_dataout_297_port, Q(8) => 
                           bus_reg_dataout_296_port, Q(7) => 
                           bus_reg_dataout_295_port, Q(6) => 
                           bus_reg_dataout_294_port, Q(5) => 
                           bus_reg_dataout_293_port, Q(4) => 
                           bus_reg_dataout_292_port, Q(3) => 
                           bus_reg_dataout_291_port, Q(2) => 
                           bus_reg_dataout_290_port, Q(1) => 
                           bus_reg_dataout_289_port, Q(0) => 
                           bus_reg_dataout_288_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_17_port);
   MUX_SELINPUT_18 : mux_N32_M1_35 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1618
                           , Y(30) => n1610, Y(29) => n1602, Y(28) => n1594, 
                           Y(27) => n1586, Y(26) => n1578, Y(25) => n1570, 
                           Y(24) => n1562, Y(23) => n1554, Y(22) => n1546, 
                           Y(21) => n1538, Y(20) => n1530, Y(19) => n1522, 
                           Y(18) => n1514, Y(17) => n1506, Y(16) => n1498, 
                           Y(15) => n1490, Y(14) => n1482, Y(13) => n1474, 
                           Y(12) => n1466, Y(11) => n1458, Y(10) => n1450, Y(9)
                           => n1442, Y(8) => n1434, Y(7) => n1426, Y(6) => 
                           n1418, Y(5) => n1410, Y(4) => n1402, Y(3) => n1394, 
                           Y(2) => n1386, Y(1) => n1378, Y(0) => n1370);
   BLOCKi_18 : reg_generic_N32_RSTVAL0_70 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_351_port, Q(30) => 
                           bus_reg_dataout_350_port, Q(29) => 
                           bus_reg_dataout_349_port, Q(28) => 
                           bus_reg_dataout_348_port, Q(27) => 
                           bus_reg_dataout_347_port, Q(26) => 
                           bus_reg_dataout_346_port, Q(25) => 
                           bus_reg_dataout_345_port, Q(24) => 
                           bus_reg_dataout_344_port, Q(23) => 
                           bus_reg_dataout_343_port, Q(22) => 
                           bus_reg_dataout_342_port, Q(21) => 
                           bus_reg_dataout_341_port, Q(20) => 
                           bus_reg_dataout_340_port, Q(19) => 
                           bus_reg_dataout_339_port, Q(18) => 
                           bus_reg_dataout_338_port, Q(17) => 
                           bus_reg_dataout_337_port, Q(16) => 
                           bus_reg_dataout_336_port, Q(15) => 
                           bus_reg_dataout_335_port, Q(14) => 
                           bus_reg_dataout_334_port, Q(13) => 
                           bus_reg_dataout_333_port, Q(12) => 
                           bus_reg_dataout_332_port, Q(11) => 
                           bus_reg_dataout_331_port, Q(10) => 
                           bus_reg_dataout_330_port, Q(9) => 
                           bus_reg_dataout_329_port, Q(8) => 
                           bus_reg_dataout_328_port, Q(7) => 
                           bus_reg_dataout_327_port, Q(6) => 
                           bus_reg_dataout_326_port, Q(5) => 
                           bus_reg_dataout_325_port, Q(4) => 
                           bus_reg_dataout_324_port, Q(3) => 
                           bus_reg_dataout_323_port, Q(2) => 
                           bus_reg_dataout_322_port, Q(1) => 
                           bus_reg_dataout_321_port, Q(0) => 
                           bus_reg_dataout_320_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_18_port);
   BLOCKi_19 : reg_generic_N32_RSTVAL0_69 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_383_port, Q(30) => 
                           bus_reg_dataout_382_port, Q(29) => 
                           bus_reg_dataout_381_port, Q(28) => 
                           bus_reg_dataout_380_port, Q(27) => 
                           bus_reg_dataout_379_port, Q(26) => 
                           bus_reg_dataout_378_port, Q(25) => 
                           bus_reg_dataout_377_port, Q(24) => 
                           bus_reg_dataout_376_port, Q(23) => 
                           bus_reg_dataout_375_port, Q(22) => 
                           bus_reg_dataout_374_port, Q(21) => 
                           bus_reg_dataout_373_port, Q(20) => 
                           bus_reg_dataout_372_port, Q(19) => 
                           bus_reg_dataout_371_port, Q(18) => 
                           bus_reg_dataout_370_port, Q(17) => 
                           bus_reg_dataout_369_port, Q(16) => 
                           bus_reg_dataout_368_port, Q(15) => 
                           bus_reg_dataout_367_port, Q(14) => 
                           bus_reg_dataout_366_port, Q(13) => 
                           bus_reg_dataout_365_port, Q(12) => 
                           bus_reg_dataout_364_port, Q(11) => 
                           bus_reg_dataout_363_port, Q(10) => 
                           bus_reg_dataout_362_port, Q(9) => 
                           bus_reg_dataout_361_port, Q(8) => 
                           bus_reg_dataout_360_port, Q(7) => 
                           bus_reg_dataout_359_port, Q(6) => 
                           bus_reg_dataout_358_port, Q(5) => 
                           bus_reg_dataout_357_port, Q(4) => 
                           bus_reg_dataout_356_port, Q(3) => 
                           bus_reg_dataout_355_port, Q(2) => 
                           bus_reg_dataout_354_port, Q(1) => 
                           bus_reg_dataout_353_port, Q(0) => 
                           bus_reg_dataout_352_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_19_port);
   MUX_SELINPUT_20 : mux_N32_M1_34 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1617
                           , Y(30) => n1609, Y(29) => n1601, Y(28) => n1593, 
                           Y(27) => n1585, Y(26) => n1577, Y(25) => n1569, 
                           Y(24) => n1561, Y(23) => n1553, Y(22) => n1545, 
                           Y(21) => n1537, Y(20) => n1529, Y(19) => n1521, 
                           Y(18) => n1513, Y(17) => n1505, Y(16) => n1497, 
                           Y(15) => n1489, Y(14) => n1481, Y(13) => n1473, 
                           Y(12) => n1465, Y(11) => n1457, Y(10) => n1449, Y(9)
                           => n1441, Y(8) => n1433, Y(7) => n1425, Y(6) => 
                           n1417, Y(5) => n1409, Y(4) => n1401, Y(3) => n1393, 
                           Y(2) => n1385, Y(1) => n1377, Y(0) => n1369);
   BLOCKi_20 : reg_generic_N32_RSTVAL0_68 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_415_port, Q(30) => 
                           bus_reg_dataout_414_port, Q(29) => 
                           bus_reg_dataout_413_port, Q(28) => 
                           bus_reg_dataout_412_port, Q(27) => 
                           bus_reg_dataout_411_port, Q(26) => 
                           bus_reg_dataout_410_port, Q(25) => 
                           bus_reg_dataout_409_port, Q(24) => 
                           bus_reg_dataout_408_port, Q(23) => 
                           bus_reg_dataout_407_port, Q(22) => 
                           bus_reg_dataout_406_port, Q(21) => 
                           bus_reg_dataout_405_port, Q(20) => 
                           bus_reg_dataout_404_port, Q(19) => 
                           bus_reg_dataout_403_port, Q(18) => 
                           bus_reg_dataout_402_port, Q(17) => 
                           bus_reg_dataout_401_port, Q(16) => 
                           bus_reg_dataout_400_port, Q(15) => 
                           bus_reg_dataout_399_port, Q(14) => 
                           bus_reg_dataout_398_port, Q(13) => 
                           bus_reg_dataout_397_port, Q(12) => 
                           bus_reg_dataout_396_port, Q(11) => 
                           bus_reg_dataout_395_port, Q(10) => 
                           bus_reg_dataout_394_port, Q(9) => 
                           bus_reg_dataout_393_port, Q(8) => 
                           bus_reg_dataout_392_port, Q(7) => 
                           bus_reg_dataout_391_port, Q(6) => 
                           bus_reg_dataout_390_port, Q(5) => 
                           bus_reg_dataout_389_port, Q(4) => 
                           bus_reg_dataout_388_port, Q(3) => 
                           bus_reg_dataout_387_port, Q(2) => 
                           bus_reg_dataout_386_port, Q(1) => 
                           bus_reg_dataout_385_port, Q(0) => 
                           bus_reg_dataout_384_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_20_port);
   BLOCKi_21 : reg_generic_N32_RSTVAL0_67 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_447_port, Q(30) => 
                           bus_reg_dataout_446_port, Q(29) => 
                           bus_reg_dataout_445_port, Q(28) => 
                           bus_reg_dataout_444_port, Q(27) => 
                           bus_reg_dataout_443_port, Q(26) => 
                           bus_reg_dataout_442_port, Q(25) => 
                           bus_reg_dataout_441_port, Q(24) => 
                           bus_reg_dataout_440_port, Q(23) => 
                           bus_reg_dataout_439_port, Q(22) => 
                           bus_reg_dataout_438_port, Q(21) => 
                           bus_reg_dataout_437_port, Q(20) => 
                           bus_reg_dataout_436_port, Q(19) => 
                           bus_reg_dataout_435_port, Q(18) => 
                           bus_reg_dataout_434_port, Q(17) => 
                           bus_reg_dataout_433_port, Q(16) => 
                           bus_reg_dataout_432_port, Q(15) => 
                           bus_reg_dataout_431_port, Q(14) => 
                           bus_reg_dataout_430_port, Q(13) => 
                           bus_reg_dataout_429_port, Q(12) => 
                           bus_reg_dataout_428_port, Q(11) => 
                           bus_reg_dataout_427_port, Q(10) => 
                           bus_reg_dataout_426_port, Q(9) => 
                           bus_reg_dataout_425_port, Q(8) => 
                           bus_reg_dataout_424_port, Q(7) => 
                           bus_reg_dataout_423_port, Q(6) => 
                           bus_reg_dataout_422_port, Q(5) => 
                           bus_reg_dataout_421_port, Q(4) => 
                           bus_reg_dataout_420_port, Q(3) => 
                           bus_reg_dataout_419_port, Q(2) => 
                           bus_reg_dataout_418_port, Q(1) => 
                           bus_reg_dataout_417_port, Q(0) => 
                           bus_reg_dataout_416_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_21_port);
   MUX_SELINPUT_22 : mux_N32_M1_33 port map( S => c_swin_masked_1bit_0_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1616
                           , Y(30) => n1608, Y(29) => n1600, Y(28) => n1592, 
                           Y(27) => n1584, Y(26) => n1576, Y(25) => n1568, 
                           Y(24) => n1560, Y(23) => n1552, Y(22) => n1544, 
                           Y(21) => n1536, Y(20) => n1528, Y(19) => n1520, 
                           Y(18) => n1512, Y(17) => n1504, Y(16) => n1496, 
                           Y(15) => n1488, Y(14) => n1480, Y(13) => n1472, 
                           Y(12) => n1464, Y(11) => n1456, Y(10) => n1448, Y(9)
                           => n1440, Y(8) => n1432, Y(7) => n1424, Y(6) => 
                           n1416, Y(5) => n1408, Y(4) => n1400, Y(3) => n1392, 
                           Y(2) => n1384, Y(1) => n1376, Y(0) => n1368);
   BLOCKi_22 : reg_generic_N32_RSTVAL0_66 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_479_port, Q(30) => 
                           bus_reg_dataout_478_port, Q(29) => 
                           bus_reg_dataout_477_port, Q(28) => 
                           bus_reg_dataout_476_port, Q(27) => 
                           bus_reg_dataout_475_port, Q(26) => 
                           bus_reg_dataout_474_port, Q(25) => 
                           bus_reg_dataout_473_port, Q(24) => 
                           bus_reg_dataout_472_port, Q(23) => 
                           bus_reg_dataout_471_port, Q(22) => 
                           bus_reg_dataout_470_port, Q(21) => 
                           bus_reg_dataout_469_port, Q(20) => 
                           bus_reg_dataout_468_port, Q(19) => 
                           bus_reg_dataout_467_port, Q(18) => 
                           bus_reg_dataout_466_port, Q(17) => 
                           bus_reg_dataout_465_port, Q(16) => 
                           bus_reg_dataout_464_port, Q(15) => 
                           bus_reg_dataout_463_port, Q(14) => 
                           bus_reg_dataout_462_port, Q(13) => 
                           bus_reg_dataout_461_port, Q(12) => 
                           bus_reg_dataout_460_port, Q(11) => 
                           bus_reg_dataout_459_port, Q(10) => 
                           bus_reg_dataout_458_port, Q(9) => 
                           bus_reg_dataout_457_port, Q(8) => 
                           bus_reg_dataout_456_port, Q(7) => 
                           bus_reg_dataout_455_port, Q(6) => 
                           bus_reg_dataout_454_port, Q(5) => 
                           bus_reg_dataout_453_port, Q(4) => 
                           bus_reg_dataout_452_port, Q(3) => 
                           bus_reg_dataout_451_port, Q(2) => 
                           bus_reg_dataout_450_port, Q(1) => 
                           bus_reg_dataout_449_port, Q(0) => 
                           bus_reg_dataout_448_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_22_port);
   BLOCKi_23 : reg_generic_N32_RSTVAL0_65 port map( D(31) => 
                           internal_inloc_data_0_31_port, D(30) => 
                           internal_inloc_data_0_30_port, D(29) => 
                           internal_inloc_data_0_29_port, D(28) => 
                           internal_inloc_data_0_28_port, D(27) => 
                           internal_inloc_data_0_27_port, D(26) => 
                           internal_inloc_data_0_26_port, D(25) => 
                           internal_inloc_data_0_25_port, D(24) => 
                           internal_inloc_data_0_24_port, D(23) => 
                           internal_inloc_data_0_23_port, D(22) => 
                           internal_inloc_data_0_22_port, D(21) => 
                           internal_inloc_data_0_21_port, D(20) => 
                           internal_inloc_data_0_20_port, D(19) => 
                           internal_inloc_data_0_19_port, D(18) => 
                           internal_inloc_data_0_18_port, D(17) => 
                           internal_inloc_data_0_17_port, D(16) => 
                           internal_inloc_data_0_16_port, D(15) => 
                           internal_inloc_data_0_15_port, D(14) => 
                           internal_inloc_data_0_14_port, D(13) => 
                           internal_inloc_data_0_13_port, D(12) => 
                           internal_inloc_data_0_12_port, D(11) => 
                           internal_inloc_data_0_11_port, D(10) => 
                           internal_inloc_data_0_10_port, D(9) => 
                           internal_inloc_data_0_9_port, D(8) => 
                           internal_inloc_data_0_8_port, D(7) => 
                           internal_inloc_data_0_7_port, D(6) => 
                           internal_inloc_data_0_6_port, D(5) => 
                           internal_inloc_data_0_5_port, D(4) => 
                           internal_inloc_data_0_4_port, D(3) => 
                           internal_inloc_data_0_3_port, D(2) => 
                           internal_inloc_data_0_2_port, D(1) => 
                           internal_inloc_data_0_1_port, D(0) => 
                           internal_inloc_data_0_0_port, Q(31) => 
                           bus_reg_dataout_511_port, Q(30) => 
                           bus_reg_dataout_510_port, Q(29) => 
                           bus_reg_dataout_509_port, Q(28) => 
                           bus_reg_dataout_508_port, Q(27) => 
                           bus_reg_dataout_507_port, Q(26) => 
                           bus_reg_dataout_506_port, Q(25) => 
                           bus_reg_dataout_505_port, Q(24) => 
                           bus_reg_dataout_504_port, Q(23) => 
                           bus_reg_dataout_503_port, Q(22) => 
                           bus_reg_dataout_502_port, Q(21) => 
                           bus_reg_dataout_501_port, Q(20) => 
                           bus_reg_dataout_500_port, Q(19) => 
                           bus_reg_dataout_499_port, Q(18) => 
                           bus_reg_dataout_498_port, Q(17) => 
                           bus_reg_dataout_497_port, Q(16) => 
                           bus_reg_dataout_496_port, Q(15) => 
                           bus_reg_dataout_495_port, Q(14) => 
                           bus_reg_dataout_494_port, Q(13) => 
                           bus_reg_dataout_493_port, Q(12) => 
                           bus_reg_dataout_492_port, Q(11) => 
                           bus_reg_dataout_491_port, Q(10) => 
                           bus_reg_dataout_490_port, Q(9) => 
                           bus_reg_dataout_489_port, Q(8) => 
                           bus_reg_dataout_488_port, Q(7) => 
                           bus_reg_dataout_487_port, Q(6) => 
                           bus_reg_dataout_486_port, Q(5) => 
                           bus_reg_dataout_485_port, Q(4) => 
                           bus_reg_dataout_484_port, Q(3) => 
                           bus_reg_dataout_483_port, Q(2) => 
                           bus_reg_dataout_482_port, Q(1) => 
                           bus_reg_dataout_481_port, Q(0) => 
                           bus_reg_dataout_480_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_23_port);
   MUX_SELINPUT_24 : mux_N32_M1_32 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1366
                           , Y(30) => n1358, Y(29) => n1350, Y(28) => n1342, 
                           Y(27) => n1334, Y(26) => n1326, Y(25) => n1318, 
                           Y(24) => n1310, Y(23) => n1302, Y(22) => n1294, 
                           Y(21) => n1286, Y(20) => n1278, Y(19) => n1270, 
                           Y(18) => n1262, Y(17) => n1254, Y(16) => n1246, 
                           Y(15) => n1238, Y(14) => n1230, Y(13) => n1222, 
                           Y(12) => n1214, Y(11) => n1206, Y(10) => n1198, Y(9)
                           => n1190, Y(8) => n1182, Y(7) => n1174, Y(6) => 
                           n1166, Y(5) => n1158, Y(4) => n1150, Y(3) => n1142, 
                           Y(2) => n1134, Y(1) => n1126, Y(0) => n1118);
   BLOCKi_24 : reg_generic_N32_RSTVAL0_64 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_543_port, Q(30) => 
                           bus_reg_dataout_542_port, Q(29) => 
                           bus_reg_dataout_541_port, Q(28) => 
                           bus_reg_dataout_540_port, Q(27) => 
                           bus_reg_dataout_539_port, Q(26) => 
                           bus_reg_dataout_538_port, Q(25) => 
                           bus_reg_dataout_537_port, Q(24) => 
                           bus_reg_dataout_536_port, Q(23) => 
                           bus_reg_dataout_535_port, Q(22) => 
                           bus_reg_dataout_534_port, Q(21) => 
                           bus_reg_dataout_533_port, Q(20) => 
                           bus_reg_dataout_532_port, Q(19) => 
                           bus_reg_dataout_531_port, Q(18) => 
                           bus_reg_dataout_530_port, Q(17) => 
                           bus_reg_dataout_529_port, Q(16) => 
                           bus_reg_dataout_528_port, Q(15) => 
                           bus_reg_dataout_527_port, Q(14) => 
                           bus_reg_dataout_526_port, Q(13) => 
                           bus_reg_dataout_525_port, Q(12) => 
                           bus_reg_dataout_524_port, Q(11) => 
                           bus_reg_dataout_523_port, Q(10) => 
                           bus_reg_dataout_522_port, Q(9) => 
                           bus_reg_dataout_521_port, Q(8) => 
                           bus_reg_dataout_520_port, Q(7) => 
                           bus_reg_dataout_519_port, Q(6) => 
                           bus_reg_dataout_518_port, Q(5) => 
                           bus_reg_dataout_517_port, Q(4) => 
                           bus_reg_dataout_516_port, Q(3) => 
                           bus_reg_dataout_515_port, Q(2) => 
                           bus_reg_dataout_514_port, Q(1) => 
                           bus_reg_dataout_513_port, Q(0) => 
                           bus_reg_dataout_512_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_24_port);
   BLOCKi_25 : reg_generic_N32_RSTVAL0_63 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_575_port, Q(30) => 
                           bus_reg_dataout_574_port, Q(29) => 
                           bus_reg_dataout_573_port, Q(28) => 
                           bus_reg_dataout_572_port, Q(27) => 
                           bus_reg_dataout_571_port, Q(26) => 
                           bus_reg_dataout_570_port, Q(25) => 
                           bus_reg_dataout_569_port, Q(24) => 
                           bus_reg_dataout_568_port, Q(23) => 
                           bus_reg_dataout_567_port, Q(22) => 
                           bus_reg_dataout_566_port, Q(21) => 
                           bus_reg_dataout_565_port, Q(20) => 
                           bus_reg_dataout_564_port, Q(19) => 
                           bus_reg_dataout_563_port, Q(18) => 
                           bus_reg_dataout_562_port, Q(17) => 
                           bus_reg_dataout_561_port, Q(16) => 
                           bus_reg_dataout_560_port, Q(15) => 
                           bus_reg_dataout_559_port, Q(14) => 
                           bus_reg_dataout_558_port, Q(13) => 
                           bus_reg_dataout_557_port, Q(12) => 
                           bus_reg_dataout_556_port, Q(11) => 
                           bus_reg_dataout_555_port, Q(10) => 
                           bus_reg_dataout_554_port, Q(9) => 
                           bus_reg_dataout_553_port, Q(8) => 
                           bus_reg_dataout_552_port, Q(7) => 
                           bus_reg_dataout_551_port, Q(6) => 
                           bus_reg_dataout_550_port, Q(5) => 
                           bus_reg_dataout_549_port, Q(4) => 
                           bus_reg_dataout_548_port, Q(3) => 
                           bus_reg_dataout_547_port, Q(2) => 
                           bus_reg_dataout_546_port, Q(1) => 
                           bus_reg_dataout_545_port, Q(0) => 
                           bus_reg_dataout_544_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_25_port);
   MUX_SELINPUT_26 : mux_N32_M1_31 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1365
                           , Y(30) => n1357, Y(29) => n1349, Y(28) => n1341, 
                           Y(27) => n1333, Y(26) => n1325, Y(25) => n1317, 
                           Y(24) => n1309, Y(23) => n1301, Y(22) => n1293, 
                           Y(21) => n1285, Y(20) => n1277, Y(19) => n1269, 
                           Y(18) => n1261, Y(17) => n1253, Y(16) => n1245, 
                           Y(15) => n1237, Y(14) => n1229, Y(13) => n1221, 
                           Y(12) => n1213, Y(11) => n1205, Y(10) => n1197, Y(9)
                           => n1189, Y(8) => n1181, Y(7) => n1173, Y(6) => 
                           n1165, Y(5) => n1157, Y(4) => n1149, Y(3) => n1141, 
                           Y(2) => n1133, Y(1) => n1125, Y(0) => n1117);
   BLOCKi_26 : reg_generic_N32_RSTVAL0_62 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_607_port, Q(30) => 
                           bus_reg_dataout_606_port, Q(29) => 
                           bus_reg_dataout_605_port, Q(28) => 
                           bus_reg_dataout_604_port, Q(27) => 
                           bus_reg_dataout_603_port, Q(26) => 
                           bus_reg_dataout_602_port, Q(25) => 
                           bus_reg_dataout_601_port, Q(24) => 
                           bus_reg_dataout_600_port, Q(23) => 
                           bus_reg_dataout_599_port, Q(22) => 
                           bus_reg_dataout_598_port, Q(21) => 
                           bus_reg_dataout_597_port, Q(20) => 
                           bus_reg_dataout_596_port, Q(19) => 
                           bus_reg_dataout_595_port, Q(18) => 
                           bus_reg_dataout_594_port, Q(17) => 
                           bus_reg_dataout_593_port, Q(16) => 
                           bus_reg_dataout_592_port, Q(15) => 
                           bus_reg_dataout_591_port, Q(14) => 
                           bus_reg_dataout_590_port, Q(13) => 
                           bus_reg_dataout_589_port, Q(12) => 
                           bus_reg_dataout_588_port, Q(11) => 
                           bus_reg_dataout_587_port, Q(10) => 
                           bus_reg_dataout_586_port, Q(9) => 
                           bus_reg_dataout_585_port, Q(8) => 
                           bus_reg_dataout_584_port, Q(7) => 
                           bus_reg_dataout_583_port, Q(6) => 
                           bus_reg_dataout_582_port, Q(5) => 
                           bus_reg_dataout_581_port, Q(4) => 
                           bus_reg_dataout_580_port, Q(3) => 
                           bus_reg_dataout_579_port, Q(2) => 
                           bus_reg_dataout_578_port, Q(1) => 
                           bus_reg_dataout_577_port, Q(0) => 
                           bus_reg_dataout_576_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_26_port);
   BLOCKi_27 : reg_generic_N32_RSTVAL0_61 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_639_port, Q(30) => 
                           bus_reg_dataout_638_port, Q(29) => 
                           bus_reg_dataout_637_port, Q(28) => 
                           bus_reg_dataout_636_port, Q(27) => 
                           bus_reg_dataout_635_port, Q(26) => 
                           bus_reg_dataout_634_port, Q(25) => 
                           bus_reg_dataout_633_port, Q(24) => 
                           bus_reg_dataout_632_port, Q(23) => 
                           bus_reg_dataout_631_port, Q(22) => 
                           bus_reg_dataout_630_port, Q(21) => 
                           bus_reg_dataout_629_port, Q(20) => 
                           bus_reg_dataout_628_port, Q(19) => 
                           bus_reg_dataout_627_port, Q(18) => 
                           bus_reg_dataout_626_port, Q(17) => 
                           bus_reg_dataout_625_port, Q(16) => 
                           bus_reg_dataout_624_port, Q(15) => 
                           bus_reg_dataout_623_port, Q(14) => 
                           bus_reg_dataout_622_port, Q(13) => 
                           bus_reg_dataout_621_port, Q(12) => 
                           bus_reg_dataout_620_port, Q(11) => 
                           bus_reg_dataout_619_port, Q(10) => 
                           bus_reg_dataout_618_port, Q(9) => 
                           bus_reg_dataout_617_port, Q(8) => 
                           bus_reg_dataout_616_port, Q(7) => 
                           bus_reg_dataout_615_port, Q(6) => 
                           bus_reg_dataout_614_port, Q(5) => 
                           bus_reg_dataout_613_port, Q(4) => 
                           bus_reg_dataout_612_port, Q(3) => 
                           bus_reg_dataout_611_port, Q(2) => 
                           bus_reg_dataout_610_port, Q(1) => 
                           bus_reg_dataout_609_port, Q(0) => 
                           bus_reg_dataout_608_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_27_port);
   MUX_SELINPUT_28 : mux_N32_M1_30 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1364
                           , Y(30) => n1356, Y(29) => n1348, Y(28) => n1340, 
                           Y(27) => n1332, Y(26) => n1324, Y(25) => n1316, 
                           Y(24) => n1308, Y(23) => n1300, Y(22) => n1292, 
                           Y(21) => n1284, Y(20) => n1276, Y(19) => n1268, 
                           Y(18) => n1260, Y(17) => n1252, Y(16) => n1244, 
                           Y(15) => n1236, Y(14) => n1228, Y(13) => n1220, 
                           Y(12) => n1212, Y(11) => n1204, Y(10) => n1196, Y(9)
                           => n1188, Y(8) => n1180, Y(7) => n1172, Y(6) => 
                           n1164, Y(5) => n1156, Y(4) => n1148, Y(3) => n1140, 
                           Y(2) => n1132, Y(1) => n1124, Y(0) => n1116);
   BLOCKi_28 : reg_generic_N32_RSTVAL0_60 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_671_port, Q(30) => 
                           bus_reg_dataout_670_port, Q(29) => 
                           bus_reg_dataout_669_port, Q(28) => 
                           bus_reg_dataout_668_port, Q(27) => 
                           bus_reg_dataout_667_port, Q(26) => 
                           bus_reg_dataout_666_port, Q(25) => 
                           bus_reg_dataout_665_port, Q(24) => 
                           bus_reg_dataout_664_port, Q(23) => 
                           bus_reg_dataout_663_port, Q(22) => 
                           bus_reg_dataout_662_port, Q(21) => 
                           bus_reg_dataout_661_port, Q(20) => 
                           bus_reg_dataout_660_port, Q(19) => 
                           bus_reg_dataout_659_port, Q(18) => 
                           bus_reg_dataout_658_port, Q(17) => 
                           bus_reg_dataout_657_port, Q(16) => 
                           bus_reg_dataout_656_port, Q(15) => 
                           bus_reg_dataout_655_port, Q(14) => 
                           bus_reg_dataout_654_port, Q(13) => 
                           bus_reg_dataout_653_port, Q(12) => 
                           bus_reg_dataout_652_port, Q(11) => 
                           bus_reg_dataout_651_port, Q(10) => 
                           bus_reg_dataout_650_port, Q(9) => 
                           bus_reg_dataout_649_port, Q(8) => 
                           bus_reg_dataout_648_port, Q(7) => 
                           bus_reg_dataout_647_port, Q(6) => 
                           bus_reg_dataout_646_port, Q(5) => 
                           bus_reg_dataout_645_port, Q(4) => 
                           bus_reg_dataout_644_port, Q(3) => 
                           bus_reg_dataout_643_port, Q(2) => 
                           bus_reg_dataout_642_port, Q(1) => 
                           bus_reg_dataout_641_port, Q(0) => 
                           bus_reg_dataout_640_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_28_port);
   BLOCKi_29 : reg_generic_N32_RSTVAL0_59 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_703_port, Q(30) => 
                           bus_reg_dataout_702_port, Q(29) => 
                           bus_reg_dataout_701_port, Q(28) => 
                           bus_reg_dataout_700_port, Q(27) => 
                           bus_reg_dataout_699_port, Q(26) => 
                           bus_reg_dataout_698_port, Q(25) => 
                           bus_reg_dataout_697_port, Q(24) => 
                           bus_reg_dataout_696_port, Q(23) => 
                           bus_reg_dataout_695_port, Q(22) => 
                           bus_reg_dataout_694_port, Q(21) => 
                           bus_reg_dataout_693_port, Q(20) => 
                           bus_reg_dataout_692_port, Q(19) => 
                           bus_reg_dataout_691_port, Q(18) => 
                           bus_reg_dataout_690_port, Q(17) => 
                           bus_reg_dataout_689_port, Q(16) => 
                           bus_reg_dataout_688_port, Q(15) => 
                           bus_reg_dataout_687_port, Q(14) => 
                           bus_reg_dataout_686_port, Q(13) => 
                           bus_reg_dataout_685_port, Q(12) => 
                           bus_reg_dataout_684_port, Q(11) => 
                           bus_reg_dataout_683_port, Q(10) => 
                           bus_reg_dataout_682_port, Q(9) => 
                           bus_reg_dataout_681_port, Q(8) => 
                           bus_reg_dataout_680_port, Q(7) => 
                           bus_reg_dataout_679_port, Q(6) => 
                           bus_reg_dataout_678_port, Q(5) => 
                           bus_reg_dataout_677_port, Q(4) => 
                           bus_reg_dataout_676_port, Q(3) => 
                           bus_reg_dataout_675_port, Q(2) => 
                           bus_reg_dataout_674_port, Q(1) => 
                           bus_reg_dataout_673_port, Q(0) => 
                           bus_reg_dataout_672_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_29_port);
   MUX_SELINPUT_30 : mux_N32_M1_29 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1363
                           , Y(30) => n1355, Y(29) => n1347, Y(28) => n1339, 
                           Y(27) => n1331, Y(26) => n1323, Y(25) => n1315, 
                           Y(24) => n1307, Y(23) => n1299, Y(22) => n1291, 
                           Y(21) => n1283, Y(20) => n1275, Y(19) => n1267, 
                           Y(18) => n1259, Y(17) => n1251, Y(16) => n1243, 
                           Y(15) => n1235, Y(14) => n1227, Y(13) => n1219, 
                           Y(12) => n1211, Y(11) => n1203, Y(10) => n1195, Y(9)
                           => n1187, Y(8) => n1179, Y(7) => n1171, Y(6) => 
                           n1163, Y(5) => n1155, Y(4) => n1147, Y(3) => n1139, 
                           Y(2) => n1131, Y(1) => n1123, Y(0) => n1115);
   BLOCKi_30 : reg_generic_N32_RSTVAL0_58 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_735_port, Q(30) => 
                           bus_reg_dataout_734_port, Q(29) => 
                           bus_reg_dataout_733_port, Q(28) => 
                           bus_reg_dataout_732_port, Q(27) => 
                           bus_reg_dataout_731_port, Q(26) => 
                           bus_reg_dataout_730_port, Q(25) => 
                           bus_reg_dataout_729_port, Q(24) => 
                           bus_reg_dataout_728_port, Q(23) => 
                           bus_reg_dataout_727_port, Q(22) => 
                           bus_reg_dataout_726_port, Q(21) => 
                           bus_reg_dataout_725_port, Q(20) => 
                           bus_reg_dataout_724_port, Q(19) => 
                           bus_reg_dataout_723_port, Q(18) => 
                           bus_reg_dataout_722_port, Q(17) => 
                           bus_reg_dataout_721_port, Q(16) => 
                           bus_reg_dataout_720_port, Q(15) => 
                           bus_reg_dataout_719_port, Q(14) => 
                           bus_reg_dataout_718_port, Q(13) => 
                           bus_reg_dataout_717_port, Q(12) => 
                           bus_reg_dataout_716_port, Q(11) => 
                           bus_reg_dataout_715_port, Q(10) => 
                           bus_reg_dataout_714_port, Q(9) => 
                           bus_reg_dataout_713_port, Q(8) => 
                           bus_reg_dataout_712_port, Q(7) => 
                           bus_reg_dataout_711_port, Q(6) => 
                           bus_reg_dataout_710_port, Q(5) => 
                           bus_reg_dataout_709_port, Q(4) => 
                           bus_reg_dataout_708_port, Q(3) => 
                           bus_reg_dataout_707_port, Q(2) => 
                           bus_reg_dataout_706_port, Q(1) => 
                           bus_reg_dataout_705_port, Q(0) => 
                           bus_reg_dataout_704_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_30_port);
   BLOCKi_31 : reg_generic_N32_RSTVAL0_57 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_767_port, Q(30) => 
                           bus_reg_dataout_766_port, Q(29) => 
                           bus_reg_dataout_765_port, Q(28) => 
                           bus_reg_dataout_764_port, Q(27) => 
                           bus_reg_dataout_763_port, Q(26) => 
                           bus_reg_dataout_762_port, Q(25) => 
                           bus_reg_dataout_761_port, Q(24) => 
                           bus_reg_dataout_760_port, Q(23) => 
                           bus_reg_dataout_759_port, Q(22) => 
                           bus_reg_dataout_758_port, Q(21) => 
                           bus_reg_dataout_757_port, Q(20) => 
                           bus_reg_dataout_756_port, Q(19) => 
                           bus_reg_dataout_755_port, Q(18) => 
                           bus_reg_dataout_754_port, Q(17) => 
                           bus_reg_dataout_753_port, Q(16) => 
                           bus_reg_dataout_752_port, Q(15) => 
                           bus_reg_dataout_751_port, Q(14) => 
                           bus_reg_dataout_750_port, Q(13) => 
                           bus_reg_dataout_749_port, Q(12) => 
                           bus_reg_dataout_748_port, Q(11) => 
                           bus_reg_dataout_747_port, Q(10) => 
                           bus_reg_dataout_746_port, Q(9) => 
                           bus_reg_dataout_745_port, Q(8) => 
                           bus_reg_dataout_744_port, Q(7) => 
                           bus_reg_dataout_743_port, Q(6) => 
                           bus_reg_dataout_742_port, Q(5) => 
                           bus_reg_dataout_741_port, Q(4) => 
                           bus_reg_dataout_740_port, Q(3) => 
                           bus_reg_dataout_739_port, Q(2) => 
                           bus_reg_dataout_738_port, Q(1) => 
                           bus_reg_dataout_737_port, Q(0) => 
                           bus_reg_dataout_736_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_31_port);
   MUX_SELINPUT_32 : mux_N32_M1_28 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1362
                           , Y(30) => n1354, Y(29) => n1346, Y(28) => n1338, 
                           Y(27) => n1330, Y(26) => n1322, Y(25) => n1314, 
                           Y(24) => n1306, Y(23) => n1298, Y(22) => n1290, 
                           Y(21) => n1282, Y(20) => n1274, Y(19) => n1266, 
                           Y(18) => n1258, Y(17) => n1250, Y(16) => n1242, 
                           Y(15) => n1234, Y(14) => n1226, Y(13) => n1218, 
                           Y(12) => n1210, Y(11) => n1202, Y(10) => n1194, Y(9)
                           => n1186, Y(8) => n1178, Y(7) => n1170, Y(6) => 
                           n1162, Y(5) => n1154, Y(4) => n1146, Y(3) => n1138, 
                           Y(2) => n1130, Y(1) => n1122, Y(0) => n1114);
   BLOCKi_32 : reg_generic_N32_RSTVAL0_56 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_799_port, Q(30) => 
                           bus_reg_dataout_798_port, Q(29) => 
                           bus_reg_dataout_797_port, Q(28) => 
                           bus_reg_dataout_796_port, Q(27) => 
                           bus_reg_dataout_795_port, Q(26) => 
                           bus_reg_dataout_794_port, Q(25) => 
                           bus_reg_dataout_793_port, Q(24) => 
                           bus_reg_dataout_792_port, Q(23) => 
                           bus_reg_dataout_791_port, Q(22) => 
                           bus_reg_dataout_790_port, Q(21) => 
                           bus_reg_dataout_789_port, Q(20) => 
                           bus_reg_dataout_788_port, Q(19) => 
                           bus_reg_dataout_787_port, Q(18) => 
                           bus_reg_dataout_786_port, Q(17) => 
                           bus_reg_dataout_785_port, Q(16) => 
                           bus_reg_dataout_784_port, Q(15) => 
                           bus_reg_dataout_783_port, Q(14) => 
                           bus_reg_dataout_782_port, Q(13) => 
                           bus_reg_dataout_781_port, Q(12) => 
                           bus_reg_dataout_780_port, Q(11) => 
                           bus_reg_dataout_779_port, Q(10) => 
                           bus_reg_dataout_778_port, Q(9) => 
                           bus_reg_dataout_777_port, Q(8) => 
                           bus_reg_dataout_776_port, Q(7) => 
                           bus_reg_dataout_775_port, Q(6) => 
                           bus_reg_dataout_774_port, Q(5) => 
                           bus_reg_dataout_773_port, Q(4) => 
                           bus_reg_dataout_772_port, Q(3) => 
                           bus_reg_dataout_771_port, Q(2) => 
                           bus_reg_dataout_770_port, Q(1) => 
                           bus_reg_dataout_769_port, Q(0) => 
                           bus_reg_dataout_768_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_32_port);
   BLOCKi_33 : reg_generic_N32_RSTVAL0_55 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_831_port, Q(30) => 
                           bus_reg_dataout_830_port, Q(29) => 
                           bus_reg_dataout_829_port, Q(28) => 
                           bus_reg_dataout_828_port, Q(27) => 
                           bus_reg_dataout_827_port, Q(26) => 
                           bus_reg_dataout_826_port, Q(25) => 
                           bus_reg_dataout_825_port, Q(24) => 
                           bus_reg_dataout_824_port, Q(23) => 
                           bus_reg_dataout_823_port, Q(22) => 
                           bus_reg_dataout_822_port, Q(21) => 
                           bus_reg_dataout_821_port, Q(20) => 
                           bus_reg_dataout_820_port, Q(19) => 
                           bus_reg_dataout_819_port, Q(18) => 
                           bus_reg_dataout_818_port, Q(17) => 
                           bus_reg_dataout_817_port, Q(16) => 
                           bus_reg_dataout_816_port, Q(15) => 
                           bus_reg_dataout_815_port, Q(14) => 
                           bus_reg_dataout_814_port, Q(13) => 
                           bus_reg_dataout_813_port, Q(12) => 
                           bus_reg_dataout_812_port, Q(11) => 
                           bus_reg_dataout_811_port, Q(10) => 
                           bus_reg_dataout_810_port, Q(9) => 
                           bus_reg_dataout_809_port, Q(8) => 
                           bus_reg_dataout_808_port, Q(7) => 
                           bus_reg_dataout_807_port, Q(6) => 
                           bus_reg_dataout_806_port, Q(5) => 
                           bus_reg_dataout_805_port, Q(4) => 
                           bus_reg_dataout_804_port, Q(3) => 
                           bus_reg_dataout_803_port, Q(2) => 
                           bus_reg_dataout_802_port, Q(1) => 
                           bus_reg_dataout_801_port, Q(0) => 
                           bus_reg_dataout_800_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_33_port);
   MUX_SELINPUT_34 : mux_N32_M1_27 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1361
                           , Y(30) => n1353, Y(29) => n1345, Y(28) => n1337, 
                           Y(27) => n1329, Y(26) => n1321, Y(25) => n1313, 
                           Y(24) => n1305, Y(23) => n1297, Y(22) => n1289, 
                           Y(21) => n1281, Y(20) => n1273, Y(19) => n1265, 
                           Y(18) => n1257, Y(17) => n1249, Y(16) => n1241, 
                           Y(15) => n1233, Y(14) => n1225, Y(13) => n1217, 
                           Y(12) => n1209, Y(11) => n1201, Y(10) => n1193, Y(9)
                           => n1185, Y(8) => n1177, Y(7) => n1169, Y(6) => 
                           n1161, Y(5) => n1153, Y(4) => n1145, Y(3) => n1137, 
                           Y(2) => n1129, Y(1) => n1121, Y(0) => n1113);
   BLOCKi_34 : reg_generic_N32_RSTVAL0_54 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_863_port, Q(30) => 
                           bus_reg_dataout_862_port, Q(29) => 
                           bus_reg_dataout_861_port, Q(28) => 
                           bus_reg_dataout_860_port, Q(27) => 
                           bus_reg_dataout_859_port, Q(26) => 
                           bus_reg_dataout_858_port, Q(25) => 
                           bus_reg_dataout_857_port, Q(24) => 
                           bus_reg_dataout_856_port, Q(23) => 
                           bus_reg_dataout_855_port, Q(22) => 
                           bus_reg_dataout_854_port, Q(21) => 
                           bus_reg_dataout_853_port, Q(20) => 
                           bus_reg_dataout_852_port, Q(19) => 
                           bus_reg_dataout_851_port, Q(18) => 
                           bus_reg_dataout_850_port, Q(17) => 
                           bus_reg_dataout_849_port, Q(16) => 
                           bus_reg_dataout_848_port, Q(15) => 
                           bus_reg_dataout_847_port, Q(14) => 
                           bus_reg_dataout_846_port, Q(13) => 
                           bus_reg_dataout_845_port, Q(12) => 
                           bus_reg_dataout_844_port, Q(11) => 
                           bus_reg_dataout_843_port, Q(10) => 
                           bus_reg_dataout_842_port, Q(9) => 
                           bus_reg_dataout_841_port, Q(8) => 
                           bus_reg_dataout_840_port, Q(7) => 
                           bus_reg_dataout_839_port, Q(6) => 
                           bus_reg_dataout_838_port, Q(5) => 
                           bus_reg_dataout_837_port, Q(4) => 
                           bus_reg_dataout_836_port, Q(3) => 
                           bus_reg_dataout_835_port, Q(2) => 
                           bus_reg_dataout_834_port, Q(1) => 
                           bus_reg_dataout_833_port, Q(0) => 
                           bus_reg_dataout_832_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_34_port);
   BLOCKi_35 : reg_generic_N32_RSTVAL0_53 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_895_port, Q(30) => 
                           bus_reg_dataout_894_port, Q(29) => 
                           bus_reg_dataout_893_port, Q(28) => 
                           bus_reg_dataout_892_port, Q(27) => 
                           bus_reg_dataout_891_port, Q(26) => 
                           bus_reg_dataout_890_port, Q(25) => 
                           bus_reg_dataout_889_port, Q(24) => 
                           bus_reg_dataout_888_port, Q(23) => 
                           bus_reg_dataout_887_port, Q(22) => 
                           bus_reg_dataout_886_port, Q(21) => 
                           bus_reg_dataout_885_port, Q(20) => 
                           bus_reg_dataout_884_port, Q(19) => 
                           bus_reg_dataout_883_port, Q(18) => 
                           bus_reg_dataout_882_port, Q(17) => 
                           bus_reg_dataout_881_port, Q(16) => 
                           bus_reg_dataout_880_port, Q(15) => 
                           bus_reg_dataout_879_port, Q(14) => 
                           bus_reg_dataout_878_port, Q(13) => 
                           bus_reg_dataout_877_port, Q(12) => 
                           bus_reg_dataout_876_port, Q(11) => 
                           bus_reg_dataout_875_port, Q(10) => 
                           bus_reg_dataout_874_port, Q(9) => 
                           bus_reg_dataout_873_port, Q(8) => 
                           bus_reg_dataout_872_port, Q(7) => 
                           bus_reg_dataout_871_port, Q(6) => 
                           bus_reg_dataout_870_port, Q(5) => 
                           bus_reg_dataout_869_port, Q(4) => 
                           bus_reg_dataout_868_port, Q(3) => 
                           bus_reg_dataout_867_port, Q(2) => 
                           bus_reg_dataout_866_port, Q(1) => 
                           bus_reg_dataout_865_port, Q(0) => 
                           bus_reg_dataout_864_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_35_port);
   MUX_SELINPUT_36 : mux_N32_M1_26 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1360
                           , Y(30) => n1352, Y(29) => n1344, Y(28) => n1336, 
                           Y(27) => n1328, Y(26) => n1320, Y(25) => n1312, 
                           Y(24) => n1304, Y(23) => n1296, Y(22) => n1288, 
                           Y(21) => n1280, Y(20) => n1272, Y(19) => n1264, 
                           Y(18) => n1256, Y(17) => n1248, Y(16) => n1240, 
                           Y(15) => n1232, Y(14) => n1224, Y(13) => n1216, 
                           Y(12) => n1208, Y(11) => n1200, Y(10) => n1192, Y(9)
                           => n1184, Y(8) => n1176, Y(7) => n1168, Y(6) => 
                           n1160, Y(5) => n1152, Y(4) => n1144, Y(3) => n1136, 
                           Y(2) => n1128, Y(1) => n1120, Y(0) => n1112);
   BLOCKi_36 : reg_generic_N32_RSTVAL0_52 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_927_port, Q(30) => 
                           bus_reg_dataout_926_port, Q(29) => 
                           bus_reg_dataout_925_port, Q(28) => 
                           bus_reg_dataout_924_port, Q(27) => 
                           bus_reg_dataout_923_port, Q(26) => 
                           bus_reg_dataout_922_port, Q(25) => 
                           bus_reg_dataout_921_port, Q(24) => 
                           bus_reg_dataout_920_port, Q(23) => 
                           bus_reg_dataout_919_port, Q(22) => 
                           bus_reg_dataout_918_port, Q(21) => 
                           bus_reg_dataout_917_port, Q(20) => 
                           bus_reg_dataout_916_port, Q(19) => 
                           bus_reg_dataout_915_port, Q(18) => 
                           bus_reg_dataout_914_port, Q(17) => 
                           bus_reg_dataout_913_port, Q(16) => 
                           bus_reg_dataout_912_port, Q(15) => 
                           bus_reg_dataout_911_port, Q(14) => 
                           bus_reg_dataout_910_port, Q(13) => 
                           bus_reg_dataout_909_port, Q(12) => 
                           bus_reg_dataout_908_port, Q(11) => 
                           bus_reg_dataout_907_port, Q(10) => 
                           bus_reg_dataout_906_port, Q(9) => 
                           bus_reg_dataout_905_port, Q(8) => 
                           bus_reg_dataout_904_port, Q(7) => 
                           bus_reg_dataout_903_port, Q(6) => 
                           bus_reg_dataout_902_port, Q(5) => 
                           bus_reg_dataout_901_port, Q(4) => 
                           bus_reg_dataout_900_port, Q(3) => 
                           bus_reg_dataout_899_port, Q(2) => 
                           bus_reg_dataout_898_port, Q(1) => 
                           bus_reg_dataout_897_port, Q(0) => 
                           bus_reg_dataout_896_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_36_port);
   BLOCKi_37 : reg_generic_N32_RSTVAL0_51 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_959_port, Q(30) => 
                           bus_reg_dataout_958_port, Q(29) => 
                           bus_reg_dataout_957_port, Q(28) => 
                           bus_reg_dataout_956_port, Q(27) => 
                           bus_reg_dataout_955_port, Q(26) => 
                           bus_reg_dataout_954_port, Q(25) => 
                           bus_reg_dataout_953_port, Q(24) => 
                           bus_reg_dataout_952_port, Q(23) => 
                           bus_reg_dataout_951_port, Q(22) => 
                           bus_reg_dataout_950_port, Q(21) => 
                           bus_reg_dataout_949_port, Q(20) => 
                           bus_reg_dataout_948_port, Q(19) => 
                           bus_reg_dataout_947_port, Q(18) => 
                           bus_reg_dataout_946_port, Q(17) => 
                           bus_reg_dataout_945_port, Q(16) => 
                           bus_reg_dataout_944_port, Q(15) => 
                           bus_reg_dataout_943_port, Q(14) => 
                           bus_reg_dataout_942_port, Q(13) => 
                           bus_reg_dataout_941_port, Q(12) => 
                           bus_reg_dataout_940_port, Q(11) => 
                           bus_reg_dataout_939_port, Q(10) => 
                           bus_reg_dataout_938_port, Q(9) => 
                           bus_reg_dataout_937_port, Q(8) => 
                           bus_reg_dataout_936_port, Q(7) => 
                           bus_reg_dataout_935_port, Q(6) => 
                           bus_reg_dataout_934_port, Q(5) => 
                           bus_reg_dataout_933_port, Q(4) => 
                           bus_reg_dataout_932_port, Q(3) => 
                           bus_reg_dataout_931_port, Q(2) => 
                           bus_reg_dataout_930_port, Q(1) => 
                           bus_reg_dataout_929_port, Q(0) => 
                           bus_reg_dataout_928_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_37_port);
   MUX_SELINPUT_38 : mux_N32_M1_25 port map( S => c_swin_masked_1bit_1_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1359
                           , Y(30) => n1351, Y(29) => n1343, Y(28) => n1335, 
                           Y(27) => n1327, Y(26) => n1319, Y(25) => n1311, 
                           Y(24) => n1303, Y(23) => n1295, Y(22) => n1287, 
                           Y(21) => n1279, Y(20) => n1271, Y(19) => n1263, 
                           Y(18) => n1255, Y(17) => n1247, Y(16) => n1239, 
                           Y(15) => n1231, Y(14) => n1223, Y(13) => n1215, 
                           Y(12) => n1207, Y(11) => n1199, Y(10) => n1191, Y(9)
                           => n1183, Y(8) => n1175, Y(7) => n1167, Y(6) => 
                           n1159, Y(5) => n1151, Y(4) => n1143, Y(3) => n1135, 
                           Y(2) => n1127, Y(1) => n1119, Y(0) => n1111);
   BLOCKi_38 : reg_generic_N32_RSTVAL0_50 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_991_port, Q(30) => 
                           bus_reg_dataout_990_port, Q(29) => 
                           bus_reg_dataout_989_port, Q(28) => 
                           bus_reg_dataout_988_port, Q(27) => 
                           bus_reg_dataout_987_port, Q(26) => 
                           bus_reg_dataout_986_port, Q(25) => 
                           bus_reg_dataout_985_port, Q(24) => 
                           bus_reg_dataout_984_port, Q(23) => 
                           bus_reg_dataout_983_port, Q(22) => 
                           bus_reg_dataout_982_port, Q(21) => 
                           bus_reg_dataout_981_port, Q(20) => 
                           bus_reg_dataout_980_port, Q(19) => 
                           bus_reg_dataout_979_port, Q(18) => 
                           bus_reg_dataout_978_port, Q(17) => 
                           bus_reg_dataout_977_port, Q(16) => 
                           bus_reg_dataout_976_port, Q(15) => 
                           bus_reg_dataout_975_port, Q(14) => 
                           bus_reg_dataout_974_port, Q(13) => 
                           bus_reg_dataout_973_port, Q(12) => 
                           bus_reg_dataout_972_port, Q(11) => 
                           bus_reg_dataout_971_port, Q(10) => 
                           bus_reg_dataout_970_port, Q(9) => 
                           bus_reg_dataout_969_port, Q(8) => 
                           bus_reg_dataout_968_port, Q(7) => 
                           bus_reg_dataout_967_port, Q(6) => 
                           bus_reg_dataout_966_port, Q(5) => 
                           bus_reg_dataout_965_port, Q(4) => 
                           bus_reg_dataout_964_port, Q(3) => 
                           bus_reg_dataout_963_port, Q(2) => 
                           bus_reg_dataout_962_port, Q(1) => 
                           bus_reg_dataout_961_port, Q(0) => 
                           bus_reg_dataout_960_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_38_port);
   BLOCKi_39 : reg_generic_N32_RSTVAL0_49 port map( D(31) => 
                           internal_inloc_data_1_31_port, D(30) => 
                           internal_inloc_data_1_30_port, D(29) => 
                           internal_inloc_data_1_29_port, D(28) => 
                           internal_inloc_data_1_28_port, D(27) => 
                           internal_inloc_data_1_27_port, D(26) => 
                           internal_inloc_data_1_26_port, D(25) => 
                           internal_inloc_data_1_25_port, D(24) => 
                           internal_inloc_data_1_24_port, D(23) => 
                           internal_inloc_data_1_23_port, D(22) => 
                           internal_inloc_data_1_22_port, D(21) => 
                           internal_inloc_data_1_21_port, D(20) => 
                           internal_inloc_data_1_20_port, D(19) => 
                           internal_inloc_data_1_19_port, D(18) => 
                           internal_inloc_data_1_18_port, D(17) => 
                           internal_inloc_data_1_17_port, D(16) => 
                           internal_inloc_data_1_16_port, D(15) => 
                           internal_inloc_data_1_15_port, D(14) => 
                           internal_inloc_data_1_14_port, D(13) => 
                           internal_inloc_data_1_13_port, D(12) => 
                           internal_inloc_data_1_12_port, D(11) => 
                           internal_inloc_data_1_11_port, D(10) => 
                           internal_inloc_data_1_10_port, D(9) => 
                           internal_inloc_data_1_9_port, D(8) => 
                           internal_inloc_data_1_8_port, D(7) => 
                           internal_inloc_data_1_7_port, D(6) => 
                           internal_inloc_data_1_6_port, D(5) => 
                           internal_inloc_data_1_5_port, D(4) => 
                           internal_inloc_data_1_4_port, D(3) => 
                           internal_inloc_data_1_3_port, D(2) => 
                           internal_inloc_data_1_2_port, D(1) => 
                           internal_inloc_data_1_1_port, D(0) => 
                           internal_inloc_data_1_0_port, Q(31) => 
                           bus_reg_dataout_1023_port, Q(30) => 
                           bus_reg_dataout_1022_port, Q(29) => 
                           bus_reg_dataout_1021_port, Q(28) => 
                           bus_reg_dataout_1020_port, Q(27) => 
                           bus_reg_dataout_1019_port, Q(26) => 
                           bus_reg_dataout_1018_port, Q(25) => 
                           bus_reg_dataout_1017_port, Q(24) => 
                           bus_reg_dataout_1016_port, Q(23) => 
                           bus_reg_dataout_1015_port, Q(22) => 
                           bus_reg_dataout_1014_port, Q(21) => 
                           bus_reg_dataout_1013_port, Q(20) => 
                           bus_reg_dataout_1012_port, Q(19) => 
                           bus_reg_dataout_1011_port, Q(18) => 
                           bus_reg_dataout_1010_port, Q(17) => 
                           bus_reg_dataout_1009_port, Q(16) => 
                           bus_reg_dataout_1008_port, Q(15) => 
                           bus_reg_dataout_1007_port, Q(14) => 
                           bus_reg_dataout_1006_port, Q(13) => 
                           bus_reg_dataout_1005_port, Q(12) => 
                           bus_reg_dataout_1004_port, Q(11) => 
                           bus_reg_dataout_1003_port, Q(10) => 
                           bus_reg_dataout_1002_port, Q(9) => 
                           bus_reg_dataout_1001_port, Q(8) => 
                           bus_reg_dataout_1000_port, Q(7) => 
                           bus_reg_dataout_999_port, Q(6) => 
                           bus_reg_dataout_998_port, Q(5) => 
                           bus_reg_dataout_997_port, Q(4) => 
                           bus_reg_dataout_996_port, Q(3) => 
                           bus_reg_dataout_995_port, Q(2) => 
                           bus_reg_dataout_994_port, Q(1) => 
                           bus_reg_dataout_993_port, Q(0) => 
                           bus_reg_dataout_992_port, Clk => CLK, Rst => RESET, 
                           Enable => en_regi_39_port);
   MUX_SELINPUT_40 : mux_N32_M1_24 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1110
                           , Y(30) => n1102, Y(29) => n1094, Y(28) => n1086, 
                           Y(27) => n1078, Y(26) => n1070, Y(25) => n1062, 
                           Y(24) => n1054, Y(23) => n1046, Y(22) => n1038, 
                           Y(21) => n1030, Y(20) => n1022, Y(19) => n1014, 
                           Y(18) => n1006, Y(17) => n998, Y(16) => n990, Y(15) 
                           => n982, Y(14) => n974, Y(13) => n966, Y(12) => n958
                           , Y(11) => n950, Y(10) => n942, Y(9) => n934, Y(8) 
                           => n926, Y(7) => n918, Y(6) => n910, Y(5) => n902, 
                           Y(4) => n894, Y(3) => n886, Y(2) => n878, Y(1) => 
                           n870, Y(0) => n862);
   BLOCKi_40 : reg_generic_N32_RSTVAL0_48 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1055_port, Q(30) => 
                           bus_reg_dataout_1054_port, Q(29) => 
                           bus_reg_dataout_1053_port, Q(28) => 
                           bus_reg_dataout_1052_port, Q(27) => 
                           bus_reg_dataout_1051_port, Q(26) => 
                           bus_reg_dataout_1050_port, Q(25) => 
                           bus_reg_dataout_1049_port, Q(24) => 
                           bus_reg_dataout_1048_port, Q(23) => 
                           bus_reg_dataout_1047_port, Q(22) => 
                           bus_reg_dataout_1046_port, Q(21) => 
                           bus_reg_dataout_1045_port, Q(20) => 
                           bus_reg_dataout_1044_port, Q(19) => 
                           bus_reg_dataout_1043_port, Q(18) => 
                           bus_reg_dataout_1042_port, Q(17) => 
                           bus_reg_dataout_1041_port, Q(16) => 
                           bus_reg_dataout_1040_port, Q(15) => 
                           bus_reg_dataout_1039_port, Q(14) => 
                           bus_reg_dataout_1038_port, Q(13) => 
                           bus_reg_dataout_1037_port, Q(12) => 
                           bus_reg_dataout_1036_port, Q(11) => 
                           bus_reg_dataout_1035_port, Q(10) => 
                           bus_reg_dataout_1034_port, Q(9) => 
                           bus_reg_dataout_1033_port, Q(8) => 
                           bus_reg_dataout_1032_port, Q(7) => 
                           bus_reg_dataout_1031_port, Q(6) => 
                           bus_reg_dataout_1030_port, Q(5) => 
                           bus_reg_dataout_1029_port, Q(4) => 
                           bus_reg_dataout_1028_port, Q(3) => 
                           bus_reg_dataout_1027_port, Q(2) => 
                           bus_reg_dataout_1026_port, Q(1) => 
                           bus_reg_dataout_1025_port, Q(0) => 
                           bus_reg_dataout_1024_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_40_port);
   BLOCKi_41 : reg_generic_N32_RSTVAL0_47 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1087_port, Q(30) => 
                           bus_reg_dataout_1086_port, Q(29) => 
                           bus_reg_dataout_1085_port, Q(28) => 
                           bus_reg_dataout_1084_port, Q(27) => 
                           bus_reg_dataout_1083_port, Q(26) => 
                           bus_reg_dataout_1082_port, Q(25) => 
                           bus_reg_dataout_1081_port, Q(24) => 
                           bus_reg_dataout_1080_port, Q(23) => 
                           bus_reg_dataout_1079_port, Q(22) => 
                           bus_reg_dataout_1078_port, Q(21) => 
                           bus_reg_dataout_1077_port, Q(20) => 
                           bus_reg_dataout_1076_port, Q(19) => 
                           bus_reg_dataout_1075_port, Q(18) => 
                           bus_reg_dataout_1074_port, Q(17) => 
                           bus_reg_dataout_1073_port, Q(16) => 
                           bus_reg_dataout_1072_port, Q(15) => 
                           bus_reg_dataout_1071_port, Q(14) => 
                           bus_reg_dataout_1070_port, Q(13) => 
                           bus_reg_dataout_1069_port, Q(12) => 
                           bus_reg_dataout_1068_port, Q(11) => 
                           bus_reg_dataout_1067_port, Q(10) => 
                           bus_reg_dataout_1066_port, Q(9) => 
                           bus_reg_dataout_1065_port, Q(8) => 
                           bus_reg_dataout_1064_port, Q(7) => 
                           bus_reg_dataout_1063_port, Q(6) => 
                           bus_reg_dataout_1062_port, Q(5) => 
                           bus_reg_dataout_1061_port, Q(4) => 
                           bus_reg_dataout_1060_port, Q(3) => 
                           bus_reg_dataout_1059_port, Q(2) => 
                           bus_reg_dataout_1058_port, Q(1) => 
                           bus_reg_dataout_1057_port, Q(0) => 
                           bus_reg_dataout_1056_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_41_port);
   MUX_SELINPUT_42 : mux_N32_M1_23 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1109
                           , Y(30) => n1101, Y(29) => n1093, Y(28) => n1085, 
                           Y(27) => n1077, Y(26) => n1069, Y(25) => n1061, 
                           Y(24) => n1053, Y(23) => n1045, Y(22) => n1037, 
                           Y(21) => n1029, Y(20) => n1021, Y(19) => n1013, 
                           Y(18) => n1005, Y(17) => n997, Y(16) => n989, Y(15) 
                           => n981, Y(14) => n973, Y(13) => n965, Y(12) => n957
                           , Y(11) => n949, Y(10) => n941, Y(9) => n933, Y(8) 
                           => n925, Y(7) => n917, Y(6) => n909, Y(5) => n901, 
                           Y(4) => n893, Y(3) => n885, Y(2) => n877, Y(1) => 
                           n869, Y(0) => n861);
   BLOCKi_42 : reg_generic_N32_RSTVAL0_46 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1119_port, Q(30) => 
                           bus_reg_dataout_1118_port, Q(29) => 
                           bus_reg_dataout_1117_port, Q(28) => 
                           bus_reg_dataout_1116_port, Q(27) => 
                           bus_reg_dataout_1115_port, Q(26) => 
                           bus_reg_dataout_1114_port, Q(25) => 
                           bus_reg_dataout_1113_port, Q(24) => 
                           bus_reg_dataout_1112_port, Q(23) => 
                           bus_reg_dataout_1111_port, Q(22) => 
                           bus_reg_dataout_1110_port, Q(21) => 
                           bus_reg_dataout_1109_port, Q(20) => 
                           bus_reg_dataout_1108_port, Q(19) => 
                           bus_reg_dataout_1107_port, Q(18) => 
                           bus_reg_dataout_1106_port, Q(17) => 
                           bus_reg_dataout_1105_port, Q(16) => 
                           bus_reg_dataout_1104_port, Q(15) => 
                           bus_reg_dataout_1103_port, Q(14) => 
                           bus_reg_dataout_1102_port, Q(13) => 
                           bus_reg_dataout_1101_port, Q(12) => 
                           bus_reg_dataout_1100_port, Q(11) => 
                           bus_reg_dataout_1099_port, Q(10) => 
                           bus_reg_dataout_1098_port, Q(9) => 
                           bus_reg_dataout_1097_port, Q(8) => 
                           bus_reg_dataout_1096_port, Q(7) => 
                           bus_reg_dataout_1095_port, Q(6) => 
                           bus_reg_dataout_1094_port, Q(5) => 
                           bus_reg_dataout_1093_port, Q(4) => 
                           bus_reg_dataout_1092_port, Q(3) => 
                           bus_reg_dataout_1091_port, Q(2) => 
                           bus_reg_dataout_1090_port, Q(1) => 
                           bus_reg_dataout_1089_port, Q(0) => 
                           bus_reg_dataout_1088_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_42_port);
   BLOCKi_43 : reg_generic_N32_RSTVAL0_45 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1151_port, Q(30) => 
                           bus_reg_dataout_1150_port, Q(29) => 
                           bus_reg_dataout_1149_port, Q(28) => 
                           bus_reg_dataout_1148_port, Q(27) => 
                           bus_reg_dataout_1147_port, Q(26) => 
                           bus_reg_dataout_1146_port, Q(25) => 
                           bus_reg_dataout_1145_port, Q(24) => 
                           bus_reg_dataout_1144_port, Q(23) => 
                           bus_reg_dataout_1143_port, Q(22) => 
                           bus_reg_dataout_1142_port, Q(21) => 
                           bus_reg_dataout_1141_port, Q(20) => 
                           bus_reg_dataout_1140_port, Q(19) => 
                           bus_reg_dataout_1139_port, Q(18) => 
                           bus_reg_dataout_1138_port, Q(17) => 
                           bus_reg_dataout_1137_port, Q(16) => 
                           bus_reg_dataout_1136_port, Q(15) => 
                           bus_reg_dataout_1135_port, Q(14) => 
                           bus_reg_dataout_1134_port, Q(13) => 
                           bus_reg_dataout_1133_port, Q(12) => 
                           bus_reg_dataout_1132_port, Q(11) => 
                           bus_reg_dataout_1131_port, Q(10) => 
                           bus_reg_dataout_1130_port, Q(9) => 
                           bus_reg_dataout_1129_port, Q(8) => 
                           bus_reg_dataout_1128_port, Q(7) => 
                           bus_reg_dataout_1127_port, Q(6) => 
                           bus_reg_dataout_1126_port, Q(5) => 
                           bus_reg_dataout_1125_port, Q(4) => 
                           bus_reg_dataout_1124_port, Q(3) => 
                           bus_reg_dataout_1123_port, Q(2) => 
                           bus_reg_dataout_1122_port, Q(1) => 
                           bus_reg_dataout_1121_port, Q(0) => 
                           bus_reg_dataout_1120_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_43_port);
   MUX_SELINPUT_44 : mux_N32_M1_22 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1108
                           , Y(30) => n1100, Y(29) => n1092, Y(28) => n1084, 
                           Y(27) => n1076, Y(26) => n1068, Y(25) => n1060, 
                           Y(24) => n1052, Y(23) => n1044, Y(22) => n1036, 
                           Y(21) => n1028, Y(20) => n1020, Y(19) => n1012, 
                           Y(18) => n1004, Y(17) => n996, Y(16) => n988, Y(15) 
                           => n980, Y(14) => n972, Y(13) => n964, Y(12) => n956
                           , Y(11) => n948, Y(10) => n940, Y(9) => n932, Y(8) 
                           => n924, Y(7) => n916, Y(6) => n908, Y(5) => n900, 
                           Y(4) => n892, Y(3) => n884, Y(2) => n876, Y(1) => 
                           n868, Y(0) => n860);
   BLOCKi_44 : reg_generic_N32_RSTVAL0_44 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1183_port, Q(30) => 
                           bus_reg_dataout_1182_port, Q(29) => 
                           bus_reg_dataout_1181_port, Q(28) => 
                           bus_reg_dataout_1180_port, Q(27) => 
                           bus_reg_dataout_1179_port, Q(26) => 
                           bus_reg_dataout_1178_port, Q(25) => 
                           bus_reg_dataout_1177_port, Q(24) => 
                           bus_reg_dataout_1176_port, Q(23) => 
                           bus_reg_dataout_1175_port, Q(22) => 
                           bus_reg_dataout_1174_port, Q(21) => 
                           bus_reg_dataout_1173_port, Q(20) => 
                           bus_reg_dataout_1172_port, Q(19) => 
                           bus_reg_dataout_1171_port, Q(18) => 
                           bus_reg_dataout_1170_port, Q(17) => 
                           bus_reg_dataout_1169_port, Q(16) => 
                           bus_reg_dataout_1168_port, Q(15) => 
                           bus_reg_dataout_1167_port, Q(14) => 
                           bus_reg_dataout_1166_port, Q(13) => 
                           bus_reg_dataout_1165_port, Q(12) => 
                           bus_reg_dataout_1164_port, Q(11) => 
                           bus_reg_dataout_1163_port, Q(10) => 
                           bus_reg_dataout_1162_port, Q(9) => 
                           bus_reg_dataout_1161_port, Q(8) => 
                           bus_reg_dataout_1160_port, Q(7) => 
                           bus_reg_dataout_1159_port, Q(6) => 
                           bus_reg_dataout_1158_port, Q(5) => 
                           bus_reg_dataout_1157_port, Q(4) => 
                           bus_reg_dataout_1156_port, Q(3) => 
                           bus_reg_dataout_1155_port, Q(2) => 
                           bus_reg_dataout_1154_port, Q(1) => 
                           bus_reg_dataout_1153_port, Q(0) => 
                           bus_reg_dataout_1152_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_44_port);
   BLOCKi_45 : reg_generic_N32_RSTVAL0_43 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1215_port, Q(30) => 
                           bus_reg_dataout_1214_port, Q(29) => 
                           bus_reg_dataout_1213_port, Q(28) => 
                           bus_reg_dataout_1212_port, Q(27) => 
                           bus_reg_dataout_1211_port, Q(26) => 
                           bus_reg_dataout_1210_port, Q(25) => 
                           bus_reg_dataout_1209_port, Q(24) => 
                           bus_reg_dataout_1208_port, Q(23) => 
                           bus_reg_dataout_1207_port, Q(22) => 
                           bus_reg_dataout_1206_port, Q(21) => 
                           bus_reg_dataout_1205_port, Q(20) => 
                           bus_reg_dataout_1204_port, Q(19) => 
                           bus_reg_dataout_1203_port, Q(18) => 
                           bus_reg_dataout_1202_port, Q(17) => 
                           bus_reg_dataout_1201_port, Q(16) => 
                           bus_reg_dataout_1200_port, Q(15) => 
                           bus_reg_dataout_1199_port, Q(14) => 
                           bus_reg_dataout_1198_port, Q(13) => 
                           bus_reg_dataout_1197_port, Q(12) => 
                           bus_reg_dataout_1196_port, Q(11) => 
                           bus_reg_dataout_1195_port, Q(10) => 
                           bus_reg_dataout_1194_port, Q(9) => 
                           bus_reg_dataout_1193_port, Q(8) => 
                           bus_reg_dataout_1192_port, Q(7) => 
                           bus_reg_dataout_1191_port, Q(6) => 
                           bus_reg_dataout_1190_port, Q(5) => 
                           bus_reg_dataout_1189_port, Q(4) => 
                           bus_reg_dataout_1188_port, Q(3) => 
                           bus_reg_dataout_1187_port, Q(2) => 
                           bus_reg_dataout_1186_port, Q(1) => 
                           bus_reg_dataout_1185_port, Q(0) => 
                           bus_reg_dataout_1184_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_45_port);
   MUX_SELINPUT_46 : mux_N32_M1_21 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1107
                           , Y(30) => n1099, Y(29) => n1091, Y(28) => n1083, 
                           Y(27) => n1075, Y(26) => n1067, Y(25) => n1059, 
                           Y(24) => n1051, Y(23) => n1043, Y(22) => n1035, 
                           Y(21) => n1027, Y(20) => n1019, Y(19) => n1011, 
                           Y(18) => n1003, Y(17) => n995, Y(16) => n987, Y(15) 
                           => n979, Y(14) => n971, Y(13) => n963, Y(12) => n955
                           , Y(11) => n947, Y(10) => n939, Y(9) => n931, Y(8) 
                           => n923, Y(7) => n915, Y(6) => n907, Y(5) => n899, 
                           Y(4) => n891, Y(3) => n883, Y(2) => n875, Y(1) => 
                           n867, Y(0) => n859);
   BLOCKi_46 : reg_generic_N32_RSTVAL0_42 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1247_port, Q(30) => 
                           bus_reg_dataout_1246_port, Q(29) => 
                           bus_reg_dataout_1245_port, Q(28) => 
                           bus_reg_dataout_1244_port, Q(27) => 
                           bus_reg_dataout_1243_port, Q(26) => 
                           bus_reg_dataout_1242_port, Q(25) => 
                           bus_reg_dataout_1241_port, Q(24) => 
                           bus_reg_dataout_1240_port, Q(23) => 
                           bus_reg_dataout_1239_port, Q(22) => 
                           bus_reg_dataout_1238_port, Q(21) => 
                           bus_reg_dataout_1237_port, Q(20) => 
                           bus_reg_dataout_1236_port, Q(19) => 
                           bus_reg_dataout_1235_port, Q(18) => 
                           bus_reg_dataout_1234_port, Q(17) => 
                           bus_reg_dataout_1233_port, Q(16) => 
                           bus_reg_dataout_1232_port, Q(15) => 
                           bus_reg_dataout_1231_port, Q(14) => 
                           bus_reg_dataout_1230_port, Q(13) => 
                           bus_reg_dataout_1229_port, Q(12) => 
                           bus_reg_dataout_1228_port, Q(11) => 
                           bus_reg_dataout_1227_port, Q(10) => 
                           bus_reg_dataout_1226_port, Q(9) => 
                           bus_reg_dataout_1225_port, Q(8) => 
                           bus_reg_dataout_1224_port, Q(7) => 
                           bus_reg_dataout_1223_port, Q(6) => 
                           bus_reg_dataout_1222_port, Q(5) => 
                           bus_reg_dataout_1221_port, Q(4) => 
                           bus_reg_dataout_1220_port, Q(3) => 
                           bus_reg_dataout_1219_port, Q(2) => 
                           bus_reg_dataout_1218_port, Q(1) => 
                           bus_reg_dataout_1217_port, Q(0) => 
                           bus_reg_dataout_1216_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_46_port);
   BLOCKi_47 : reg_generic_N32_RSTVAL0_41 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1279_port, Q(30) => 
                           bus_reg_dataout_1278_port, Q(29) => 
                           bus_reg_dataout_1277_port, Q(28) => 
                           bus_reg_dataout_1276_port, Q(27) => 
                           bus_reg_dataout_1275_port, Q(26) => 
                           bus_reg_dataout_1274_port, Q(25) => 
                           bus_reg_dataout_1273_port, Q(24) => 
                           bus_reg_dataout_1272_port, Q(23) => 
                           bus_reg_dataout_1271_port, Q(22) => 
                           bus_reg_dataout_1270_port, Q(21) => 
                           bus_reg_dataout_1269_port, Q(20) => 
                           bus_reg_dataout_1268_port, Q(19) => 
                           bus_reg_dataout_1267_port, Q(18) => 
                           bus_reg_dataout_1266_port, Q(17) => 
                           bus_reg_dataout_1265_port, Q(16) => 
                           bus_reg_dataout_1264_port, Q(15) => 
                           bus_reg_dataout_1263_port, Q(14) => 
                           bus_reg_dataout_1262_port, Q(13) => 
                           bus_reg_dataout_1261_port, Q(12) => 
                           bus_reg_dataout_1260_port, Q(11) => 
                           bus_reg_dataout_1259_port, Q(10) => 
                           bus_reg_dataout_1258_port, Q(9) => 
                           bus_reg_dataout_1257_port, Q(8) => 
                           bus_reg_dataout_1256_port, Q(7) => 
                           bus_reg_dataout_1255_port, Q(6) => 
                           bus_reg_dataout_1254_port, Q(5) => 
                           bus_reg_dataout_1253_port, Q(4) => 
                           bus_reg_dataout_1252_port, Q(3) => 
                           bus_reg_dataout_1251_port, Q(2) => 
                           bus_reg_dataout_1250_port, Q(1) => 
                           bus_reg_dataout_1249_port, Q(0) => 
                           bus_reg_dataout_1248_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_47_port);
   MUX_SELINPUT_48 : mux_N32_M1_20 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1106
                           , Y(30) => n1098, Y(29) => n1090, Y(28) => n1082, 
                           Y(27) => n1074, Y(26) => n1066, Y(25) => n1058, 
                           Y(24) => n1050, Y(23) => n1042, Y(22) => n1034, 
                           Y(21) => n1026, Y(20) => n1018, Y(19) => n1010, 
                           Y(18) => n1002, Y(17) => n994, Y(16) => n986, Y(15) 
                           => n978, Y(14) => n970, Y(13) => n962, Y(12) => n954
                           , Y(11) => n946, Y(10) => n938, Y(9) => n930, Y(8) 
                           => n922, Y(7) => n914, Y(6) => n906, Y(5) => n898, 
                           Y(4) => n890, Y(3) => n882, Y(2) => n874, Y(1) => 
                           n866, Y(0) => n858);
   BLOCKi_48 : reg_generic_N32_RSTVAL0_40 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1311_port, Q(30) => 
                           bus_reg_dataout_1310_port, Q(29) => 
                           bus_reg_dataout_1309_port, Q(28) => 
                           bus_reg_dataout_1308_port, Q(27) => 
                           bus_reg_dataout_1307_port, Q(26) => 
                           bus_reg_dataout_1306_port, Q(25) => 
                           bus_reg_dataout_1305_port, Q(24) => 
                           bus_reg_dataout_1304_port, Q(23) => 
                           bus_reg_dataout_1303_port, Q(22) => 
                           bus_reg_dataout_1302_port, Q(21) => 
                           bus_reg_dataout_1301_port, Q(20) => 
                           bus_reg_dataout_1300_port, Q(19) => 
                           bus_reg_dataout_1299_port, Q(18) => 
                           bus_reg_dataout_1298_port, Q(17) => 
                           bus_reg_dataout_1297_port, Q(16) => 
                           bus_reg_dataout_1296_port, Q(15) => 
                           bus_reg_dataout_1295_port, Q(14) => 
                           bus_reg_dataout_1294_port, Q(13) => 
                           bus_reg_dataout_1293_port, Q(12) => 
                           bus_reg_dataout_1292_port, Q(11) => 
                           bus_reg_dataout_1291_port, Q(10) => 
                           bus_reg_dataout_1290_port, Q(9) => 
                           bus_reg_dataout_1289_port, Q(8) => 
                           bus_reg_dataout_1288_port, Q(7) => 
                           bus_reg_dataout_1287_port, Q(6) => 
                           bus_reg_dataout_1286_port, Q(5) => 
                           bus_reg_dataout_1285_port, Q(4) => 
                           bus_reg_dataout_1284_port, Q(3) => 
                           bus_reg_dataout_1283_port, Q(2) => 
                           bus_reg_dataout_1282_port, Q(1) => 
                           bus_reg_dataout_1281_port, Q(0) => 
                           bus_reg_dataout_1280_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_48_port);
   BLOCKi_49 : reg_generic_N32_RSTVAL0_39 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1343_port, Q(30) => 
                           bus_reg_dataout_1342_port, Q(29) => 
                           bus_reg_dataout_1341_port, Q(28) => 
                           bus_reg_dataout_1340_port, Q(27) => 
                           bus_reg_dataout_1339_port, Q(26) => 
                           bus_reg_dataout_1338_port, Q(25) => 
                           bus_reg_dataout_1337_port, Q(24) => 
                           bus_reg_dataout_1336_port, Q(23) => 
                           bus_reg_dataout_1335_port, Q(22) => 
                           bus_reg_dataout_1334_port, Q(21) => 
                           bus_reg_dataout_1333_port, Q(20) => 
                           bus_reg_dataout_1332_port, Q(19) => 
                           bus_reg_dataout_1331_port, Q(18) => 
                           bus_reg_dataout_1330_port, Q(17) => 
                           bus_reg_dataout_1329_port, Q(16) => 
                           bus_reg_dataout_1328_port, Q(15) => 
                           bus_reg_dataout_1327_port, Q(14) => 
                           bus_reg_dataout_1326_port, Q(13) => 
                           bus_reg_dataout_1325_port, Q(12) => 
                           bus_reg_dataout_1324_port, Q(11) => 
                           bus_reg_dataout_1323_port, Q(10) => 
                           bus_reg_dataout_1322_port, Q(9) => 
                           bus_reg_dataout_1321_port, Q(8) => 
                           bus_reg_dataout_1320_port, Q(7) => 
                           bus_reg_dataout_1319_port, Q(6) => 
                           bus_reg_dataout_1318_port, Q(5) => 
                           bus_reg_dataout_1317_port, Q(4) => 
                           bus_reg_dataout_1316_port, Q(3) => 
                           bus_reg_dataout_1315_port, Q(2) => 
                           bus_reg_dataout_1314_port, Q(1) => 
                           bus_reg_dataout_1313_port, Q(0) => 
                           bus_reg_dataout_1312_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_49_port);
   MUX_SELINPUT_50 : mux_N32_M1_19 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1105
                           , Y(30) => n1097, Y(29) => n1089, Y(28) => n1081, 
                           Y(27) => n1073, Y(26) => n1065, Y(25) => n1057, 
                           Y(24) => n1049, Y(23) => n1041, Y(22) => n1033, 
                           Y(21) => n1025, Y(20) => n1017, Y(19) => n1009, 
                           Y(18) => n1001, Y(17) => n993, Y(16) => n985, Y(15) 
                           => n977, Y(14) => n969, Y(13) => n961, Y(12) => n953
                           , Y(11) => n945, Y(10) => n937, Y(9) => n929, Y(8) 
                           => n921, Y(7) => n913, Y(6) => n905, Y(5) => n897, 
                           Y(4) => n889, Y(3) => n881, Y(2) => n873, Y(1) => 
                           n865, Y(0) => n857);
   BLOCKi_50 : reg_generic_N32_RSTVAL0_38 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1375_port, Q(30) => 
                           bus_reg_dataout_1374_port, Q(29) => 
                           bus_reg_dataout_1373_port, Q(28) => 
                           bus_reg_dataout_1372_port, Q(27) => 
                           bus_reg_dataout_1371_port, Q(26) => 
                           bus_reg_dataout_1370_port, Q(25) => 
                           bus_reg_dataout_1369_port, Q(24) => 
                           bus_reg_dataout_1368_port, Q(23) => 
                           bus_reg_dataout_1367_port, Q(22) => 
                           bus_reg_dataout_1366_port, Q(21) => 
                           bus_reg_dataout_1365_port, Q(20) => 
                           bus_reg_dataout_1364_port, Q(19) => 
                           bus_reg_dataout_1363_port, Q(18) => 
                           bus_reg_dataout_1362_port, Q(17) => 
                           bus_reg_dataout_1361_port, Q(16) => 
                           bus_reg_dataout_1360_port, Q(15) => 
                           bus_reg_dataout_1359_port, Q(14) => 
                           bus_reg_dataout_1358_port, Q(13) => 
                           bus_reg_dataout_1357_port, Q(12) => 
                           bus_reg_dataout_1356_port, Q(11) => 
                           bus_reg_dataout_1355_port, Q(10) => 
                           bus_reg_dataout_1354_port, Q(9) => 
                           bus_reg_dataout_1353_port, Q(8) => 
                           bus_reg_dataout_1352_port, Q(7) => 
                           bus_reg_dataout_1351_port, Q(6) => 
                           bus_reg_dataout_1350_port, Q(5) => 
                           bus_reg_dataout_1349_port, Q(4) => 
                           bus_reg_dataout_1348_port, Q(3) => 
                           bus_reg_dataout_1347_port, Q(2) => 
                           bus_reg_dataout_1346_port, Q(1) => 
                           bus_reg_dataout_1345_port, Q(0) => 
                           bus_reg_dataout_1344_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_50_port);
   BLOCKi_51 : reg_generic_N32_RSTVAL0_37 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1407_port, Q(30) => 
                           bus_reg_dataout_1406_port, Q(29) => 
                           bus_reg_dataout_1405_port, Q(28) => 
                           bus_reg_dataout_1404_port, Q(27) => 
                           bus_reg_dataout_1403_port, Q(26) => 
                           bus_reg_dataout_1402_port, Q(25) => 
                           bus_reg_dataout_1401_port, Q(24) => 
                           bus_reg_dataout_1400_port, Q(23) => 
                           bus_reg_dataout_1399_port, Q(22) => 
                           bus_reg_dataout_1398_port, Q(21) => 
                           bus_reg_dataout_1397_port, Q(20) => 
                           bus_reg_dataout_1396_port, Q(19) => 
                           bus_reg_dataout_1395_port, Q(18) => 
                           bus_reg_dataout_1394_port, Q(17) => 
                           bus_reg_dataout_1393_port, Q(16) => 
                           bus_reg_dataout_1392_port, Q(15) => 
                           bus_reg_dataout_1391_port, Q(14) => 
                           bus_reg_dataout_1390_port, Q(13) => 
                           bus_reg_dataout_1389_port, Q(12) => 
                           bus_reg_dataout_1388_port, Q(11) => 
                           bus_reg_dataout_1387_port, Q(10) => 
                           bus_reg_dataout_1386_port, Q(9) => 
                           bus_reg_dataout_1385_port, Q(8) => 
                           bus_reg_dataout_1384_port, Q(7) => 
                           bus_reg_dataout_1383_port, Q(6) => 
                           bus_reg_dataout_1382_port, Q(5) => 
                           bus_reg_dataout_1381_port, Q(4) => 
                           bus_reg_dataout_1380_port, Q(3) => 
                           bus_reg_dataout_1379_port, Q(2) => 
                           bus_reg_dataout_1378_port, Q(1) => 
                           bus_reg_dataout_1377_port, Q(0) => 
                           bus_reg_dataout_1376_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_51_port);
   MUX_SELINPUT_52 : mux_N32_M1_18 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1104
                           , Y(30) => n1096, Y(29) => n1088, Y(28) => n1080, 
                           Y(27) => n1072, Y(26) => n1064, Y(25) => n1056, 
                           Y(24) => n1048, Y(23) => n1040, Y(22) => n1032, 
                           Y(21) => n1024, Y(20) => n1016, Y(19) => n1008, 
                           Y(18) => n1000, Y(17) => n992, Y(16) => n984, Y(15) 
                           => n976, Y(14) => n968, Y(13) => n960, Y(12) => n952
                           , Y(11) => n944, Y(10) => n936, Y(9) => n928, Y(8) 
                           => n920, Y(7) => n912, Y(6) => n904, Y(5) => n896, 
                           Y(4) => n888, Y(3) => n880, Y(2) => n872, Y(1) => 
                           n864, Y(0) => n856);
   BLOCKi_52 : reg_generic_N32_RSTVAL0_36 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1439_port, Q(30) => 
                           bus_reg_dataout_1438_port, Q(29) => 
                           bus_reg_dataout_1437_port, Q(28) => 
                           bus_reg_dataout_1436_port, Q(27) => 
                           bus_reg_dataout_1435_port, Q(26) => 
                           bus_reg_dataout_1434_port, Q(25) => 
                           bus_reg_dataout_1433_port, Q(24) => 
                           bus_reg_dataout_1432_port, Q(23) => 
                           bus_reg_dataout_1431_port, Q(22) => 
                           bus_reg_dataout_1430_port, Q(21) => 
                           bus_reg_dataout_1429_port, Q(20) => 
                           bus_reg_dataout_1428_port, Q(19) => 
                           bus_reg_dataout_1427_port, Q(18) => 
                           bus_reg_dataout_1426_port, Q(17) => 
                           bus_reg_dataout_1425_port, Q(16) => 
                           bus_reg_dataout_1424_port, Q(15) => 
                           bus_reg_dataout_1423_port, Q(14) => 
                           bus_reg_dataout_1422_port, Q(13) => 
                           bus_reg_dataout_1421_port, Q(12) => 
                           bus_reg_dataout_1420_port, Q(11) => 
                           bus_reg_dataout_1419_port, Q(10) => 
                           bus_reg_dataout_1418_port, Q(9) => 
                           bus_reg_dataout_1417_port, Q(8) => 
                           bus_reg_dataout_1416_port, Q(7) => 
                           bus_reg_dataout_1415_port, Q(6) => 
                           bus_reg_dataout_1414_port, Q(5) => 
                           bus_reg_dataout_1413_port, Q(4) => 
                           bus_reg_dataout_1412_port, Q(3) => 
                           bus_reg_dataout_1411_port, Q(2) => 
                           bus_reg_dataout_1410_port, Q(1) => 
                           bus_reg_dataout_1409_port, Q(0) => 
                           bus_reg_dataout_1408_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_52_port);
   BLOCKi_53 : reg_generic_N32_RSTVAL0_35 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1471_port, Q(30) => 
                           bus_reg_dataout_1470_port, Q(29) => 
                           bus_reg_dataout_1469_port, Q(28) => 
                           bus_reg_dataout_1468_port, Q(27) => 
                           bus_reg_dataout_1467_port, Q(26) => 
                           bus_reg_dataout_1466_port, Q(25) => 
                           bus_reg_dataout_1465_port, Q(24) => 
                           bus_reg_dataout_1464_port, Q(23) => 
                           bus_reg_dataout_1463_port, Q(22) => 
                           bus_reg_dataout_1462_port, Q(21) => 
                           bus_reg_dataout_1461_port, Q(20) => 
                           bus_reg_dataout_1460_port, Q(19) => 
                           bus_reg_dataout_1459_port, Q(18) => 
                           bus_reg_dataout_1458_port, Q(17) => 
                           bus_reg_dataout_1457_port, Q(16) => 
                           bus_reg_dataout_1456_port, Q(15) => 
                           bus_reg_dataout_1455_port, Q(14) => 
                           bus_reg_dataout_1454_port, Q(13) => 
                           bus_reg_dataout_1453_port, Q(12) => 
                           bus_reg_dataout_1452_port, Q(11) => 
                           bus_reg_dataout_1451_port, Q(10) => 
                           bus_reg_dataout_1450_port, Q(9) => 
                           bus_reg_dataout_1449_port, Q(8) => 
                           bus_reg_dataout_1448_port, Q(7) => 
                           bus_reg_dataout_1447_port, Q(6) => 
                           bus_reg_dataout_1446_port, Q(5) => 
                           bus_reg_dataout_1445_port, Q(4) => 
                           bus_reg_dataout_1444_port, Q(3) => 
                           bus_reg_dataout_1443_port, Q(2) => 
                           bus_reg_dataout_1442_port, Q(1) => 
                           bus_reg_dataout_1441_port, Q(0) => 
                           bus_reg_dataout_1440_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_53_port);
   MUX_SELINPUT_54 : mux_N32_M1_17 port map( S => c_swin_masked_1bit_2_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n1103
                           , Y(30) => n1095, Y(29) => n1087, Y(28) => n1079, 
                           Y(27) => n1071, Y(26) => n1063, Y(25) => n1055, 
                           Y(24) => n1047, Y(23) => n1039, Y(22) => n1031, 
                           Y(21) => n1023, Y(20) => n1015, Y(19) => n1007, 
                           Y(18) => n999, Y(17) => n991, Y(16) => n983, Y(15) 
                           => n975, Y(14) => n967, Y(13) => n959, Y(12) => n951
                           , Y(11) => n943, Y(10) => n935, Y(9) => n927, Y(8) 
                           => n919, Y(7) => n911, Y(6) => n903, Y(5) => n895, 
                           Y(4) => n887, Y(3) => n879, Y(2) => n871, Y(1) => 
                           n863, Y(0) => n855);
   BLOCKi_54 : reg_generic_N32_RSTVAL0_34 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1503_port, Q(30) => 
                           bus_reg_dataout_1502_port, Q(29) => 
                           bus_reg_dataout_1501_port, Q(28) => 
                           bus_reg_dataout_1500_port, Q(27) => 
                           bus_reg_dataout_1499_port, Q(26) => 
                           bus_reg_dataout_1498_port, Q(25) => 
                           bus_reg_dataout_1497_port, Q(24) => 
                           bus_reg_dataout_1496_port, Q(23) => 
                           bus_reg_dataout_1495_port, Q(22) => 
                           bus_reg_dataout_1494_port, Q(21) => 
                           bus_reg_dataout_1493_port, Q(20) => 
                           bus_reg_dataout_1492_port, Q(19) => 
                           bus_reg_dataout_1491_port, Q(18) => 
                           bus_reg_dataout_1490_port, Q(17) => 
                           bus_reg_dataout_1489_port, Q(16) => 
                           bus_reg_dataout_1488_port, Q(15) => 
                           bus_reg_dataout_1487_port, Q(14) => 
                           bus_reg_dataout_1486_port, Q(13) => 
                           bus_reg_dataout_1485_port, Q(12) => 
                           bus_reg_dataout_1484_port, Q(11) => 
                           bus_reg_dataout_1483_port, Q(10) => 
                           bus_reg_dataout_1482_port, Q(9) => 
                           bus_reg_dataout_1481_port, Q(8) => 
                           bus_reg_dataout_1480_port, Q(7) => 
                           bus_reg_dataout_1479_port, Q(6) => 
                           bus_reg_dataout_1478_port, Q(5) => 
                           bus_reg_dataout_1477_port, Q(4) => 
                           bus_reg_dataout_1476_port, Q(3) => 
                           bus_reg_dataout_1475_port, Q(2) => 
                           bus_reg_dataout_1474_port, Q(1) => 
                           bus_reg_dataout_1473_port, Q(0) => 
                           bus_reg_dataout_1472_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_54_port);
   BLOCKi_55 : reg_generic_N32_RSTVAL0_33 port map( D(31) => 
                           internal_inloc_data_2_31_port, D(30) => 
                           internal_inloc_data_2_30_port, D(29) => 
                           internal_inloc_data_2_29_port, D(28) => 
                           internal_inloc_data_2_28_port, D(27) => 
                           internal_inloc_data_2_27_port, D(26) => 
                           internal_inloc_data_2_26_port, D(25) => 
                           internal_inloc_data_2_25_port, D(24) => 
                           internal_inloc_data_2_24_port, D(23) => 
                           internal_inloc_data_2_23_port, D(22) => 
                           internal_inloc_data_2_22_port, D(21) => 
                           internal_inloc_data_2_21_port, D(20) => 
                           internal_inloc_data_2_20_port, D(19) => 
                           internal_inloc_data_2_19_port, D(18) => 
                           internal_inloc_data_2_18_port, D(17) => 
                           internal_inloc_data_2_17_port, D(16) => 
                           internal_inloc_data_2_16_port, D(15) => 
                           internal_inloc_data_2_15_port, D(14) => 
                           internal_inloc_data_2_14_port, D(13) => 
                           internal_inloc_data_2_13_port, D(12) => 
                           internal_inloc_data_2_12_port, D(11) => 
                           internal_inloc_data_2_11_port, D(10) => 
                           internal_inloc_data_2_10_port, D(9) => 
                           internal_inloc_data_2_9_port, D(8) => 
                           internal_inloc_data_2_8_port, D(7) => 
                           internal_inloc_data_2_7_port, D(6) => 
                           internal_inloc_data_2_6_port, D(5) => 
                           internal_inloc_data_2_5_port, D(4) => 
                           internal_inloc_data_2_4_port, D(3) => 
                           internal_inloc_data_2_3_port, D(2) => 
                           internal_inloc_data_2_2_port, D(1) => 
                           internal_inloc_data_2_1_port, D(0) => 
                           internal_inloc_data_2_0_port, Q(31) => 
                           bus_reg_dataout_1535_port, Q(30) => 
                           bus_reg_dataout_1534_port, Q(29) => 
                           bus_reg_dataout_1533_port, Q(28) => 
                           bus_reg_dataout_1532_port, Q(27) => 
                           bus_reg_dataout_1531_port, Q(26) => 
                           bus_reg_dataout_1530_port, Q(25) => 
                           bus_reg_dataout_1529_port, Q(24) => 
                           bus_reg_dataout_1528_port, Q(23) => 
                           bus_reg_dataout_1527_port, Q(22) => 
                           bus_reg_dataout_1526_port, Q(21) => 
                           bus_reg_dataout_1525_port, Q(20) => 
                           bus_reg_dataout_1524_port, Q(19) => 
                           bus_reg_dataout_1523_port, Q(18) => 
                           bus_reg_dataout_1522_port, Q(17) => 
                           bus_reg_dataout_1521_port, Q(16) => 
                           bus_reg_dataout_1520_port, Q(15) => 
                           bus_reg_dataout_1519_port, Q(14) => 
                           bus_reg_dataout_1518_port, Q(13) => 
                           bus_reg_dataout_1517_port, Q(12) => 
                           bus_reg_dataout_1516_port, Q(11) => 
                           bus_reg_dataout_1515_port, Q(10) => 
                           bus_reg_dataout_1514_port, Q(9) => 
                           bus_reg_dataout_1513_port, Q(8) => 
                           bus_reg_dataout_1512_port, Q(7) => 
                           bus_reg_dataout_1511_port, Q(6) => 
                           bus_reg_dataout_1510_port, Q(5) => 
                           bus_reg_dataout_1509_port, Q(4) => 
                           bus_reg_dataout_1508_port, Q(3) => 
                           bus_reg_dataout_1507_port, Q(2) => 
                           bus_reg_dataout_1506_port, Q(1) => 
                           bus_reg_dataout_1505_port, Q(0) => 
                           bus_reg_dataout_1504_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_55_port);
   MUX_SELINPUT_56 : mux_N32_M1_16 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n854,
                           Y(30) => n846, Y(29) => n838, Y(28) => n830, Y(27) 
                           => n822, Y(26) => n814, Y(25) => n806, Y(24) => n798
                           , Y(23) => n790, Y(22) => n782, Y(21) => n774, Y(20)
                           => n766, Y(19) => n758, Y(18) => n750, Y(17) => n742
                           , Y(16) => n734, Y(15) => n726, Y(14) => n718, Y(13)
                           => n710, Y(12) => n702, Y(11) => n694, Y(10) => n686
                           , Y(9) => n678, Y(8) => n670, Y(7) => n662, Y(6) => 
                           n654, Y(5) => n646, Y(4) => n638, Y(3) => n630, Y(2)
                           => n622, Y(1) => n614, Y(0) => n606);
   BLOCKi_56 : reg_generic_N32_RSTVAL0_32 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1567_port, Q(30) => 
                           bus_reg_dataout_1566_port, Q(29) => 
                           bus_reg_dataout_1565_port, Q(28) => 
                           bus_reg_dataout_1564_port, Q(27) => 
                           bus_reg_dataout_1563_port, Q(26) => 
                           bus_reg_dataout_1562_port, Q(25) => 
                           bus_reg_dataout_1561_port, Q(24) => 
                           bus_reg_dataout_1560_port, Q(23) => 
                           bus_reg_dataout_1559_port, Q(22) => 
                           bus_reg_dataout_1558_port, Q(21) => 
                           bus_reg_dataout_1557_port, Q(20) => 
                           bus_reg_dataout_1556_port, Q(19) => 
                           bus_reg_dataout_1555_port, Q(18) => 
                           bus_reg_dataout_1554_port, Q(17) => 
                           bus_reg_dataout_1553_port, Q(16) => 
                           bus_reg_dataout_1552_port, Q(15) => 
                           bus_reg_dataout_1551_port, Q(14) => 
                           bus_reg_dataout_1550_port, Q(13) => 
                           bus_reg_dataout_1549_port, Q(12) => 
                           bus_reg_dataout_1548_port, Q(11) => 
                           bus_reg_dataout_1547_port, Q(10) => 
                           bus_reg_dataout_1546_port, Q(9) => 
                           bus_reg_dataout_1545_port, Q(8) => 
                           bus_reg_dataout_1544_port, Q(7) => 
                           bus_reg_dataout_1543_port, Q(6) => 
                           bus_reg_dataout_1542_port, Q(5) => 
                           bus_reg_dataout_1541_port, Q(4) => 
                           bus_reg_dataout_1540_port, Q(3) => 
                           bus_reg_dataout_1539_port, Q(2) => 
                           bus_reg_dataout_1538_port, Q(1) => 
                           bus_reg_dataout_1537_port, Q(0) => 
                           bus_reg_dataout_1536_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_56_port);
   BLOCKi_57 : reg_generic_N32_RSTVAL0_31 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1599_port, Q(30) => 
                           bus_reg_dataout_1598_port, Q(29) => 
                           bus_reg_dataout_1597_port, Q(28) => 
                           bus_reg_dataout_1596_port, Q(27) => 
                           bus_reg_dataout_1595_port, Q(26) => 
                           bus_reg_dataout_1594_port, Q(25) => 
                           bus_reg_dataout_1593_port, Q(24) => 
                           bus_reg_dataout_1592_port, Q(23) => 
                           bus_reg_dataout_1591_port, Q(22) => 
                           bus_reg_dataout_1590_port, Q(21) => 
                           bus_reg_dataout_1589_port, Q(20) => 
                           bus_reg_dataout_1588_port, Q(19) => 
                           bus_reg_dataout_1587_port, Q(18) => 
                           bus_reg_dataout_1586_port, Q(17) => 
                           bus_reg_dataout_1585_port, Q(16) => 
                           bus_reg_dataout_1584_port, Q(15) => 
                           bus_reg_dataout_1583_port, Q(14) => 
                           bus_reg_dataout_1582_port, Q(13) => 
                           bus_reg_dataout_1581_port, Q(12) => 
                           bus_reg_dataout_1580_port, Q(11) => 
                           bus_reg_dataout_1579_port, Q(10) => 
                           bus_reg_dataout_1578_port, Q(9) => 
                           bus_reg_dataout_1577_port, Q(8) => 
                           bus_reg_dataout_1576_port, Q(7) => 
                           bus_reg_dataout_1575_port, Q(6) => 
                           bus_reg_dataout_1574_port, Q(5) => 
                           bus_reg_dataout_1573_port, Q(4) => 
                           bus_reg_dataout_1572_port, Q(3) => 
                           bus_reg_dataout_1571_port, Q(2) => 
                           bus_reg_dataout_1570_port, Q(1) => 
                           bus_reg_dataout_1569_port, Q(0) => 
                           bus_reg_dataout_1568_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_57_port);
   MUX_SELINPUT_58 : mux_N32_M1_15 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n853,
                           Y(30) => n845, Y(29) => n837, Y(28) => n829, Y(27) 
                           => n821, Y(26) => n813, Y(25) => n805, Y(24) => n797
                           , Y(23) => n789, Y(22) => n781, Y(21) => n773, Y(20)
                           => n765, Y(19) => n757, Y(18) => n749, Y(17) => n741
                           , Y(16) => n733, Y(15) => n725, Y(14) => n717, Y(13)
                           => n709, Y(12) => n701, Y(11) => n693, Y(10) => n685
                           , Y(9) => n677, Y(8) => n669, Y(7) => n661, Y(6) => 
                           n653, Y(5) => n645, Y(4) => n637, Y(3) => n629, Y(2)
                           => n621, Y(1) => n613, Y(0) => n605);
   BLOCKi_58 : reg_generic_N32_RSTVAL0_30 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1631_port, Q(30) => 
                           bus_reg_dataout_1630_port, Q(29) => 
                           bus_reg_dataout_1629_port, Q(28) => 
                           bus_reg_dataout_1628_port, Q(27) => 
                           bus_reg_dataout_1627_port, Q(26) => 
                           bus_reg_dataout_1626_port, Q(25) => 
                           bus_reg_dataout_1625_port, Q(24) => 
                           bus_reg_dataout_1624_port, Q(23) => 
                           bus_reg_dataout_1623_port, Q(22) => 
                           bus_reg_dataout_1622_port, Q(21) => 
                           bus_reg_dataout_1621_port, Q(20) => 
                           bus_reg_dataout_1620_port, Q(19) => 
                           bus_reg_dataout_1619_port, Q(18) => 
                           bus_reg_dataout_1618_port, Q(17) => 
                           bus_reg_dataout_1617_port, Q(16) => 
                           bus_reg_dataout_1616_port, Q(15) => 
                           bus_reg_dataout_1615_port, Q(14) => 
                           bus_reg_dataout_1614_port, Q(13) => 
                           bus_reg_dataout_1613_port, Q(12) => 
                           bus_reg_dataout_1612_port, Q(11) => 
                           bus_reg_dataout_1611_port, Q(10) => 
                           bus_reg_dataout_1610_port, Q(9) => 
                           bus_reg_dataout_1609_port, Q(8) => 
                           bus_reg_dataout_1608_port, Q(7) => 
                           bus_reg_dataout_1607_port, Q(6) => 
                           bus_reg_dataout_1606_port, Q(5) => 
                           bus_reg_dataout_1605_port, Q(4) => 
                           bus_reg_dataout_1604_port, Q(3) => 
                           bus_reg_dataout_1603_port, Q(2) => 
                           bus_reg_dataout_1602_port, Q(1) => 
                           bus_reg_dataout_1601_port, Q(0) => 
                           bus_reg_dataout_1600_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_58_port);
   BLOCKi_59 : reg_generic_N32_RSTVAL0_29 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1663_port, Q(30) => 
                           bus_reg_dataout_1662_port, Q(29) => 
                           bus_reg_dataout_1661_port, Q(28) => 
                           bus_reg_dataout_1660_port, Q(27) => 
                           bus_reg_dataout_1659_port, Q(26) => 
                           bus_reg_dataout_1658_port, Q(25) => 
                           bus_reg_dataout_1657_port, Q(24) => 
                           bus_reg_dataout_1656_port, Q(23) => 
                           bus_reg_dataout_1655_port, Q(22) => 
                           bus_reg_dataout_1654_port, Q(21) => 
                           bus_reg_dataout_1653_port, Q(20) => 
                           bus_reg_dataout_1652_port, Q(19) => 
                           bus_reg_dataout_1651_port, Q(18) => 
                           bus_reg_dataout_1650_port, Q(17) => 
                           bus_reg_dataout_1649_port, Q(16) => 
                           bus_reg_dataout_1648_port, Q(15) => 
                           bus_reg_dataout_1647_port, Q(14) => 
                           bus_reg_dataout_1646_port, Q(13) => 
                           bus_reg_dataout_1645_port, Q(12) => 
                           bus_reg_dataout_1644_port, Q(11) => 
                           bus_reg_dataout_1643_port, Q(10) => 
                           bus_reg_dataout_1642_port, Q(9) => 
                           bus_reg_dataout_1641_port, Q(8) => 
                           bus_reg_dataout_1640_port, Q(7) => 
                           bus_reg_dataout_1639_port, Q(6) => 
                           bus_reg_dataout_1638_port, Q(5) => 
                           bus_reg_dataout_1637_port, Q(4) => 
                           bus_reg_dataout_1636_port, Q(3) => 
                           bus_reg_dataout_1635_port, Q(2) => 
                           bus_reg_dataout_1634_port, Q(1) => 
                           bus_reg_dataout_1633_port, Q(0) => 
                           bus_reg_dataout_1632_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_59_port);
   MUX_SELINPUT_60 : mux_N32_M1_14 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n852,
                           Y(30) => n844, Y(29) => n836, Y(28) => n828, Y(27) 
                           => n820, Y(26) => n812, Y(25) => n804, Y(24) => n796
                           , Y(23) => n788, Y(22) => n780, Y(21) => n772, Y(20)
                           => n764, Y(19) => n756, Y(18) => n748, Y(17) => n740
                           , Y(16) => n732, Y(15) => n724, Y(14) => n716, Y(13)
                           => n708, Y(12) => n700, Y(11) => n692, Y(10) => n684
                           , Y(9) => n676, Y(8) => n668, Y(7) => n660, Y(6) => 
                           n652, Y(5) => n644, Y(4) => n636, Y(3) => n628, Y(2)
                           => n620, Y(1) => n612, Y(0) => n604);
   BLOCKi_60 : reg_generic_N32_RSTVAL0_28 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1695_port, Q(30) => 
                           bus_reg_dataout_1694_port, Q(29) => 
                           bus_reg_dataout_1693_port, Q(28) => 
                           bus_reg_dataout_1692_port, Q(27) => 
                           bus_reg_dataout_1691_port, Q(26) => 
                           bus_reg_dataout_1690_port, Q(25) => 
                           bus_reg_dataout_1689_port, Q(24) => 
                           bus_reg_dataout_1688_port, Q(23) => 
                           bus_reg_dataout_1687_port, Q(22) => 
                           bus_reg_dataout_1686_port, Q(21) => 
                           bus_reg_dataout_1685_port, Q(20) => 
                           bus_reg_dataout_1684_port, Q(19) => 
                           bus_reg_dataout_1683_port, Q(18) => 
                           bus_reg_dataout_1682_port, Q(17) => 
                           bus_reg_dataout_1681_port, Q(16) => 
                           bus_reg_dataout_1680_port, Q(15) => 
                           bus_reg_dataout_1679_port, Q(14) => 
                           bus_reg_dataout_1678_port, Q(13) => 
                           bus_reg_dataout_1677_port, Q(12) => 
                           bus_reg_dataout_1676_port, Q(11) => 
                           bus_reg_dataout_1675_port, Q(10) => 
                           bus_reg_dataout_1674_port, Q(9) => 
                           bus_reg_dataout_1673_port, Q(8) => 
                           bus_reg_dataout_1672_port, Q(7) => 
                           bus_reg_dataout_1671_port, Q(6) => 
                           bus_reg_dataout_1670_port, Q(5) => 
                           bus_reg_dataout_1669_port, Q(4) => 
                           bus_reg_dataout_1668_port, Q(3) => 
                           bus_reg_dataout_1667_port, Q(2) => 
                           bus_reg_dataout_1666_port, Q(1) => 
                           bus_reg_dataout_1665_port, Q(0) => 
                           bus_reg_dataout_1664_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_60_port);
   BLOCKi_61 : reg_generic_N32_RSTVAL0_27 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1727_port, Q(30) => 
                           bus_reg_dataout_1726_port, Q(29) => 
                           bus_reg_dataout_1725_port, Q(28) => 
                           bus_reg_dataout_1724_port, Q(27) => 
                           bus_reg_dataout_1723_port, Q(26) => 
                           bus_reg_dataout_1722_port, Q(25) => 
                           bus_reg_dataout_1721_port, Q(24) => 
                           bus_reg_dataout_1720_port, Q(23) => 
                           bus_reg_dataout_1719_port, Q(22) => 
                           bus_reg_dataout_1718_port, Q(21) => 
                           bus_reg_dataout_1717_port, Q(20) => 
                           bus_reg_dataout_1716_port, Q(19) => 
                           bus_reg_dataout_1715_port, Q(18) => 
                           bus_reg_dataout_1714_port, Q(17) => 
                           bus_reg_dataout_1713_port, Q(16) => 
                           bus_reg_dataout_1712_port, Q(15) => 
                           bus_reg_dataout_1711_port, Q(14) => 
                           bus_reg_dataout_1710_port, Q(13) => 
                           bus_reg_dataout_1709_port, Q(12) => 
                           bus_reg_dataout_1708_port, Q(11) => 
                           bus_reg_dataout_1707_port, Q(10) => 
                           bus_reg_dataout_1706_port, Q(9) => 
                           bus_reg_dataout_1705_port, Q(8) => 
                           bus_reg_dataout_1704_port, Q(7) => 
                           bus_reg_dataout_1703_port, Q(6) => 
                           bus_reg_dataout_1702_port, Q(5) => 
                           bus_reg_dataout_1701_port, Q(4) => 
                           bus_reg_dataout_1700_port, Q(3) => 
                           bus_reg_dataout_1699_port, Q(2) => 
                           bus_reg_dataout_1698_port, Q(1) => 
                           bus_reg_dataout_1697_port, Q(0) => 
                           bus_reg_dataout_1696_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_61_port);
   MUX_SELINPUT_62 : mux_N32_M1_13 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n851,
                           Y(30) => n843, Y(29) => n835, Y(28) => n827, Y(27) 
                           => n819, Y(26) => n811, Y(25) => n803, Y(24) => n795
                           , Y(23) => n787, Y(22) => n779, Y(21) => n771, Y(20)
                           => n763, Y(19) => n755, Y(18) => n747, Y(17) => n739
                           , Y(16) => n731, Y(15) => n723, Y(14) => n715, Y(13)
                           => n707, Y(12) => n699, Y(11) => n691, Y(10) => n683
                           , Y(9) => n675, Y(8) => n667, Y(7) => n659, Y(6) => 
                           n651, Y(5) => n643, Y(4) => n635, Y(3) => n627, Y(2)
                           => n619, Y(1) => n611, Y(0) => n603);
   BLOCKi_62 : reg_generic_N32_RSTVAL0_26 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1759_port, Q(30) => 
                           bus_reg_dataout_1758_port, Q(29) => 
                           bus_reg_dataout_1757_port, Q(28) => 
                           bus_reg_dataout_1756_port, Q(27) => 
                           bus_reg_dataout_1755_port, Q(26) => 
                           bus_reg_dataout_1754_port, Q(25) => 
                           bus_reg_dataout_1753_port, Q(24) => 
                           bus_reg_dataout_1752_port, Q(23) => 
                           bus_reg_dataout_1751_port, Q(22) => 
                           bus_reg_dataout_1750_port, Q(21) => 
                           bus_reg_dataout_1749_port, Q(20) => 
                           bus_reg_dataout_1748_port, Q(19) => 
                           bus_reg_dataout_1747_port, Q(18) => 
                           bus_reg_dataout_1746_port, Q(17) => 
                           bus_reg_dataout_1745_port, Q(16) => 
                           bus_reg_dataout_1744_port, Q(15) => 
                           bus_reg_dataout_1743_port, Q(14) => 
                           bus_reg_dataout_1742_port, Q(13) => 
                           bus_reg_dataout_1741_port, Q(12) => 
                           bus_reg_dataout_1740_port, Q(11) => 
                           bus_reg_dataout_1739_port, Q(10) => 
                           bus_reg_dataout_1738_port, Q(9) => 
                           bus_reg_dataout_1737_port, Q(8) => 
                           bus_reg_dataout_1736_port, Q(7) => 
                           bus_reg_dataout_1735_port, Q(6) => 
                           bus_reg_dataout_1734_port, Q(5) => 
                           bus_reg_dataout_1733_port, Q(4) => 
                           bus_reg_dataout_1732_port, Q(3) => 
                           bus_reg_dataout_1731_port, Q(2) => 
                           bus_reg_dataout_1730_port, Q(1) => 
                           bus_reg_dataout_1729_port, Q(0) => 
                           bus_reg_dataout_1728_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_62_port);
   BLOCKi_63 : reg_generic_N32_RSTVAL0_25 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1791_port, Q(30) => 
                           bus_reg_dataout_1790_port, Q(29) => 
                           bus_reg_dataout_1789_port, Q(28) => 
                           bus_reg_dataout_1788_port, Q(27) => 
                           bus_reg_dataout_1787_port, Q(26) => 
                           bus_reg_dataout_1786_port, Q(25) => 
                           bus_reg_dataout_1785_port, Q(24) => 
                           bus_reg_dataout_1784_port, Q(23) => 
                           bus_reg_dataout_1783_port, Q(22) => 
                           bus_reg_dataout_1782_port, Q(21) => 
                           bus_reg_dataout_1781_port, Q(20) => 
                           bus_reg_dataout_1780_port, Q(19) => 
                           bus_reg_dataout_1779_port, Q(18) => 
                           bus_reg_dataout_1778_port, Q(17) => 
                           bus_reg_dataout_1777_port, Q(16) => 
                           bus_reg_dataout_1776_port, Q(15) => 
                           bus_reg_dataout_1775_port, Q(14) => 
                           bus_reg_dataout_1774_port, Q(13) => 
                           bus_reg_dataout_1773_port, Q(12) => 
                           bus_reg_dataout_1772_port, Q(11) => 
                           bus_reg_dataout_1771_port, Q(10) => 
                           bus_reg_dataout_1770_port, Q(9) => 
                           bus_reg_dataout_1769_port, Q(8) => 
                           bus_reg_dataout_1768_port, Q(7) => 
                           bus_reg_dataout_1767_port, Q(6) => 
                           bus_reg_dataout_1766_port, Q(5) => 
                           bus_reg_dataout_1765_port, Q(4) => 
                           bus_reg_dataout_1764_port, Q(3) => 
                           bus_reg_dataout_1763_port, Q(2) => 
                           bus_reg_dataout_1762_port, Q(1) => 
                           bus_reg_dataout_1761_port, Q(0) => 
                           bus_reg_dataout_1760_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_63_port);
   MUX_SELINPUT_64 : mux_N32_M1_12 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n850,
                           Y(30) => n842, Y(29) => n834, Y(28) => n826, Y(27) 
                           => n818, Y(26) => n810, Y(25) => n802, Y(24) => n794
                           , Y(23) => n786, Y(22) => n778, Y(21) => n770, Y(20)
                           => n762, Y(19) => n754, Y(18) => n746, Y(17) => n738
                           , Y(16) => n730, Y(15) => n722, Y(14) => n714, Y(13)
                           => n706, Y(12) => n698, Y(11) => n690, Y(10) => n682
                           , Y(9) => n674, Y(8) => n666, Y(7) => n658, Y(6) => 
                           n650, Y(5) => n642, Y(4) => n634, Y(3) => n626, Y(2)
                           => n618, Y(1) => n610, Y(0) => n602);
   BLOCKi_64 : reg_generic_N32_RSTVAL0_24 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1823_port, Q(30) => 
                           bus_reg_dataout_1822_port, Q(29) => 
                           bus_reg_dataout_1821_port, Q(28) => 
                           bus_reg_dataout_1820_port, Q(27) => 
                           bus_reg_dataout_1819_port, Q(26) => 
                           bus_reg_dataout_1818_port, Q(25) => 
                           bus_reg_dataout_1817_port, Q(24) => 
                           bus_reg_dataout_1816_port, Q(23) => 
                           bus_reg_dataout_1815_port, Q(22) => 
                           bus_reg_dataout_1814_port, Q(21) => 
                           bus_reg_dataout_1813_port, Q(20) => 
                           bus_reg_dataout_1812_port, Q(19) => 
                           bus_reg_dataout_1811_port, Q(18) => 
                           bus_reg_dataout_1810_port, Q(17) => 
                           bus_reg_dataout_1809_port, Q(16) => 
                           bus_reg_dataout_1808_port, Q(15) => 
                           bus_reg_dataout_1807_port, Q(14) => 
                           bus_reg_dataout_1806_port, Q(13) => 
                           bus_reg_dataout_1805_port, Q(12) => 
                           bus_reg_dataout_1804_port, Q(11) => 
                           bus_reg_dataout_1803_port, Q(10) => 
                           bus_reg_dataout_1802_port, Q(9) => 
                           bus_reg_dataout_1801_port, Q(8) => 
                           bus_reg_dataout_1800_port, Q(7) => 
                           bus_reg_dataout_1799_port, Q(6) => 
                           bus_reg_dataout_1798_port, Q(5) => 
                           bus_reg_dataout_1797_port, Q(4) => 
                           bus_reg_dataout_1796_port, Q(3) => 
                           bus_reg_dataout_1795_port, Q(2) => 
                           bus_reg_dataout_1794_port, Q(1) => 
                           bus_reg_dataout_1793_port, Q(0) => 
                           bus_reg_dataout_1792_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_64_port);
   BLOCKi_65 : reg_generic_N32_RSTVAL0_23 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1855_port, Q(30) => 
                           bus_reg_dataout_1854_port, Q(29) => 
                           bus_reg_dataout_1853_port, Q(28) => 
                           bus_reg_dataout_1852_port, Q(27) => 
                           bus_reg_dataout_1851_port, Q(26) => 
                           bus_reg_dataout_1850_port, Q(25) => 
                           bus_reg_dataout_1849_port, Q(24) => 
                           bus_reg_dataout_1848_port, Q(23) => 
                           bus_reg_dataout_1847_port, Q(22) => 
                           bus_reg_dataout_1846_port, Q(21) => 
                           bus_reg_dataout_1845_port, Q(20) => 
                           bus_reg_dataout_1844_port, Q(19) => 
                           bus_reg_dataout_1843_port, Q(18) => 
                           bus_reg_dataout_1842_port, Q(17) => 
                           bus_reg_dataout_1841_port, Q(16) => 
                           bus_reg_dataout_1840_port, Q(15) => 
                           bus_reg_dataout_1839_port, Q(14) => 
                           bus_reg_dataout_1838_port, Q(13) => 
                           bus_reg_dataout_1837_port, Q(12) => 
                           bus_reg_dataout_1836_port, Q(11) => 
                           bus_reg_dataout_1835_port, Q(10) => 
                           bus_reg_dataout_1834_port, Q(9) => 
                           bus_reg_dataout_1833_port, Q(8) => 
                           bus_reg_dataout_1832_port, Q(7) => 
                           bus_reg_dataout_1831_port, Q(6) => 
                           bus_reg_dataout_1830_port, Q(5) => 
                           bus_reg_dataout_1829_port, Q(4) => 
                           bus_reg_dataout_1828_port, Q(3) => 
                           bus_reg_dataout_1827_port, Q(2) => 
                           bus_reg_dataout_1826_port, Q(1) => 
                           bus_reg_dataout_1825_port, Q(0) => 
                           bus_reg_dataout_1824_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_65_port);
   MUX_SELINPUT_66 : mux_N32_M1_11 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n849,
                           Y(30) => n841, Y(29) => n833, Y(28) => n825, Y(27) 
                           => n817, Y(26) => n809, Y(25) => n801, Y(24) => n793
                           , Y(23) => n785, Y(22) => n777, Y(21) => n769, Y(20)
                           => n761, Y(19) => n753, Y(18) => n745, Y(17) => n737
                           , Y(16) => n729, Y(15) => n721, Y(14) => n713, Y(13)
                           => n705, Y(12) => n697, Y(11) => n689, Y(10) => n681
                           , Y(9) => n673, Y(8) => n665, Y(7) => n657, Y(6) => 
                           n649, Y(5) => n641, Y(4) => n633, Y(3) => n625, Y(2)
                           => n617, Y(1) => n609, Y(0) => n601);
   BLOCKi_66 : reg_generic_N32_RSTVAL0_22 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1887_port, Q(30) => 
                           bus_reg_dataout_1886_port, Q(29) => 
                           bus_reg_dataout_1885_port, Q(28) => 
                           bus_reg_dataout_1884_port, Q(27) => 
                           bus_reg_dataout_1883_port, Q(26) => 
                           bus_reg_dataout_1882_port, Q(25) => 
                           bus_reg_dataout_1881_port, Q(24) => 
                           bus_reg_dataout_1880_port, Q(23) => 
                           bus_reg_dataout_1879_port, Q(22) => 
                           bus_reg_dataout_1878_port, Q(21) => 
                           bus_reg_dataout_1877_port, Q(20) => 
                           bus_reg_dataout_1876_port, Q(19) => 
                           bus_reg_dataout_1875_port, Q(18) => 
                           bus_reg_dataout_1874_port, Q(17) => 
                           bus_reg_dataout_1873_port, Q(16) => 
                           bus_reg_dataout_1872_port, Q(15) => 
                           bus_reg_dataout_1871_port, Q(14) => 
                           bus_reg_dataout_1870_port, Q(13) => 
                           bus_reg_dataout_1869_port, Q(12) => 
                           bus_reg_dataout_1868_port, Q(11) => 
                           bus_reg_dataout_1867_port, Q(10) => 
                           bus_reg_dataout_1866_port, Q(9) => 
                           bus_reg_dataout_1865_port, Q(8) => 
                           bus_reg_dataout_1864_port, Q(7) => 
                           bus_reg_dataout_1863_port, Q(6) => 
                           bus_reg_dataout_1862_port, Q(5) => 
                           bus_reg_dataout_1861_port, Q(4) => 
                           bus_reg_dataout_1860_port, Q(3) => 
                           bus_reg_dataout_1859_port, Q(2) => 
                           bus_reg_dataout_1858_port, Q(1) => 
                           bus_reg_dataout_1857_port, Q(0) => 
                           bus_reg_dataout_1856_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_66_port);
   BLOCKi_67 : reg_generic_N32_RSTVAL0_21 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1919_port, Q(30) => 
                           bus_reg_dataout_1918_port, Q(29) => 
                           bus_reg_dataout_1917_port, Q(28) => 
                           bus_reg_dataout_1916_port, Q(27) => 
                           bus_reg_dataout_1915_port, Q(26) => 
                           bus_reg_dataout_1914_port, Q(25) => 
                           bus_reg_dataout_1913_port, Q(24) => 
                           bus_reg_dataout_1912_port, Q(23) => 
                           bus_reg_dataout_1911_port, Q(22) => 
                           bus_reg_dataout_1910_port, Q(21) => 
                           bus_reg_dataout_1909_port, Q(20) => 
                           bus_reg_dataout_1908_port, Q(19) => 
                           bus_reg_dataout_1907_port, Q(18) => 
                           bus_reg_dataout_1906_port, Q(17) => 
                           bus_reg_dataout_1905_port, Q(16) => 
                           bus_reg_dataout_1904_port, Q(15) => 
                           bus_reg_dataout_1903_port, Q(14) => 
                           bus_reg_dataout_1902_port, Q(13) => 
                           bus_reg_dataout_1901_port, Q(12) => 
                           bus_reg_dataout_1900_port, Q(11) => 
                           bus_reg_dataout_1899_port, Q(10) => 
                           bus_reg_dataout_1898_port, Q(9) => 
                           bus_reg_dataout_1897_port, Q(8) => 
                           bus_reg_dataout_1896_port, Q(7) => 
                           bus_reg_dataout_1895_port, Q(6) => 
                           bus_reg_dataout_1894_port, Q(5) => 
                           bus_reg_dataout_1893_port, Q(4) => 
                           bus_reg_dataout_1892_port, Q(3) => 
                           bus_reg_dataout_1891_port, Q(2) => 
                           bus_reg_dataout_1890_port, Q(1) => 
                           bus_reg_dataout_1889_port, Q(0) => 
                           bus_reg_dataout_1888_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_67_port);
   MUX_SELINPUT_68 : mux_N32_M1_10 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n848,
                           Y(30) => n840, Y(29) => n832, Y(28) => n824, Y(27) 
                           => n816, Y(26) => n808, Y(25) => n800, Y(24) => n792
                           , Y(23) => n784, Y(22) => n776, Y(21) => n768, Y(20)
                           => n760, Y(19) => n752, Y(18) => n744, Y(17) => n736
                           , Y(16) => n728, Y(15) => n720, Y(14) => n712, Y(13)
                           => n704, Y(12) => n696, Y(11) => n688, Y(10) => n680
                           , Y(9) => n672, Y(8) => n664, Y(7) => n656, Y(6) => 
                           n648, Y(5) => n640, Y(4) => n632, Y(3) => n624, Y(2)
                           => n616, Y(1) => n608, Y(0) => n600);
   BLOCKi_68 : reg_generic_N32_RSTVAL0_20 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1951_port, Q(30) => 
                           bus_reg_dataout_1950_port, Q(29) => 
                           bus_reg_dataout_1949_port, Q(28) => 
                           bus_reg_dataout_1948_port, Q(27) => 
                           bus_reg_dataout_1947_port, Q(26) => 
                           bus_reg_dataout_1946_port, Q(25) => 
                           bus_reg_dataout_1945_port, Q(24) => 
                           bus_reg_dataout_1944_port, Q(23) => 
                           bus_reg_dataout_1943_port, Q(22) => 
                           bus_reg_dataout_1942_port, Q(21) => 
                           bus_reg_dataout_1941_port, Q(20) => 
                           bus_reg_dataout_1940_port, Q(19) => 
                           bus_reg_dataout_1939_port, Q(18) => 
                           bus_reg_dataout_1938_port, Q(17) => 
                           bus_reg_dataout_1937_port, Q(16) => 
                           bus_reg_dataout_1936_port, Q(15) => 
                           bus_reg_dataout_1935_port, Q(14) => 
                           bus_reg_dataout_1934_port, Q(13) => 
                           bus_reg_dataout_1933_port, Q(12) => 
                           bus_reg_dataout_1932_port, Q(11) => 
                           bus_reg_dataout_1931_port, Q(10) => 
                           bus_reg_dataout_1930_port, Q(9) => 
                           bus_reg_dataout_1929_port, Q(8) => 
                           bus_reg_dataout_1928_port, Q(7) => 
                           bus_reg_dataout_1927_port, Q(6) => 
                           bus_reg_dataout_1926_port, Q(5) => 
                           bus_reg_dataout_1925_port, Q(4) => 
                           bus_reg_dataout_1924_port, Q(3) => 
                           bus_reg_dataout_1923_port, Q(2) => 
                           bus_reg_dataout_1922_port, Q(1) => 
                           bus_reg_dataout_1921_port, Q(0) => 
                           bus_reg_dataout_1920_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_68_port);
   BLOCKi_69 : reg_generic_N32_RSTVAL0_19 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_1983_port, Q(30) => 
                           bus_reg_dataout_1982_port, Q(29) => 
                           bus_reg_dataout_1981_port, Q(28) => 
                           bus_reg_dataout_1980_port, Q(27) => 
                           bus_reg_dataout_1979_port, Q(26) => 
                           bus_reg_dataout_1978_port, Q(25) => 
                           bus_reg_dataout_1977_port, Q(24) => 
                           bus_reg_dataout_1976_port, Q(23) => 
                           bus_reg_dataout_1975_port, Q(22) => 
                           bus_reg_dataout_1974_port, Q(21) => 
                           bus_reg_dataout_1973_port, Q(20) => 
                           bus_reg_dataout_1972_port, Q(19) => 
                           bus_reg_dataout_1971_port, Q(18) => 
                           bus_reg_dataout_1970_port, Q(17) => 
                           bus_reg_dataout_1969_port, Q(16) => 
                           bus_reg_dataout_1968_port, Q(15) => 
                           bus_reg_dataout_1967_port, Q(14) => 
                           bus_reg_dataout_1966_port, Q(13) => 
                           bus_reg_dataout_1965_port, Q(12) => 
                           bus_reg_dataout_1964_port, Q(11) => 
                           bus_reg_dataout_1963_port, Q(10) => 
                           bus_reg_dataout_1962_port, Q(9) => 
                           bus_reg_dataout_1961_port, Q(8) => 
                           bus_reg_dataout_1960_port, Q(7) => 
                           bus_reg_dataout_1959_port, Q(6) => 
                           bus_reg_dataout_1958_port, Q(5) => 
                           bus_reg_dataout_1957_port, Q(4) => 
                           bus_reg_dataout_1956_port, Q(3) => 
                           bus_reg_dataout_1955_port, Q(2) => 
                           bus_reg_dataout_1954_port, Q(1) => 
                           bus_reg_dataout_1953_port, Q(0) => 
                           bus_reg_dataout_1952_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_69_port);
   MUX_SELINPUT_70 : mux_N32_M1_9 port map( S => c_swin_masked_1bit_3_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n847,
                           Y(30) => n839, Y(29) => n831, Y(28) => n823, Y(27) 
                           => n815, Y(26) => n807, Y(25) => n799, Y(24) => n791
                           , Y(23) => n783, Y(22) => n775, Y(21) => n767, Y(20)
                           => n759, Y(19) => n751, Y(18) => n743, Y(17) => n735
                           , Y(16) => n727, Y(15) => n719, Y(14) => n711, Y(13)
                           => n703, Y(12) => n695, Y(11) => n687, Y(10) => n679
                           , Y(9) => n671, Y(8) => n663, Y(7) => n655, Y(6) => 
                           n647, Y(5) => n639, Y(4) => n631, Y(3) => n623, Y(2)
                           => n615, Y(1) => n607, Y(0) => n599);
   BLOCKi_70 : reg_generic_N32_RSTVAL0_18 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_2015_port, Q(30) => 
                           bus_reg_dataout_2014_port, Q(29) => 
                           bus_reg_dataout_2013_port, Q(28) => 
                           bus_reg_dataout_2012_port, Q(27) => 
                           bus_reg_dataout_2011_port, Q(26) => 
                           bus_reg_dataout_2010_port, Q(25) => 
                           bus_reg_dataout_2009_port, Q(24) => 
                           bus_reg_dataout_2008_port, Q(23) => 
                           bus_reg_dataout_2007_port, Q(22) => 
                           bus_reg_dataout_2006_port, Q(21) => 
                           bus_reg_dataout_2005_port, Q(20) => 
                           bus_reg_dataout_2004_port, Q(19) => 
                           bus_reg_dataout_2003_port, Q(18) => 
                           bus_reg_dataout_2002_port, Q(17) => 
                           bus_reg_dataout_2001_port, Q(16) => 
                           bus_reg_dataout_2000_port, Q(15) => 
                           bus_reg_dataout_1999_port, Q(14) => 
                           bus_reg_dataout_1998_port, Q(13) => 
                           bus_reg_dataout_1997_port, Q(12) => 
                           bus_reg_dataout_1996_port, Q(11) => 
                           bus_reg_dataout_1995_port, Q(10) => 
                           bus_reg_dataout_1994_port, Q(9) => 
                           bus_reg_dataout_1993_port, Q(8) => 
                           bus_reg_dataout_1992_port, Q(7) => 
                           bus_reg_dataout_1991_port, Q(6) => 
                           bus_reg_dataout_1990_port, Q(5) => 
                           bus_reg_dataout_1989_port, Q(4) => 
                           bus_reg_dataout_1988_port, Q(3) => 
                           bus_reg_dataout_1987_port, Q(2) => 
                           bus_reg_dataout_1986_port, Q(1) => 
                           bus_reg_dataout_1985_port, Q(0) => 
                           bus_reg_dataout_1984_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_70_port);
   BLOCKi_71 : reg_generic_N32_RSTVAL0_17 port map( D(31) => 
                           internal_inloc_data_3_31_port, D(30) => 
                           internal_inloc_data_3_30_port, D(29) => 
                           internal_inloc_data_3_29_port, D(28) => 
                           internal_inloc_data_3_28_port, D(27) => 
                           internal_inloc_data_3_27_port, D(26) => 
                           internal_inloc_data_3_26_port, D(25) => 
                           internal_inloc_data_3_25_port, D(24) => 
                           internal_inloc_data_3_24_port, D(23) => 
                           internal_inloc_data_3_23_port, D(22) => 
                           internal_inloc_data_3_22_port, D(21) => 
                           internal_inloc_data_3_21_port, D(20) => 
                           internal_inloc_data_3_20_port, D(19) => 
                           internal_inloc_data_3_19_port, D(18) => 
                           internal_inloc_data_3_18_port, D(17) => 
                           internal_inloc_data_3_17_port, D(16) => 
                           internal_inloc_data_3_16_port, D(15) => 
                           internal_inloc_data_3_15_port, D(14) => 
                           internal_inloc_data_3_14_port, D(13) => 
                           internal_inloc_data_3_13_port, D(12) => 
                           internal_inloc_data_3_12_port, D(11) => 
                           internal_inloc_data_3_11_port, D(10) => 
                           internal_inloc_data_3_10_port, D(9) => 
                           internal_inloc_data_3_9_port, D(8) => 
                           internal_inloc_data_3_8_port, D(7) => 
                           internal_inloc_data_3_7_port, D(6) => 
                           internal_inloc_data_3_6_port, D(5) => 
                           internal_inloc_data_3_5_port, D(4) => 
                           internal_inloc_data_3_4_port, D(3) => 
                           internal_inloc_data_3_3_port, D(2) => 
                           internal_inloc_data_3_2_port, D(1) => 
                           internal_inloc_data_3_1_port, D(0) => 
                           internal_inloc_data_3_0_port, Q(31) => 
                           bus_reg_dataout_2047_port, Q(30) => 
                           bus_reg_dataout_2046_port, Q(29) => 
                           bus_reg_dataout_2045_port, Q(28) => 
                           bus_reg_dataout_2044_port, Q(27) => 
                           bus_reg_dataout_2043_port, Q(26) => 
                           bus_reg_dataout_2042_port, Q(25) => 
                           bus_reg_dataout_2041_port, Q(24) => 
                           bus_reg_dataout_2040_port, Q(23) => 
                           bus_reg_dataout_2039_port, Q(22) => 
                           bus_reg_dataout_2038_port, Q(21) => 
                           bus_reg_dataout_2037_port, Q(20) => 
                           bus_reg_dataout_2036_port, Q(19) => 
                           bus_reg_dataout_2035_port, Q(18) => 
                           bus_reg_dataout_2034_port, Q(17) => 
                           bus_reg_dataout_2033_port, Q(16) => 
                           bus_reg_dataout_2032_port, Q(15) => 
                           bus_reg_dataout_2031_port, Q(14) => 
                           bus_reg_dataout_2030_port, Q(13) => 
                           bus_reg_dataout_2029_port, Q(12) => 
                           bus_reg_dataout_2028_port, Q(11) => 
                           bus_reg_dataout_2027_port, Q(10) => 
                           bus_reg_dataout_2026_port, Q(9) => 
                           bus_reg_dataout_2025_port, Q(8) => 
                           bus_reg_dataout_2024_port, Q(7) => 
                           bus_reg_dataout_2023_port, Q(6) => 
                           bus_reg_dataout_2022_port, Q(5) => 
                           bus_reg_dataout_2021_port, Q(4) => 
                           bus_reg_dataout_2020_port, Q(3) => 
                           bus_reg_dataout_2019_port, Q(2) => 
                           bus_reg_dataout_2018_port, Q(1) => 
                           bus_reg_dataout_2017_port, Q(0) => 
                           bus_reg_dataout_2016_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_71_port);
   MUX_SELINPUT_72 : mux_N32_M1_8 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n598,
                           Y(30) => n590, Y(29) => n582, Y(28) => n574, Y(27) 
                           => n566, Y(26) => n558, Y(25) => n550, Y(24) => n542
                           , Y(23) => n534, Y(22) => n526, Y(21) => n518, Y(20)
                           => n510, Y(19) => n502, Y(18) => n494, Y(17) => n486
                           , Y(16) => n478, Y(15) => n470, Y(14) => n462, Y(13)
                           => n454, Y(12) => n446, Y(11) => n438, Y(10) => n430
                           , Y(9) => n422, Y(8) => n414, Y(7) => n406, Y(6) => 
                           n398, Y(5) => n390, Y(4) => n382, Y(3) => n374, Y(2)
                           => n366, Y(1) => n358, Y(0) => n350);
   BLOCKi_72 : reg_generic_N32_RSTVAL0_16 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2079_port, Q(30) => 
                           bus_reg_dataout_2078_port, Q(29) => 
                           bus_reg_dataout_2077_port, Q(28) => 
                           bus_reg_dataout_2076_port, Q(27) => 
                           bus_reg_dataout_2075_port, Q(26) => 
                           bus_reg_dataout_2074_port, Q(25) => 
                           bus_reg_dataout_2073_port, Q(24) => 
                           bus_reg_dataout_2072_port, Q(23) => 
                           bus_reg_dataout_2071_port, Q(22) => 
                           bus_reg_dataout_2070_port, Q(21) => 
                           bus_reg_dataout_2069_port, Q(20) => 
                           bus_reg_dataout_2068_port, Q(19) => 
                           bus_reg_dataout_2067_port, Q(18) => 
                           bus_reg_dataout_2066_port, Q(17) => 
                           bus_reg_dataout_2065_port, Q(16) => 
                           bus_reg_dataout_2064_port, Q(15) => 
                           bus_reg_dataout_2063_port, Q(14) => 
                           bus_reg_dataout_2062_port, Q(13) => 
                           bus_reg_dataout_2061_port, Q(12) => 
                           bus_reg_dataout_2060_port, Q(11) => 
                           bus_reg_dataout_2059_port, Q(10) => 
                           bus_reg_dataout_2058_port, Q(9) => 
                           bus_reg_dataout_2057_port, Q(8) => 
                           bus_reg_dataout_2056_port, Q(7) => 
                           bus_reg_dataout_2055_port, Q(6) => 
                           bus_reg_dataout_2054_port, Q(5) => 
                           bus_reg_dataout_2053_port, Q(4) => 
                           bus_reg_dataout_2052_port, Q(3) => 
                           bus_reg_dataout_2051_port, Q(2) => 
                           bus_reg_dataout_2050_port, Q(1) => 
                           bus_reg_dataout_2049_port, Q(0) => 
                           bus_reg_dataout_2048_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_72_port);
   BLOCKi_73 : reg_generic_N32_RSTVAL0_15 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2111_port, Q(30) => 
                           bus_reg_dataout_2110_port, Q(29) => 
                           bus_reg_dataout_2109_port, Q(28) => 
                           bus_reg_dataout_2108_port, Q(27) => 
                           bus_reg_dataout_2107_port, Q(26) => 
                           bus_reg_dataout_2106_port, Q(25) => 
                           bus_reg_dataout_2105_port, Q(24) => 
                           bus_reg_dataout_2104_port, Q(23) => 
                           bus_reg_dataout_2103_port, Q(22) => 
                           bus_reg_dataout_2102_port, Q(21) => 
                           bus_reg_dataout_2101_port, Q(20) => 
                           bus_reg_dataout_2100_port, Q(19) => 
                           bus_reg_dataout_2099_port, Q(18) => 
                           bus_reg_dataout_2098_port, Q(17) => 
                           bus_reg_dataout_2097_port, Q(16) => 
                           bus_reg_dataout_2096_port, Q(15) => 
                           bus_reg_dataout_2095_port, Q(14) => 
                           bus_reg_dataout_2094_port, Q(13) => 
                           bus_reg_dataout_2093_port, Q(12) => 
                           bus_reg_dataout_2092_port, Q(11) => 
                           bus_reg_dataout_2091_port, Q(10) => 
                           bus_reg_dataout_2090_port, Q(9) => 
                           bus_reg_dataout_2089_port, Q(8) => 
                           bus_reg_dataout_2088_port, Q(7) => 
                           bus_reg_dataout_2087_port, Q(6) => 
                           bus_reg_dataout_2086_port, Q(5) => 
                           bus_reg_dataout_2085_port, Q(4) => 
                           bus_reg_dataout_2084_port, Q(3) => 
                           bus_reg_dataout_2083_port, Q(2) => 
                           bus_reg_dataout_2082_port, Q(1) => 
                           bus_reg_dataout_2081_port, Q(0) => 
                           bus_reg_dataout_2080_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_73_port);
   MUX_SELINPUT_74 : mux_N32_M1_7 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n597,
                           Y(30) => n589, Y(29) => n581, Y(28) => n573, Y(27) 
                           => n565, Y(26) => n557, Y(25) => n549, Y(24) => n541
                           , Y(23) => n533, Y(22) => n525, Y(21) => n517, Y(20)
                           => n509, Y(19) => n501, Y(18) => n493, Y(17) => n485
                           , Y(16) => n477, Y(15) => n469, Y(14) => n461, Y(13)
                           => n453, Y(12) => n445, Y(11) => n437, Y(10) => n429
                           , Y(9) => n421, Y(8) => n413, Y(7) => n405, Y(6) => 
                           n397, Y(5) => n389, Y(4) => n381, Y(3) => n373, Y(2)
                           => n365, Y(1) => n357, Y(0) => n349);
   BLOCKi_74 : reg_generic_N32_RSTVAL0_14 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2143_port, Q(30) => 
                           bus_reg_dataout_2142_port, Q(29) => 
                           bus_reg_dataout_2141_port, Q(28) => 
                           bus_reg_dataout_2140_port, Q(27) => 
                           bus_reg_dataout_2139_port, Q(26) => 
                           bus_reg_dataout_2138_port, Q(25) => 
                           bus_reg_dataout_2137_port, Q(24) => 
                           bus_reg_dataout_2136_port, Q(23) => 
                           bus_reg_dataout_2135_port, Q(22) => 
                           bus_reg_dataout_2134_port, Q(21) => 
                           bus_reg_dataout_2133_port, Q(20) => 
                           bus_reg_dataout_2132_port, Q(19) => 
                           bus_reg_dataout_2131_port, Q(18) => 
                           bus_reg_dataout_2130_port, Q(17) => 
                           bus_reg_dataout_2129_port, Q(16) => 
                           bus_reg_dataout_2128_port, Q(15) => 
                           bus_reg_dataout_2127_port, Q(14) => 
                           bus_reg_dataout_2126_port, Q(13) => 
                           bus_reg_dataout_2125_port, Q(12) => 
                           bus_reg_dataout_2124_port, Q(11) => 
                           bus_reg_dataout_2123_port, Q(10) => 
                           bus_reg_dataout_2122_port, Q(9) => 
                           bus_reg_dataout_2121_port, Q(8) => 
                           bus_reg_dataout_2120_port, Q(7) => 
                           bus_reg_dataout_2119_port, Q(6) => 
                           bus_reg_dataout_2118_port, Q(5) => 
                           bus_reg_dataout_2117_port, Q(4) => 
                           bus_reg_dataout_2116_port, Q(3) => 
                           bus_reg_dataout_2115_port, Q(2) => 
                           bus_reg_dataout_2114_port, Q(1) => 
                           bus_reg_dataout_2113_port, Q(0) => 
                           bus_reg_dataout_2112_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_74_port);
   BLOCKi_75 : reg_generic_N32_RSTVAL0_13 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2175_port, Q(30) => 
                           bus_reg_dataout_2174_port, Q(29) => 
                           bus_reg_dataout_2173_port, Q(28) => 
                           bus_reg_dataout_2172_port, Q(27) => 
                           bus_reg_dataout_2171_port, Q(26) => 
                           bus_reg_dataout_2170_port, Q(25) => 
                           bus_reg_dataout_2169_port, Q(24) => 
                           bus_reg_dataout_2168_port, Q(23) => 
                           bus_reg_dataout_2167_port, Q(22) => 
                           bus_reg_dataout_2166_port, Q(21) => 
                           bus_reg_dataout_2165_port, Q(20) => 
                           bus_reg_dataout_2164_port, Q(19) => 
                           bus_reg_dataout_2163_port, Q(18) => 
                           bus_reg_dataout_2162_port, Q(17) => 
                           bus_reg_dataout_2161_port, Q(16) => 
                           bus_reg_dataout_2160_port, Q(15) => 
                           bus_reg_dataout_2159_port, Q(14) => 
                           bus_reg_dataout_2158_port, Q(13) => 
                           bus_reg_dataout_2157_port, Q(12) => 
                           bus_reg_dataout_2156_port, Q(11) => 
                           bus_reg_dataout_2155_port, Q(10) => 
                           bus_reg_dataout_2154_port, Q(9) => 
                           bus_reg_dataout_2153_port, Q(8) => 
                           bus_reg_dataout_2152_port, Q(7) => 
                           bus_reg_dataout_2151_port, Q(6) => 
                           bus_reg_dataout_2150_port, Q(5) => 
                           bus_reg_dataout_2149_port, Q(4) => 
                           bus_reg_dataout_2148_port, Q(3) => 
                           bus_reg_dataout_2147_port, Q(2) => 
                           bus_reg_dataout_2146_port, Q(1) => 
                           bus_reg_dataout_2145_port, Q(0) => 
                           bus_reg_dataout_2144_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_75_port);
   MUX_SELINPUT_76 : mux_N32_M1_6 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n596,
                           Y(30) => n588, Y(29) => n580, Y(28) => n572, Y(27) 
                           => n564, Y(26) => n556, Y(25) => n548, Y(24) => n540
                           , Y(23) => n532, Y(22) => n524, Y(21) => n516, Y(20)
                           => n508, Y(19) => n500, Y(18) => n492, Y(17) => n484
                           , Y(16) => n476, Y(15) => n468, Y(14) => n460, Y(13)
                           => n452, Y(12) => n444, Y(11) => n436, Y(10) => n428
                           , Y(9) => n420, Y(8) => n412, Y(7) => n404, Y(6) => 
                           n396, Y(5) => n388, Y(4) => n380, Y(3) => n372, Y(2)
                           => n364, Y(1) => n356, Y(0) => n348);
   BLOCKi_76 : reg_generic_N32_RSTVAL0_12 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2207_port, Q(30) => 
                           bus_reg_dataout_2206_port, Q(29) => 
                           bus_reg_dataout_2205_port, Q(28) => 
                           bus_reg_dataout_2204_port, Q(27) => 
                           bus_reg_dataout_2203_port, Q(26) => 
                           bus_reg_dataout_2202_port, Q(25) => 
                           bus_reg_dataout_2201_port, Q(24) => 
                           bus_reg_dataout_2200_port, Q(23) => 
                           bus_reg_dataout_2199_port, Q(22) => 
                           bus_reg_dataout_2198_port, Q(21) => 
                           bus_reg_dataout_2197_port, Q(20) => 
                           bus_reg_dataout_2196_port, Q(19) => 
                           bus_reg_dataout_2195_port, Q(18) => 
                           bus_reg_dataout_2194_port, Q(17) => 
                           bus_reg_dataout_2193_port, Q(16) => 
                           bus_reg_dataout_2192_port, Q(15) => 
                           bus_reg_dataout_2191_port, Q(14) => 
                           bus_reg_dataout_2190_port, Q(13) => 
                           bus_reg_dataout_2189_port, Q(12) => 
                           bus_reg_dataout_2188_port, Q(11) => 
                           bus_reg_dataout_2187_port, Q(10) => 
                           bus_reg_dataout_2186_port, Q(9) => 
                           bus_reg_dataout_2185_port, Q(8) => 
                           bus_reg_dataout_2184_port, Q(7) => 
                           bus_reg_dataout_2183_port, Q(6) => 
                           bus_reg_dataout_2182_port, Q(5) => 
                           bus_reg_dataout_2181_port, Q(4) => 
                           bus_reg_dataout_2180_port, Q(3) => 
                           bus_reg_dataout_2179_port, Q(2) => 
                           bus_reg_dataout_2178_port, Q(1) => 
                           bus_reg_dataout_2177_port, Q(0) => 
                           bus_reg_dataout_2176_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_76_port);
   BLOCKi_77 : reg_generic_N32_RSTVAL0_11 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2239_port, Q(30) => 
                           bus_reg_dataout_2238_port, Q(29) => 
                           bus_reg_dataout_2237_port, Q(28) => 
                           bus_reg_dataout_2236_port, Q(27) => 
                           bus_reg_dataout_2235_port, Q(26) => 
                           bus_reg_dataout_2234_port, Q(25) => 
                           bus_reg_dataout_2233_port, Q(24) => 
                           bus_reg_dataout_2232_port, Q(23) => 
                           bus_reg_dataout_2231_port, Q(22) => 
                           bus_reg_dataout_2230_port, Q(21) => 
                           bus_reg_dataout_2229_port, Q(20) => 
                           bus_reg_dataout_2228_port, Q(19) => 
                           bus_reg_dataout_2227_port, Q(18) => 
                           bus_reg_dataout_2226_port, Q(17) => 
                           bus_reg_dataout_2225_port, Q(16) => 
                           bus_reg_dataout_2224_port, Q(15) => 
                           bus_reg_dataout_2223_port, Q(14) => 
                           bus_reg_dataout_2222_port, Q(13) => 
                           bus_reg_dataout_2221_port, Q(12) => 
                           bus_reg_dataout_2220_port, Q(11) => 
                           bus_reg_dataout_2219_port, Q(10) => 
                           bus_reg_dataout_2218_port, Q(9) => 
                           bus_reg_dataout_2217_port, Q(8) => 
                           bus_reg_dataout_2216_port, Q(7) => 
                           bus_reg_dataout_2215_port, Q(6) => 
                           bus_reg_dataout_2214_port, Q(5) => 
                           bus_reg_dataout_2213_port, Q(4) => 
                           bus_reg_dataout_2212_port, Q(3) => 
                           bus_reg_dataout_2211_port, Q(2) => 
                           bus_reg_dataout_2210_port, Q(1) => 
                           bus_reg_dataout_2209_port, Q(0) => 
                           bus_reg_dataout_2208_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_77_port);
   MUX_SELINPUT_78 : mux_N32_M1_5 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n595,
                           Y(30) => n587, Y(29) => n579, Y(28) => n571, Y(27) 
                           => n563, Y(26) => n555, Y(25) => n547, Y(24) => n539
                           , Y(23) => n531, Y(22) => n523, Y(21) => n515, Y(20)
                           => n507, Y(19) => n499, Y(18) => n491, Y(17) => n483
                           , Y(16) => n475, Y(15) => n467, Y(14) => n459, Y(13)
                           => n451, Y(12) => n443, Y(11) => n435, Y(10) => n427
                           , Y(9) => n419, Y(8) => n411, Y(7) => n403, Y(6) => 
                           n395, Y(5) => n387, Y(4) => n379, Y(3) => n371, Y(2)
                           => n363, Y(1) => n355, Y(0) => n347);
   BLOCKi_78 : reg_generic_N32_RSTVAL0_10 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2271_port, Q(30) => 
                           bus_reg_dataout_2270_port, Q(29) => 
                           bus_reg_dataout_2269_port, Q(28) => 
                           bus_reg_dataout_2268_port, Q(27) => 
                           bus_reg_dataout_2267_port, Q(26) => 
                           bus_reg_dataout_2266_port, Q(25) => 
                           bus_reg_dataout_2265_port, Q(24) => 
                           bus_reg_dataout_2264_port, Q(23) => 
                           bus_reg_dataout_2263_port, Q(22) => 
                           bus_reg_dataout_2262_port, Q(21) => 
                           bus_reg_dataout_2261_port, Q(20) => 
                           bus_reg_dataout_2260_port, Q(19) => 
                           bus_reg_dataout_2259_port, Q(18) => 
                           bus_reg_dataout_2258_port, Q(17) => 
                           bus_reg_dataout_2257_port, Q(16) => 
                           bus_reg_dataout_2256_port, Q(15) => 
                           bus_reg_dataout_2255_port, Q(14) => 
                           bus_reg_dataout_2254_port, Q(13) => 
                           bus_reg_dataout_2253_port, Q(12) => 
                           bus_reg_dataout_2252_port, Q(11) => 
                           bus_reg_dataout_2251_port, Q(10) => 
                           bus_reg_dataout_2250_port, Q(9) => 
                           bus_reg_dataout_2249_port, Q(8) => 
                           bus_reg_dataout_2248_port, Q(7) => 
                           bus_reg_dataout_2247_port, Q(6) => 
                           bus_reg_dataout_2246_port, Q(5) => 
                           bus_reg_dataout_2245_port, Q(4) => 
                           bus_reg_dataout_2244_port, Q(3) => 
                           bus_reg_dataout_2243_port, Q(2) => 
                           bus_reg_dataout_2242_port, Q(1) => 
                           bus_reg_dataout_2241_port, Q(0) => 
                           bus_reg_dataout_2240_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_78_port);
   BLOCKi_79 : reg_generic_N32_RSTVAL0_9 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2303_port, Q(30) => 
                           bus_reg_dataout_2302_port, Q(29) => 
                           bus_reg_dataout_2301_port, Q(28) => 
                           bus_reg_dataout_2300_port, Q(27) => 
                           bus_reg_dataout_2299_port, Q(26) => 
                           bus_reg_dataout_2298_port, Q(25) => 
                           bus_reg_dataout_2297_port, Q(24) => 
                           bus_reg_dataout_2296_port, Q(23) => 
                           bus_reg_dataout_2295_port, Q(22) => 
                           bus_reg_dataout_2294_port, Q(21) => 
                           bus_reg_dataout_2293_port, Q(20) => 
                           bus_reg_dataout_2292_port, Q(19) => 
                           bus_reg_dataout_2291_port, Q(18) => 
                           bus_reg_dataout_2290_port, Q(17) => 
                           bus_reg_dataout_2289_port, Q(16) => 
                           bus_reg_dataout_2288_port, Q(15) => 
                           bus_reg_dataout_2287_port, Q(14) => 
                           bus_reg_dataout_2286_port, Q(13) => 
                           bus_reg_dataout_2285_port, Q(12) => 
                           bus_reg_dataout_2284_port, Q(11) => 
                           bus_reg_dataout_2283_port, Q(10) => 
                           bus_reg_dataout_2282_port, Q(9) => 
                           bus_reg_dataout_2281_port, Q(8) => 
                           bus_reg_dataout_2280_port, Q(7) => 
                           bus_reg_dataout_2279_port, Q(6) => 
                           bus_reg_dataout_2278_port, Q(5) => 
                           bus_reg_dataout_2277_port, Q(4) => 
                           bus_reg_dataout_2276_port, Q(3) => 
                           bus_reg_dataout_2275_port, Q(2) => 
                           bus_reg_dataout_2274_port, Q(1) => 
                           bus_reg_dataout_2273_port, Q(0) => 
                           bus_reg_dataout_2272_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_79_port);
   MUX_SELINPUT_80 : mux_N32_M1_4 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n594,
                           Y(30) => n586, Y(29) => n578, Y(28) => n570, Y(27) 
                           => n562, Y(26) => n554, Y(25) => n546, Y(24) => n538
                           , Y(23) => n530, Y(22) => n522, Y(21) => n514, Y(20)
                           => n506, Y(19) => n498, Y(18) => n490, Y(17) => n482
                           , Y(16) => n474, Y(15) => n466, Y(14) => n458, Y(13)
                           => n450, Y(12) => n442, Y(11) => n434, Y(10) => n426
                           , Y(9) => n418, Y(8) => n410, Y(7) => n402, Y(6) => 
                           n394, Y(5) => n386, Y(4) => n378, Y(3) => n370, Y(2)
                           => n362, Y(1) => n354, Y(0) => n346);
   BLOCKi_80 : reg_generic_N32_RSTVAL0_8 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2335_port, Q(30) => 
                           bus_reg_dataout_2334_port, Q(29) => 
                           bus_reg_dataout_2333_port, Q(28) => 
                           bus_reg_dataout_2332_port, Q(27) => 
                           bus_reg_dataout_2331_port, Q(26) => 
                           bus_reg_dataout_2330_port, Q(25) => 
                           bus_reg_dataout_2329_port, Q(24) => 
                           bus_reg_dataout_2328_port, Q(23) => 
                           bus_reg_dataout_2327_port, Q(22) => 
                           bus_reg_dataout_2326_port, Q(21) => 
                           bus_reg_dataout_2325_port, Q(20) => 
                           bus_reg_dataout_2324_port, Q(19) => 
                           bus_reg_dataout_2323_port, Q(18) => 
                           bus_reg_dataout_2322_port, Q(17) => 
                           bus_reg_dataout_2321_port, Q(16) => 
                           bus_reg_dataout_2320_port, Q(15) => 
                           bus_reg_dataout_2319_port, Q(14) => 
                           bus_reg_dataout_2318_port, Q(13) => 
                           bus_reg_dataout_2317_port, Q(12) => 
                           bus_reg_dataout_2316_port, Q(11) => 
                           bus_reg_dataout_2315_port, Q(10) => 
                           bus_reg_dataout_2314_port, Q(9) => 
                           bus_reg_dataout_2313_port, Q(8) => 
                           bus_reg_dataout_2312_port, Q(7) => 
                           bus_reg_dataout_2311_port, Q(6) => 
                           bus_reg_dataout_2310_port, Q(5) => 
                           bus_reg_dataout_2309_port, Q(4) => 
                           bus_reg_dataout_2308_port, Q(3) => 
                           bus_reg_dataout_2307_port, Q(2) => 
                           bus_reg_dataout_2306_port, Q(1) => 
                           bus_reg_dataout_2305_port, Q(0) => 
                           bus_reg_dataout_2304_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_80_port);
   BLOCKi_81 : reg_generic_N32_RSTVAL0_7 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2367_port, Q(30) => 
                           bus_reg_dataout_2366_port, Q(29) => 
                           bus_reg_dataout_2365_port, Q(28) => 
                           bus_reg_dataout_2364_port, Q(27) => 
                           bus_reg_dataout_2363_port, Q(26) => 
                           bus_reg_dataout_2362_port, Q(25) => 
                           bus_reg_dataout_2361_port, Q(24) => 
                           bus_reg_dataout_2360_port, Q(23) => 
                           bus_reg_dataout_2359_port, Q(22) => 
                           bus_reg_dataout_2358_port, Q(21) => 
                           bus_reg_dataout_2357_port, Q(20) => 
                           bus_reg_dataout_2356_port, Q(19) => 
                           bus_reg_dataout_2355_port, Q(18) => 
                           bus_reg_dataout_2354_port, Q(17) => 
                           bus_reg_dataout_2353_port, Q(16) => 
                           bus_reg_dataout_2352_port, Q(15) => 
                           bus_reg_dataout_2351_port, Q(14) => 
                           bus_reg_dataout_2350_port, Q(13) => 
                           bus_reg_dataout_2349_port, Q(12) => 
                           bus_reg_dataout_2348_port, Q(11) => 
                           bus_reg_dataout_2347_port, Q(10) => 
                           bus_reg_dataout_2346_port, Q(9) => 
                           bus_reg_dataout_2345_port, Q(8) => 
                           bus_reg_dataout_2344_port, Q(7) => 
                           bus_reg_dataout_2343_port, Q(6) => 
                           bus_reg_dataout_2342_port, Q(5) => 
                           bus_reg_dataout_2341_port, Q(4) => 
                           bus_reg_dataout_2340_port, Q(3) => 
                           bus_reg_dataout_2339_port, Q(2) => 
                           bus_reg_dataout_2338_port, Q(1) => 
                           bus_reg_dataout_2337_port, Q(0) => 
                           bus_reg_dataout_2336_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_81_port);
   MUX_SELINPUT_82 : mux_N32_M1_3 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n593,
                           Y(30) => n585, Y(29) => n577, Y(28) => n569, Y(27) 
                           => n561, Y(26) => n553, Y(25) => n545, Y(24) => n537
                           , Y(23) => n529, Y(22) => n521, Y(21) => n513, Y(20)
                           => n505, Y(19) => n497, Y(18) => n489, Y(17) => n481
                           , Y(16) => n473, Y(15) => n465, Y(14) => n457, Y(13)
                           => n449, Y(12) => n441, Y(11) => n433, Y(10) => n425
                           , Y(9) => n417, Y(8) => n409, Y(7) => n401, Y(6) => 
                           n393, Y(5) => n385, Y(4) => n377, Y(3) => n369, Y(2)
                           => n361, Y(1) => n353, Y(0) => n345);
   BLOCKi_82 : reg_generic_N32_RSTVAL0_6 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2399_port, Q(30) => 
                           bus_reg_dataout_2398_port, Q(29) => 
                           bus_reg_dataout_2397_port, Q(28) => 
                           bus_reg_dataout_2396_port, Q(27) => 
                           bus_reg_dataout_2395_port, Q(26) => 
                           bus_reg_dataout_2394_port, Q(25) => 
                           bus_reg_dataout_2393_port, Q(24) => 
                           bus_reg_dataout_2392_port, Q(23) => 
                           bus_reg_dataout_2391_port, Q(22) => 
                           bus_reg_dataout_2390_port, Q(21) => 
                           bus_reg_dataout_2389_port, Q(20) => 
                           bus_reg_dataout_2388_port, Q(19) => 
                           bus_reg_dataout_2387_port, Q(18) => 
                           bus_reg_dataout_2386_port, Q(17) => 
                           bus_reg_dataout_2385_port, Q(16) => 
                           bus_reg_dataout_2384_port, Q(15) => 
                           bus_reg_dataout_2383_port, Q(14) => 
                           bus_reg_dataout_2382_port, Q(13) => 
                           bus_reg_dataout_2381_port, Q(12) => 
                           bus_reg_dataout_2380_port, Q(11) => 
                           bus_reg_dataout_2379_port, Q(10) => 
                           bus_reg_dataout_2378_port, Q(9) => 
                           bus_reg_dataout_2377_port, Q(8) => 
                           bus_reg_dataout_2376_port, Q(7) => 
                           bus_reg_dataout_2375_port, Q(6) => 
                           bus_reg_dataout_2374_port, Q(5) => 
                           bus_reg_dataout_2373_port, Q(4) => 
                           bus_reg_dataout_2372_port, Q(3) => 
                           bus_reg_dataout_2371_port, Q(2) => 
                           bus_reg_dataout_2370_port, Q(1) => 
                           bus_reg_dataout_2369_port, Q(0) => 
                           bus_reg_dataout_2368_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_82_port);
   BLOCKi_83 : reg_generic_N32_RSTVAL0_5 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2431_port, Q(30) => 
                           bus_reg_dataout_2430_port, Q(29) => 
                           bus_reg_dataout_2429_port, Q(28) => 
                           bus_reg_dataout_2428_port, Q(27) => 
                           bus_reg_dataout_2427_port, Q(26) => 
                           bus_reg_dataout_2426_port, Q(25) => 
                           bus_reg_dataout_2425_port, Q(24) => 
                           bus_reg_dataout_2424_port, Q(23) => 
                           bus_reg_dataout_2423_port, Q(22) => 
                           bus_reg_dataout_2422_port, Q(21) => 
                           bus_reg_dataout_2421_port, Q(20) => 
                           bus_reg_dataout_2420_port, Q(19) => 
                           bus_reg_dataout_2419_port, Q(18) => 
                           bus_reg_dataout_2418_port, Q(17) => 
                           bus_reg_dataout_2417_port, Q(16) => 
                           bus_reg_dataout_2416_port, Q(15) => 
                           bus_reg_dataout_2415_port, Q(14) => 
                           bus_reg_dataout_2414_port, Q(13) => 
                           bus_reg_dataout_2413_port, Q(12) => 
                           bus_reg_dataout_2412_port, Q(11) => 
                           bus_reg_dataout_2411_port, Q(10) => 
                           bus_reg_dataout_2410_port, Q(9) => 
                           bus_reg_dataout_2409_port, Q(8) => 
                           bus_reg_dataout_2408_port, Q(7) => 
                           bus_reg_dataout_2407_port, Q(6) => 
                           bus_reg_dataout_2406_port, Q(5) => 
                           bus_reg_dataout_2405_port, Q(4) => 
                           bus_reg_dataout_2404_port, Q(3) => 
                           bus_reg_dataout_2403_port, Q(2) => 
                           bus_reg_dataout_2402_port, Q(1) => 
                           bus_reg_dataout_2401_port, Q(0) => 
                           bus_reg_dataout_2400_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_83_port);
   MUX_SELINPUT_84 : mux_N32_M1_2 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n592,
                           Y(30) => n584, Y(29) => n576, Y(28) => n568, Y(27) 
                           => n560, Y(26) => n552, Y(25) => n544, Y(24) => n536
                           , Y(23) => n528, Y(22) => n520, Y(21) => n512, Y(20)
                           => n504, Y(19) => n496, Y(18) => n488, Y(17) => n480
                           , Y(16) => n472, Y(15) => n464, Y(14) => n456, Y(13)
                           => n448, Y(12) => n440, Y(11) => n432, Y(10) => n424
                           , Y(9) => n416, Y(8) => n408, Y(7) => n400, Y(6) => 
                           n392, Y(5) => n384, Y(4) => n376, Y(3) => n368, Y(2)
                           => n360, Y(1) => n352, Y(0) => n344);
   BLOCKi_84 : reg_generic_N32_RSTVAL0_4 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2463_port, Q(30) => 
                           bus_reg_dataout_2462_port, Q(29) => 
                           bus_reg_dataout_2461_port, Q(28) => 
                           bus_reg_dataout_2460_port, Q(27) => 
                           bus_reg_dataout_2459_port, Q(26) => 
                           bus_reg_dataout_2458_port, Q(25) => 
                           bus_reg_dataout_2457_port, Q(24) => 
                           bus_reg_dataout_2456_port, Q(23) => 
                           bus_reg_dataout_2455_port, Q(22) => 
                           bus_reg_dataout_2454_port, Q(21) => 
                           bus_reg_dataout_2453_port, Q(20) => 
                           bus_reg_dataout_2452_port, Q(19) => 
                           bus_reg_dataout_2451_port, Q(18) => 
                           bus_reg_dataout_2450_port, Q(17) => 
                           bus_reg_dataout_2449_port, Q(16) => 
                           bus_reg_dataout_2448_port, Q(15) => 
                           bus_reg_dataout_2447_port, Q(14) => 
                           bus_reg_dataout_2446_port, Q(13) => 
                           bus_reg_dataout_2445_port, Q(12) => 
                           bus_reg_dataout_2444_port, Q(11) => 
                           bus_reg_dataout_2443_port, Q(10) => 
                           bus_reg_dataout_2442_port, Q(9) => 
                           bus_reg_dataout_2441_port, Q(8) => 
                           bus_reg_dataout_2440_port, Q(7) => 
                           bus_reg_dataout_2439_port, Q(6) => 
                           bus_reg_dataout_2438_port, Q(5) => 
                           bus_reg_dataout_2437_port, Q(4) => 
                           bus_reg_dataout_2436_port, Q(3) => 
                           bus_reg_dataout_2435_port, Q(2) => 
                           bus_reg_dataout_2434_port, Q(1) => 
                           bus_reg_dataout_2433_port, Q(0) => 
                           bus_reg_dataout_2432_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_84_port);
   BLOCKi_85 : reg_generic_N32_RSTVAL0_3 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2495_port, Q(30) => 
                           bus_reg_dataout_2494_port, Q(29) => 
                           bus_reg_dataout_2493_port, Q(28) => 
                           bus_reg_dataout_2492_port, Q(27) => 
                           bus_reg_dataout_2491_port, Q(26) => 
                           bus_reg_dataout_2490_port, Q(25) => 
                           bus_reg_dataout_2489_port, Q(24) => 
                           bus_reg_dataout_2488_port, Q(23) => 
                           bus_reg_dataout_2487_port, Q(22) => 
                           bus_reg_dataout_2486_port, Q(21) => 
                           bus_reg_dataout_2485_port, Q(20) => 
                           bus_reg_dataout_2484_port, Q(19) => 
                           bus_reg_dataout_2483_port, Q(18) => 
                           bus_reg_dataout_2482_port, Q(17) => 
                           bus_reg_dataout_2481_port, Q(16) => 
                           bus_reg_dataout_2480_port, Q(15) => 
                           bus_reg_dataout_2479_port, Q(14) => 
                           bus_reg_dataout_2478_port, Q(13) => 
                           bus_reg_dataout_2477_port, Q(12) => 
                           bus_reg_dataout_2476_port, Q(11) => 
                           bus_reg_dataout_2475_port, Q(10) => 
                           bus_reg_dataout_2474_port, Q(9) => 
                           bus_reg_dataout_2473_port, Q(8) => 
                           bus_reg_dataout_2472_port, Q(7) => 
                           bus_reg_dataout_2471_port, Q(6) => 
                           bus_reg_dataout_2470_port, Q(5) => 
                           bus_reg_dataout_2469_port, Q(4) => 
                           bus_reg_dataout_2468_port, Q(3) => 
                           bus_reg_dataout_2467_port, Q(2) => 
                           bus_reg_dataout_2466_port, Q(1) => 
                           bus_reg_dataout_2465_port, Q(0) => 
                           bus_reg_dataout_2464_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_85_port);
   MUX_SELINPUT_86 : mux_N32_M1_1 port map( S => c_swin_masked_1bit_4_0_port, 
                           Q(63) => BUS_FROMEM(31), Q(62) => BUS_FROMEM(30), 
                           Q(61) => BUS_FROMEM(29), Q(60) => BUS_FROMEM(28), 
                           Q(59) => BUS_FROMEM(27), Q(58) => BUS_FROMEM(26), 
                           Q(57) => BUS_FROMEM(25), Q(56) => BUS_FROMEM(24), 
                           Q(55) => BUS_FROMEM(23), Q(54) => BUS_FROMEM(22), 
                           Q(53) => BUS_FROMEM(21), Q(52) => BUS_FROMEM(20), 
                           Q(51) => BUS_FROMEM(19), Q(50) => BUS_FROMEM(18), 
                           Q(49) => BUS_FROMEM(17), Q(48) => BUS_FROMEM(16), 
                           Q(47) => BUS_FROMEM(15), Q(46) => BUS_FROMEM(14), 
                           Q(45) => BUS_FROMEM(13), Q(44) => BUS_FROMEM(12), 
                           Q(43) => BUS_FROMEM(11), Q(42) => BUS_FROMEM(10), 
                           Q(41) => BUS_FROMEM(9), Q(40) => BUS_FROMEM(8), 
                           Q(39) => BUS_FROMEM(7), Q(38) => BUS_FROMEM(6), 
                           Q(37) => BUS_FROMEM(5), Q(36) => BUS_FROMEM(4), 
                           Q(35) => BUS_FROMEM(3), Q(34) => BUS_FROMEM(2), 
                           Q(33) => BUS_FROMEM(1), Q(32) => BUS_FROMEM(0), 
                           Q(31) => DATAIN(31), Q(30) => DATAIN(30), Q(29) => 
                           DATAIN(29), Q(28) => DATAIN(28), Q(27) => DATAIN(27)
                           , Q(26) => DATAIN(26), Q(25) => DATAIN(25), Q(24) =>
                           DATAIN(24), Q(23) => DATAIN(23), Q(22) => DATAIN(22)
                           , Q(21) => DATAIN(21), Q(20) => DATAIN(20), Q(19) =>
                           DATAIN(19), Q(18) => DATAIN(18), Q(17) => DATAIN(17)
                           , Q(16) => DATAIN(16), Q(15) => DATAIN(15), Q(14) =>
                           DATAIN(14), Q(13) => DATAIN(13), Q(12) => DATAIN(12)
                           , Q(11) => DATAIN(11), Q(10) => DATAIN(10), Q(9) => 
                           DATAIN(9), Q(8) => DATAIN(8), Q(7) => DATAIN(7), 
                           Q(6) => DATAIN(6), Q(5) => DATAIN(5), Q(4) => 
                           DATAIN(4), Q(3) => DATAIN(3), Q(2) => DATAIN(2), 
                           Q(1) => DATAIN(1), Q(0) => DATAIN(0), Y(31) => n591,
                           Y(30) => n583, Y(29) => n575, Y(28) => n567, Y(27) 
                           => n559, Y(26) => n551, Y(25) => n543, Y(24) => n535
                           , Y(23) => n527, Y(22) => n519, Y(21) => n511, Y(20)
                           => n503, Y(19) => n495, Y(18) => n487, Y(17) => n479
                           , Y(16) => n471, Y(15) => n463, Y(14) => n455, Y(13)
                           => n447, Y(12) => n439, Y(11) => n431, Y(10) => n423
                           , Y(9) => n415, Y(8) => n407, Y(7) => n399, Y(6) => 
                           n391, Y(5) => n383, Y(4) => n375, Y(3) => n367, Y(2)
                           => n359, Y(1) => n351, Y(0) => n343);
   BLOCKi_86 : reg_generic_N32_RSTVAL0_2 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2527_port, Q(30) => 
                           bus_reg_dataout_2526_port, Q(29) => 
                           bus_reg_dataout_2525_port, Q(28) => 
                           bus_reg_dataout_2524_port, Q(27) => 
                           bus_reg_dataout_2523_port, Q(26) => 
                           bus_reg_dataout_2522_port, Q(25) => 
                           bus_reg_dataout_2521_port, Q(24) => 
                           bus_reg_dataout_2520_port, Q(23) => 
                           bus_reg_dataout_2519_port, Q(22) => 
                           bus_reg_dataout_2518_port, Q(21) => 
                           bus_reg_dataout_2517_port, Q(20) => 
                           bus_reg_dataout_2516_port, Q(19) => 
                           bus_reg_dataout_2515_port, Q(18) => 
                           bus_reg_dataout_2514_port, Q(17) => 
                           bus_reg_dataout_2513_port, Q(16) => 
                           bus_reg_dataout_2512_port, Q(15) => 
                           bus_reg_dataout_2511_port, Q(14) => 
                           bus_reg_dataout_2510_port, Q(13) => 
                           bus_reg_dataout_2509_port, Q(12) => 
                           bus_reg_dataout_2508_port, Q(11) => 
                           bus_reg_dataout_2507_port, Q(10) => 
                           bus_reg_dataout_2506_port, Q(9) => 
                           bus_reg_dataout_2505_port, Q(8) => 
                           bus_reg_dataout_2504_port, Q(7) => 
                           bus_reg_dataout_2503_port, Q(6) => 
                           bus_reg_dataout_2502_port, Q(5) => 
                           bus_reg_dataout_2501_port, Q(4) => 
                           bus_reg_dataout_2500_port, Q(3) => 
                           bus_reg_dataout_2499_port, Q(2) => 
                           bus_reg_dataout_2498_port, Q(1) => 
                           bus_reg_dataout_2497_port, Q(0) => 
                           bus_reg_dataout_2496_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_86_port);
   BLOCKi_87 : reg_generic_N32_RSTVAL0_1 port map( D(31) => 
                           internal_inloc_data_4_31_port, D(30) => 
                           internal_inloc_data_4_30_port, D(29) => 
                           internal_inloc_data_4_29_port, D(28) => 
                           internal_inloc_data_4_28_port, D(27) => 
                           internal_inloc_data_4_27_port, D(26) => 
                           internal_inloc_data_4_26_port, D(25) => 
                           internal_inloc_data_4_25_port, D(24) => 
                           internal_inloc_data_4_24_port, D(23) => 
                           internal_inloc_data_4_23_port, D(22) => 
                           internal_inloc_data_4_22_port, D(21) => 
                           internal_inloc_data_4_21_port, D(20) => 
                           internal_inloc_data_4_20_port, D(19) => 
                           internal_inloc_data_4_19_port, D(18) => 
                           internal_inloc_data_4_18_port, D(17) => 
                           internal_inloc_data_4_17_port, D(16) => 
                           internal_inloc_data_4_16_port, D(15) => 
                           internal_inloc_data_4_15_port, D(14) => 
                           internal_inloc_data_4_14_port, D(13) => 
                           internal_inloc_data_4_13_port, D(12) => 
                           internal_inloc_data_4_12_port, D(11) => 
                           internal_inloc_data_4_11_port, D(10) => 
                           internal_inloc_data_4_10_port, D(9) => 
                           internal_inloc_data_4_9_port, D(8) => 
                           internal_inloc_data_4_8_port, D(7) => 
                           internal_inloc_data_4_7_port, D(6) => 
                           internal_inloc_data_4_6_port, D(5) => 
                           internal_inloc_data_4_5_port, D(4) => 
                           internal_inloc_data_4_4_port, D(3) => 
                           internal_inloc_data_4_3_port, D(2) => 
                           internal_inloc_data_4_2_port, D(1) => 
                           internal_inloc_data_4_1_port, D(0) => 
                           internal_inloc_data_4_0_port, Q(31) => 
                           bus_reg_dataout_2559_port, Q(30) => 
                           bus_reg_dataout_2558_port, Q(29) => 
                           bus_reg_dataout_2557_port, Q(28) => 
                           bus_reg_dataout_2556_port, Q(27) => 
                           bus_reg_dataout_2555_port, Q(26) => 
                           bus_reg_dataout_2554_port, Q(25) => 
                           bus_reg_dataout_2553_port, Q(24) => 
                           bus_reg_dataout_2552_port, Q(23) => 
                           bus_reg_dataout_2551_port, Q(22) => 
                           bus_reg_dataout_2550_port, Q(21) => 
                           bus_reg_dataout_2549_port, Q(20) => 
                           bus_reg_dataout_2548_port, Q(19) => 
                           bus_reg_dataout_2547_port, Q(18) => 
                           bus_reg_dataout_2546_port, Q(17) => 
                           bus_reg_dataout_2545_port, Q(16) => 
                           bus_reg_dataout_2544_port, Q(15) => 
                           bus_reg_dataout_2543_port, Q(14) => 
                           bus_reg_dataout_2542_port, Q(13) => 
                           bus_reg_dataout_2541_port, Q(12) => 
                           bus_reg_dataout_2540_port, Q(11) => 
                           bus_reg_dataout_2539_port, Q(10) => 
                           bus_reg_dataout_2538_port, Q(9) => 
                           bus_reg_dataout_2537_port, Q(8) => 
                           bus_reg_dataout_2536_port, Q(7) => 
                           bus_reg_dataout_2535_port, Q(6) => 
                           bus_reg_dataout_2534_port, Q(5) => 
                           bus_reg_dataout_2533_port, Q(4) => 
                           bus_reg_dataout_2532_port, Q(3) => 
                           bus_reg_dataout_2531_port, Q(2) => 
                           bus_reg_dataout_2530_port, Q(1) => 
                           bus_reg_dataout_2529_port, Q(0) => 
                           bus_reg_dataout_2528_port, Clk => CLK, Rst => RESET,
                           Enable => en_regi_87_port);
   DEC : decoder_N5 port map( Q(4) => ADD_WR(4), Q(3) => ADD_WR(3), Q(2) => 
                           ADD_WR(2), Q(1) => ADD_WR(1), Q(0) => ADD_WR(0), 
                           Y(31) => dec_output_31_port, Y(30) => 
                           dec_output_30_port, Y(29) => dec_output_29_port, 
                           Y(28) => dec_output_28_port, Y(27) => 
                           dec_output_27_port, Y(26) => dec_output_26_port, 
                           Y(25) => dec_output_25_port, Y(24) => 
                           dec_output_24_port, Y(23) => dec_output_23_port, 
                           Y(22) => dec_output_22_port, Y(21) => 
                           dec_output_21_port, Y(20) => dec_output_20_port, 
                           Y(19) => dec_output_19_port, Y(18) => 
                           dec_output_18_port, Y(17) => dec_output_17_port, 
                           Y(16) => dec_output_16_port, Y(15) => 
                           dec_output_15_port, Y(14) => dec_output_14_port, 
                           Y(13) => dec_output_13_port, Y(12) => 
                           dec_output_12_port, Y(11) => dec_output_11_port, 
                           Y(10) => dec_output_10_port, Y(9) => 
                           dec_output_9_port, Y(8) => dec_output_8_port, Y(7) 
                           => dec_output_7_port, Y(6) => dec_output_6_port, 
                           Y(5) => dec_output_5_port, Y(4) => dec_output_4_port
                           , Y(3) => dec_output_3_port, Y(2) => 
                           dec_output_2_port, Y(1) => dec_output_1_port, Y(0) 
                           => dec_output_0_port);
   ConnMtx : connection_mtx_M8_N8_F5 port map( dec(31) => 
                           dec_out_with_wen_31_port, dec(30) => 
                           dec_out_with_wen_30_port, dec(29) => 
                           dec_out_with_wen_29_port, dec(28) => 
                           dec_out_with_wen_28_port, dec(27) => 
                           dec_out_with_wen_27_port, dec(26) => 
                           dec_out_with_wen_26_port, dec(25) => 
                           dec_out_with_wen_25_port, dec(24) => 
                           dec_out_with_wen_24_port, dec(23) => 
                           dec_out_with_wen_23_port, dec(22) => 
                           dec_out_with_wen_22_port, dec(21) => 
                           dec_out_with_wen_21_port, dec(20) => 
                           dec_out_with_wen_20_port, dec(19) => 
                           dec_out_with_wen_19_port, dec(18) => 
                           dec_out_with_wen_18_port, dec(17) => 
                           dec_out_with_wen_17_port, dec(16) => 
                           dec_out_with_wen_16_port, dec(15) => 
                           dec_out_with_wen_15_port, dec(14) => 
                           dec_out_with_wen_14_port, dec(13) => 
                           dec_out_with_wen_13_port, dec(12) => 
                           dec_out_with_wen_12_port, dec(11) => 
                           dec_out_with_wen_11_port, dec(10) => 
                           dec_out_with_wen_10_port, dec(9) => 
                           dec_out_with_wen_9_port, dec(8) => 
                           dec_out_with_wen_8_port, dec(7) => 
                           dec_out_with_wen_7_port, dec(6) => 
                           dec_out_with_wen_6_port, dec(5) => 
                           dec_out_with_wen_5_port, dec(4) => 
                           dec_out_with_wen_4_port, dec(3) => 
                           dec_out_with_wen_3_port, dec(2) => 
                           dec_out_with_wen_2_port, dec(1) => 
                           dec_out_with_wen_1_port, dec(0) => 
                           dec_out_with_wen_0_port, addr_pop(15) => 
                           fill_address_ext_15_port, addr_pop(14) => 
                           fill_address_ext_14_port, addr_pop(13) => 
                           fill_address_ext_13_port, addr_pop(12) => 
                           fill_address_ext_12_port, addr_pop(11) => 
                           fill_address_ext_11_port, addr_pop(10) => 
                           fill_address_ext_10_port, addr_pop(9) => 
                           fill_address_ext_9_port, addr_pop(8) => 
                           fill_address_ext_8_port, addr_pop(7) => 
                           fill_address_ext_7_port, addr_pop(6) => 
                           fill_address_ext_6_port, addr_pop(5) => 
                           fill_address_ext_5_port, addr_pop(4) => 
                           fill_address_ext_4_port, addr_pop(3) => 
                           fill_address_ext_3_port, addr_pop(2) => 
                           fill_address_ext_2_port, addr_pop(1) => 
                           fill_address_ext_1_port, addr_pop(0) => 
                           fill_address_ext_0_port, win(4) => c_win_4_port, 
                           win(3) => c_win_3_port, win(2) => c_win_2_port, 
                           win(1) => c_win_1_port, win(0) => c_win_0_port, 
                           swp(4) => c_swin_masked_1bit_4_0_port, swp(3) => 
                           c_swin_masked_1bit_3_0_port, swp(2) => 
                           c_swin_masked_1bit_2_0_port, swp(1) => 
                           c_swin_masked_1bit_1_0_port, swp(0) => 
                           c_swin_masked_1bit_0_0_port, sel(87) => 
                           en_regi_87_port, sel(86) => en_regi_86_port, sel(85)
                           => en_regi_85_port, sel(84) => en_regi_84_port, 
                           sel(83) => en_regi_83_port, sel(82) => 
                           en_regi_82_port, sel(81) => en_regi_81_port, sel(80)
                           => en_regi_80_port, sel(79) => en_regi_79_port, 
                           sel(78) => en_regi_78_port, sel(77) => 
                           en_regi_77_port, sel(76) => en_regi_76_port, sel(75)
                           => en_regi_75_port, sel(74) => en_regi_74_port, 
                           sel(73) => en_regi_73_port, sel(72) => 
                           en_regi_72_port, sel(71) => en_regi_71_port, sel(70)
                           => en_regi_70_port, sel(69) => en_regi_69_port, 
                           sel(68) => en_regi_68_port, sel(67) => 
                           en_regi_67_port, sel(66) => en_regi_66_port, sel(65)
                           => en_regi_65_port, sel(64) => en_regi_64_port, 
                           sel(63) => en_regi_63_port, sel(62) => 
                           en_regi_62_port, sel(61) => en_regi_61_port, sel(60)
                           => en_regi_60_port, sel(59) => en_regi_59_port, 
                           sel(58) => en_regi_58_port, sel(57) => 
                           en_regi_57_port, sel(56) => en_regi_56_port, sel(55)
                           => en_regi_55_port, sel(54) => en_regi_54_port, 
                           sel(53) => en_regi_53_port, sel(52) => 
                           en_regi_52_port, sel(51) => en_regi_51_port, sel(50)
                           => en_regi_50_port, sel(49) => en_regi_49_port, 
                           sel(48) => en_regi_48_port, sel(47) => 
                           en_regi_47_port, sel(46) => en_regi_46_port, sel(45)
                           => en_regi_45_port, sel(44) => en_regi_44_port, 
                           sel(43) => en_regi_43_port, sel(42) => 
                           en_regi_42_port, sel(41) => en_regi_41_port, sel(40)
                           => en_regi_40_port, sel(39) => en_regi_39_port, 
                           sel(38) => en_regi_38_port, sel(37) => 
                           en_regi_37_port, sel(36) => en_regi_36_port, sel(35)
                           => en_regi_35_port, sel(34) => en_regi_34_port, 
                           sel(33) => en_regi_33_port, sel(32) => 
                           en_regi_32_port, sel(31) => en_regi_31_port, sel(30)
                           => en_regi_30_port, sel(29) => en_regi_29_port, 
                           sel(28) => en_regi_28_port, sel(27) => 
                           en_regi_27_port, sel(26) => en_regi_26_port, sel(25)
                           => en_regi_25_port, sel(24) => en_regi_24_port, 
                           sel(23) => en_regi_23_port, sel(22) => 
                           en_regi_22_port, sel(21) => en_regi_21_port, sel(20)
                           => en_regi_20_port, sel(19) => en_regi_19_port, 
                           sel(18) => en_regi_18_port, sel(17) => 
                           en_regi_17_port, sel(16) => en_regi_16_port, sel(15)
                           => en_regi_15_port, sel(14) => en_regi_14_port, 
                           sel(13) => en_regi_13_port, sel(12) => 
                           en_regi_12_port, sel(11) => en_regi_11_port, sel(10)
                           => en_regi_10_port, sel(9) => en_regi_9_port, sel(8)
                           => en_regi_8_port, sel(7) => en_regi_7_port, sel(6) 
                           => en_regi_6_port, sel(5) => en_regi_5_port, sel(4) 
                           => en_regi_4_port, sel(3) => en_regi_3_port, sel(2) 
                           => en_regi_2_port, sel(1) => en_regi_1_port, sel(0) 
                           => en_regi_0_port);
   SWP_NEXT_CALC : nwin_calc_F5_1 port map( c_win(4) => c_swin_4_port, c_win(3)
                           => c_swin_3_port, c_win(2) => c_swin_2_port, 
                           c_win(1) => c_swin_1_port, c_win(0) => c_swin_0_port
                           , sel(1) => donespill_donefill_encoding_1_port, 
                           sel(0) => donespill_donefill_encoding_0_port, 
                           n_win(4) => next_swp_4_port, n_win(3) => 
                           next_swp_3_port, n_win(2) => next_swp_2_port, 
                           n_win(1) => next_swp_1_port, n_win(0) => 
                           next_swp_0_port);
   SWP : reg_generic_N5_RSTVAL1_1 port map( D(4) => next_swp_4_port, D(3) => 
                           next_swp_3_port, D(2) => next_swp_2_port, D(1) => 
                           next_swp_1_port, D(0) => next_swp_0_port, Q(4) => 
                           c_swin_4_port, Q(3) => c_swin_3_port, Q(2) => 
                           c_swin_2_port, Q(1) => c_swin_1_port, Q(0) => 
                           c_swin_0_port, Clk => CLK, Rst => RESET, Enable => 
                           X_Logic1_port);
   EQ_CHECK : equal_check_N5_0 port map( A(4) => c_win_2_port, A(3) => 
                           c_win_1_port, A(2) => c_win_0_port, A(1) => 
                           c_win_4_port, A(0) => c_win_3_port, B(4) => 
                           c_swin_4_port, B(3) => c_swin_3_port, B(2) => 
                           c_swin_2_port, B(1) => c_swin_1_port, B(0) => 
                           c_swin_0_port, EQUAL => spilleq);
   SELBLOCK_INLOC : in_loc_selblock_NBIT_DATA32_N8_F5 port map( regs(2559) => 
                           bus_reg_dataout_2559_port, regs(2558) => 
                           bus_reg_dataout_2558_port, regs(2557) => 
                           bus_reg_dataout_2557_port, regs(2556) => 
                           bus_reg_dataout_2556_port, regs(2555) => 
                           bus_reg_dataout_2555_port, regs(2554) => 
                           bus_reg_dataout_2554_port, regs(2553) => 
                           bus_reg_dataout_2553_port, regs(2552) => 
                           bus_reg_dataout_2552_port, regs(2551) => 
                           bus_reg_dataout_2551_port, regs(2550) => 
                           bus_reg_dataout_2550_port, regs(2549) => 
                           bus_reg_dataout_2549_port, regs(2548) => 
                           bus_reg_dataout_2548_port, regs(2547) => 
                           bus_reg_dataout_2547_port, regs(2546) => 
                           bus_reg_dataout_2546_port, regs(2545) => 
                           bus_reg_dataout_2545_port, regs(2544) => 
                           bus_reg_dataout_2544_port, regs(2543) => 
                           bus_reg_dataout_2543_port, regs(2542) => 
                           bus_reg_dataout_2542_port, regs(2541) => 
                           bus_reg_dataout_2541_port, regs(2540) => 
                           bus_reg_dataout_2540_port, regs(2539) => 
                           bus_reg_dataout_2539_port, regs(2538) => 
                           bus_reg_dataout_2538_port, regs(2537) => 
                           bus_reg_dataout_2537_port, regs(2536) => 
                           bus_reg_dataout_2536_port, regs(2535) => 
                           bus_reg_dataout_2535_port, regs(2534) => 
                           bus_reg_dataout_2534_port, regs(2533) => 
                           bus_reg_dataout_2533_port, regs(2532) => 
                           bus_reg_dataout_2532_port, regs(2531) => 
                           bus_reg_dataout_2531_port, regs(2530) => 
                           bus_reg_dataout_2530_port, regs(2529) => 
                           bus_reg_dataout_2529_port, regs(2528) => 
                           bus_reg_dataout_2528_port, regs(2527) => 
                           bus_reg_dataout_2527_port, regs(2526) => 
                           bus_reg_dataout_2526_port, regs(2525) => 
                           bus_reg_dataout_2525_port, regs(2524) => 
                           bus_reg_dataout_2524_port, regs(2523) => 
                           bus_reg_dataout_2523_port, regs(2522) => 
                           bus_reg_dataout_2522_port, regs(2521) => 
                           bus_reg_dataout_2521_port, regs(2520) => 
                           bus_reg_dataout_2520_port, regs(2519) => 
                           bus_reg_dataout_2519_port, regs(2518) => 
                           bus_reg_dataout_2518_port, regs(2517) => 
                           bus_reg_dataout_2517_port, regs(2516) => 
                           bus_reg_dataout_2516_port, regs(2515) => 
                           bus_reg_dataout_2515_port, regs(2514) => 
                           bus_reg_dataout_2514_port, regs(2513) => 
                           bus_reg_dataout_2513_port, regs(2512) => 
                           bus_reg_dataout_2512_port, regs(2511) => 
                           bus_reg_dataout_2511_port, regs(2510) => 
                           bus_reg_dataout_2510_port, regs(2509) => 
                           bus_reg_dataout_2509_port, regs(2508) => 
                           bus_reg_dataout_2508_port, regs(2507) => 
                           bus_reg_dataout_2507_port, regs(2506) => 
                           bus_reg_dataout_2506_port, regs(2505) => 
                           bus_reg_dataout_2505_port, regs(2504) => 
                           bus_reg_dataout_2504_port, regs(2503) => 
                           bus_reg_dataout_2503_port, regs(2502) => 
                           bus_reg_dataout_2502_port, regs(2501) => 
                           bus_reg_dataout_2501_port, regs(2500) => 
                           bus_reg_dataout_2500_port, regs(2499) => 
                           bus_reg_dataout_2499_port, regs(2498) => 
                           bus_reg_dataout_2498_port, regs(2497) => 
                           bus_reg_dataout_2497_port, regs(2496) => 
                           bus_reg_dataout_2496_port, regs(2495) => 
                           bus_reg_dataout_2495_port, regs(2494) => 
                           bus_reg_dataout_2494_port, regs(2493) => 
                           bus_reg_dataout_2493_port, regs(2492) => 
                           bus_reg_dataout_2492_port, regs(2491) => 
                           bus_reg_dataout_2491_port, regs(2490) => 
                           bus_reg_dataout_2490_port, regs(2489) => 
                           bus_reg_dataout_2489_port, regs(2488) => 
                           bus_reg_dataout_2488_port, regs(2487) => 
                           bus_reg_dataout_2487_port, regs(2486) => 
                           bus_reg_dataout_2486_port, regs(2485) => 
                           bus_reg_dataout_2485_port, regs(2484) => 
                           bus_reg_dataout_2484_port, regs(2483) => 
                           bus_reg_dataout_2483_port, regs(2482) => 
                           bus_reg_dataout_2482_port, regs(2481) => 
                           bus_reg_dataout_2481_port, regs(2480) => 
                           bus_reg_dataout_2480_port, regs(2479) => 
                           bus_reg_dataout_2479_port, regs(2478) => 
                           bus_reg_dataout_2478_port, regs(2477) => 
                           bus_reg_dataout_2477_port, regs(2476) => 
                           bus_reg_dataout_2476_port, regs(2475) => 
                           bus_reg_dataout_2475_port, regs(2474) => 
                           bus_reg_dataout_2474_port, regs(2473) => 
                           bus_reg_dataout_2473_port, regs(2472) => 
                           bus_reg_dataout_2472_port, regs(2471) => 
                           bus_reg_dataout_2471_port, regs(2470) => 
                           bus_reg_dataout_2470_port, regs(2469) => 
                           bus_reg_dataout_2469_port, regs(2468) => 
                           bus_reg_dataout_2468_port, regs(2467) => 
                           bus_reg_dataout_2467_port, regs(2466) => 
                           bus_reg_dataout_2466_port, regs(2465) => 
                           bus_reg_dataout_2465_port, regs(2464) => 
                           bus_reg_dataout_2464_port, regs(2463) => 
                           bus_reg_dataout_2463_port, regs(2462) => 
                           bus_reg_dataout_2462_port, regs(2461) => 
                           bus_reg_dataout_2461_port, regs(2460) => 
                           bus_reg_dataout_2460_port, regs(2459) => 
                           bus_reg_dataout_2459_port, regs(2458) => 
                           bus_reg_dataout_2458_port, regs(2457) => 
                           bus_reg_dataout_2457_port, regs(2456) => 
                           bus_reg_dataout_2456_port, regs(2455) => 
                           bus_reg_dataout_2455_port, regs(2454) => 
                           bus_reg_dataout_2454_port, regs(2453) => 
                           bus_reg_dataout_2453_port, regs(2452) => 
                           bus_reg_dataout_2452_port, regs(2451) => 
                           bus_reg_dataout_2451_port, regs(2450) => 
                           bus_reg_dataout_2450_port, regs(2449) => 
                           bus_reg_dataout_2449_port, regs(2448) => 
                           bus_reg_dataout_2448_port, regs(2447) => 
                           bus_reg_dataout_2447_port, regs(2446) => 
                           bus_reg_dataout_2446_port, regs(2445) => 
                           bus_reg_dataout_2445_port, regs(2444) => 
                           bus_reg_dataout_2444_port, regs(2443) => 
                           bus_reg_dataout_2443_port, regs(2442) => 
                           bus_reg_dataout_2442_port, regs(2441) => 
                           bus_reg_dataout_2441_port, regs(2440) => 
                           bus_reg_dataout_2440_port, regs(2439) => 
                           bus_reg_dataout_2439_port, regs(2438) => 
                           bus_reg_dataout_2438_port, regs(2437) => 
                           bus_reg_dataout_2437_port, regs(2436) => 
                           bus_reg_dataout_2436_port, regs(2435) => 
                           bus_reg_dataout_2435_port, regs(2434) => 
                           bus_reg_dataout_2434_port, regs(2433) => 
                           bus_reg_dataout_2433_port, regs(2432) => 
                           bus_reg_dataout_2432_port, regs(2431) => 
                           bus_reg_dataout_2431_port, regs(2430) => 
                           bus_reg_dataout_2430_port, regs(2429) => 
                           bus_reg_dataout_2429_port, regs(2428) => 
                           bus_reg_dataout_2428_port, regs(2427) => 
                           bus_reg_dataout_2427_port, regs(2426) => 
                           bus_reg_dataout_2426_port, regs(2425) => 
                           bus_reg_dataout_2425_port, regs(2424) => 
                           bus_reg_dataout_2424_port, regs(2423) => 
                           bus_reg_dataout_2423_port, regs(2422) => 
                           bus_reg_dataout_2422_port, regs(2421) => 
                           bus_reg_dataout_2421_port, regs(2420) => 
                           bus_reg_dataout_2420_port, regs(2419) => 
                           bus_reg_dataout_2419_port, regs(2418) => 
                           bus_reg_dataout_2418_port, regs(2417) => 
                           bus_reg_dataout_2417_port, regs(2416) => 
                           bus_reg_dataout_2416_port, regs(2415) => 
                           bus_reg_dataout_2415_port, regs(2414) => 
                           bus_reg_dataout_2414_port, regs(2413) => 
                           bus_reg_dataout_2413_port, regs(2412) => 
                           bus_reg_dataout_2412_port, regs(2411) => 
                           bus_reg_dataout_2411_port, regs(2410) => 
                           bus_reg_dataout_2410_port, regs(2409) => 
                           bus_reg_dataout_2409_port, regs(2408) => 
                           bus_reg_dataout_2408_port, regs(2407) => 
                           bus_reg_dataout_2407_port, regs(2406) => 
                           bus_reg_dataout_2406_port, regs(2405) => 
                           bus_reg_dataout_2405_port, regs(2404) => 
                           bus_reg_dataout_2404_port, regs(2403) => 
                           bus_reg_dataout_2403_port, regs(2402) => 
                           bus_reg_dataout_2402_port, regs(2401) => 
                           bus_reg_dataout_2401_port, regs(2400) => 
                           bus_reg_dataout_2400_port, regs(2399) => 
                           bus_reg_dataout_2399_port, regs(2398) => 
                           bus_reg_dataout_2398_port, regs(2397) => 
                           bus_reg_dataout_2397_port, regs(2396) => 
                           bus_reg_dataout_2396_port, regs(2395) => 
                           bus_reg_dataout_2395_port, regs(2394) => 
                           bus_reg_dataout_2394_port, regs(2393) => 
                           bus_reg_dataout_2393_port, regs(2392) => 
                           bus_reg_dataout_2392_port, regs(2391) => 
                           bus_reg_dataout_2391_port, regs(2390) => 
                           bus_reg_dataout_2390_port, regs(2389) => 
                           bus_reg_dataout_2389_port, regs(2388) => 
                           bus_reg_dataout_2388_port, regs(2387) => 
                           bus_reg_dataout_2387_port, regs(2386) => 
                           bus_reg_dataout_2386_port, regs(2385) => 
                           bus_reg_dataout_2385_port, regs(2384) => 
                           bus_reg_dataout_2384_port, regs(2383) => 
                           bus_reg_dataout_2383_port, regs(2382) => 
                           bus_reg_dataout_2382_port, regs(2381) => 
                           bus_reg_dataout_2381_port, regs(2380) => 
                           bus_reg_dataout_2380_port, regs(2379) => 
                           bus_reg_dataout_2379_port, regs(2378) => 
                           bus_reg_dataout_2378_port, regs(2377) => 
                           bus_reg_dataout_2377_port, regs(2376) => 
                           bus_reg_dataout_2376_port, regs(2375) => 
                           bus_reg_dataout_2375_port, regs(2374) => 
                           bus_reg_dataout_2374_port, regs(2373) => 
                           bus_reg_dataout_2373_port, regs(2372) => 
                           bus_reg_dataout_2372_port, regs(2371) => 
                           bus_reg_dataout_2371_port, regs(2370) => 
                           bus_reg_dataout_2370_port, regs(2369) => 
                           bus_reg_dataout_2369_port, regs(2368) => 
                           bus_reg_dataout_2368_port, regs(2367) => 
                           bus_reg_dataout_2367_port, regs(2366) => 
                           bus_reg_dataout_2366_port, regs(2365) => 
                           bus_reg_dataout_2365_port, regs(2364) => 
                           bus_reg_dataout_2364_port, regs(2363) => 
                           bus_reg_dataout_2363_port, regs(2362) => 
                           bus_reg_dataout_2362_port, regs(2361) => 
                           bus_reg_dataout_2361_port, regs(2360) => 
                           bus_reg_dataout_2360_port, regs(2359) => 
                           bus_reg_dataout_2359_port, regs(2358) => 
                           bus_reg_dataout_2358_port, regs(2357) => 
                           bus_reg_dataout_2357_port, regs(2356) => 
                           bus_reg_dataout_2356_port, regs(2355) => 
                           bus_reg_dataout_2355_port, regs(2354) => 
                           bus_reg_dataout_2354_port, regs(2353) => 
                           bus_reg_dataout_2353_port, regs(2352) => 
                           bus_reg_dataout_2352_port, regs(2351) => 
                           bus_reg_dataout_2351_port, regs(2350) => 
                           bus_reg_dataout_2350_port, regs(2349) => 
                           bus_reg_dataout_2349_port, regs(2348) => 
                           bus_reg_dataout_2348_port, regs(2347) => 
                           bus_reg_dataout_2347_port, regs(2346) => 
                           bus_reg_dataout_2346_port, regs(2345) => 
                           bus_reg_dataout_2345_port, regs(2344) => 
                           bus_reg_dataout_2344_port, regs(2343) => 
                           bus_reg_dataout_2343_port, regs(2342) => 
                           bus_reg_dataout_2342_port, regs(2341) => 
                           bus_reg_dataout_2341_port, regs(2340) => 
                           bus_reg_dataout_2340_port, regs(2339) => 
                           bus_reg_dataout_2339_port, regs(2338) => 
                           bus_reg_dataout_2338_port, regs(2337) => 
                           bus_reg_dataout_2337_port, regs(2336) => 
                           bus_reg_dataout_2336_port, regs(2335) => 
                           bus_reg_dataout_2335_port, regs(2334) => 
                           bus_reg_dataout_2334_port, regs(2333) => 
                           bus_reg_dataout_2333_port, regs(2332) => 
                           bus_reg_dataout_2332_port, regs(2331) => 
                           bus_reg_dataout_2331_port, regs(2330) => 
                           bus_reg_dataout_2330_port, regs(2329) => 
                           bus_reg_dataout_2329_port, regs(2328) => 
                           bus_reg_dataout_2328_port, regs(2327) => 
                           bus_reg_dataout_2327_port, regs(2326) => 
                           bus_reg_dataout_2326_port, regs(2325) => 
                           bus_reg_dataout_2325_port, regs(2324) => 
                           bus_reg_dataout_2324_port, regs(2323) => 
                           bus_reg_dataout_2323_port, regs(2322) => 
                           bus_reg_dataout_2322_port, regs(2321) => 
                           bus_reg_dataout_2321_port, regs(2320) => 
                           bus_reg_dataout_2320_port, regs(2319) => 
                           bus_reg_dataout_2319_port, regs(2318) => 
                           bus_reg_dataout_2318_port, regs(2317) => 
                           bus_reg_dataout_2317_port, regs(2316) => 
                           bus_reg_dataout_2316_port, regs(2315) => 
                           bus_reg_dataout_2315_port, regs(2314) => 
                           bus_reg_dataout_2314_port, regs(2313) => 
                           bus_reg_dataout_2313_port, regs(2312) => 
                           bus_reg_dataout_2312_port, regs(2311) => 
                           bus_reg_dataout_2311_port, regs(2310) => 
                           bus_reg_dataout_2310_port, regs(2309) => 
                           bus_reg_dataout_2309_port, regs(2308) => 
                           bus_reg_dataout_2308_port, regs(2307) => 
                           bus_reg_dataout_2307_port, regs(2306) => 
                           bus_reg_dataout_2306_port, regs(2305) => 
                           bus_reg_dataout_2305_port, regs(2304) => 
                           bus_reg_dataout_2304_port, regs(2303) => 
                           bus_reg_dataout_2303_port, regs(2302) => 
                           bus_reg_dataout_2302_port, regs(2301) => 
                           bus_reg_dataout_2301_port, regs(2300) => 
                           bus_reg_dataout_2300_port, regs(2299) => 
                           bus_reg_dataout_2299_port, regs(2298) => 
                           bus_reg_dataout_2298_port, regs(2297) => 
                           bus_reg_dataout_2297_port, regs(2296) => 
                           bus_reg_dataout_2296_port, regs(2295) => 
                           bus_reg_dataout_2295_port, regs(2294) => 
                           bus_reg_dataout_2294_port, regs(2293) => 
                           bus_reg_dataout_2293_port, regs(2292) => 
                           bus_reg_dataout_2292_port, regs(2291) => 
                           bus_reg_dataout_2291_port, regs(2290) => 
                           bus_reg_dataout_2290_port, regs(2289) => 
                           bus_reg_dataout_2289_port, regs(2288) => 
                           bus_reg_dataout_2288_port, regs(2287) => 
                           bus_reg_dataout_2287_port, regs(2286) => 
                           bus_reg_dataout_2286_port, regs(2285) => 
                           bus_reg_dataout_2285_port, regs(2284) => 
                           bus_reg_dataout_2284_port, regs(2283) => 
                           bus_reg_dataout_2283_port, regs(2282) => 
                           bus_reg_dataout_2282_port, regs(2281) => 
                           bus_reg_dataout_2281_port, regs(2280) => 
                           bus_reg_dataout_2280_port, regs(2279) => 
                           bus_reg_dataout_2279_port, regs(2278) => 
                           bus_reg_dataout_2278_port, regs(2277) => 
                           bus_reg_dataout_2277_port, regs(2276) => 
                           bus_reg_dataout_2276_port, regs(2275) => 
                           bus_reg_dataout_2275_port, regs(2274) => 
                           bus_reg_dataout_2274_port, regs(2273) => 
                           bus_reg_dataout_2273_port, regs(2272) => 
                           bus_reg_dataout_2272_port, regs(2271) => 
                           bus_reg_dataout_2271_port, regs(2270) => 
                           bus_reg_dataout_2270_port, regs(2269) => 
                           bus_reg_dataout_2269_port, regs(2268) => 
                           bus_reg_dataout_2268_port, regs(2267) => 
                           bus_reg_dataout_2267_port, regs(2266) => 
                           bus_reg_dataout_2266_port, regs(2265) => 
                           bus_reg_dataout_2265_port, regs(2264) => 
                           bus_reg_dataout_2264_port, regs(2263) => 
                           bus_reg_dataout_2263_port, regs(2262) => 
                           bus_reg_dataout_2262_port, regs(2261) => 
                           bus_reg_dataout_2261_port, regs(2260) => 
                           bus_reg_dataout_2260_port, regs(2259) => 
                           bus_reg_dataout_2259_port, regs(2258) => 
                           bus_reg_dataout_2258_port, regs(2257) => 
                           bus_reg_dataout_2257_port, regs(2256) => 
                           bus_reg_dataout_2256_port, regs(2255) => 
                           bus_reg_dataout_2255_port, regs(2254) => 
                           bus_reg_dataout_2254_port, regs(2253) => 
                           bus_reg_dataout_2253_port, regs(2252) => 
                           bus_reg_dataout_2252_port, regs(2251) => 
                           bus_reg_dataout_2251_port, regs(2250) => 
                           bus_reg_dataout_2250_port, regs(2249) => 
                           bus_reg_dataout_2249_port, regs(2248) => 
                           bus_reg_dataout_2248_port, regs(2247) => 
                           bus_reg_dataout_2247_port, regs(2246) => 
                           bus_reg_dataout_2246_port, regs(2245) => 
                           bus_reg_dataout_2245_port, regs(2244) => 
                           bus_reg_dataout_2244_port, regs(2243) => 
                           bus_reg_dataout_2243_port, regs(2242) => 
                           bus_reg_dataout_2242_port, regs(2241) => 
                           bus_reg_dataout_2241_port, regs(2240) => 
                           bus_reg_dataout_2240_port, regs(2239) => 
                           bus_reg_dataout_2239_port, regs(2238) => 
                           bus_reg_dataout_2238_port, regs(2237) => 
                           bus_reg_dataout_2237_port, regs(2236) => 
                           bus_reg_dataout_2236_port, regs(2235) => 
                           bus_reg_dataout_2235_port, regs(2234) => 
                           bus_reg_dataout_2234_port, regs(2233) => 
                           bus_reg_dataout_2233_port, regs(2232) => 
                           bus_reg_dataout_2232_port, regs(2231) => 
                           bus_reg_dataout_2231_port, regs(2230) => 
                           bus_reg_dataout_2230_port, regs(2229) => 
                           bus_reg_dataout_2229_port, regs(2228) => 
                           bus_reg_dataout_2228_port, regs(2227) => 
                           bus_reg_dataout_2227_port, regs(2226) => 
                           bus_reg_dataout_2226_port, regs(2225) => 
                           bus_reg_dataout_2225_port, regs(2224) => 
                           bus_reg_dataout_2224_port, regs(2223) => 
                           bus_reg_dataout_2223_port, regs(2222) => 
                           bus_reg_dataout_2222_port, regs(2221) => 
                           bus_reg_dataout_2221_port, regs(2220) => 
                           bus_reg_dataout_2220_port, regs(2219) => 
                           bus_reg_dataout_2219_port, regs(2218) => 
                           bus_reg_dataout_2218_port, regs(2217) => 
                           bus_reg_dataout_2217_port, regs(2216) => 
                           bus_reg_dataout_2216_port, regs(2215) => 
                           bus_reg_dataout_2215_port, regs(2214) => 
                           bus_reg_dataout_2214_port, regs(2213) => 
                           bus_reg_dataout_2213_port, regs(2212) => 
                           bus_reg_dataout_2212_port, regs(2211) => 
                           bus_reg_dataout_2211_port, regs(2210) => 
                           bus_reg_dataout_2210_port, regs(2209) => 
                           bus_reg_dataout_2209_port, regs(2208) => 
                           bus_reg_dataout_2208_port, regs(2207) => 
                           bus_reg_dataout_2207_port, regs(2206) => 
                           bus_reg_dataout_2206_port, regs(2205) => 
                           bus_reg_dataout_2205_port, regs(2204) => 
                           bus_reg_dataout_2204_port, regs(2203) => 
                           bus_reg_dataout_2203_port, regs(2202) => 
                           bus_reg_dataout_2202_port, regs(2201) => 
                           bus_reg_dataout_2201_port, regs(2200) => 
                           bus_reg_dataout_2200_port, regs(2199) => 
                           bus_reg_dataout_2199_port, regs(2198) => 
                           bus_reg_dataout_2198_port, regs(2197) => 
                           bus_reg_dataout_2197_port, regs(2196) => 
                           bus_reg_dataout_2196_port, regs(2195) => 
                           bus_reg_dataout_2195_port, regs(2194) => 
                           bus_reg_dataout_2194_port, regs(2193) => 
                           bus_reg_dataout_2193_port, regs(2192) => 
                           bus_reg_dataout_2192_port, regs(2191) => 
                           bus_reg_dataout_2191_port, regs(2190) => 
                           bus_reg_dataout_2190_port, regs(2189) => 
                           bus_reg_dataout_2189_port, regs(2188) => 
                           bus_reg_dataout_2188_port, regs(2187) => 
                           bus_reg_dataout_2187_port, regs(2186) => 
                           bus_reg_dataout_2186_port, regs(2185) => 
                           bus_reg_dataout_2185_port, regs(2184) => 
                           bus_reg_dataout_2184_port, regs(2183) => 
                           bus_reg_dataout_2183_port, regs(2182) => 
                           bus_reg_dataout_2182_port, regs(2181) => 
                           bus_reg_dataout_2181_port, regs(2180) => 
                           bus_reg_dataout_2180_port, regs(2179) => 
                           bus_reg_dataout_2179_port, regs(2178) => 
                           bus_reg_dataout_2178_port, regs(2177) => 
                           bus_reg_dataout_2177_port, regs(2176) => 
                           bus_reg_dataout_2176_port, regs(2175) => 
                           bus_reg_dataout_2175_port, regs(2174) => 
                           bus_reg_dataout_2174_port, regs(2173) => 
                           bus_reg_dataout_2173_port, regs(2172) => 
                           bus_reg_dataout_2172_port, regs(2171) => 
                           bus_reg_dataout_2171_port, regs(2170) => 
                           bus_reg_dataout_2170_port, regs(2169) => 
                           bus_reg_dataout_2169_port, regs(2168) => 
                           bus_reg_dataout_2168_port, regs(2167) => 
                           bus_reg_dataout_2167_port, regs(2166) => 
                           bus_reg_dataout_2166_port, regs(2165) => 
                           bus_reg_dataout_2165_port, regs(2164) => 
                           bus_reg_dataout_2164_port, regs(2163) => 
                           bus_reg_dataout_2163_port, regs(2162) => 
                           bus_reg_dataout_2162_port, regs(2161) => 
                           bus_reg_dataout_2161_port, regs(2160) => 
                           bus_reg_dataout_2160_port, regs(2159) => 
                           bus_reg_dataout_2159_port, regs(2158) => 
                           bus_reg_dataout_2158_port, regs(2157) => 
                           bus_reg_dataout_2157_port, regs(2156) => 
                           bus_reg_dataout_2156_port, regs(2155) => 
                           bus_reg_dataout_2155_port, regs(2154) => 
                           bus_reg_dataout_2154_port, regs(2153) => 
                           bus_reg_dataout_2153_port, regs(2152) => 
                           bus_reg_dataout_2152_port, regs(2151) => 
                           bus_reg_dataout_2151_port, regs(2150) => 
                           bus_reg_dataout_2150_port, regs(2149) => 
                           bus_reg_dataout_2149_port, regs(2148) => 
                           bus_reg_dataout_2148_port, regs(2147) => 
                           bus_reg_dataout_2147_port, regs(2146) => 
                           bus_reg_dataout_2146_port, regs(2145) => 
                           bus_reg_dataout_2145_port, regs(2144) => 
                           bus_reg_dataout_2144_port, regs(2143) => 
                           bus_reg_dataout_2143_port, regs(2142) => 
                           bus_reg_dataout_2142_port, regs(2141) => 
                           bus_reg_dataout_2141_port, regs(2140) => 
                           bus_reg_dataout_2140_port, regs(2139) => 
                           bus_reg_dataout_2139_port, regs(2138) => 
                           bus_reg_dataout_2138_port, regs(2137) => 
                           bus_reg_dataout_2137_port, regs(2136) => 
                           bus_reg_dataout_2136_port, regs(2135) => 
                           bus_reg_dataout_2135_port, regs(2134) => 
                           bus_reg_dataout_2134_port, regs(2133) => 
                           bus_reg_dataout_2133_port, regs(2132) => 
                           bus_reg_dataout_2132_port, regs(2131) => 
                           bus_reg_dataout_2131_port, regs(2130) => 
                           bus_reg_dataout_2130_port, regs(2129) => 
                           bus_reg_dataout_2129_port, regs(2128) => 
                           bus_reg_dataout_2128_port, regs(2127) => 
                           bus_reg_dataout_2127_port, regs(2126) => 
                           bus_reg_dataout_2126_port, regs(2125) => 
                           bus_reg_dataout_2125_port, regs(2124) => 
                           bus_reg_dataout_2124_port, regs(2123) => 
                           bus_reg_dataout_2123_port, regs(2122) => 
                           bus_reg_dataout_2122_port, regs(2121) => 
                           bus_reg_dataout_2121_port, regs(2120) => 
                           bus_reg_dataout_2120_port, regs(2119) => 
                           bus_reg_dataout_2119_port, regs(2118) => 
                           bus_reg_dataout_2118_port, regs(2117) => 
                           bus_reg_dataout_2117_port, regs(2116) => 
                           bus_reg_dataout_2116_port, regs(2115) => 
                           bus_reg_dataout_2115_port, regs(2114) => 
                           bus_reg_dataout_2114_port, regs(2113) => 
                           bus_reg_dataout_2113_port, regs(2112) => 
                           bus_reg_dataout_2112_port, regs(2111) => 
                           bus_reg_dataout_2111_port, regs(2110) => 
                           bus_reg_dataout_2110_port, regs(2109) => 
                           bus_reg_dataout_2109_port, regs(2108) => 
                           bus_reg_dataout_2108_port, regs(2107) => 
                           bus_reg_dataout_2107_port, regs(2106) => 
                           bus_reg_dataout_2106_port, regs(2105) => 
                           bus_reg_dataout_2105_port, regs(2104) => 
                           bus_reg_dataout_2104_port, regs(2103) => 
                           bus_reg_dataout_2103_port, regs(2102) => 
                           bus_reg_dataout_2102_port, regs(2101) => 
                           bus_reg_dataout_2101_port, regs(2100) => 
                           bus_reg_dataout_2100_port, regs(2099) => 
                           bus_reg_dataout_2099_port, regs(2098) => 
                           bus_reg_dataout_2098_port, regs(2097) => 
                           bus_reg_dataout_2097_port, regs(2096) => 
                           bus_reg_dataout_2096_port, regs(2095) => 
                           bus_reg_dataout_2095_port, regs(2094) => 
                           bus_reg_dataout_2094_port, regs(2093) => 
                           bus_reg_dataout_2093_port, regs(2092) => 
                           bus_reg_dataout_2092_port, regs(2091) => 
                           bus_reg_dataout_2091_port, regs(2090) => 
                           bus_reg_dataout_2090_port, regs(2089) => 
                           bus_reg_dataout_2089_port, regs(2088) => 
                           bus_reg_dataout_2088_port, regs(2087) => 
                           bus_reg_dataout_2087_port, regs(2086) => 
                           bus_reg_dataout_2086_port, regs(2085) => 
                           bus_reg_dataout_2085_port, regs(2084) => 
                           bus_reg_dataout_2084_port, regs(2083) => 
                           bus_reg_dataout_2083_port, regs(2082) => 
                           bus_reg_dataout_2082_port, regs(2081) => 
                           bus_reg_dataout_2081_port, regs(2080) => 
                           bus_reg_dataout_2080_port, regs(2079) => 
                           bus_reg_dataout_2079_port, regs(2078) => 
                           bus_reg_dataout_2078_port, regs(2077) => 
                           bus_reg_dataout_2077_port, regs(2076) => 
                           bus_reg_dataout_2076_port, regs(2075) => 
                           bus_reg_dataout_2075_port, regs(2074) => 
                           bus_reg_dataout_2074_port, regs(2073) => 
                           bus_reg_dataout_2073_port, regs(2072) => 
                           bus_reg_dataout_2072_port, regs(2071) => 
                           bus_reg_dataout_2071_port, regs(2070) => 
                           bus_reg_dataout_2070_port, regs(2069) => 
                           bus_reg_dataout_2069_port, regs(2068) => 
                           bus_reg_dataout_2068_port, regs(2067) => 
                           bus_reg_dataout_2067_port, regs(2066) => 
                           bus_reg_dataout_2066_port, regs(2065) => 
                           bus_reg_dataout_2065_port, regs(2064) => 
                           bus_reg_dataout_2064_port, regs(2063) => 
                           bus_reg_dataout_2063_port, regs(2062) => 
                           bus_reg_dataout_2062_port, regs(2061) => 
                           bus_reg_dataout_2061_port, regs(2060) => 
                           bus_reg_dataout_2060_port, regs(2059) => 
                           bus_reg_dataout_2059_port, regs(2058) => 
                           bus_reg_dataout_2058_port, regs(2057) => 
                           bus_reg_dataout_2057_port, regs(2056) => 
                           bus_reg_dataout_2056_port, regs(2055) => 
                           bus_reg_dataout_2055_port, regs(2054) => 
                           bus_reg_dataout_2054_port, regs(2053) => 
                           bus_reg_dataout_2053_port, regs(2052) => 
                           bus_reg_dataout_2052_port, regs(2051) => 
                           bus_reg_dataout_2051_port, regs(2050) => 
                           bus_reg_dataout_2050_port, regs(2049) => 
                           bus_reg_dataout_2049_port, regs(2048) => 
                           bus_reg_dataout_2048_port, regs(2047) => 
                           bus_reg_dataout_2047_port, regs(2046) => 
                           bus_reg_dataout_2046_port, regs(2045) => 
                           bus_reg_dataout_2045_port, regs(2044) => 
                           bus_reg_dataout_2044_port, regs(2043) => 
                           bus_reg_dataout_2043_port, regs(2042) => 
                           bus_reg_dataout_2042_port, regs(2041) => 
                           bus_reg_dataout_2041_port, regs(2040) => 
                           bus_reg_dataout_2040_port, regs(2039) => 
                           bus_reg_dataout_2039_port, regs(2038) => 
                           bus_reg_dataout_2038_port, regs(2037) => 
                           bus_reg_dataout_2037_port, regs(2036) => 
                           bus_reg_dataout_2036_port, regs(2035) => 
                           bus_reg_dataout_2035_port, regs(2034) => 
                           bus_reg_dataout_2034_port, regs(2033) => 
                           bus_reg_dataout_2033_port, regs(2032) => 
                           bus_reg_dataout_2032_port, regs(2031) => 
                           bus_reg_dataout_2031_port, regs(2030) => 
                           bus_reg_dataout_2030_port, regs(2029) => 
                           bus_reg_dataout_2029_port, regs(2028) => 
                           bus_reg_dataout_2028_port, regs(2027) => 
                           bus_reg_dataout_2027_port, regs(2026) => 
                           bus_reg_dataout_2026_port, regs(2025) => 
                           bus_reg_dataout_2025_port, regs(2024) => 
                           bus_reg_dataout_2024_port, regs(2023) => 
                           bus_reg_dataout_2023_port, regs(2022) => 
                           bus_reg_dataout_2022_port, regs(2021) => 
                           bus_reg_dataout_2021_port, regs(2020) => 
                           bus_reg_dataout_2020_port, regs(2019) => 
                           bus_reg_dataout_2019_port, regs(2018) => 
                           bus_reg_dataout_2018_port, regs(2017) => 
                           bus_reg_dataout_2017_port, regs(2016) => 
                           bus_reg_dataout_2016_port, regs(2015) => 
                           bus_reg_dataout_2015_port, regs(2014) => 
                           bus_reg_dataout_2014_port, regs(2013) => 
                           bus_reg_dataout_2013_port, regs(2012) => 
                           bus_reg_dataout_2012_port, regs(2011) => 
                           bus_reg_dataout_2011_port, regs(2010) => 
                           bus_reg_dataout_2010_port, regs(2009) => 
                           bus_reg_dataout_2009_port, regs(2008) => 
                           bus_reg_dataout_2008_port, regs(2007) => 
                           bus_reg_dataout_2007_port, regs(2006) => 
                           bus_reg_dataout_2006_port, regs(2005) => 
                           bus_reg_dataout_2005_port, regs(2004) => 
                           bus_reg_dataout_2004_port, regs(2003) => 
                           bus_reg_dataout_2003_port, regs(2002) => 
                           bus_reg_dataout_2002_port, regs(2001) => 
                           bus_reg_dataout_2001_port, regs(2000) => 
                           bus_reg_dataout_2000_port, regs(1999) => 
                           bus_reg_dataout_1999_port, regs(1998) => 
                           bus_reg_dataout_1998_port, regs(1997) => 
                           bus_reg_dataout_1997_port, regs(1996) => 
                           bus_reg_dataout_1996_port, regs(1995) => 
                           bus_reg_dataout_1995_port, regs(1994) => 
                           bus_reg_dataout_1994_port, regs(1993) => 
                           bus_reg_dataout_1993_port, regs(1992) => 
                           bus_reg_dataout_1992_port, regs(1991) => 
                           bus_reg_dataout_1991_port, regs(1990) => 
                           bus_reg_dataout_1990_port, regs(1989) => 
                           bus_reg_dataout_1989_port, regs(1988) => 
                           bus_reg_dataout_1988_port, regs(1987) => 
                           bus_reg_dataout_1987_port, regs(1986) => 
                           bus_reg_dataout_1986_port, regs(1985) => 
                           bus_reg_dataout_1985_port, regs(1984) => 
                           bus_reg_dataout_1984_port, regs(1983) => 
                           bus_reg_dataout_1983_port, regs(1982) => 
                           bus_reg_dataout_1982_port, regs(1981) => 
                           bus_reg_dataout_1981_port, regs(1980) => 
                           bus_reg_dataout_1980_port, regs(1979) => 
                           bus_reg_dataout_1979_port, regs(1978) => 
                           bus_reg_dataout_1978_port, regs(1977) => 
                           bus_reg_dataout_1977_port, regs(1976) => 
                           bus_reg_dataout_1976_port, regs(1975) => 
                           bus_reg_dataout_1975_port, regs(1974) => 
                           bus_reg_dataout_1974_port, regs(1973) => 
                           bus_reg_dataout_1973_port, regs(1972) => 
                           bus_reg_dataout_1972_port, regs(1971) => 
                           bus_reg_dataout_1971_port, regs(1970) => 
                           bus_reg_dataout_1970_port, regs(1969) => 
                           bus_reg_dataout_1969_port, regs(1968) => 
                           bus_reg_dataout_1968_port, regs(1967) => 
                           bus_reg_dataout_1967_port, regs(1966) => 
                           bus_reg_dataout_1966_port, regs(1965) => 
                           bus_reg_dataout_1965_port, regs(1964) => 
                           bus_reg_dataout_1964_port, regs(1963) => 
                           bus_reg_dataout_1963_port, regs(1962) => 
                           bus_reg_dataout_1962_port, regs(1961) => 
                           bus_reg_dataout_1961_port, regs(1960) => 
                           bus_reg_dataout_1960_port, regs(1959) => 
                           bus_reg_dataout_1959_port, regs(1958) => 
                           bus_reg_dataout_1958_port, regs(1957) => 
                           bus_reg_dataout_1957_port, regs(1956) => 
                           bus_reg_dataout_1956_port, regs(1955) => 
                           bus_reg_dataout_1955_port, regs(1954) => 
                           bus_reg_dataout_1954_port, regs(1953) => 
                           bus_reg_dataout_1953_port, regs(1952) => 
                           bus_reg_dataout_1952_port, regs(1951) => 
                           bus_reg_dataout_1951_port, regs(1950) => 
                           bus_reg_dataout_1950_port, regs(1949) => 
                           bus_reg_dataout_1949_port, regs(1948) => 
                           bus_reg_dataout_1948_port, regs(1947) => 
                           bus_reg_dataout_1947_port, regs(1946) => 
                           bus_reg_dataout_1946_port, regs(1945) => 
                           bus_reg_dataout_1945_port, regs(1944) => 
                           bus_reg_dataout_1944_port, regs(1943) => 
                           bus_reg_dataout_1943_port, regs(1942) => 
                           bus_reg_dataout_1942_port, regs(1941) => 
                           bus_reg_dataout_1941_port, regs(1940) => 
                           bus_reg_dataout_1940_port, regs(1939) => 
                           bus_reg_dataout_1939_port, regs(1938) => 
                           bus_reg_dataout_1938_port, regs(1937) => 
                           bus_reg_dataout_1937_port, regs(1936) => 
                           bus_reg_dataout_1936_port, regs(1935) => 
                           bus_reg_dataout_1935_port, regs(1934) => 
                           bus_reg_dataout_1934_port, regs(1933) => 
                           bus_reg_dataout_1933_port, regs(1932) => 
                           bus_reg_dataout_1932_port, regs(1931) => 
                           bus_reg_dataout_1931_port, regs(1930) => 
                           bus_reg_dataout_1930_port, regs(1929) => 
                           bus_reg_dataout_1929_port, regs(1928) => 
                           bus_reg_dataout_1928_port, regs(1927) => 
                           bus_reg_dataout_1927_port, regs(1926) => 
                           bus_reg_dataout_1926_port, regs(1925) => 
                           bus_reg_dataout_1925_port, regs(1924) => 
                           bus_reg_dataout_1924_port, regs(1923) => 
                           bus_reg_dataout_1923_port, regs(1922) => 
                           bus_reg_dataout_1922_port, regs(1921) => 
                           bus_reg_dataout_1921_port, regs(1920) => 
                           bus_reg_dataout_1920_port, regs(1919) => 
                           bus_reg_dataout_1919_port, regs(1918) => 
                           bus_reg_dataout_1918_port, regs(1917) => 
                           bus_reg_dataout_1917_port, regs(1916) => 
                           bus_reg_dataout_1916_port, regs(1915) => 
                           bus_reg_dataout_1915_port, regs(1914) => 
                           bus_reg_dataout_1914_port, regs(1913) => 
                           bus_reg_dataout_1913_port, regs(1912) => 
                           bus_reg_dataout_1912_port, regs(1911) => 
                           bus_reg_dataout_1911_port, regs(1910) => 
                           bus_reg_dataout_1910_port, regs(1909) => 
                           bus_reg_dataout_1909_port, regs(1908) => 
                           bus_reg_dataout_1908_port, regs(1907) => 
                           bus_reg_dataout_1907_port, regs(1906) => 
                           bus_reg_dataout_1906_port, regs(1905) => 
                           bus_reg_dataout_1905_port, regs(1904) => 
                           bus_reg_dataout_1904_port, regs(1903) => 
                           bus_reg_dataout_1903_port, regs(1902) => 
                           bus_reg_dataout_1902_port, regs(1901) => 
                           bus_reg_dataout_1901_port, regs(1900) => 
                           bus_reg_dataout_1900_port, regs(1899) => 
                           bus_reg_dataout_1899_port, regs(1898) => 
                           bus_reg_dataout_1898_port, regs(1897) => 
                           bus_reg_dataout_1897_port, regs(1896) => 
                           bus_reg_dataout_1896_port, regs(1895) => 
                           bus_reg_dataout_1895_port, regs(1894) => 
                           bus_reg_dataout_1894_port, regs(1893) => 
                           bus_reg_dataout_1893_port, regs(1892) => 
                           bus_reg_dataout_1892_port, regs(1891) => 
                           bus_reg_dataout_1891_port, regs(1890) => 
                           bus_reg_dataout_1890_port, regs(1889) => 
                           bus_reg_dataout_1889_port, regs(1888) => 
                           bus_reg_dataout_1888_port, regs(1887) => 
                           bus_reg_dataout_1887_port, regs(1886) => 
                           bus_reg_dataout_1886_port, regs(1885) => 
                           bus_reg_dataout_1885_port, regs(1884) => 
                           bus_reg_dataout_1884_port, regs(1883) => 
                           bus_reg_dataout_1883_port, regs(1882) => 
                           bus_reg_dataout_1882_port, regs(1881) => 
                           bus_reg_dataout_1881_port, regs(1880) => 
                           bus_reg_dataout_1880_port, regs(1879) => 
                           bus_reg_dataout_1879_port, regs(1878) => 
                           bus_reg_dataout_1878_port, regs(1877) => 
                           bus_reg_dataout_1877_port, regs(1876) => 
                           bus_reg_dataout_1876_port, regs(1875) => 
                           bus_reg_dataout_1875_port, regs(1874) => 
                           bus_reg_dataout_1874_port, regs(1873) => 
                           bus_reg_dataout_1873_port, regs(1872) => 
                           bus_reg_dataout_1872_port, regs(1871) => 
                           bus_reg_dataout_1871_port, regs(1870) => 
                           bus_reg_dataout_1870_port, regs(1869) => 
                           bus_reg_dataout_1869_port, regs(1868) => 
                           bus_reg_dataout_1868_port, regs(1867) => 
                           bus_reg_dataout_1867_port, regs(1866) => 
                           bus_reg_dataout_1866_port, regs(1865) => 
                           bus_reg_dataout_1865_port, regs(1864) => 
                           bus_reg_dataout_1864_port, regs(1863) => 
                           bus_reg_dataout_1863_port, regs(1862) => 
                           bus_reg_dataout_1862_port, regs(1861) => 
                           bus_reg_dataout_1861_port, regs(1860) => 
                           bus_reg_dataout_1860_port, regs(1859) => 
                           bus_reg_dataout_1859_port, regs(1858) => 
                           bus_reg_dataout_1858_port, regs(1857) => 
                           bus_reg_dataout_1857_port, regs(1856) => 
                           bus_reg_dataout_1856_port, regs(1855) => 
                           bus_reg_dataout_1855_port, regs(1854) => 
                           bus_reg_dataout_1854_port, regs(1853) => 
                           bus_reg_dataout_1853_port, regs(1852) => 
                           bus_reg_dataout_1852_port, regs(1851) => 
                           bus_reg_dataout_1851_port, regs(1850) => 
                           bus_reg_dataout_1850_port, regs(1849) => 
                           bus_reg_dataout_1849_port, regs(1848) => 
                           bus_reg_dataout_1848_port, regs(1847) => 
                           bus_reg_dataout_1847_port, regs(1846) => 
                           bus_reg_dataout_1846_port, regs(1845) => 
                           bus_reg_dataout_1845_port, regs(1844) => 
                           bus_reg_dataout_1844_port, regs(1843) => 
                           bus_reg_dataout_1843_port, regs(1842) => 
                           bus_reg_dataout_1842_port, regs(1841) => 
                           bus_reg_dataout_1841_port, regs(1840) => 
                           bus_reg_dataout_1840_port, regs(1839) => 
                           bus_reg_dataout_1839_port, regs(1838) => 
                           bus_reg_dataout_1838_port, regs(1837) => 
                           bus_reg_dataout_1837_port, regs(1836) => 
                           bus_reg_dataout_1836_port, regs(1835) => 
                           bus_reg_dataout_1835_port, regs(1834) => 
                           bus_reg_dataout_1834_port, regs(1833) => 
                           bus_reg_dataout_1833_port, regs(1832) => 
                           bus_reg_dataout_1832_port, regs(1831) => 
                           bus_reg_dataout_1831_port, regs(1830) => 
                           bus_reg_dataout_1830_port, regs(1829) => 
                           bus_reg_dataout_1829_port, regs(1828) => 
                           bus_reg_dataout_1828_port, regs(1827) => 
                           bus_reg_dataout_1827_port, regs(1826) => 
                           bus_reg_dataout_1826_port, regs(1825) => 
                           bus_reg_dataout_1825_port, regs(1824) => 
                           bus_reg_dataout_1824_port, regs(1823) => 
                           bus_reg_dataout_1823_port, regs(1822) => 
                           bus_reg_dataout_1822_port, regs(1821) => 
                           bus_reg_dataout_1821_port, regs(1820) => 
                           bus_reg_dataout_1820_port, regs(1819) => 
                           bus_reg_dataout_1819_port, regs(1818) => 
                           bus_reg_dataout_1818_port, regs(1817) => 
                           bus_reg_dataout_1817_port, regs(1816) => 
                           bus_reg_dataout_1816_port, regs(1815) => 
                           bus_reg_dataout_1815_port, regs(1814) => 
                           bus_reg_dataout_1814_port, regs(1813) => 
                           bus_reg_dataout_1813_port, regs(1812) => 
                           bus_reg_dataout_1812_port, regs(1811) => 
                           bus_reg_dataout_1811_port, regs(1810) => 
                           bus_reg_dataout_1810_port, regs(1809) => 
                           bus_reg_dataout_1809_port, regs(1808) => 
                           bus_reg_dataout_1808_port, regs(1807) => 
                           bus_reg_dataout_1807_port, regs(1806) => 
                           bus_reg_dataout_1806_port, regs(1805) => 
                           bus_reg_dataout_1805_port, regs(1804) => 
                           bus_reg_dataout_1804_port, regs(1803) => 
                           bus_reg_dataout_1803_port, regs(1802) => 
                           bus_reg_dataout_1802_port, regs(1801) => 
                           bus_reg_dataout_1801_port, regs(1800) => 
                           bus_reg_dataout_1800_port, regs(1799) => 
                           bus_reg_dataout_1799_port, regs(1798) => 
                           bus_reg_dataout_1798_port, regs(1797) => 
                           bus_reg_dataout_1797_port, regs(1796) => 
                           bus_reg_dataout_1796_port, regs(1795) => 
                           bus_reg_dataout_1795_port, regs(1794) => 
                           bus_reg_dataout_1794_port, regs(1793) => 
                           bus_reg_dataout_1793_port, regs(1792) => 
                           bus_reg_dataout_1792_port, regs(1791) => 
                           bus_reg_dataout_1791_port, regs(1790) => 
                           bus_reg_dataout_1790_port, regs(1789) => 
                           bus_reg_dataout_1789_port, regs(1788) => 
                           bus_reg_dataout_1788_port, regs(1787) => 
                           bus_reg_dataout_1787_port, regs(1786) => 
                           bus_reg_dataout_1786_port, regs(1785) => 
                           bus_reg_dataout_1785_port, regs(1784) => 
                           bus_reg_dataout_1784_port, regs(1783) => 
                           bus_reg_dataout_1783_port, regs(1782) => 
                           bus_reg_dataout_1782_port, regs(1781) => 
                           bus_reg_dataout_1781_port, regs(1780) => 
                           bus_reg_dataout_1780_port, regs(1779) => 
                           bus_reg_dataout_1779_port, regs(1778) => 
                           bus_reg_dataout_1778_port, regs(1777) => 
                           bus_reg_dataout_1777_port, regs(1776) => 
                           bus_reg_dataout_1776_port, regs(1775) => 
                           bus_reg_dataout_1775_port, regs(1774) => 
                           bus_reg_dataout_1774_port, regs(1773) => 
                           bus_reg_dataout_1773_port, regs(1772) => 
                           bus_reg_dataout_1772_port, regs(1771) => 
                           bus_reg_dataout_1771_port, regs(1770) => 
                           bus_reg_dataout_1770_port, regs(1769) => 
                           bus_reg_dataout_1769_port, regs(1768) => 
                           bus_reg_dataout_1768_port, regs(1767) => 
                           bus_reg_dataout_1767_port, regs(1766) => 
                           bus_reg_dataout_1766_port, regs(1765) => 
                           bus_reg_dataout_1765_port, regs(1764) => 
                           bus_reg_dataout_1764_port, regs(1763) => 
                           bus_reg_dataout_1763_port, regs(1762) => 
                           bus_reg_dataout_1762_port, regs(1761) => 
                           bus_reg_dataout_1761_port, regs(1760) => 
                           bus_reg_dataout_1760_port, regs(1759) => 
                           bus_reg_dataout_1759_port, regs(1758) => 
                           bus_reg_dataout_1758_port, regs(1757) => 
                           bus_reg_dataout_1757_port, regs(1756) => 
                           bus_reg_dataout_1756_port, regs(1755) => 
                           bus_reg_dataout_1755_port, regs(1754) => 
                           bus_reg_dataout_1754_port, regs(1753) => 
                           bus_reg_dataout_1753_port, regs(1752) => 
                           bus_reg_dataout_1752_port, regs(1751) => 
                           bus_reg_dataout_1751_port, regs(1750) => 
                           bus_reg_dataout_1750_port, regs(1749) => 
                           bus_reg_dataout_1749_port, regs(1748) => 
                           bus_reg_dataout_1748_port, regs(1747) => 
                           bus_reg_dataout_1747_port, regs(1746) => 
                           bus_reg_dataout_1746_port, regs(1745) => 
                           bus_reg_dataout_1745_port, regs(1744) => 
                           bus_reg_dataout_1744_port, regs(1743) => 
                           bus_reg_dataout_1743_port, regs(1742) => 
                           bus_reg_dataout_1742_port, regs(1741) => 
                           bus_reg_dataout_1741_port, regs(1740) => 
                           bus_reg_dataout_1740_port, regs(1739) => 
                           bus_reg_dataout_1739_port, regs(1738) => 
                           bus_reg_dataout_1738_port, regs(1737) => 
                           bus_reg_dataout_1737_port, regs(1736) => 
                           bus_reg_dataout_1736_port, regs(1735) => 
                           bus_reg_dataout_1735_port, regs(1734) => 
                           bus_reg_dataout_1734_port, regs(1733) => 
                           bus_reg_dataout_1733_port, regs(1732) => 
                           bus_reg_dataout_1732_port, regs(1731) => 
                           bus_reg_dataout_1731_port, regs(1730) => 
                           bus_reg_dataout_1730_port, regs(1729) => 
                           bus_reg_dataout_1729_port, regs(1728) => 
                           bus_reg_dataout_1728_port, regs(1727) => 
                           bus_reg_dataout_1727_port, regs(1726) => 
                           bus_reg_dataout_1726_port, regs(1725) => 
                           bus_reg_dataout_1725_port, regs(1724) => 
                           bus_reg_dataout_1724_port, regs(1723) => 
                           bus_reg_dataout_1723_port, regs(1722) => 
                           bus_reg_dataout_1722_port, regs(1721) => 
                           bus_reg_dataout_1721_port, regs(1720) => 
                           bus_reg_dataout_1720_port, regs(1719) => 
                           bus_reg_dataout_1719_port, regs(1718) => 
                           bus_reg_dataout_1718_port, regs(1717) => 
                           bus_reg_dataout_1717_port, regs(1716) => 
                           bus_reg_dataout_1716_port, regs(1715) => 
                           bus_reg_dataout_1715_port, regs(1714) => 
                           bus_reg_dataout_1714_port, regs(1713) => 
                           bus_reg_dataout_1713_port, regs(1712) => 
                           bus_reg_dataout_1712_port, regs(1711) => 
                           bus_reg_dataout_1711_port, regs(1710) => 
                           bus_reg_dataout_1710_port, regs(1709) => 
                           bus_reg_dataout_1709_port, regs(1708) => 
                           bus_reg_dataout_1708_port, regs(1707) => 
                           bus_reg_dataout_1707_port, regs(1706) => 
                           bus_reg_dataout_1706_port, regs(1705) => 
                           bus_reg_dataout_1705_port, regs(1704) => 
                           bus_reg_dataout_1704_port, regs(1703) => 
                           bus_reg_dataout_1703_port, regs(1702) => 
                           bus_reg_dataout_1702_port, regs(1701) => 
                           bus_reg_dataout_1701_port, regs(1700) => 
                           bus_reg_dataout_1700_port, regs(1699) => 
                           bus_reg_dataout_1699_port, regs(1698) => 
                           bus_reg_dataout_1698_port, regs(1697) => 
                           bus_reg_dataout_1697_port, regs(1696) => 
                           bus_reg_dataout_1696_port, regs(1695) => 
                           bus_reg_dataout_1695_port, regs(1694) => 
                           bus_reg_dataout_1694_port, regs(1693) => 
                           bus_reg_dataout_1693_port, regs(1692) => 
                           bus_reg_dataout_1692_port, regs(1691) => 
                           bus_reg_dataout_1691_port, regs(1690) => 
                           bus_reg_dataout_1690_port, regs(1689) => 
                           bus_reg_dataout_1689_port, regs(1688) => 
                           bus_reg_dataout_1688_port, regs(1687) => 
                           bus_reg_dataout_1687_port, regs(1686) => 
                           bus_reg_dataout_1686_port, regs(1685) => 
                           bus_reg_dataout_1685_port, regs(1684) => 
                           bus_reg_dataout_1684_port, regs(1683) => 
                           bus_reg_dataout_1683_port, regs(1682) => 
                           bus_reg_dataout_1682_port, regs(1681) => 
                           bus_reg_dataout_1681_port, regs(1680) => 
                           bus_reg_dataout_1680_port, regs(1679) => 
                           bus_reg_dataout_1679_port, regs(1678) => 
                           bus_reg_dataout_1678_port, regs(1677) => 
                           bus_reg_dataout_1677_port, regs(1676) => 
                           bus_reg_dataout_1676_port, regs(1675) => 
                           bus_reg_dataout_1675_port, regs(1674) => 
                           bus_reg_dataout_1674_port, regs(1673) => 
                           bus_reg_dataout_1673_port, regs(1672) => 
                           bus_reg_dataout_1672_port, regs(1671) => 
                           bus_reg_dataout_1671_port, regs(1670) => 
                           bus_reg_dataout_1670_port, regs(1669) => 
                           bus_reg_dataout_1669_port, regs(1668) => 
                           bus_reg_dataout_1668_port, regs(1667) => 
                           bus_reg_dataout_1667_port, regs(1666) => 
                           bus_reg_dataout_1666_port, regs(1665) => 
                           bus_reg_dataout_1665_port, regs(1664) => 
                           bus_reg_dataout_1664_port, regs(1663) => 
                           bus_reg_dataout_1663_port, regs(1662) => 
                           bus_reg_dataout_1662_port, regs(1661) => 
                           bus_reg_dataout_1661_port, regs(1660) => 
                           bus_reg_dataout_1660_port, regs(1659) => 
                           bus_reg_dataout_1659_port, regs(1658) => 
                           bus_reg_dataout_1658_port, regs(1657) => 
                           bus_reg_dataout_1657_port, regs(1656) => 
                           bus_reg_dataout_1656_port, regs(1655) => 
                           bus_reg_dataout_1655_port, regs(1654) => 
                           bus_reg_dataout_1654_port, regs(1653) => 
                           bus_reg_dataout_1653_port, regs(1652) => 
                           bus_reg_dataout_1652_port, regs(1651) => 
                           bus_reg_dataout_1651_port, regs(1650) => 
                           bus_reg_dataout_1650_port, regs(1649) => 
                           bus_reg_dataout_1649_port, regs(1648) => 
                           bus_reg_dataout_1648_port, regs(1647) => 
                           bus_reg_dataout_1647_port, regs(1646) => 
                           bus_reg_dataout_1646_port, regs(1645) => 
                           bus_reg_dataout_1645_port, regs(1644) => 
                           bus_reg_dataout_1644_port, regs(1643) => 
                           bus_reg_dataout_1643_port, regs(1642) => 
                           bus_reg_dataout_1642_port, regs(1641) => 
                           bus_reg_dataout_1641_port, regs(1640) => 
                           bus_reg_dataout_1640_port, regs(1639) => 
                           bus_reg_dataout_1639_port, regs(1638) => 
                           bus_reg_dataout_1638_port, regs(1637) => 
                           bus_reg_dataout_1637_port, regs(1636) => 
                           bus_reg_dataout_1636_port, regs(1635) => 
                           bus_reg_dataout_1635_port, regs(1634) => 
                           bus_reg_dataout_1634_port, regs(1633) => 
                           bus_reg_dataout_1633_port, regs(1632) => 
                           bus_reg_dataout_1632_port, regs(1631) => 
                           bus_reg_dataout_1631_port, regs(1630) => 
                           bus_reg_dataout_1630_port, regs(1629) => 
                           bus_reg_dataout_1629_port, regs(1628) => 
                           bus_reg_dataout_1628_port, regs(1627) => 
                           bus_reg_dataout_1627_port, regs(1626) => 
                           bus_reg_dataout_1626_port, regs(1625) => 
                           bus_reg_dataout_1625_port, regs(1624) => 
                           bus_reg_dataout_1624_port, regs(1623) => 
                           bus_reg_dataout_1623_port, regs(1622) => 
                           bus_reg_dataout_1622_port, regs(1621) => 
                           bus_reg_dataout_1621_port, regs(1620) => 
                           bus_reg_dataout_1620_port, regs(1619) => 
                           bus_reg_dataout_1619_port, regs(1618) => 
                           bus_reg_dataout_1618_port, regs(1617) => 
                           bus_reg_dataout_1617_port, regs(1616) => 
                           bus_reg_dataout_1616_port, regs(1615) => 
                           bus_reg_dataout_1615_port, regs(1614) => 
                           bus_reg_dataout_1614_port, regs(1613) => 
                           bus_reg_dataout_1613_port, regs(1612) => 
                           bus_reg_dataout_1612_port, regs(1611) => 
                           bus_reg_dataout_1611_port, regs(1610) => 
                           bus_reg_dataout_1610_port, regs(1609) => 
                           bus_reg_dataout_1609_port, regs(1608) => 
                           bus_reg_dataout_1608_port, regs(1607) => 
                           bus_reg_dataout_1607_port, regs(1606) => 
                           bus_reg_dataout_1606_port, regs(1605) => 
                           bus_reg_dataout_1605_port, regs(1604) => 
                           bus_reg_dataout_1604_port, regs(1603) => 
                           bus_reg_dataout_1603_port, regs(1602) => 
                           bus_reg_dataout_1602_port, regs(1601) => 
                           bus_reg_dataout_1601_port, regs(1600) => 
                           bus_reg_dataout_1600_port, regs(1599) => 
                           bus_reg_dataout_1599_port, regs(1598) => 
                           bus_reg_dataout_1598_port, regs(1597) => 
                           bus_reg_dataout_1597_port, regs(1596) => 
                           bus_reg_dataout_1596_port, regs(1595) => 
                           bus_reg_dataout_1595_port, regs(1594) => 
                           bus_reg_dataout_1594_port, regs(1593) => 
                           bus_reg_dataout_1593_port, regs(1592) => 
                           bus_reg_dataout_1592_port, regs(1591) => 
                           bus_reg_dataout_1591_port, regs(1590) => 
                           bus_reg_dataout_1590_port, regs(1589) => 
                           bus_reg_dataout_1589_port, regs(1588) => 
                           bus_reg_dataout_1588_port, regs(1587) => 
                           bus_reg_dataout_1587_port, regs(1586) => 
                           bus_reg_dataout_1586_port, regs(1585) => 
                           bus_reg_dataout_1585_port, regs(1584) => 
                           bus_reg_dataout_1584_port, regs(1583) => 
                           bus_reg_dataout_1583_port, regs(1582) => 
                           bus_reg_dataout_1582_port, regs(1581) => 
                           bus_reg_dataout_1581_port, regs(1580) => 
                           bus_reg_dataout_1580_port, regs(1579) => 
                           bus_reg_dataout_1579_port, regs(1578) => 
                           bus_reg_dataout_1578_port, regs(1577) => 
                           bus_reg_dataout_1577_port, regs(1576) => 
                           bus_reg_dataout_1576_port, regs(1575) => 
                           bus_reg_dataout_1575_port, regs(1574) => 
                           bus_reg_dataout_1574_port, regs(1573) => 
                           bus_reg_dataout_1573_port, regs(1572) => 
                           bus_reg_dataout_1572_port, regs(1571) => 
                           bus_reg_dataout_1571_port, regs(1570) => 
                           bus_reg_dataout_1570_port, regs(1569) => 
                           bus_reg_dataout_1569_port, regs(1568) => 
                           bus_reg_dataout_1568_port, regs(1567) => 
                           bus_reg_dataout_1567_port, regs(1566) => 
                           bus_reg_dataout_1566_port, regs(1565) => 
                           bus_reg_dataout_1565_port, regs(1564) => 
                           bus_reg_dataout_1564_port, regs(1563) => 
                           bus_reg_dataout_1563_port, regs(1562) => 
                           bus_reg_dataout_1562_port, regs(1561) => 
                           bus_reg_dataout_1561_port, regs(1560) => 
                           bus_reg_dataout_1560_port, regs(1559) => 
                           bus_reg_dataout_1559_port, regs(1558) => 
                           bus_reg_dataout_1558_port, regs(1557) => 
                           bus_reg_dataout_1557_port, regs(1556) => 
                           bus_reg_dataout_1556_port, regs(1555) => 
                           bus_reg_dataout_1555_port, regs(1554) => 
                           bus_reg_dataout_1554_port, regs(1553) => 
                           bus_reg_dataout_1553_port, regs(1552) => 
                           bus_reg_dataout_1552_port, regs(1551) => 
                           bus_reg_dataout_1551_port, regs(1550) => 
                           bus_reg_dataout_1550_port, regs(1549) => 
                           bus_reg_dataout_1549_port, regs(1548) => 
                           bus_reg_dataout_1548_port, regs(1547) => 
                           bus_reg_dataout_1547_port, regs(1546) => 
                           bus_reg_dataout_1546_port, regs(1545) => 
                           bus_reg_dataout_1545_port, regs(1544) => 
                           bus_reg_dataout_1544_port, regs(1543) => 
                           bus_reg_dataout_1543_port, regs(1542) => 
                           bus_reg_dataout_1542_port, regs(1541) => 
                           bus_reg_dataout_1541_port, regs(1540) => 
                           bus_reg_dataout_1540_port, regs(1539) => 
                           bus_reg_dataout_1539_port, regs(1538) => 
                           bus_reg_dataout_1538_port, regs(1537) => 
                           bus_reg_dataout_1537_port, regs(1536) => 
                           bus_reg_dataout_1536_port, regs(1535) => 
                           bus_reg_dataout_1535_port, regs(1534) => 
                           bus_reg_dataout_1534_port, regs(1533) => 
                           bus_reg_dataout_1533_port, regs(1532) => 
                           bus_reg_dataout_1532_port, regs(1531) => 
                           bus_reg_dataout_1531_port, regs(1530) => 
                           bus_reg_dataout_1530_port, regs(1529) => 
                           bus_reg_dataout_1529_port, regs(1528) => 
                           bus_reg_dataout_1528_port, regs(1527) => 
                           bus_reg_dataout_1527_port, regs(1526) => 
                           bus_reg_dataout_1526_port, regs(1525) => 
                           bus_reg_dataout_1525_port, regs(1524) => 
                           bus_reg_dataout_1524_port, regs(1523) => 
                           bus_reg_dataout_1523_port, regs(1522) => 
                           bus_reg_dataout_1522_port, regs(1521) => 
                           bus_reg_dataout_1521_port, regs(1520) => 
                           bus_reg_dataout_1520_port, regs(1519) => 
                           bus_reg_dataout_1519_port, regs(1518) => 
                           bus_reg_dataout_1518_port, regs(1517) => 
                           bus_reg_dataout_1517_port, regs(1516) => 
                           bus_reg_dataout_1516_port, regs(1515) => 
                           bus_reg_dataout_1515_port, regs(1514) => 
                           bus_reg_dataout_1514_port, regs(1513) => 
                           bus_reg_dataout_1513_port, regs(1512) => 
                           bus_reg_dataout_1512_port, regs(1511) => 
                           bus_reg_dataout_1511_port, regs(1510) => 
                           bus_reg_dataout_1510_port, regs(1509) => 
                           bus_reg_dataout_1509_port, regs(1508) => 
                           bus_reg_dataout_1508_port, regs(1507) => 
                           bus_reg_dataout_1507_port, regs(1506) => 
                           bus_reg_dataout_1506_port, regs(1505) => 
                           bus_reg_dataout_1505_port, regs(1504) => 
                           bus_reg_dataout_1504_port, regs(1503) => 
                           bus_reg_dataout_1503_port, regs(1502) => 
                           bus_reg_dataout_1502_port, regs(1501) => 
                           bus_reg_dataout_1501_port, regs(1500) => 
                           bus_reg_dataout_1500_port, regs(1499) => 
                           bus_reg_dataout_1499_port, regs(1498) => 
                           bus_reg_dataout_1498_port, regs(1497) => 
                           bus_reg_dataout_1497_port, regs(1496) => 
                           bus_reg_dataout_1496_port, regs(1495) => 
                           bus_reg_dataout_1495_port, regs(1494) => 
                           bus_reg_dataout_1494_port, regs(1493) => 
                           bus_reg_dataout_1493_port, regs(1492) => 
                           bus_reg_dataout_1492_port, regs(1491) => 
                           bus_reg_dataout_1491_port, regs(1490) => 
                           bus_reg_dataout_1490_port, regs(1489) => 
                           bus_reg_dataout_1489_port, regs(1488) => 
                           bus_reg_dataout_1488_port, regs(1487) => 
                           bus_reg_dataout_1487_port, regs(1486) => 
                           bus_reg_dataout_1486_port, regs(1485) => 
                           bus_reg_dataout_1485_port, regs(1484) => 
                           bus_reg_dataout_1484_port, regs(1483) => 
                           bus_reg_dataout_1483_port, regs(1482) => 
                           bus_reg_dataout_1482_port, regs(1481) => 
                           bus_reg_dataout_1481_port, regs(1480) => 
                           bus_reg_dataout_1480_port, regs(1479) => 
                           bus_reg_dataout_1479_port, regs(1478) => 
                           bus_reg_dataout_1478_port, regs(1477) => 
                           bus_reg_dataout_1477_port, regs(1476) => 
                           bus_reg_dataout_1476_port, regs(1475) => 
                           bus_reg_dataout_1475_port, regs(1474) => 
                           bus_reg_dataout_1474_port, regs(1473) => 
                           bus_reg_dataout_1473_port, regs(1472) => 
                           bus_reg_dataout_1472_port, regs(1471) => 
                           bus_reg_dataout_1471_port, regs(1470) => 
                           bus_reg_dataout_1470_port, regs(1469) => 
                           bus_reg_dataout_1469_port, regs(1468) => 
                           bus_reg_dataout_1468_port, regs(1467) => 
                           bus_reg_dataout_1467_port, regs(1466) => 
                           bus_reg_dataout_1466_port, regs(1465) => 
                           bus_reg_dataout_1465_port, regs(1464) => 
                           bus_reg_dataout_1464_port, regs(1463) => 
                           bus_reg_dataout_1463_port, regs(1462) => 
                           bus_reg_dataout_1462_port, regs(1461) => 
                           bus_reg_dataout_1461_port, regs(1460) => 
                           bus_reg_dataout_1460_port, regs(1459) => 
                           bus_reg_dataout_1459_port, regs(1458) => 
                           bus_reg_dataout_1458_port, regs(1457) => 
                           bus_reg_dataout_1457_port, regs(1456) => 
                           bus_reg_dataout_1456_port, regs(1455) => 
                           bus_reg_dataout_1455_port, regs(1454) => 
                           bus_reg_dataout_1454_port, regs(1453) => 
                           bus_reg_dataout_1453_port, regs(1452) => 
                           bus_reg_dataout_1452_port, regs(1451) => 
                           bus_reg_dataout_1451_port, regs(1450) => 
                           bus_reg_dataout_1450_port, regs(1449) => 
                           bus_reg_dataout_1449_port, regs(1448) => 
                           bus_reg_dataout_1448_port, regs(1447) => 
                           bus_reg_dataout_1447_port, regs(1446) => 
                           bus_reg_dataout_1446_port, regs(1445) => 
                           bus_reg_dataout_1445_port, regs(1444) => 
                           bus_reg_dataout_1444_port, regs(1443) => 
                           bus_reg_dataout_1443_port, regs(1442) => 
                           bus_reg_dataout_1442_port, regs(1441) => 
                           bus_reg_dataout_1441_port, regs(1440) => 
                           bus_reg_dataout_1440_port, regs(1439) => 
                           bus_reg_dataout_1439_port, regs(1438) => 
                           bus_reg_dataout_1438_port, regs(1437) => 
                           bus_reg_dataout_1437_port, regs(1436) => 
                           bus_reg_dataout_1436_port, regs(1435) => 
                           bus_reg_dataout_1435_port, regs(1434) => 
                           bus_reg_dataout_1434_port, regs(1433) => 
                           bus_reg_dataout_1433_port, regs(1432) => 
                           bus_reg_dataout_1432_port, regs(1431) => 
                           bus_reg_dataout_1431_port, regs(1430) => 
                           bus_reg_dataout_1430_port, regs(1429) => 
                           bus_reg_dataout_1429_port, regs(1428) => 
                           bus_reg_dataout_1428_port, regs(1427) => 
                           bus_reg_dataout_1427_port, regs(1426) => 
                           bus_reg_dataout_1426_port, regs(1425) => 
                           bus_reg_dataout_1425_port, regs(1424) => 
                           bus_reg_dataout_1424_port, regs(1423) => 
                           bus_reg_dataout_1423_port, regs(1422) => 
                           bus_reg_dataout_1422_port, regs(1421) => 
                           bus_reg_dataout_1421_port, regs(1420) => 
                           bus_reg_dataout_1420_port, regs(1419) => 
                           bus_reg_dataout_1419_port, regs(1418) => 
                           bus_reg_dataout_1418_port, regs(1417) => 
                           bus_reg_dataout_1417_port, regs(1416) => 
                           bus_reg_dataout_1416_port, regs(1415) => 
                           bus_reg_dataout_1415_port, regs(1414) => 
                           bus_reg_dataout_1414_port, regs(1413) => 
                           bus_reg_dataout_1413_port, regs(1412) => 
                           bus_reg_dataout_1412_port, regs(1411) => 
                           bus_reg_dataout_1411_port, regs(1410) => 
                           bus_reg_dataout_1410_port, regs(1409) => 
                           bus_reg_dataout_1409_port, regs(1408) => 
                           bus_reg_dataout_1408_port, regs(1407) => 
                           bus_reg_dataout_1407_port, regs(1406) => 
                           bus_reg_dataout_1406_port, regs(1405) => 
                           bus_reg_dataout_1405_port, regs(1404) => 
                           bus_reg_dataout_1404_port, regs(1403) => 
                           bus_reg_dataout_1403_port, regs(1402) => 
                           bus_reg_dataout_1402_port, regs(1401) => 
                           bus_reg_dataout_1401_port, regs(1400) => 
                           bus_reg_dataout_1400_port, regs(1399) => 
                           bus_reg_dataout_1399_port, regs(1398) => 
                           bus_reg_dataout_1398_port, regs(1397) => 
                           bus_reg_dataout_1397_port, regs(1396) => 
                           bus_reg_dataout_1396_port, regs(1395) => 
                           bus_reg_dataout_1395_port, regs(1394) => 
                           bus_reg_dataout_1394_port, regs(1393) => 
                           bus_reg_dataout_1393_port, regs(1392) => 
                           bus_reg_dataout_1392_port, regs(1391) => 
                           bus_reg_dataout_1391_port, regs(1390) => 
                           bus_reg_dataout_1390_port, regs(1389) => 
                           bus_reg_dataout_1389_port, regs(1388) => 
                           bus_reg_dataout_1388_port, regs(1387) => 
                           bus_reg_dataout_1387_port, regs(1386) => 
                           bus_reg_dataout_1386_port, regs(1385) => 
                           bus_reg_dataout_1385_port, regs(1384) => 
                           bus_reg_dataout_1384_port, regs(1383) => 
                           bus_reg_dataout_1383_port, regs(1382) => 
                           bus_reg_dataout_1382_port, regs(1381) => 
                           bus_reg_dataout_1381_port, regs(1380) => 
                           bus_reg_dataout_1380_port, regs(1379) => 
                           bus_reg_dataout_1379_port, regs(1378) => 
                           bus_reg_dataout_1378_port, regs(1377) => 
                           bus_reg_dataout_1377_port, regs(1376) => 
                           bus_reg_dataout_1376_port, regs(1375) => 
                           bus_reg_dataout_1375_port, regs(1374) => 
                           bus_reg_dataout_1374_port, regs(1373) => 
                           bus_reg_dataout_1373_port, regs(1372) => 
                           bus_reg_dataout_1372_port, regs(1371) => 
                           bus_reg_dataout_1371_port, regs(1370) => 
                           bus_reg_dataout_1370_port, regs(1369) => 
                           bus_reg_dataout_1369_port, regs(1368) => 
                           bus_reg_dataout_1368_port, regs(1367) => 
                           bus_reg_dataout_1367_port, regs(1366) => 
                           bus_reg_dataout_1366_port, regs(1365) => 
                           bus_reg_dataout_1365_port, regs(1364) => 
                           bus_reg_dataout_1364_port, regs(1363) => 
                           bus_reg_dataout_1363_port, regs(1362) => 
                           bus_reg_dataout_1362_port, regs(1361) => 
                           bus_reg_dataout_1361_port, regs(1360) => 
                           bus_reg_dataout_1360_port, regs(1359) => 
                           bus_reg_dataout_1359_port, regs(1358) => 
                           bus_reg_dataout_1358_port, regs(1357) => 
                           bus_reg_dataout_1357_port, regs(1356) => 
                           bus_reg_dataout_1356_port, regs(1355) => 
                           bus_reg_dataout_1355_port, regs(1354) => 
                           bus_reg_dataout_1354_port, regs(1353) => 
                           bus_reg_dataout_1353_port, regs(1352) => 
                           bus_reg_dataout_1352_port, regs(1351) => 
                           bus_reg_dataout_1351_port, regs(1350) => 
                           bus_reg_dataout_1350_port, regs(1349) => 
                           bus_reg_dataout_1349_port, regs(1348) => 
                           bus_reg_dataout_1348_port, regs(1347) => 
                           bus_reg_dataout_1347_port, regs(1346) => 
                           bus_reg_dataout_1346_port, regs(1345) => 
                           bus_reg_dataout_1345_port, regs(1344) => 
                           bus_reg_dataout_1344_port, regs(1343) => 
                           bus_reg_dataout_1343_port, regs(1342) => 
                           bus_reg_dataout_1342_port, regs(1341) => 
                           bus_reg_dataout_1341_port, regs(1340) => 
                           bus_reg_dataout_1340_port, regs(1339) => 
                           bus_reg_dataout_1339_port, regs(1338) => 
                           bus_reg_dataout_1338_port, regs(1337) => 
                           bus_reg_dataout_1337_port, regs(1336) => 
                           bus_reg_dataout_1336_port, regs(1335) => 
                           bus_reg_dataout_1335_port, regs(1334) => 
                           bus_reg_dataout_1334_port, regs(1333) => 
                           bus_reg_dataout_1333_port, regs(1332) => 
                           bus_reg_dataout_1332_port, regs(1331) => 
                           bus_reg_dataout_1331_port, regs(1330) => 
                           bus_reg_dataout_1330_port, regs(1329) => 
                           bus_reg_dataout_1329_port, regs(1328) => 
                           bus_reg_dataout_1328_port, regs(1327) => 
                           bus_reg_dataout_1327_port, regs(1326) => 
                           bus_reg_dataout_1326_port, regs(1325) => 
                           bus_reg_dataout_1325_port, regs(1324) => 
                           bus_reg_dataout_1324_port, regs(1323) => 
                           bus_reg_dataout_1323_port, regs(1322) => 
                           bus_reg_dataout_1322_port, regs(1321) => 
                           bus_reg_dataout_1321_port, regs(1320) => 
                           bus_reg_dataout_1320_port, regs(1319) => 
                           bus_reg_dataout_1319_port, regs(1318) => 
                           bus_reg_dataout_1318_port, regs(1317) => 
                           bus_reg_dataout_1317_port, regs(1316) => 
                           bus_reg_dataout_1316_port, regs(1315) => 
                           bus_reg_dataout_1315_port, regs(1314) => 
                           bus_reg_dataout_1314_port, regs(1313) => 
                           bus_reg_dataout_1313_port, regs(1312) => 
                           bus_reg_dataout_1312_port, regs(1311) => 
                           bus_reg_dataout_1311_port, regs(1310) => 
                           bus_reg_dataout_1310_port, regs(1309) => 
                           bus_reg_dataout_1309_port, regs(1308) => 
                           bus_reg_dataout_1308_port, regs(1307) => 
                           bus_reg_dataout_1307_port, regs(1306) => 
                           bus_reg_dataout_1306_port, regs(1305) => 
                           bus_reg_dataout_1305_port, regs(1304) => 
                           bus_reg_dataout_1304_port, regs(1303) => 
                           bus_reg_dataout_1303_port, regs(1302) => 
                           bus_reg_dataout_1302_port, regs(1301) => 
                           bus_reg_dataout_1301_port, regs(1300) => 
                           bus_reg_dataout_1300_port, regs(1299) => 
                           bus_reg_dataout_1299_port, regs(1298) => 
                           bus_reg_dataout_1298_port, regs(1297) => 
                           bus_reg_dataout_1297_port, regs(1296) => 
                           bus_reg_dataout_1296_port, regs(1295) => 
                           bus_reg_dataout_1295_port, regs(1294) => 
                           bus_reg_dataout_1294_port, regs(1293) => 
                           bus_reg_dataout_1293_port, regs(1292) => 
                           bus_reg_dataout_1292_port, regs(1291) => 
                           bus_reg_dataout_1291_port, regs(1290) => 
                           bus_reg_dataout_1290_port, regs(1289) => 
                           bus_reg_dataout_1289_port, regs(1288) => 
                           bus_reg_dataout_1288_port, regs(1287) => 
                           bus_reg_dataout_1287_port, regs(1286) => 
                           bus_reg_dataout_1286_port, regs(1285) => 
                           bus_reg_dataout_1285_port, regs(1284) => 
                           bus_reg_dataout_1284_port, regs(1283) => 
                           bus_reg_dataout_1283_port, regs(1282) => 
                           bus_reg_dataout_1282_port, regs(1281) => 
                           bus_reg_dataout_1281_port, regs(1280) => 
                           bus_reg_dataout_1280_port, regs(1279) => 
                           bus_reg_dataout_1279_port, regs(1278) => 
                           bus_reg_dataout_1278_port, regs(1277) => 
                           bus_reg_dataout_1277_port, regs(1276) => 
                           bus_reg_dataout_1276_port, regs(1275) => 
                           bus_reg_dataout_1275_port, regs(1274) => 
                           bus_reg_dataout_1274_port, regs(1273) => 
                           bus_reg_dataout_1273_port, regs(1272) => 
                           bus_reg_dataout_1272_port, regs(1271) => 
                           bus_reg_dataout_1271_port, regs(1270) => 
                           bus_reg_dataout_1270_port, regs(1269) => 
                           bus_reg_dataout_1269_port, regs(1268) => 
                           bus_reg_dataout_1268_port, regs(1267) => 
                           bus_reg_dataout_1267_port, regs(1266) => 
                           bus_reg_dataout_1266_port, regs(1265) => 
                           bus_reg_dataout_1265_port, regs(1264) => 
                           bus_reg_dataout_1264_port, regs(1263) => 
                           bus_reg_dataout_1263_port, regs(1262) => 
                           bus_reg_dataout_1262_port, regs(1261) => 
                           bus_reg_dataout_1261_port, regs(1260) => 
                           bus_reg_dataout_1260_port, regs(1259) => 
                           bus_reg_dataout_1259_port, regs(1258) => 
                           bus_reg_dataout_1258_port, regs(1257) => 
                           bus_reg_dataout_1257_port, regs(1256) => 
                           bus_reg_dataout_1256_port, regs(1255) => 
                           bus_reg_dataout_1255_port, regs(1254) => 
                           bus_reg_dataout_1254_port, regs(1253) => 
                           bus_reg_dataout_1253_port, regs(1252) => 
                           bus_reg_dataout_1252_port, regs(1251) => 
                           bus_reg_dataout_1251_port, regs(1250) => 
                           bus_reg_dataout_1250_port, regs(1249) => 
                           bus_reg_dataout_1249_port, regs(1248) => 
                           bus_reg_dataout_1248_port, regs(1247) => 
                           bus_reg_dataout_1247_port, regs(1246) => 
                           bus_reg_dataout_1246_port, regs(1245) => 
                           bus_reg_dataout_1245_port, regs(1244) => 
                           bus_reg_dataout_1244_port, regs(1243) => 
                           bus_reg_dataout_1243_port, regs(1242) => 
                           bus_reg_dataout_1242_port, regs(1241) => 
                           bus_reg_dataout_1241_port, regs(1240) => 
                           bus_reg_dataout_1240_port, regs(1239) => 
                           bus_reg_dataout_1239_port, regs(1238) => 
                           bus_reg_dataout_1238_port, regs(1237) => 
                           bus_reg_dataout_1237_port, regs(1236) => 
                           bus_reg_dataout_1236_port, regs(1235) => 
                           bus_reg_dataout_1235_port, regs(1234) => 
                           bus_reg_dataout_1234_port, regs(1233) => 
                           bus_reg_dataout_1233_port, regs(1232) => 
                           bus_reg_dataout_1232_port, regs(1231) => 
                           bus_reg_dataout_1231_port, regs(1230) => 
                           bus_reg_dataout_1230_port, regs(1229) => 
                           bus_reg_dataout_1229_port, regs(1228) => 
                           bus_reg_dataout_1228_port, regs(1227) => 
                           bus_reg_dataout_1227_port, regs(1226) => 
                           bus_reg_dataout_1226_port, regs(1225) => 
                           bus_reg_dataout_1225_port, regs(1224) => 
                           bus_reg_dataout_1224_port, regs(1223) => 
                           bus_reg_dataout_1223_port, regs(1222) => 
                           bus_reg_dataout_1222_port, regs(1221) => 
                           bus_reg_dataout_1221_port, regs(1220) => 
                           bus_reg_dataout_1220_port, regs(1219) => 
                           bus_reg_dataout_1219_port, regs(1218) => 
                           bus_reg_dataout_1218_port, regs(1217) => 
                           bus_reg_dataout_1217_port, regs(1216) => 
                           bus_reg_dataout_1216_port, regs(1215) => 
                           bus_reg_dataout_1215_port, regs(1214) => 
                           bus_reg_dataout_1214_port, regs(1213) => 
                           bus_reg_dataout_1213_port, regs(1212) => 
                           bus_reg_dataout_1212_port, regs(1211) => 
                           bus_reg_dataout_1211_port, regs(1210) => 
                           bus_reg_dataout_1210_port, regs(1209) => 
                           bus_reg_dataout_1209_port, regs(1208) => 
                           bus_reg_dataout_1208_port, regs(1207) => 
                           bus_reg_dataout_1207_port, regs(1206) => 
                           bus_reg_dataout_1206_port, regs(1205) => 
                           bus_reg_dataout_1205_port, regs(1204) => 
                           bus_reg_dataout_1204_port, regs(1203) => 
                           bus_reg_dataout_1203_port, regs(1202) => 
                           bus_reg_dataout_1202_port, regs(1201) => 
                           bus_reg_dataout_1201_port, regs(1200) => 
                           bus_reg_dataout_1200_port, regs(1199) => 
                           bus_reg_dataout_1199_port, regs(1198) => 
                           bus_reg_dataout_1198_port, regs(1197) => 
                           bus_reg_dataout_1197_port, regs(1196) => 
                           bus_reg_dataout_1196_port, regs(1195) => 
                           bus_reg_dataout_1195_port, regs(1194) => 
                           bus_reg_dataout_1194_port, regs(1193) => 
                           bus_reg_dataout_1193_port, regs(1192) => 
                           bus_reg_dataout_1192_port, regs(1191) => 
                           bus_reg_dataout_1191_port, regs(1190) => 
                           bus_reg_dataout_1190_port, regs(1189) => 
                           bus_reg_dataout_1189_port, regs(1188) => 
                           bus_reg_dataout_1188_port, regs(1187) => 
                           bus_reg_dataout_1187_port, regs(1186) => 
                           bus_reg_dataout_1186_port, regs(1185) => 
                           bus_reg_dataout_1185_port, regs(1184) => 
                           bus_reg_dataout_1184_port, regs(1183) => 
                           bus_reg_dataout_1183_port, regs(1182) => 
                           bus_reg_dataout_1182_port, regs(1181) => 
                           bus_reg_dataout_1181_port, regs(1180) => 
                           bus_reg_dataout_1180_port, regs(1179) => 
                           bus_reg_dataout_1179_port, regs(1178) => 
                           bus_reg_dataout_1178_port, regs(1177) => 
                           bus_reg_dataout_1177_port, regs(1176) => 
                           bus_reg_dataout_1176_port, regs(1175) => 
                           bus_reg_dataout_1175_port, regs(1174) => 
                           bus_reg_dataout_1174_port, regs(1173) => 
                           bus_reg_dataout_1173_port, regs(1172) => 
                           bus_reg_dataout_1172_port, regs(1171) => 
                           bus_reg_dataout_1171_port, regs(1170) => 
                           bus_reg_dataout_1170_port, regs(1169) => 
                           bus_reg_dataout_1169_port, regs(1168) => 
                           bus_reg_dataout_1168_port, regs(1167) => 
                           bus_reg_dataout_1167_port, regs(1166) => 
                           bus_reg_dataout_1166_port, regs(1165) => 
                           bus_reg_dataout_1165_port, regs(1164) => 
                           bus_reg_dataout_1164_port, regs(1163) => 
                           bus_reg_dataout_1163_port, regs(1162) => 
                           bus_reg_dataout_1162_port, regs(1161) => 
                           bus_reg_dataout_1161_port, regs(1160) => 
                           bus_reg_dataout_1160_port, regs(1159) => 
                           bus_reg_dataout_1159_port, regs(1158) => 
                           bus_reg_dataout_1158_port, regs(1157) => 
                           bus_reg_dataout_1157_port, regs(1156) => 
                           bus_reg_dataout_1156_port, regs(1155) => 
                           bus_reg_dataout_1155_port, regs(1154) => 
                           bus_reg_dataout_1154_port, regs(1153) => 
                           bus_reg_dataout_1153_port, regs(1152) => 
                           bus_reg_dataout_1152_port, regs(1151) => 
                           bus_reg_dataout_1151_port, regs(1150) => 
                           bus_reg_dataout_1150_port, regs(1149) => 
                           bus_reg_dataout_1149_port, regs(1148) => 
                           bus_reg_dataout_1148_port, regs(1147) => 
                           bus_reg_dataout_1147_port, regs(1146) => 
                           bus_reg_dataout_1146_port, regs(1145) => 
                           bus_reg_dataout_1145_port, regs(1144) => 
                           bus_reg_dataout_1144_port, regs(1143) => 
                           bus_reg_dataout_1143_port, regs(1142) => 
                           bus_reg_dataout_1142_port, regs(1141) => 
                           bus_reg_dataout_1141_port, regs(1140) => 
                           bus_reg_dataout_1140_port, regs(1139) => 
                           bus_reg_dataout_1139_port, regs(1138) => 
                           bus_reg_dataout_1138_port, regs(1137) => 
                           bus_reg_dataout_1137_port, regs(1136) => 
                           bus_reg_dataout_1136_port, regs(1135) => 
                           bus_reg_dataout_1135_port, regs(1134) => 
                           bus_reg_dataout_1134_port, regs(1133) => 
                           bus_reg_dataout_1133_port, regs(1132) => 
                           bus_reg_dataout_1132_port, regs(1131) => 
                           bus_reg_dataout_1131_port, regs(1130) => 
                           bus_reg_dataout_1130_port, regs(1129) => 
                           bus_reg_dataout_1129_port, regs(1128) => 
                           bus_reg_dataout_1128_port, regs(1127) => 
                           bus_reg_dataout_1127_port, regs(1126) => 
                           bus_reg_dataout_1126_port, regs(1125) => 
                           bus_reg_dataout_1125_port, regs(1124) => 
                           bus_reg_dataout_1124_port, regs(1123) => 
                           bus_reg_dataout_1123_port, regs(1122) => 
                           bus_reg_dataout_1122_port, regs(1121) => 
                           bus_reg_dataout_1121_port, regs(1120) => 
                           bus_reg_dataout_1120_port, regs(1119) => 
                           bus_reg_dataout_1119_port, regs(1118) => 
                           bus_reg_dataout_1118_port, regs(1117) => 
                           bus_reg_dataout_1117_port, regs(1116) => 
                           bus_reg_dataout_1116_port, regs(1115) => 
                           bus_reg_dataout_1115_port, regs(1114) => 
                           bus_reg_dataout_1114_port, regs(1113) => 
                           bus_reg_dataout_1113_port, regs(1112) => 
                           bus_reg_dataout_1112_port, regs(1111) => 
                           bus_reg_dataout_1111_port, regs(1110) => 
                           bus_reg_dataout_1110_port, regs(1109) => 
                           bus_reg_dataout_1109_port, regs(1108) => 
                           bus_reg_dataout_1108_port, regs(1107) => 
                           bus_reg_dataout_1107_port, regs(1106) => 
                           bus_reg_dataout_1106_port, regs(1105) => 
                           bus_reg_dataout_1105_port, regs(1104) => 
                           bus_reg_dataout_1104_port, regs(1103) => 
                           bus_reg_dataout_1103_port, regs(1102) => 
                           bus_reg_dataout_1102_port, regs(1101) => 
                           bus_reg_dataout_1101_port, regs(1100) => 
                           bus_reg_dataout_1100_port, regs(1099) => 
                           bus_reg_dataout_1099_port, regs(1098) => 
                           bus_reg_dataout_1098_port, regs(1097) => 
                           bus_reg_dataout_1097_port, regs(1096) => 
                           bus_reg_dataout_1096_port, regs(1095) => 
                           bus_reg_dataout_1095_port, regs(1094) => 
                           bus_reg_dataout_1094_port, regs(1093) => 
                           bus_reg_dataout_1093_port, regs(1092) => 
                           bus_reg_dataout_1092_port, regs(1091) => 
                           bus_reg_dataout_1091_port, regs(1090) => 
                           bus_reg_dataout_1090_port, regs(1089) => 
                           bus_reg_dataout_1089_port, regs(1088) => 
                           bus_reg_dataout_1088_port, regs(1087) => 
                           bus_reg_dataout_1087_port, regs(1086) => 
                           bus_reg_dataout_1086_port, regs(1085) => 
                           bus_reg_dataout_1085_port, regs(1084) => 
                           bus_reg_dataout_1084_port, regs(1083) => 
                           bus_reg_dataout_1083_port, regs(1082) => 
                           bus_reg_dataout_1082_port, regs(1081) => 
                           bus_reg_dataout_1081_port, regs(1080) => 
                           bus_reg_dataout_1080_port, regs(1079) => 
                           bus_reg_dataout_1079_port, regs(1078) => 
                           bus_reg_dataout_1078_port, regs(1077) => 
                           bus_reg_dataout_1077_port, regs(1076) => 
                           bus_reg_dataout_1076_port, regs(1075) => 
                           bus_reg_dataout_1075_port, regs(1074) => 
                           bus_reg_dataout_1074_port, regs(1073) => 
                           bus_reg_dataout_1073_port, regs(1072) => 
                           bus_reg_dataout_1072_port, regs(1071) => 
                           bus_reg_dataout_1071_port, regs(1070) => 
                           bus_reg_dataout_1070_port, regs(1069) => 
                           bus_reg_dataout_1069_port, regs(1068) => 
                           bus_reg_dataout_1068_port, regs(1067) => 
                           bus_reg_dataout_1067_port, regs(1066) => 
                           bus_reg_dataout_1066_port, regs(1065) => 
                           bus_reg_dataout_1065_port, regs(1064) => 
                           bus_reg_dataout_1064_port, regs(1063) => 
                           bus_reg_dataout_1063_port, regs(1062) => 
                           bus_reg_dataout_1062_port, regs(1061) => 
                           bus_reg_dataout_1061_port, regs(1060) => 
                           bus_reg_dataout_1060_port, regs(1059) => 
                           bus_reg_dataout_1059_port, regs(1058) => 
                           bus_reg_dataout_1058_port, regs(1057) => 
                           bus_reg_dataout_1057_port, regs(1056) => 
                           bus_reg_dataout_1056_port, regs(1055) => 
                           bus_reg_dataout_1055_port, regs(1054) => 
                           bus_reg_dataout_1054_port, regs(1053) => 
                           bus_reg_dataout_1053_port, regs(1052) => 
                           bus_reg_dataout_1052_port, regs(1051) => 
                           bus_reg_dataout_1051_port, regs(1050) => 
                           bus_reg_dataout_1050_port, regs(1049) => 
                           bus_reg_dataout_1049_port, regs(1048) => 
                           bus_reg_dataout_1048_port, regs(1047) => 
                           bus_reg_dataout_1047_port, regs(1046) => 
                           bus_reg_dataout_1046_port, regs(1045) => 
                           bus_reg_dataout_1045_port, regs(1044) => 
                           bus_reg_dataout_1044_port, regs(1043) => 
                           bus_reg_dataout_1043_port, regs(1042) => 
                           bus_reg_dataout_1042_port, regs(1041) => 
                           bus_reg_dataout_1041_port, regs(1040) => 
                           bus_reg_dataout_1040_port, regs(1039) => 
                           bus_reg_dataout_1039_port, regs(1038) => 
                           bus_reg_dataout_1038_port, regs(1037) => 
                           bus_reg_dataout_1037_port, regs(1036) => 
                           bus_reg_dataout_1036_port, regs(1035) => 
                           bus_reg_dataout_1035_port, regs(1034) => 
                           bus_reg_dataout_1034_port, regs(1033) => 
                           bus_reg_dataout_1033_port, regs(1032) => 
                           bus_reg_dataout_1032_port, regs(1031) => 
                           bus_reg_dataout_1031_port, regs(1030) => 
                           bus_reg_dataout_1030_port, regs(1029) => 
                           bus_reg_dataout_1029_port, regs(1028) => 
                           bus_reg_dataout_1028_port, regs(1027) => 
                           bus_reg_dataout_1027_port, regs(1026) => 
                           bus_reg_dataout_1026_port, regs(1025) => 
                           bus_reg_dataout_1025_port, regs(1024) => 
                           bus_reg_dataout_1024_port, regs(1023) => 
                           bus_reg_dataout_1023_port, regs(1022) => 
                           bus_reg_dataout_1022_port, regs(1021) => 
                           bus_reg_dataout_1021_port, regs(1020) => 
                           bus_reg_dataout_1020_port, regs(1019) => 
                           bus_reg_dataout_1019_port, regs(1018) => 
                           bus_reg_dataout_1018_port, regs(1017) => 
                           bus_reg_dataout_1017_port, regs(1016) => 
                           bus_reg_dataout_1016_port, regs(1015) => 
                           bus_reg_dataout_1015_port, regs(1014) => 
                           bus_reg_dataout_1014_port, regs(1013) => 
                           bus_reg_dataout_1013_port, regs(1012) => 
                           bus_reg_dataout_1012_port, regs(1011) => 
                           bus_reg_dataout_1011_port, regs(1010) => 
                           bus_reg_dataout_1010_port, regs(1009) => 
                           bus_reg_dataout_1009_port, regs(1008) => 
                           bus_reg_dataout_1008_port, regs(1007) => 
                           bus_reg_dataout_1007_port, regs(1006) => 
                           bus_reg_dataout_1006_port, regs(1005) => 
                           bus_reg_dataout_1005_port, regs(1004) => 
                           bus_reg_dataout_1004_port, regs(1003) => 
                           bus_reg_dataout_1003_port, regs(1002) => 
                           bus_reg_dataout_1002_port, regs(1001) => 
                           bus_reg_dataout_1001_port, regs(1000) => 
                           bus_reg_dataout_1000_port, regs(999) => 
                           bus_reg_dataout_999_port, regs(998) => 
                           bus_reg_dataout_998_port, regs(997) => 
                           bus_reg_dataout_997_port, regs(996) => 
                           bus_reg_dataout_996_port, regs(995) => 
                           bus_reg_dataout_995_port, regs(994) => 
                           bus_reg_dataout_994_port, regs(993) => 
                           bus_reg_dataout_993_port, regs(992) => 
                           bus_reg_dataout_992_port, regs(991) => 
                           bus_reg_dataout_991_port, regs(990) => 
                           bus_reg_dataout_990_port, regs(989) => 
                           bus_reg_dataout_989_port, regs(988) => 
                           bus_reg_dataout_988_port, regs(987) => 
                           bus_reg_dataout_987_port, regs(986) => 
                           bus_reg_dataout_986_port, regs(985) => 
                           bus_reg_dataout_985_port, regs(984) => 
                           bus_reg_dataout_984_port, regs(983) => 
                           bus_reg_dataout_983_port, regs(982) => 
                           bus_reg_dataout_982_port, regs(981) => 
                           bus_reg_dataout_981_port, regs(980) => 
                           bus_reg_dataout_980_port, regs(979) => 
                           bus_reg_dataout_979_port, regs(978) => 
                           bus_reg_dataout_978_port, regs(977) => 
                           bus_reg_dataout_977_port, regs(976) => 
                           bus_reg_dataout_976_port, regs(975) => 
                           bus_reg_dataout_975_port, regs(974) => 
                           bus_reg_dataout_974_port, regs(973) => 
                           bus_reg_dataout_973_port, regs(972) => 
                           bus_reg_dataout_972_port, regs(971) => 
                           bus_reg_dataout_971_port, regs(970) => 
                           bus_reg_dataout_970_port, regs(969) => 
                           bus_reg_dataout_969_port, regs(968) => 
                           bus_reg_dataout_968_port, regs(967) => 
                           bus_reg_dataout_967_port, regs(966) => 
                           bus_reg_dataout_966_port, regs(965) => 
                           bus_reg_dataout_965_port, regs(964) => 
                           bus_reg_dataout_964_port, regs(963) => 
                           bus_reg_dataout_963_port, regs(962) => 
                           bus_reg_dataout_962_port, regs(961) => 
                           bus_reg_dataout_961_port, regs(960) => 
                           bus_reg_dataout_960_port, regs(959) => 
                           bus_reg_dataout_959_port, regs(958) => 
                           bus_reg_dataout_958_port, regs(957) => 
                           bus_reg_dataout_957_port, regs(956) => 
                           bus_reg_dataout_956_port, regs(955) => 
                           bus_reg_dataout_955_port, regs(954) => 
                           bus_reg_dataout_954_port, regs(953) => 
                           bus_reg_dataout_953_port, regs(952) => 
                           bus_reg_dataout_952_port, regs(951) => 
                           bus_reg_dataout_951_port, regs(950) => 
                           bus_reg_dataout_950_port, regs(949) => 
                           bus_reg_dataout_949_port, regs(948) => 
                           bus_reg_dataout_948_port, regs(947) => 
                           bus_reg_dataout_947_port, regs(946) => 
                           bus_reg_dataout_946_port, regs(945) => 
                           bus_reg_dataout_945_port, regs(944) => 
                           bus_reg_dataout_944_port, regs(943) => 
                           bus_reg_dataout_943_port, regs(942) => 
                           bus_reg_dataout_942_port, regs(941) => 
                           bus_reg_dataout_941_port, regs(940) => 
                           bus_reg_dataout_940_port, regs(939) => 
                           bus_reg_dataout_939_port, regs(938) => 
                           bus_reg_dataout_938_port, regs(937) => 
                           bus_reg_dataout_937_port, regs(936) => 
                           bus_reg_dataout_936_port, regs(935) => 
                           bus_reg_dataout_935_port, regs(934) => 
                           bus_reg_dataout_934_port, regs(933) => 
                           bus_reg_dataout_933_port, regs(932) => 
                           bus_reg_dataout_932_port, regs(931) => 
                           bus_reg_dataout_931_port, regs(930) => 
                           bus_reg_dataout_930_port, regs(929) => 
                           bus_reg_dataout_929_port, regs(928) => 
                           bus_reg_dataout_928_port, regs(927) => 
                           bus_reg_dataout_927_port, regs(926) => 
                           bus_reg_dataout_926_port, regs(925) => 
                           bus_reg_dataout_925_port, regs(924) => 
                           bus_reg_dataout_924_port, regs(923) => 
                           bus_reg_dataout_923_port, regs(922) => 
                           bus_reg_dataout_922_port, regs(921) => 
                           bus_reg_dataout_921_port, regs(920) => 
                           bus_reg_dataout_920_port, regs(919) => 
                           bus_reg_dataout_919_port, regs(918) => 
                           bus_reg_dataout_918_port, regs(917) => 
                           bus_reg_dataout_917_port, regs(916) => 
                           bus_reg_dataout_916_port, regs(915) => 
                           bus_reg_dataout_915_port, regs(914) => 
                           bus_reg_dataout_914_port, regs(913) => 
                           bus_reg_dataout_913_port, regs(912) => 
                           bus_reg_dataout_912_port, regs(911) => 
                           bus_reg_dataout_911_port, regs(910) => 
                           bus_reg_dataout_910_port, regs(909) => 
                           bus_reg_dataout_909_port, regs(908) => 
                           bus_reg_dataout_908_port, regs(907) => 
                           bus_reg_dataout_907_port, regs(906) => 
                           bus_reg_dataout_906_port, regs(905) => 
                           bus_reg_dataout_905_port, regs(904) => 
                           bus_reg_dataout_904_port, regs(903) => 
                           bus_reg_dataout_903_port, regs(902) => 
                           bus_reg_dataout_902_port, regs(901) => 
                           bus_reg_dataout_901_port, regs(900) => 
                           bus_reg_dataout_900_port, regs(899) => 
                           bus_reg_dataout_899_port, regs(898) => 
                           bus_reg_dataout_898_port, regs(897) => 
                           bus_reg_dataout_897_port, regs(896) => 
                           bus_reg_dataout_896_port, regs(895) => 
                           bus_reg_dataout_895_port, regs(894) => 
                           bus_reg_dataout_894_port, regs(893) => 
                           bus_reg_dataout_893_port, regs(892) => 
                           bus_reg_dataout_892_port, regs(891) => 
                           bus_reg_dataout_891_port, regs(890) => 
                           bus_reg_dataout_890_port, regs(889) => 
                           bus_reg_dataout_889_port, regs(888) => 
                           bus_reg_dataout_888_port, regs(887) => 
                           bus_reg_dataout_887_port, regs(886) => 
                           bus_reg_dataout_886_port, regs(885) => 
                           bus_reg_dataout_885_port, regs(884) => 
                           bus_reg_dataout_884_port, regs(883) => 
                           bus_reg_dataout_883_port, regs(882) => 
                           bus_reg_dataout_882_port, regs(881) => 
                           bus_reg_dataout_881_port, regs(880) => 
                           bus_reg_dataout_880_port, regs(879) => 
                           bus_reg_dataout_879_port, regs(878) => 
                           bus_reg_dataout_878_port, regs(877) => 
                           bus_reg_dataout_877_port, regs(876) => 
                           bus_reg_dataout_876_port, regs(875) => 
                           bus_reg_dataout_875_port, regs(874) => 
                           bus_reg_dataout_874_port, regs(873) => 
                           bus_reg_dataout_873_port, regs(872) => 
                           bus_reg_dataout_872_port, regs(871) => 
                           bus_reg_dataout_871_port, regs(870) => 
                           bus_reg_dataout_870_port, regs(869) => 
                           bus_reg_dataout_869_port, regs(868) => 
                           bus_reg_dataout_868_port, regs(867) => 
                           bus_reg_dataout_867_port, regs(866) => 
                           bus_reg_dataout_866_port, regs(865) => 
                           bus_reg_dataout_865_port, regs(864) => 
                           bus_reg_dataout_864_port, regs(863) => 
                           bus_reg_dataout_863_port, regs(862) => 
                           bus_reg_dataout_862_port, regs(861) => 
                           bus_reg_dataout_861_port, regs(860) => 
                           bus_reg_dataout_860_port, regs(859) => 
                           bus_reg_dataout_859_port, regs(858) => 
                           bus_reg_dataout_858_port, regs(857) => 
                           bus_reg_dataout_857_port, regs(856) => 
                           bus_reg_dataout_856_port, regs(855) => 
                           bus_reg_dataout_855_port, regs(854) => 
                           bus_reg_dataout_854_port, regs(853) => 
                           bus_reg_dataout_853_port, regs(852) => 
                           bus_reg_dataout_852_port, regs(851) => 
                           bus_reg_dataout_851_port, regs(850) => 
                           bus_reg_dataout_850_port, regs(849) => 
                           bus_reg_dataout_849_port, regs(848) => 
                           bus_reg_dataout_848_port, regs(847) => 
                           bus_reg_dataout_847_port, regs(846) => 
                           bus_reg_dataout_846_port, regs(845) => 
                           bus_reg_dataout_845_port, regs(844) => 
                           bus_reg_dataout_844_port, regs(843) => 
                           bus_reg_dataout_843_port, regs(842) => 
                           bus_reg_dataout_842_port, regs(841) => 
                           bus_reg_dataout_841_port, regs(840) => 
                           bus_reg_dataout_840_port, regs(839) => 
                           bus_reg_dataout_839_port, regs(838) => 
                           bus_reg_dataout_838_port, regs(837) => 
                           bus_reg_dataout_837_port, regs(836) => 
                           bus_reg_dataout_836_port, regs(835) => 
                           bus_reg_dataout_835_port, regs(834) => 
                           bus_reg_dataout_834_port, regs(833) => 
                           bus_reg_dataout_833_port, regs(832) => 
                           bus_reg_dataout_832_port, regs(831) => 
                           bus_reg_dataout_831_port, regs(830) => 
                           bus_reg_dataout_830_port, regs(829) => 
                           bus_reg_dataout_829_port, regs(828) => 
                           bus_reg_dataout_828_port, regs(827) => 
                           bus_reg_dataout_827_port, regs(826) => 
                           bus_reg_dataout_826_port, regs(825) => 
                           bus_reg_dataout_825_port, regs(824) => 
                           bus_reg_dataout_824_port, regs(823) => 
                           bus_reg_dataout_823_port, regs(822) => 
                           bus_reg_dataout_822_port, regs(821) => 
                           bus_reg_dataout_821_port, regs(820) => 
                           bus_reg_dataout_820_port, regs(819) => 
                           bus_reg_dataout_819_port, regs(818) => 
                           bus_reg_dataout_818_port, regs(817) => 
                           bus_reg_dataout_817_port, regs(816) => 
                           bus_reg_dataout_816_port, regs(815) => 
                           bus_reg_dataout_815_port, regs(814) => 
                           bus_reg_dataout_814_port, regs(813) => 
                           bus_reg_dataout_813_port, regs(812) => 
                           bus_reg_dataout_812_port, regs(811) => 
                           bus_reg_dataout_811_port, regs(810) => 
                           bus_reg_dataout_810_port, regs(809) => 
                           bus_reg_dataout_809_port, regs(808) => 
                           bus_reg_dataout_808_port, regs(807) => 
                           bus_reg_dataout_807_port, regs(806) => 
                           bus_reg_dataout_806_port, regs(805) => 
                           bus_reg_dataout_805_port, regs(804) => 
                           bus_reg_dataout_804_port, regs(803) => 
                           bus_reg_dataout_803_port, regs(802) => 
                           bus_reg_dataout_802_port, regs(801) => 
                           bus_reg_dataout_801_port, regs(800) => 
                           bus_reg_dataout_800_port, regs(799) => 
                           bus_reg_dataout_799_port, regs(798) => 
                           bus_reg_dataout_798_port, regs(797) => 
                           bus_reg_dataout_797_port, regs(796) => 
                           bus_reg_dataout_796_port, regs(795) => 
                           bus_reg_dataout_795_port, regs(794) => 
                           bus_reg_dataout_794_port, regs(793) => 
                           bus_reg_dataout_793_port, regs(792) => 
                           bus_reg_dataout_792_port, regs(791) => 
                           bus_reg_dataout_791_port, regs(790) => 
                           bus_reg_dataout_790_port, regs(789) => 
                           bus_reg_dataout_789_port, regs(788) => 
                           bus_reg_dataout_788_port, regs(787) => 
                           bus_reg_dataout_787_port, regs(786) => 
                           bus_reg_dataout_786_port, regs(785) => 
                           bus_reg_dataout_785_port, regs(784) => 
                           bus_reg_dataout_784_port, regs(783) => 
                           bus_reg_dataout_783_port, regs(782) => 
                           bus_reg_dataout_782_port, regs(781) => 
                           bus_reg_dataout_781_port, regs(780) => 
                           bus_reg_dataout_780_port, regs(779) => 
                           bus_reg_dataout_779_port, regs(778) => 
                           bus_reg_dataout_778_port, regs(777) => 
                           bus_reg_dataout_777_port, regs(776) => 
                           bus_reg_dataout_776_port, regs(775) => 
                           bus_reg_dataout_775_port, regs(774) => 
                           bus_reg_dataout_774_port, regs(773) => 
                           bus_reg_dataout_773_port, regs(772) => 
                           bus_reg_dataout_772_port, regs(771) => 
                           bus_reg_dataout_771_port, regs(770) => 
                           bus_reg_dataout_770_port, regs(769) => 
                           bus_reg_dataout_769_port, regs(768) => 
                           bus_reg_dataout_768_port, regs(767) => 
                           bus_reg_dataout_767_port, regs(766) => 
                           bus_reg_dataout_766_port, regs(765) => 
                           bus_reg_dataout_765_port, regs(764) => 
                           bus_reg_dataout_764_port, regs(763) => 
                           bus_reg_dataout_763_port, regs(762) => 
                           bus_reg_dataout_762_port, regs(761) => 
                           bus_reg_dataout_761_port, regs(760) => 
                           bus_reg_dataout_760_port, regs(759) => 
                           bus_reg_dataout_759_port, regs(758) => 
                           bus_reg_dataout_758_port, regs(757) => 
                           bus_reg_dataout_757_port, regs(756) => 
                           bus_reg_dataout_756_port, regs(755) => 
                           bus_reg_dataout_755_port, regs(754) => 
                           bus_reg_dataout_754_port, regs(753) => 
                           bus_reg_dataout_753_port, regs(752) => 
                           bus_reg_dataout_752_port, regs(751) => 
                           bus_reg_dataout_751_port, regs(750) => 
                           bus_reg_dataout_750_port, regs(749) => 
                           bus_reg_dataout_749_port, regs(748) => 
                           bus_reg_dataout_748_port, regs(747) => 
                           bus_reg_dataout_747_port, regs(746) => 
                           bus_reg_dataout_746_port, regs(745) => 
                           bus_reg_dataout_745_port, regs(744) => 
                           bus_reg_dataout_744_port, regs(743) => 
                           bus_reg_dataout_743_port, regs(742) => 
                           bus_reg_dataout_742_port, regs(741) => 
                           bus_reg_dataout_741_port, regs(740) => 
                           bus_reg_dataout_740_port, regs(739) => 
                           bus_reg_dataout_739_port, regs(738) => 
                           bus_reg_dataout_738_port, regs(737) => 
                           bus_reg_dataout_737_port, regs(736) => 
                           bus_reg_dataout_736_port, regs(735) => 
                           bus_reg_dataout_735_port, regs(734) => 
                           bus_reg_dataout_734_port, regs(733) => 
                           bus_reg_dataout_733_port, regs(732) => 
                           bus_reg_dataout_732_port, regs(731) => 
                           bus_reg_dataout_731_port, regs(730) => 
                           bus_reg_dataout_730_port, regs(729) => 
                           bus_reg_dataout_729_port, regs(728) => 
                           bus_reg_dataout_728_port, regs(727) => 
                           bus_reg_dataout_727_port, regs(726) => 
                           bus_reg_dataout_726_port, regs(725) => 
                           bus_reg_dataout_725_port, regs(724) => 
                           bus_reg_dataout_724_port, regs(723) => 
                           bus_reg_dataout_723_port, regs(722) => 
                           bus_reg_dataout_722_port, regs(721) => 
                           bus_reg_dataout_721_port, regs(720) => 
                           bus_reg_dataout_720_port, regs(719) => 
                           bus_reg_dataout_719_port, regs(718) => 
                           bus_reg_dataout_718_port, regs(717) => 
                           bus_reg_dataout_717_port, regs(716) => 
                           bus_reg_dataout_716_port, regs(715) => 
                           bus_reg_dataout_715_port, regs(714) => 
                           bus_reg_dataout_714_port, regs(713) => 
                           bus_reg_dataout_713_port, regs(712) => 
                           bus_reg_dataout_712_port, regs(711) => 
                           bus_reg_dataout_711_port, regs(710) => 
                           bus_reg_dataout_710_port, regs(709) => 
                           bus_reg_dataout_709_port, regs(708) => 
                           bus_reg_dataout_708_port, regs(707) => 
                           bus_reg_dataout_707_port, regs(706) => 
                           bus_reg_dataout_706_port, regs(705) => 
                           bus_reg_dataout_705_port, regs(704) => 
                           bus_reg_dataout_704_port, regs(703) => 
                           bus_reg_dataout_703_port, regs(702) => 
                           bus_reg_dataout_702_port, regs(701) => 
                           bus_reg_dataout_701_port, regs(700) => 
                           bus_reg_dataout_700_port, regs(699) => 
                           bus_reg_dataout_699_port, regs(698) => 
                           bus_reg_dataout_698_port, regs(697) => 
                           bus_reg_dataout_697_port, regs(696) => 
                           bus_reg_dataout_696_port, regs(695) => 
                           bus_reg_dataout_695_port, regs(694) => 
                           bus_reg_dataout_694_port, regs(693) => 
                           bus_reg_dataout_693_port, regs(692) => 
                           bus_reg_dataout_692_port, regs(691) => 
                           bus_reg_dataout_691_port, regs(690) => 
                           bus_reg_dataout_690_port, regs(689) => 
                           bus_reg_dataout_689_port, regs(688) => 
                           bus_reg_dataout_688_port, regs(687) => 
                           bus_reg_dataout_687_port, regs(686) => 
                           bus_reg_dataout_686_port, regs(685) => 
                           bus_reg_dataout_685_port, regs(684) => 
                           bus_reg_dataout_684_port, regs(683) => 
                           bus_reg_dataout_683_port, regs(682) => 
                           bus_reg_dataout_682_port, regs(681) => 
                           bus_reg_dataout_681_port, regs(680) => 
                           bus_reg_dataout_680_port, regs(679) => 
                           bus_reg_dataout_679_port, regs(678) => 
                           bus_reg_dataout_678_port, regs(677) => 
                           bus_reg_dataout_677_port, regs(676) => 
                           bus_reg_dataout_676_port, regs(675) => 
                           bus_reg_dataout_675_port, regs(674) => 
                           bus_reg_dataout_674_port, regs(673) => 
                           bus_reg_dataout_673_port, regs(672) => 
                           bus_reg_dataout_672_port, regs(671) => 
                           bus_reg_dataout_671_port, regs(670) => 
                           bus_reg_dataout_670_port, regs(669) => 
                           bus_reg_dataout_669_port, regs(668) => 
                           bus_reg_dataout_668_port, regs(667) => 
                           bus_reg_dataout_667_port, regs(666) => 
                           bus_reg_dataout_666_port, regs(665) => 
                           bus_reg_dataout_665_port, regs(664) => 
                           bus_reg_dataout_664_port, regs(663) => 
                           bus_reg_dataout_663_port, regs(662) => 
                           bus_reg_dataout_662_port, regs(661) => 
                           bus_reg_dataout_661_port, regs(660) => 
                           bus_reg_dataout_660_port, regs(659) => 
                           bus_reg_dataout_659_port, regs(658) => 
                           bus_reg_dataout_658_port, regs(657) => 
                           bus_reg_dataout_657_port, regs(656) => 
                           bus_reg_dataout_656_port, regs(655) => 
                           bus_reg_dataout_655_port, regs(654) => 
                           bus_reg_dataout_654_port, regs(653) => 
                           bus_reg_dataout_653_port, regs(652) => 
                           bus_reg_dataout_652_port, regs(651) => 
                           bus_reg_dataout_651_port, regs(650) => 
                           bus_reg_dataout_650_port, regs(649) => 
                           bus_reg_dataout_649_port, regs(648) => 
                           bus_reg_dataout_648_port, regs(647) => 
                           bus_reg_dataout_647_port, regs(646) => 
                           bus_reg_dataout_646_port, regs(645) => 
                           bus_reg_dataout_645_port, regs(644) => 
                           bus_reg_dataout_644_port, regs(643) => 
                           bus_reg_dataout_643_port, regs(642) => 
                           bus_reg_dataout_642_port, regs(641) => 
                           bus_reg_dataout_641_port, regs(640) => 
                           bus_reg_dataout_640_port, regs(639) => 
                           bus_reg_dataout_639_port, regs(638) => 
                           bus_reg_dataout_638_port, regs(637) => 
                           bus_reg_dataout_637_port, regs(636) => 
                           bus_reg_dataout_636_port, regs(635) => 
                           bus_reg_dataout_635_port, regs(634) => 
                           bus_reg_dataout_634_port, regs(633) => 
                           bus_reg_dataout_633_port, regs(632) => 
                           bus_reg_dataout_632_port, regs(631) => 
                           bus_reg_dataout_631_port, regs(630) => 
                           bus_reg_dataout_630_port, regs(629) => 
                           bus_reg_dataout_629_port, regs(628) => 
                           bus_reg_dataout_628_port, regs(627) => 
                           bus_reg_dataout_627_port, regs(626) => 
                           bus_reg_dataout_626_port, regs(625) => 
                           bus_reg_dataout_625_port, regs(624) => 
                           bus_reg_dataout_624_port, regs(623) => 
                           bus_reg_dataout_623_port, regs(622) => 
                           bus_reg_dataout_622_port, regs(621) => 
                           bus_reg_dataout_621_port, regs(620) => 
                           bus_reg_dataout_620_port, regs(619) => 
                           bus_reg_dataout_619_port, regs(618) => 
                           bus_reg_dataout_618_port, regs(617) => 
                           bus_reg_dataout_617_port, regs(616) => 
                           bus_reg_dataout_616_port, regs(615) => 
                           bus_reg_dataout_615_port, regs(614) => 
                           bus_reg_dataout_614_port, regs(613) => 
                           bus_reg_dataout_613_port, regs(612) => 
                           bus_reg_dataout_612_port, regs(611) => 
                           bus_reg_dataout_611_port, regs(610) => 
                           bus_reg_dataout_610_port, regs(609) => 
                           bus_reg_dataout_609_port, regs(608) => 
                           bus_reg_dataout_608_port, regs(607) => 
                           bus_reg_dataout_607_port, regs(606) => 
                           bus_reg_dataout_606_port, regs(605) => 
                           bus_reg_dataout_605_port, regs(604) => 
                           bus_reg_dataout_604_port, regs(603) => 
                           bus_reg_dataout_603_port, regs(602) => 
                           bus_reg_dataout_602_port, regs(601) => 
                           bus_reg_dataout_601_port, regs(600) => 
                           bus_reg_dataout_600_port, regs(599) => 
                           bus_reg_dataout_599_port, regs(598) => 
                           bus_reg_dataout_598_port, regs(597) => 
                           bus_reg_dataout_597_port, regs(596) => 
                           bus_reg_dataout_596_port, regs(595) => 
                           bus_reg_dataout_595_port, regs(594) => 
                           bus_reg_dataout_594_port, regs(593) => 
                           bus_reg_dataout_593_port, regs(592) => 
                           bus_reg_dataout_592_port, regs(591) => 
                           bus_reg_dataout_591_port, regs(590) => 
                           bus_reg_dataout_590_port, regs(589) => 
                           bus_reg_dataout_589_port, regs(588) => 
                           bus_reg_dataout_588_port, regs(587) => 
                           bus_reg_dataout_587_port, regs(586) => 
                           bus_reg_dataout_586_port, regs(585) => 
                           bus_reg_dataout_585_port, regs(584) => 
                           bus_reg_dataout_584_port, regs(583) => 
                           bus_reg_dataout_583_port, regs(582) => 
                           bus_reg_dataout_582_port, regs(581) => 
                           bus_reg_dataout_581_port, regs(580) => 
                           bus_reg_dataout_580_port, regs(579) => 
                           bus_reg_dataout_579_port, regs(578) => 
                           bus_reg_dataout_578_port, regs(577) => 
                           bus_reg_dataout_577_port, regs(576) => 
                           bus_reg_dataout_576_port, regs(575) => 
                           bus_reg_dataout_575_port, regs(574) => 
                           bus_reg_dataout_574_port, regs(573) => 
                           bus_reg_dataout_573_port, regs(572) => 
                           bus_reg_dataout_572_port, regs(571) => 
                           bus_reg_dataout_571_port, regs(570) => 
                           bus_reg_dataout_570_port, regs(569) => 
                           bus_reg_dataout_569_port, regs(568) => 
                           bus_reg_dataout_568_port, regs(567) => 
                           bus_reg_dataout_567_port, regs(566) => 
                           bus_reg_dataout_566_port, regs(565) => 
                           bus_reg_dataout_565_port, regs(564) => 
                           bus_reg_dataout_564_port, regs(563) => 
                           bus_reg_dataout_563_port, regs(562) => 
                           bus_reg_dataout_562_port, regs(561) => 
                           bus_reg_dataout_561_port, regs(560) => 
                           bus_reg_dataout_560_port, regs(559) => 
                           bus_reg_dataout_559_port, regs(558) => 
                           bus_reg_dataout_558_port, regs(557) => 
                           bus_reg_dataout_557_port, regs(556) => 
                           bus_reg_dataout_556_port, regs(555) => 
                           bus_reg_dataout_555_port, regs(554) => 
                           bus_reg_dataout_554_port, regs(553) => 
                           bus_reg_dataout_553_port, regs(552) => 
                           bus_reg_dataout_552_port, regs(551) => 
                           bus_reg_dataout_551_port, regs(550) => 
                           bus_reg_dataout_550_port, regs(549) => 
                           bus_reg_dataout_549_port, regs(548) => 
                           bus_reg_dataout_548_port, regs(547) => 
                           bus_reg_dataout_547_port, regs(546) => 
                           bus_reg_dataout_546_port, regs(545) => 
                           bus_reg_dataout_545_port, regs(544) => 
                           bus_reg_dataout_544_port, regs(543) => 
                           bus_reg_dataout_543_port, regs(542) => 
                           bus_reg_dataout_542_port, regs(541) => 
                           bus_reg_dataout_541_port, regs(540) => 
                           bus_reg_dataout_540_port, regs(539) => 
                           bus_reg_dataout_539_port, regs(538) => 
                           bus_reg_dataout_538_port, regs(537) => 
                           bus_reg_dataout_537_port, regs(536) => 
                           bus_reg_dataout_536_port, regs(535) => 
                           bus_reg_dataout_535_port, regs(534) => 
                           bus_reg_dataout_534_port, regs(533) => 
                           bus_reg_dataout_533_port, regs(532) => 
                           bus_reg_dataout_532_port, regs(531) => 
                           bus_reg_dataout_531_port, regs(530) => 
                           bus_reg_dataout_530_port, regs(529) => 
                           bus_reg_dataout_529_port, regs(528) => 
                           bus_reg_dataout_528_port, regs(527) => 
                           bus_reg_dataout_527_port, regs(526) => 
                           bus_reg_dataout_526_port, regs(525) => 
                           bus_reg_dataout_525_port, regs(524) => 
                           bus_reg_dataout_524_port, regs(523) => 
                           bus_reg_dataout_523_port, regs(522) => 
                           bus_reg_dataout_522_port, regs(521) => 
                           bus_reg_dataout_521_port, regs(520) => 
                           bus_reg_dataout_520_port, regs(519) => 
                           bus_reg_dataout_519_port, regs(518) => 
                           bus_reg_dataout_518_port, regs(517) => 
                           bus_reg_dataout_517_port, regs(516) => 
                           bus_reg_dataout_516_port, regs(515) => 
                           bus_reg_dataout_515_port, regs(514) => 
                           bus_reg_dataout_514_port, regs(513) => 
                           bus_reg_dataout_513_port, regs(512) => 
                           bus_reg_dataout_512_port, regs(511) => 
                           bus_reg_dataout_511_port, regs(510) => 
                           bus_reg_dataout_510_port, regs(509) => 
                           bus_reg_dataout_509_port, regs(508) => 
                           bus_reg_dataout_508_port, regs(507) => 
                           bus_reg_dataout_507_port, regs(506) => 
                           bus_reg_dataout_506_port, regs(505) => 
                           bus_reg_dataout_505_port, regs(504) => 
                           bus_reg_dataout_504_port, regs(503) => 
                           bus_reg_dataout_503_port, regs(502) => 
                           bus_reg_dataout_502_port, regs(501) => 
                           bus_reg_dataout_501_port, regs(500) => 
                           bus_reg_dataout_500_port, regs(499) => 
                           bus_reg_dataout_499_port, regs(498) => 
                           bus_reg_dataout_498_port, regs(497) => 
                           bus_reg_dataout_497_port, regs(496) => 
                           bus_reg_dataout_496_port, regs(495) => 
                           bus_reg_dataout_495_port, regs(494) => 
                           bus_reg_dataout_494_port, regs(493) => 
                           bus_reg_dataout_493_port, regs(492) => 
                           bus_reg_dataout_492_port, regs(491) => 
                           bus_reg_dataout_491_port, regs(490) => 
                           bus_reg_dataout_490_port, regs(489) => 
                           bus_reg_dataout_489_port, regs(488) => 
                           bus_reg_dataout_488_port, regs(487) => 
                           bus_reg_dataout_487_port, regs(486) => 
                           bus_reg_dataout_486_port, regs(485) => 
                           bus_reg_dataout_485_port, regs(484) => 
                           bus_reg_dataout_484_port, regs(483) => 
                           bus_reg_dataout_483_port, regs(482) => 
                           bus_reg_dataout_482_port, regs(481) => 
                           bus_reg_dataout_481_port, regs(480) => 
                           bus_reg_dataout_480_port, regs(479) => 
                           bus_reg_dataout_479_port, regs(478) => 
                           bus_reg_dataout_478_port, regs(477) => 
                           bus_reg_dataout_477_port, regs(476) => 
                           bus_reg_dataout_476_port, regs(475) => 
                           bus_reg_dataout_475_port, regs(474) => 
                           bus_reg_dataout_474_port, regs(473) => 
                           bus_reg_dataout_473_port, regs(472) => 
                           bus_reg_dataout_472_port, regs(471) => 
                           bus_reg_dataout_471_port, regs(470) => 
                           bus_reg_dataout_470_port, regs(469) => 
                           bus_reg_dataout_469_port, regs(468) => 
                           bus_reg_dataout_468_port, regs(467) => 
                           bus_reg_dataout_467_port, regs(466) => 
                           bus_reg_dataout_466_port, regs(465) => 
                           bus_reg_dataout_465_port, regs(464) => 
                           bus_reg_dataout_464_port, regs(463) => 
                           bus_reg_dataout_463_port, regs(462) => 
                           bus_reg_dataout_462_port, regs(461) => 
                           bus_reg_dataout_461_port, regs(460) => 
                           bus_reg_dataout_460_port, regs(459) => 
                           bus_reg_dataout_459_port, regs(458) => 
                           bus_reg_dataout_458_port, regs(457) => 
                           bus_reg_dataout_457_port, regs(456) => 
                           bus_reg_dataout_456_port, regs(455) => 
                           bus_reg_dataout_455_port, regs(454) => 
                           bus_reg_dataout_454_port, regs(453) => 
                           bus_reg_dataout_453_port, regs(452) => 
                           bus_reg_dataout_452_port, regs(451) => 
                           bus_reg_dataout_451_port, regs(450) => 
                           bus_reg_dataout_450_port, regs(449) => 
                           bus_reg_dataout_449_port, regs(448) => 
                           bus_reg_dataout_448_port, regs(447) => 
                           bus_reg_dataout_447_port, regs(446) => 
                           bus_reg_dataout_446_port, regs(445) => 
                           bus_reg_dataout_445_port, regs(444) => 
                           bus_reg_dataout_444_port, regs(443) => 
                           bus_reg_dataout_443_port, regs(442) => 
                           bus_reg_dataout_442_port, regs(441) => 
                           bus_reg_dataout_441_port, regs(440) => 
                           bus_reg_dataout_440_port, regs(439) => 
                           bus_reg_dataout_439_port, regs(438) => 
                           bus_reg_dataout_438_port, regs(437) => 
                           bus_reg_dataout_437_port, regs(436) => 
                           bus_reg_dataout_436_port, regs(435) => 
                           bus_reg_dataout_435_port, regs(434) => 
                           bus_reg_dataout_434_port, regs(433) => 
                           bus_reg_dataout_433_port, regs(432) => 
                           bus_reg_dataout_432_port, regs(431) => 
                           bus_reg_dataout_431_port, regs(430) => 
                           bus_reg_dataout_430_port, regs(429) => 
                           bus_reg_dataout_429_port, regs(428) => 
                           bus_reg_dataout_428_port, regs(427) => 
                           bus_reg_dataout_427_port, regs(426) => 
                           bus_reg_dataout_426_port, regs(425) => 
                           bus_reg_dataout_425_port, regs(424) => 
                           bus_reg_dataout_424_port, regs(423) => 
                           bus_reg_dataout_423_port, regs(422) => 
                           bus_reg_dataout_422_port, regs(421) => 
                           bus_reg_dataout_421_port, regs(420) => 
                           bus_reg_dataout_420_port, regs(419) => 
                           bus_reg_dataout_419_port, regs(418) => 
                           bus_reg_dataout_418_port, regs(417) => 
                           bus_reg_dataout_417_port, regs(416) => 
                           bus_reg_dataout_416_port, regs(415) => 
                           bus_reg_dataout_415_port, regs(414) => 
                           bus_reg_dataout_414_port, regs(413) => 
                           bus_reg_dataout_413_port, regs(412) => 
                           bus_reg_dataout_412_port, regs(411) => 
                           bus_reg_dataout_411_port, regs(410) => 
                           bus_reg_dataout_410_port, regs(409) => 
                           bus_reg_dataout_409_port, regs(408) => 
                           bus_reg_dataout_408_port, regs(407) => 
                           bus_reg_dataout_407_port, regs(406) => 
                           bus_reg_dataout_406_port, regs(405) => 
                           bus_reg_dataout_405_port, regs(404) => 
                           bus_reg_dataout_404_port, regs(403) => 
                           bus_reg_dataout_403_port, regs(402) => 
                           bus_reg_dataout_402_port, regs(401) => 
                           bus_reg_dataout_401_port, regs(400) => 
                           bus_reg_dataout_400_port, regs(399) => 
                           bus_reg_dataout_399_port, regs(398) => 
                           bus_reg_dataout_398_port, regs(397) => 
                           bus_reg_dataout_397_port, regs(396) => 
                           bus_reg_dataout_396_port, regs(395) => 
                           bus_reg_dataout_395_port, regs(394) => 
                           bus_reg_dataout_394_port, regs(393) => 
                           bus_reg_dataout_393_port, regs(392) => 
                           bus_reg_dataout_392_port, regs(391) => 
                           bus_reg_dataout_391_port, regs(390) => 
                           bus_reg_dataout_390_port, regs(389) => 
                           bus_reg_dataout_389_port, regs(388) => 
                           bus_reg_dataout_388_port, regs(387) => 
                           bus_reg_dataout_387_port, regs(386) => 
                           bus_reg_dataout_386_port, regs(385) => 
                           bus_reg_dataout_385_port, regs(384) => 
                           bus_reg_dataout_384_port, regs(383) => 
                           bus_reg_dataout_383_port, regs(382) => 
                           bus_reg_dataout_382_port, regs(381) => 
                           bus_reg_dataout_381_port, regs(380) => 
                           bus_reg_dataout_380_port, regs(379) => 
                           bus_reg_dataout_379_port, regs(378) => 
                           bus_reg_dataout_378_port, regs(377) => 
                           bus_reg_dataout_377_port, regs(376) => 
                           bus_reg_dataout_376_port, regs(375) => 
                           bus_reg_dataout_375_port, regs(374) => 
                           bus_reg_dataout_374_port, regs(373) => 
                           bus_reg_dataout_373_port, regs(372) => 
                           bus_reg_dataout_372_port, regs(371) => 
                           bus_reg_dataout_371_port, regs(370) => 
                           bus_reg_dataout_370_port, regs(369) => 
                           bus_reg_dataout_369_port, regs(368) => 
                           bus_reg_dataout_368_port, regs(367) => 
                           bus_reg_dataout_367_port, regs(366) => 
                           bus_reg_dataout_366_port, regs(365) => 
                           bus_reg_dataout_365_port, regs(364) => 
                           bus_reg_dataout_364_port, regs(363) => 
                           bus_reg_dataout_363_port, regs(362) => 
                           bus_reg_dataout_362_port, regs(361) => 
                           bus_reg_dataout_361_port, regs(360) => 
                           bus_reg_dataout_360_port, regs(359) => 
                           bus_reg_dataout_359_port, regs(358) => 
                           bus_reg_dataout_358_port, regs(357) => 
                           bus_reg_dataout_357_port, regs(356) => 
                           bus_reg_dataout_356_port, regs(355) => 
                           bus_reg_dataout_355_port, regs(354) => 
                           bus_reg_dataout_354_port, regs(353) => 
                           bus_reg_dataout_353_port, regs(352) => 
                           bus_reg_dataout_352_port, regs(351) => 
                           bus_reg_dataout_351_port, regs(350) => 
                           bus_reg_dataout_350_port, regs(349) => 
                           bus_reg_dataout_349_port, regs(348) => 
                           bus_reg_dataout_348_port, regs(347) => 
                           bus_reg_dataout_347_port, regs(346) => 
                           bus_reg_dataout_346_port, regs(345) => 
                           bus_reg_dataout_345_port, regs(344) => 
                           bus_reg_dataout_344_port, regs(343) => 
                           bus_reg_dataout_343_port, regs(342) => 
                           bus_reg_dataout_342_port, regs(341) => 
                           bus_reg_dataout_341_port, regs(340) => 
                           bus_reg_dataout_340_port, regs(339) => 
                           bus_reg_dataout_339_port, regs(338) => 
                           bus_reg_dataout_338_port, regs(337) => 
                           bus_reg_dataout_337_port, regs(336) => 
                           bus_reg_dataout_336_port, regs(335) => 
                           bus_reg_dataout_335_port, regs(334) => 
                           bus_reg_dataout_334_port, regs(333) => 
                           bus_reg_dataout_333_port, regs(332) => 
                           bus_reg_dataout_332_port, regs(331) => 
                           bus_reg_dataout_331_port, regs(330) => 
                           bus_reg_dataout_330_port, regs(329) => 
                           bus_reg_dataout_329_port, regs(328) => 
                           bus_reg_dataout_328_port, regs(327) => 
                           bus_reg_dataout_327_port, regs(326) => 
                           bus_reg_dataout_326_port, regs(325) => 
                           bus_reg_dataout_325_port, regs(324) => 
                           bus_reg_dataout_324_port, regs(323) => 
                           bus_reg_dataout_323_port, regs(322) => 
                           bus_reg_dataout_322_port, regs(321) => 
                           bus_reg_dataout_321_port, regs(320) => 
                           bus_reg_dataout_320_port, regs(319) => 
                           bus_reg_dataout_319_port, regs(318) => 
                           bus_reg_dataout_318_port, regs(317) => 
                           bus_reg_dataout_317_port, regs(316) => 
                           bus_reg_dataout_316_port, regs(315) => 
                           bus_reg_dataout_315_port, regs(314) => 
                           bus_reg_dataout_314_port, regs(313) => 
                           bus_reg_dataout_313_port, regs(312) => 
                           bus_reg_dataout_312_port, regs(311) => 
                           bus_reg_dataout_311_port, regs(310) => 
                           bus_reg_dataout_310_port, regs(309) => 
                           bus_reg_dataout_309_port, regs(308) => 
                           bus_reg_dataout_308_port, regs(307) => 
                           bus_reg_dataout_307_port, regs(306) => 
                           bus_reg_dataout_306_port, regs(305) => 
                           bus_reg_dataout_305_port, regs(304) => 
                           bus_reg_dataout_304_port, regs(303) => 
                           bus_reg_dataout_303_port, regs(302) => 
                           bus_reg_dataout_302_port, regs(301) => 
                           bus_reg_dataout_301_port, regs(300) => 
                           bus_reg_dataout_300_port, regs(299) => 
                           bus_reg_dataout_299_port, regs(298) => 
                           bus_reg_dataout_298_port, regs(297) => 
                           bus_reg_dataout_297_port, regs(296) => 
                           bus_reg_dataout_296_port, regs(295) => 
                           bus_reg_dataout_295_port, regs(294) => 
                           bus_reg_dataout_294_port, regs(293) => 
                           bus_reg_dataout_293_port, regs(292) => 
                           bus_reg_dataout_292_port, regs(291) => 
                           bus_reg_dataout_291_port, regs(290) => 
                           bus_reg_dataout_290_port, regs(289) => 
                           bus_reg_dataout_289_port, regs(288) => 
                           bus_reg_dataout_288_port, regs(287) => 
                           bus_reg_dataout_287_port, regs(286) => 
                           bus_reg_dataout_286_port, regs(285) => 
                           bus_reg_dataout_285_port, regs(284) => 
                           bus_reg_dataout_284_port, regs(283) => 
                           bus_reg_dataout_283_port, regs(282) => 
                           bus_reg_dataout_282_port, regs(281) => 
                           bus_reg_dataout_281_port, regs(280) => 
                           bus_reg_dataout_280_port, regs(279) => 
                           bus_reg_dataout_279_port, regs(278) => 
                           bus_reg_dataout_278_port, regs(277) => 
                           bus_reg_dataout_277_port, regs(276) => 
                           bus_reg_dataout_276_port, regs(275) => 
                           bus_reg_dataout_275_port, regs(274) => 
                           bus_reg_dataout_274_port, regs(273) => 
                           bus_reg_dataout_273_port, regs(272) => 
                           bus_reg_dataout_272_port, regs(271) => 
                           bus_reg_dataout_271_port, regs(270) => 
                           bus_reg_dataout_270_port, regs(269) => 
                           bus_reg_dataout_269_port, regs(268) => 
                           bus_reg_dataout_268_port, regs(267) => 
                           bus_reg_dataout_267_port, regs(266) => 
                           bus_reg_dataout_266_port, regs(265) => 
                           bus_reg_dataout_265_port, regs(264) => 
                           bus_reg_dataout_264_port, regs(263) => 
                           bus_reg_dataout_263_port, regs(262) => 
                           bus_reg_dataout_262_port, regs(261) => 
                           bus_reg_dataout_261_port, regs(260) => 
                           bus_reg_dataout_260_port, regs(259) => 
                           bus_reg_dataout_259_port, regs(258) => 
                           bus_reg_dataout_258_port, regs(257) => 
                           bus_reg_dataout_257_port, regs(256) => 
                           bus_reg_dataout_256_port, regs(255) => 
                           bus_reg_dataout_255_port, regs(254) => 
                           bus_reg_dataout_254_port, regs(253) => 
                           bus_reg_dataout_253_port, regs(252) => 
                           bus_reg_dataout_252_port, regs(251) => 
                           bus_reg_dataout_251_port, regs(250) => 
                           bus_reg_dataout_250_port, regs(249) => 
                           bus_reg_dataout_249_port, regs(248) => 
                           bus_reg_dataout_248_port, regs(247) => 
                           bus_reg_dataout_247_port, regs(246) => 
                           bus_reg_dataout_246_port, regs(245) => 
                           bus_reg_dataout_245_port, regs(244) => 
                           bus_reg_dataout_244_port, regs(243) => 
                           bus_reg_dataout_243_port, regs(242) => 
                           bus_reg_dataout_242_port, regs(241) => 
                           bus_reg_dataout_241_port, regs(240) => 
                           bus_reg_dataout_240_port, regs(239) => 
                           bus_reg_dataout_239_port, regs(238) => 
                           bus_reg_dataout_238_port, regs(237) => 
                           bus_reg_dataout_237_port, regs(236) => 
                           bus_reg_dataout_236_port, regs(235) => 
                           bus_reg_dataout_235_port, regs(234) => 
                           bus_reg_dataout_234_port, regs(233) => 
                           bus_reg_dataout_233_port, regs(232) => 
                           bus_reg_dataout_232_port, regs(231) => 
                           bus_reg_dataout_231_port, regs(230) => 
                           bus_reg_dataout_230_port, regs(229) => 
                           bus_reg_dataout_229_port, regs(228) => 
                           bus_reg_dataout_228_port, regs(227) => 
                           bus_reg_dataout_227_port, regs(226) => 
                           bus_reg_dataout_226_port, regs(225) => 
                           bus_reg_dataout_225_port, regs(224) => 
                           bus_reg_dataout_224_port, regs(223) => 
                           bus_reg_dataout_223_port, regs(222) => 
                           bus_reg_dataout_222_port, regs(221) => 
                           bus_reg_dataout_221_port, regs(220) => 
                           bus_reg_dataout_220_port, regs(219) => 
                           bus_reg_dataout_219_port, regs(218) => 
                           bus_reg_dataout_218_port, regs(217) => 
                           bus_reg_dataout_217_port, regs(216) => 
                           bus_reg_dataout_216_port, regs(215) => 
                           bus_reg_dataout_215_port, regs(214) => 
                           bus_reg_dataout_214_port, regs(213) => 
                           bus_reg_dataout_213_port, regs(212) => 
                           bus_reg_dataout_212_port, regs(211) => 
                           bus_reg_dataout_211_port, regs(210) => 
                           bus_reg_dataout_210_port, regs(209) => 
                           bus_reg_dataout_209_port, regs(208) => 
                           bus_reg_dataout_208_port, regs(207) => 
                           bus_reg_dataout_207_port, regs(206) => 
                           bus_reg_dataout_206_port, regs(205) => 
                           bus_reg_dataout_205_port, regs(204) => 
                           bus_reg_dataout_204_port, regs(203) => 
                           bus_reg_dataout_203_port, regs(202) => 
                           bus_reg_dataout_202_port, regs(201) => 
                           bus_reg_dataout_201_port, regs(200) => 
                           bus_reg_dataout_200_port, regs(199) => 
                           bus_reg_dataout_199_port, regs(198) => 
                           bus_reg_dataout_198_port, regs(197) => 
                           bus_reg_dataout_197_port, regs(196) => 
                           bus_reg_dataout_196_port, regs(195) => 
                           bus_reg_dataout_195_port, regs(194) => 
                           bus_reg_dataout_194_port, regs(193) => 
                           bus_reg_dataout_193_port, regs(192) => 
                           bus_reg_dataout_192_port, regs(191) => 
                           bus_reg_dataout_191_port, regs(190) => 
                           bus_reg_dataout_190_port, regs(189) => 
                           bus_reg_dataout_189_port, regs(188) => 
                           bus_reg_dataout_188_port, regs(187) => 
                           bus_reg_dataout_187_port, regs(186) => 
                           bus_reg_dataout_186_port, regs(185) => 
                           bus_reg_dataout_185_port, regs(184) => 
                           bus_reg_dataout_184_port, regs(183) => 
                           bus_reg_dataout_183_port, regs(182) => 
                           bus_reg_dataout_182_port, regs(181) => 
                           bus_reg_dataout_181_port, regs(180) => 
                           bus_reg_dataout_180_port, regs(179) => 
                           bus_reg_dataout_179_port, regs(178) => 
                           bus_reg_dataout_178_port, regs(177) => 
                           bus_reg_dataout_177_port, regs(176) => 
                           bus_reg_dataout_176_port, regs(175) => 
                           bus_reg_dataout_175_port, regs(174) => 
                           bus_reg_dataout_174_port, regs(173) => 
                           bus_reg_dataout_173_port, regs(172) => 
                           bus_reg_dataout_172_port, regs(171) => 
                           bus_reg_dataout_171_port, regs(170) => 
                           bus_reg_dataout_170_port, regs(169) => 
                           bus_reg_dataout_169_port, regs(168) => 
                           bus_reg_dataout_168_port, regs(167) => 
                           bus_reg_dataout_167_port, regs(166) => 
                           bus_reg_dataout_166_port, regs(165) => 
                           bus_reg_dataout_165_port, regs(164) => 
                           bus_reg_dataout_164_port, regs(163) => 
                           bus_reg_dataout_163_port, regs(162) => 
                           bus_reg_dataout_162_port, regs(161) => 
                           bus_reg_dataout_161_port, regs(160) => 
                           bus_reg_dataout_160_port, regs(159) => 
                           bus_reg_dataout_159_port, regs(158) => 
                           bus_reg_dataout_158_port, regs(157) => 
                           bus_reg_dataout_157_port, regs(156) => 
                           bus_reg_dataout_156_port, regs(155) => 
                           bus_reg_dataout_155_port, regs(154) => 
                           bus_reg_dataout_154_port, regs(153) => 
                           bus_reg_dataout_153_port, regs(152) => 
                           bus_reg_dataout_152_port, regs(151) => 
                           bus_reg_dataout_151_port, regs(150) => 
                           bus_reg_dataout_150_port, regs(149) => 
                           bus_reg_dataout_149_port, regs(148) => 
                           bus_reg_dataout_148_port, regs(147) => 
                           bus_reg_dataout_147_port, regs(146) => 
                           bus_reg_dataout_146_port, regs(145) => 
                           bus_reg_dataout_145_port, regs(144) => 
                           bus_reg_dataout_144_port, regs(143) => 
                           bus_reg_dataout_143_port, regs(142) => 
                           bus_reg_dataout_142_port, regs(141) => 
                           bus_reg_dataout_141_port, regs(140) => 
                           bus_reg_dataout_140_port, regs(139) => 
                           bus_reg_dataout_139_port, regs(138) => 
                           bus_reg_dataout_138_port, regs(137) => 
                           bus_reg_dataout_137_port, regs(136) => 
                           bus_reg_dataout_136_port, regs(135) => 
                           bus_reg_dataout_135_port, regs(134) => 
                           bus_reg_dataout_134_port, regs(133) => 
                           bus_reg_dataout_133_port, regs(132) => 
                           bus_reg_dataout_132_port, regs(131) => 
                           bus_reg_dataout_131_port, regs(130) => 
                           bus_reg_dataout_130_port, regs(129) => 
                           bus_reg_dataout_129_port, regs(128) => 
                           bus_reg_dataout_128_port, regs(127) => 
                           bus_reg_dataout_127_port, regs(126) => 
                           bus_reg_dataout_126_port, regs(125) => 
                           bus_reg_dataout_125_port, regs(124) => 
                           bus_reg_dataout_124_port, regs(123) => 
                           bus_reg_dataout_123_port, regs(122) => 
                           bus_reg_dataout_122_port, regs(121) => 
                           bus_reg_dataout_121_port, regs(120) => 
                           bus_reg_dataout_120_port, regs(119) => 
                           bus_reg_dataout_119_port, regs(118) => 
                           bus_reg_dataout_118_port, regs(117) => 
                           bus_reg_dataout_117_port, regs(116) => 
                           bus_reg_dataout_116_port, regs(115) => 
                           bus_reg_dataout_115_port, regs(114) => 
                           bus_reg_dataout_114_port, regs(113) => 
                           bus_reg_dataout_113_port, regs(112) => 
                           bus_reg_dataout_112_port, regs(111) => 
                           bus_reg_dataout_111_port, regs(110) => 
                           bus_reg_dataout_110_port, regs(109) => 
                           bus_reg_dataout_109_port, regs(108) => 
                           bus_reg_dataout_108_port, regs(107) => 
                           bus_reg_dataout_107_port, regs(106) => 
                           bus_reg_dataout_106_port, regs(105) => 
                           bus_reg_dataout_105_port, regs(104) => 
                           bus_reg_dataout_104_port, regs(103) => 
                           bus_reg_dataout_103_port, regs(102) => 
                           bus_reg_dataout_102_port, regs(101) => 
                           bus_reg_dataout_101_port, regs(100) => 
                           bus_reg_dataout_100_port, regs(99) => 
                           bus_reg_dataout_99_port, regs(98) => 
                           bus_reg_dataout_98_port, regs(97) => 
                           bus_reg_dataout_97_port, regs(96) => 
                           bus_reg_dataout_96_port, regs(95) => 
                           bus_reg_dataout_95_port, regs(94) => 
                           bus_reg_dataout_94_port, regs(93) => 
                           bus_reg_dataout_93_port, regs(92) => 
                           bus_reg_dataout_92_port, regs(91) => 
                           bus_reg_dataout_91_port, regs(90) => 
                           bus_reg_dataout_90_port, regs(89) => 
                           bus_reg_dataout_89_port, regs(88) => 
                           bus_reg_dataout_88_port, regs(87) => 
                           bus_reg_dataout_87_port, regs(86) => 
                           bus_reg_dataout_86_port, regs(85) => 
                           bus_reg_dataout_85_port, regs(84) => 
                           bus_reg_dataout_84_port, regs(83) => 
                           bus_reg_dataout_83_port, regs(82) => 
                           bus_reg_dataout_82_port, regs(81) => 
                           bus_reg_dataout_81_port, regs(80) => 
                           bus_reg_dataout_80_port, regs(79) => 
                           bus_reg_dataout_79_port, regs(78) => 
                           bus_reg_dataout_78_port, regs(77) => 
                           bus_reg_dataout_77_port, regs(76) => 
                           bus_reg_dataout_76_port, regs(75) => 
                           bus_reg_dataout_75_port, regs(74) => 
                           bus_reg_dataout_74_port, regs(73) => 
                           bus_reg_dataout_73_port, regs(72) => 
                           bus_reg_dataout_72_port, regs(71) => 
                           bus_reg_dataout_71_port, regs(70) => 
                           bus_reg_dataout_70_port, regs(69) => 
                           bus_reg_dataout_69_port, regs(68) => 
                           bus_reg_dataout_68_port, regs(67) => 
                           bus_reg_dataout_67_port, regs(66) => 
                           bus_reg_dataout_66_port, regs(65) => 
                           bus_reg_dataout_65_port, regs(64) => 
                           bus_reg_dataout_64_port, regs(63) => 
                           bus_reg_dataout_63_port, regs(62) => 
                           bus_reg_dataout_62_port, regs(61) => 
                           bus_reg_dataout_61_port, regs(60) => 
                           bus_reg_dataout_60_port, regs(59) => 
                           bus_reg_dataout_59_port, regs(58) => 
                           bus_reg_dataout_58_port, regs(57) => 
                           bus_reg_dataout_57_port, regs(56) => 
                           bus_reg_dataout_56_port, regs(55) => 
                           bus_reg_dataout_55_port, regs(54) => 
                           bus_reg_dataout_54_port, regs(53) => 
                           bus_reg_dataout_53_port, regs(52) => 
                           bus_reg_dataout_52_port, regs(51) => 
                           bus_reg_dataout_51_port, regs(50) => 
                           bus_reg_dataout_50_port, regs(49) => 
                           bus_reg_dataout_49_port, regs(48) => 
                           bus_reg_dataout_48_port, regs(47) => 
                           bus_reg_dataout_47_port, regs(46) => 
                           bus_reg_dataout_46_port, regs(45) => 
                           bus_reg_dataout_45_port, regs(44) => 
                           bus_reg_dataout_44_port, regs(43) => 
                           bus_reg_dataout_43_port, regs(42) => 
                           bus_reg_dataout_42_port, regs(41) => 
                           bus_reg_dataout_41_port, regs(40) => 
                           bus_reg_dataout_40_port, regs(39) => 
                           bus_reg_dataout_39_port, regs(38) => 
                           bus_reg_dataout_38_port, regs(37) => 
                           bus_reg_dataout_37_port, regs(36) => 
                           bus_reg_dataout_36_port, regs(35) => 
                           bus_reg_dataout_35_port, regs(34) => 
                           bus_reg_dataout_34_port, regs(33) => 
                           bus_reg_dataout_33_port, regs(32) => 
                           bus_reg_dataout_32_port, regs(31) => 
                           bus_reg_dataout_31_port, regs(30) => 
                           bus_reg_dataout_30_port, regs(29) => 
                           bus_reg_dataout_29_port, regs(28) => 
                           bus_reg_dataout_28_port, regs(27) => 
                           bus_reg_dataout_27_port, regs(26) => 
                           bus_reg_dataout_26_port, regs(25) => 
                           bus_reg_dataout_25_port, regs(24) => 
                           bus_reg_dataout_24_port, regs(23) => 
                           bus_reg_dataout_23_port, regs(22) => 
                           bus_reg_dataout_22_port, regs(21) => 
                           bus_reg_dataout_21_port, regs(20) => 
                           bus_reg_dataout_20_port, regs(19) => 
                           bus_reg_dataout_19_port, regs(18) => 
                           bus_reg_dataout_18_port, regs(17) => 
                           bus_reg_dataout_17_port, regs(16) => 
                           bus_reg_dataout_16_port, regs(15) => 
                           bus_reg_dataout_15_port, regs(14) => 
                           bus_reg_dataout_14_port, regs(13) => 
                           bus_reg_dataout_13_port, regs(12) => 
                           bus_reg_dataout_12_port, regs(11) => 
                           bus_reg_dataout_11_port, regs(10) => 
                           bus_reg_dataout_10_port, regs(9) => 
                           bus_reg_dataout_9_port, regs(8) => 
                           bus_reg_dataout_8_port, regs(7) => 
                           bus_reg_dataout_7_port, regs(6) => 
                           bus_reg_dataout_6_port, regs(5) => 
                           bus_reg_dataout_5_port, regs(4) => 
                           bus_reg_dataout_4_port, regs(3) => 
                           bus_reg_dataout_3_port, regs(2) => 
                           bus_reg_dataout_2_port, regs(1) => 
                           bus_reg_dataout_1_port, regs(0) => 
                           bus_reg_dataout_0_port, win(4) => c_swin_4_port, 
                           win(3) => c_swin_3_port, win(2) => c_swin_2_port, 
                           win(1) => c_swin_1_port, win(0) => c_swin_0_port, 
                           curr_proc_regs(511) => 
                           bus_sel_savedwin_data_511_port, curr_proc_regs(510) 
                           => bus_sel_savedwin_data_510_port, 
                           curr_proc_regs(509) => 
                           bus_sel_savedwin_data_509_port, curr_proc_regs(508) 
                           => bus_sel_savedwin_data_508_port, 
                           curr_proc_regs(507) => 
                           bus_sel_savedwin_data_507_port, curr_proc_regs(506) 
                           => bus_sel_savedwin_data_506_port, 
                           curr_proc_regs(505) => 
                           bus_sel_savedwin_data_505_port, curr_proc_regs(504) 
                           => bus_sel_savedwin_data_504_port, 
                           curr_proc_regs(503) => 
                           bus_sel_savedwin_data_503_port, curr_proc_regs(502) 
                           => bus_sel_savedwin_data_502_port, 
                           curr_proc_regs(501) => 
                           bus_sel_savedwin_data_501_port, curr_proc_regs(500) 
                           => bus_sel_savedwin_data_500_port, 
                           curr_proc_regs(499) => 
                           bus_sel_savedwin_data_499_port, curr_proc_regs(498) 
                           => bus_sel_savedwin_data_498_port, 
                           curr_proc_regs(497) => 
                           bus_sel_savedwin_data_497_port, curr_proc_regs(496) 
                           => bus_sel_savedwin_data_496_port, 
                           curr_proc_regs(495) => 
                           bus_sel_savedwin_data_495_port, curr_proc_regs(494) 
                           => bus_sel_savedwin_data_494_port, 
                           curr_proc_regs(493) => 
                           bus_sel_savedwin_data_493_port, curr_proc_regs(492) 
                           => bus_sel_savedwin_data_492_port, 
                           curr_proc_regs(491) => 
                           bus_sel_savedwin_data_491_port, curr_proc_regs(490) 
                           => bus_sel_savedwin_data_490_port, 
                           curr_proc_regs(489) => 
                           bus_sel_savedwin_data_489_port, curr_proc_regs(488) 
                           => bus_sel_savedwin_data_488_port, 
                           curr_proc_regs(487) => 
                           bus_sel_savedwin_data_487_port, curr_proc_regs(486) 
                           => bus_sel_savedwin_data_486_port, 
                           curr_proc_regs(485) => 
                           bus_sel_savedwin_data_485_port, curr_proc_regs(484) 
                           => bus_sel_savedwin_data_484_port, 
                           curr_proc_regs(483) => 
                           bus_sel_savedwin_data_483_port, curr_proc_regs(482) 
                           => bus_sel_savedwin_data_482_port, 
                           curr_proc_regs(481) => 
                           bus_sel_savedwin_data_481_port, curr_proc_regs(480) 
                           => bus_sel_savedwin_data_480_port, 
                           curr_proc_regs(479) => 
                           bus_sel_savedwin_data_479_port, curr_proc_regs(478) 
                           => bus_sel_savedwin_data_478_port, 
                           curr_proc_regs(477) => 
                           bus_sel_savedwin_data_477_port, curr_proc_regs(476) 
                           => bus_sel_savedwin_data_476_port, 
                           curr_proc_regs(475) => 
                           bus_sel_savedwin_data_475_port, curr_proc_regs(474) 
                           => bus_sel_savedwin_data_474_port, 
                           curr_proc_regs(473) => 
                           bus_sel_savedwin_data_473_port, curr_proc_regs(472) 
                           => bus_sel_savedwin_data_472_port, 
                           curr_proc_regs(471) => 
                           bus_sel_savedwin_data_471_port, curr_proc_regs(470) 
                           => bus_sel_savedwin_data_470_port, 
                           curr_proc_regs(469) => 
                           bus_sel_savedwin_data_469_port, curr_proc_regs(468) 
                           => bus_sel_savedwin_data_468_port, 
                           curr_proc_regs(467) => 
                           bus_sel_savedwin_data_467_port, curr_proc_regs(466) 
                           => bus_sel_savedwin_data_466_port, 
                           curr_proc_regs(465) => 
                           bus_sel_savedwin_data_465_port, curr_proc_regs(464) 
                           => bus_sel_savedwin_data_464_port, 
                           curr_proc_regs(463) => 
                           bus_sel_savedwin_data_463_port, curr_proc_regs(462) 
                           => bus_sel_savedwin_data_462_port, 
                           curr_proc_regs(461) => 
                           bus_sel_savedwin_data_461_port, curr_proc_regs(460) 
                           => bus_sel_savedwin_data_460_port, 
                           curr_proc_regs(459) => 
                           bus_sel_savedwin_data_459_port, curr_proc_regs(458) 
                           => bus_sel_savedwin_data_458_port, 
                           curr_proc_regs(457) => 
                           bus_sel_savedwin_data_457_port, curr_proc_regs(456) 
                           => bus_sel_savedwin_data_456_port, 
                           curr_proc_regs(455) => 
                           bus_sel_savedwin_data_455_port, curr_proc_regs(454) 
                           => bus_sel_savedwin_data_454_port, 
                           curr_proc_regs(453) => 
                           bus_sel_savedwin_data_453_port, curr_proc_regs(452) 
                           => bus_sel_savedwin_data_452_port, 
                           curr_proc_regs(451) => 
                           bus_sel_savedwin_data_451_port, curr_proc_regs(450) 
                           => bus_sel_savedwin_data_450_port, 
                           curr_proc_regs(449) => 
                           bus_sel_savedwin_data_449_port, curr_proc_regs(448) 
                           => bus_sel_savedwin_data_448_port, 
                           curr_proc_regs(447) => 
                           bus_sel_savedwin_data_447_port, curr_proc_regs(446) 
                           => bus_sel_savedwin_data_446_port, 
                           curr_proc_regs(445) => 
                           bus_sel_savedwin_data_445_port, curr_proc_regs(444) 
                           => bus_sel_savedwin_data_444_port, 
                           curr_proc_regs(443) => 
                           bus_sel_savedwin_data_443_port, curr_proc_regs(442) 
                           => bus_sel_savedwin_data_442_port, 
                           curr_proc_regs(441) => 
                           bus_sel_savedwin_data_441_port, curr_proc_regs(440) 
                           => bus_sel_savedwin_data_440_port, 
                           curr_proc_regs(439) => 
                           bus_sel_savedwin_data_439_port, curr_proc_regs(438) 
                           => bus_sel_savedwin_data_438_port, 
                           curr_proc_regs(437) => 
                           bus_sel_savedwin_data_437_port, curr_proc_regs(436) 
                           => bus_sel_savedwin_data_436_port, 
                           curr_proc_regs(435) => 
                           bus_sel_savedwin_data_435_port, curr_proc_regs(434) 
                           => bus_sel_savedwin_data_434_port, 
                           curr_proc_regs(433) => 
                           bus_sel_savedwin_data_433_port, curr_proc_regs(432) 
                           => bus_sel_savedwin_data_432_port, 
                           curr_proc_regs(431) => 
                           bus_sel_savedwin_data_431_port, curr_proc_regs(430) 
                           => bus_sel_savedwin_data_430_port, 
                           curr_proc_regs(429) => 
                           bus_sel_savedwin_data_429_port, curr_proc_regs(428) 
                           => bus_sel_savedwin_data_428_port, 
                           curr_proc_regs(427) => 
                           bus_sel_savedwin_data_427_port, curr_proc_regs(426) 
                           => bus_sel_savedwin_data_426_port, 
                           curr_proc_regs(425) => 
                           bus_sel_savedwin_data_425_port, curr_proc_regs(424) 
                           => bus_sel_savedwin_data_424_port, 
                           curr_proc_regs(423) => 
                           bus_sel_savedwin_data_423_port, curr_proc_regs(422) 
                           => bus_sel_savedwin_data_422_port, 
                           curr_proc_regs(421) => 
                           bus_sel_savedwin_data_421_port, curr_proc_regs(420) 
                           => bus_sel_savedwin_data_420_port, 
                           curr_proc_regs(419) => 
                           bus_sel_savedwin_data_419_port, curr_proc_regs(418) 
                           => bus_sel_savedwin_data_418_port, 
                           curr_proc_regs(417) => 
                           bus_sel_savedwin_data_417_port, curr_proc_regs(416) 
                           => bus_sel_savedwin_data_416_port, 
                           curr_proc_regs(415) => 
                           bus_sel_savedwin_data_415_port, curr_proc_regs(414) 
                           => bus_sel_savedwin_data_414_port, 
                           curr_proc_regs(413) => 
                           bus_sel_savedwin_data_413_port, curr_proc_regs(412) 
                           => bus_sel_savedwin_data_412_port, 
                           curr_proc_regs(411) => 
                           bus_sel_savedwin_data_411_port, curr_proc_regs(410) 
                           => bus_sel_savedwin_data_410_port, 
                           curr_proc_regs(409) => 
                           bus_sel_savedwin_data_409_port, curr_proc_regs(408) 
                           => bus_sel_savedwin_data_408_port, 
                           curr_proc_regs(407) => 
                           bus_sel_savedwin_data_407_port, curr_proc_regs(406) 
                           => bus_sel_savedwin_data_406_port, 
                           curr_proc_regs(405) => 
                           bus_sel_savedwin_data_405_port, curr_proc_regs(404) 
                           => bus_sel_savedwin_data_404_port, 
                           curr_proc_regs(403) => 
                           bus_sel_savedwin_data_403_port, curr_proc_regs(402) 
                           => bus_sel_savedwin_data_402_port, 
                           curr_proc_regs(401) => 
                           bus_sel_savedwin_data_401_port, curr_proc_regs(400) 
                           => bus_sel_savedwin_data_400_port, 
                           curr_proc_regs(399) => 
                           bus_sel_savedwin_data_399_port, curr_proc_regs(398) 
                           => bus_sel_savedwin_data_398_port, 
                           curr_proc_regs(397) => 
                           bus_sel_savedwin_data_397_port, curr_proc_regs(396) 
                           => bus_sel_savedwin_data_396_port, 
                           curr_proc_regs(395) => 
                           bus_sel_savedwin_data_395_port, curr_proc_regs(394) 
                           => bus_sel_savedwin_data_394_port, 
                           curr_proc_regs(393) => 
                           bus_sel_savedwin_data_393_port, curr_proc_regs(392) 
                           => bus_sel_savedwin_data_392_port, 
                           curr_proc_regs(391) => 
                           bus_sel_savedwin_data_391_port, curr_proc_regs(390) 
                           => bus_sel_savedwin_data_390_port, 
                           curr_proc_regs(389) => 
                           bus_sel_savedwin_data_389_port, curr_proc_regs(388) 
                           => bus_sel_savedwin_data_388_port, 
                           curr_proc_regs(387) => 
                           bus_sel_savedwin_data_387_port, curr_proc_regs(386) 
                           => bus_sel_savedwin_data_386_port, 
                           curr_proc_regs(385) => 
                           bus_sel_savedwin_data_385_port, curr_proc_regs(384) 
                           => bus_sel_savedwin_data_384_port, 
                           curr_proc_regs(383) => 
                           bus_sel_savedwin_data_383_port, curr_proc_regs(382) 
                           => bus_sel_savedwin_data_382_port, 
                           curr_proc_regs(381) => 
                           bus_sel_savedwin_data_381_port, curr_proc_regs(380) 
                           => bus_sel_savedwin_data_380_port, 
                           curr_proc_regs(379) => 
                           bus_sel_savedwin_data_379_port, curr_proc_regs(378) 
                           => bus_sel_savedwin_data_378_port, 
                           curr_proc_regs(377) => 
                           bus_sel_savedwin_data_377_port, curr_proc_regs(376) 
                           => bus_sel_savedwin_data_376_port, 
                           curr_proc_regs(375) => 
                           bus_sel_savedwin_data_375_port, curr_proc_regs(374) 
                           => bus_sel_savedwin_data_374_port, 
                           curr_proc_regs(373) => 
                           bus_sel_savedwin_data_373_port, curr_proc_regs(372) 
                           => bus_sel_savedwin_data_372_port, 
                           curr_proc_regs(371) => 
                           bus_sel_savedwin_data_371_port, curr_proc_regs(370) 
                           => bus_sel_savedwin_data_370_port, 
                           curr_proc_regs(369) => 
                           bus_sel_savedwin_data_369_port, curr_proc_regs(368) 
                           => bus_sel_savedwin_data_368_port, 
                           curr_proc_regs(367) => 
                           bus_sel_savedwin_data_367_port, curr_proc_regs(366) 
                           => bus_sel_savedwin_data_366_port, 
                           curr_proc_regs(365) => 
                           bus_sel_savedwin_data_365_port, curr_proc_regs(364) 
                           => bus_sel_savedwin_data_364_port, 
                           curr_proc_regs(363) => 
                           bus_sel_savedwin_data_363_port, curr_proc_regs(362) 
                           => bus_sel_savedwin_data_362_port, 
                           curr_proc_regs(361) => 
                           bus_sel_savedwin_data_361_port, curr_proc_regs(360) 
                           => bus_sel_savedwin_data_360_port, 
                           curr_proc_regs(359) => 
                           bus_sel_savedwin_data_359_port, curr_proc_regs(358) 
                           => bus_sel_savedwin_data_358_port, 
                           curr_proc_regs(357) => 
                           bus_sel_savedwin_data_357_port, curr_proc_regs(356) 
                           => bus_sel_savedwin_data_356_port, 
                           curr_proc_regs(355) => 
                           bus_sel_savedwin_data_355_port, curr_proc_regs(354) 
                           => bus_sel_savedwin_data_354_port, 
                           curr_proc_regs(353) => 
                           bus_sel_savedwin_data_353_port, curr_proc_regs(352) 
                           => bus_sel_savedwin_data_352_port, 
                           curr_proc_regs(351) => 
                           bus_sel_savedwin_data_351_port, curr_proc_regs(350) 
                           => bus_sel_savedwin_data_350_port, 
                           curr_proc_regs(349) => 
                           bus_sel_savedwin_data_349_port, curr_proc_regs(348) 
                           => bus_sel_savedwin_data_348_port, 
                           curr_proc_regs(347) => 
                           bus_sel_savedwin_data_347_port, curr_proc_regs(346) 
                           => bus_sel_savedwin_data_346_port, 
                           curr_proc_regs(345) => 
                           bus_sel_savedwin_data_345_port, curr_proc_regs(344) 
                           => bus_sel_savedwin_data_344_port, 
                           curr_proc_regs(343) => 
                           bus_sel_savedwin_data_343_port, curr_proc_regs(342) 
                           => bus_sel_savedwin_data_342_port, 
                           curr_proc_regs(341) => 
                           bus_sel_savedwin_data_341_port, curr_proc_regs(340) 
                           => bus_sel_savedwin_data_340_port, 
                           curr_proc_regs(339) => 
                           bus_sel_savedwin_data_339_port, curr_proc_regs(338) 
                           => bus_sel_savedwin_data_338_port, 
                           curr_proc_regs(337) => 
                           bus_sel_savedwin_data_337_port, curr_proc_regs(336) 
                           => bus_sel_savedwin_data_336_port, 
                           curr_proc_regs(335) => 
                           bus_sel_savedwin_data_335_port, curr_proc_regs(334) 
                           => bus_sel_savedwin_data_334_port, 
                           curr_proc_regs(333) => 
                           bus_sel_savedwin_data_333_port, curr_proc_regs(332) 
                           => bus_sel_savedwin_data_332_port, 
                           curr_proc_regs(331) => 
                           bus_sel_savedwin_data_331_port, curr_proc_regs(330) 
                           => bus_sel_savedwin_data_330_port, 
                           curr_proc_regs(329) => 
                           bus_sel_savedwin_data_329_port, curr_proc_regs(328) 
                           => bus_sel_savedwin_data_328_port, 
                           curr_proc_regs(327) => 
                           bus_sel_savedwin_data_327_port, curr_proc_regs(326) 
                           => bus_sel_savedwin_data_326_port, 
                           curr_proc_regs(325) => 
                           bus_sel_savedwin_data_325_port, curr_proc_regs(324) 
                           => bus_sel_savedwin_data_324_port, 
                           curr_proc_regs(323) => 
                           bus_sel_savedwin_data_323_port, curr_proc_regs(322) 
                           => bus_sel_savedwin_data_322_port, 
                           curr_proc_regs(321) => 
                           bus_sel_savedwin_data_321_port, curr_proc_regs(320) 
                           => bus_sel_savedwin_data_320_port, 
                           curr_proc_regs(319) => 
                           bus_sel_savedwin_data_319_port, curr_proc_regs(318) 
                           => bus_sel_savedwin_data_318_port, 
                           curr_proc_regs(317) => 
                           bus_sel_savedwin_data_317_port, curr_proc_regs(316) 
                           => bus_sel_savedwin_data_316_port, 
                           curr_proc_regs(315) => 
                           bus_sel_savedwin_data_315_port, curr_proc_regs(314) 
                           => bus_sel_savedwin_data_314_port, 
                           curr_proc_regs(313) => 
                           bus_sel_savedwin_data_313_port, curr_proc_regs(312) 
                           => bus_sel_savedwin_data_312_port, 
                           curr_proc_regs(311) => 
                           bus_sel_savedwin_data_311_port, curr_proc_regs(310) 
                           => bus_sel_savedwin_data_310_port, 
                           curr_proc_regs(309) => 
                           bus_sel_savedwin_data_309_port, curr_proc_regs(308) 
                           => bus_sel_savedwin_data_308_port, 
                           curr_proc_regs(307) => 
                           bus_sel_savedwin_data_307_port, curr_proc_regs(306) 
                           => bus_sel_savedwin_data_306_port, 
                           curr_proc_regs(305) => 
                           bus_sel_savedwin_data_305_port, curr_proc_regs(304) 
                           => bus_sel_savedwin_data_304_port, 
                           curr_proc_regs(303) => 
                           bus_sel_savedwin_data_303_port, curr_proc_regs(302) 
                           => bus_sel_savedwin_data_302_port, 
                           curr_proc_regs(301) => 
                           bus_sel_savedwin_data_301_port, curr_proc_regs(300) 
                           => bus_sel_savedwin_data_300_port, 
                           curr_proc_regs(299) => 
                           bus_sel_savedwin_data_299_port, curr_proc_regs(298) 
                           => bus_sel_savedwin_data_298_port, 
                           curr_proc_regs(297) => 
                           bus_sel_savedwin_data_297_port, curr_proc_regs(296) 
                           => bus_sel_savedwin_data_296_port, 
                           curr_proc_regs(295) => 
                           bus_sel_savedwin_data_295_port, curr_proc_regs(294) 
                           => bus_sel_savedwin_data_294_port, 
                           curr_proc_regs(293) => 
                           bus_sel_savedwin_data_293_port, curr_proc_regs(292) 
                           => bus_sel_savedwin_data_292_port, 
                           curr_proc_regs(291) => 
                           bus_sel_savedwin_data_291_port, curr_proc_regs(290) 
                           => bus_sel_savedwin_data_290_port, 
                           curr_proc_regs(289) => 
                           bus_sel_savedwin_data_289_port, curr_proc_regs(288) 
                           => bus_sel_savedwin_data_288_port, 
                           curr_proc_regs(287) => 
                           bus_sel_savedwin_data_287_port, curr_proc_regs(286) 
                           => bus_sel_savedwin_data_286_port, 
                           curr_proc_regs(285) => 
                           bus_sel_savedwin_data_285_port, curr_proc_regs(284) 
                           => bus_sel_savedwin_data_284_port, 
                           curr_proc_regs(283) => 
                           bus_sel_savedwin_data_283_port, curr_proc_regs(282) 
                           => bus_sel_savedwin_data_282_port, 
                           curr_proc_regs(281) => 
                           bus_sel_savedwin_data_281_port, curr_proc_regs(280) 
                           => bus_sel_savedwin_data_280_port, 
                           curr_proc_regs(279) => 
                           bus_sel_savedwin_data_279_port, curr_proc_regs(278) 
                           => bus_sel_savedwin_data_278_port, 
                           curr_proc_regs(277) => 
                           bus_sel_savedwin_data_277_port, curr_proc_regs(276) 
                           => bus_sel_savedwin_data_276_port, 
                           curr_proc_regs(275) => 
                           bus_sel_savedwin_data_275_port, curr_proc_regs(274) 
                           => bus_sel_savedwin_data_274_port, 
                           curr_proc_regs(273) => 
                           bus_sel_savedwin_data_273_port, curr_proc_regs(272) 
                           => bus_sel_savedwin_data_272_port, 
                           curr_proc_regs(271) => 
                           bus_sel_savedwin_data_271_port, curr_proc_regs(270) 
                           => bus_sel_savedwin_data_270_port, 
                           curr_proc_regs(269) => 
                           bus_sel_savedwin_data_269_port, curr_proc_regs(268) 
                           => bus_sel_savedwin_data_268_port, 
                           curr_proc_regs(267) => 
                           bus_sel_savedwin_data_267_port, curr_proc_regs(266) 
                           => bus_sel_savedwin_data_266_port, 
                           curr_proc_regs(265) => 
                           bus_sel_savedwin_data_265_port, curr_proc_regs(264) 
                           => bus_sel_savedwin_data_264_port, 
                           curr_proc_regs(263) => 
                           bus_sel_savedwin_data_263_port, curr_proc_regs(262) 
                           => bus_sel_savedwin_data_262_port, 
                           curr_proc_regs(261) => 
                           bus_sel_savedwin_data_261_port, curr_proc_regs(260) 
                           => bus_sel_savedwin_data_260_port, 
                           curr_proc_regs(259) => 
                           bus_sel_savedwin_data_259_port, curr_proc_regs(258) 
                           => bus_sel_savedwin_data_258_port, 
                           curr_proc_regs(257) => 
                           bus_sel_savedwin_data_257_port, curr_proc_regs(256) 
                           => bus_sel_savedwin_data_256_port, 
                           curr_proc_regs(255) => 
                           bus_sel_savedwin_data_255_port, curr_proc_regs(254) 
                           => bus_sel_savedwin_data_254_port, 
                           curr_proc_regs(253) => 
                           bus_sel_savedwin_data_253_port, curr_proc_regs(252) 
                           => bus_sel_savedwin_data_252_port, 
                           curr_proc_regs(251) => 
                           bus_sel_savedwin_data_251_port, curr_proc_regs(250) 
                           => bus_sel_savedwin_data_250_port, 
                           curr_proc_regs(249) => 
                           bus_sel_savedwin_data_249_port, curr_proc_regs(248) 
                           => bus_sel_savedwin_data_248_port, 
                           curr_proc_regs(247) => 
                           bus_sel_savedwin_data_247_port, curr_proc_regs(246) 
                           => bus_sel_savedwin_data_246_port, 
                           curr_proc_regs(245) => 
                           bus_sel_savedwin_data_245_port, curr_proc_regs(244) 
                           => bus_sel_savedwin_data_244_port, 
                           curr_proc_regs(243) => 
                           bus_sel_savedwin_data_243_port, curr_proc_regs(242) 
                           => bus_sel_savedwin_data_242_port, 
                           curr_proc_regs(241) => 
                           bus_sel_savedwin_data_241_port, curr_proc_regs(240) 
                           => bus_sel_savedwin_data_240_port, 
                           curr_proc_regs(239) => 
                           bus_sel_savedwin_data_239_port, curr_proc_regs(238) 
                           => bus_sel_savedwin_data_238_port, 
                           curr_proc_regs(237) => 
                           bus_sel_savedwin_data_237_port, curr_proc_regs(236) 
                           => bus_sel_savedwin_data_236_port, 
                           curr_proc_regs(235) => 
                           bus_sel_savedwin_data_235_port, curr_proc_regs(234) 
                           => bus_sel_savedwin_data_234_port, 
                           curr_proc_regs(233) => 
                           bus_sel_savedwin_data_233_port, curr_proc_regs(232) 
                           => bus_sel_savedwin_data_232_port, 
                           curr_proc_regs(231) => 
                           bus_sel_savedwin_data_231_port, curr_proc_regs(230) 
                           => bus_sel_savedwin_data_230_port, 
                           curr_proc_regs(229) => 
                           bus_sel_savedwin_data_229_port, curr_proc_regs(228) 
                           => bus_sel_savedwin_data_228_port, 
                           curr_proc_regs(227) => 
                           bus_sel_savedwin_data_227_port, curr_proc_regs(226) 
                           => bus_sel_savedwin_data_226_port, 
                           curr_proc_regs(225) => 
                           bus_sel_savedwin_data_225_port, curr_proc_regs(224) 
                           => bus_sel_savedwin_data_224_port, 
                           curr_proc_regs(223) => 
                           bus_sel_savedwin_data_223_port, curr_proc_regs(222) 
                           => bus_sel_savedwin_data_222_port, 
                           curr_proc_regs(221) => 
                           bus_sel_savedwin_data_221_port, curr_proc_regs(220) 
                           => bus_sel_savedwin_data_220_port, 
                           curr_proc_regs(219) => 
                           bus_sel_savedwin_data_219_port, curr_proc_regs(218) 
                           => bus_sel_savedwin_data_218_port, 
                           curr_proc_regs(217) => 
                           bus_sel_savedwin_data_217_port, curr_proc_regs(216) 
                           => bus_sel_savedwin_data_216_port, 
                           curr_proc_regs(215) => 
                           bus_sel_savedwin_data_215_port, curr_proc_regs(214) 
                           => bus_sel_savedwin_data_214_port, 
                           curr_proc_regs(213) => 
                           bus_sel_savedwin_data_213_port, curr_proc_regs(212) 
                           => bus_sel_savedwin_data_212_port, 
                           curr_proc_regs(211) => 
                           bus_sel_savedwin_data_211_port, curr_proc_regs(210) 
                           => bus_sel_savedwin_data_210_port, 
                           curr_proc_regs(209) => 
                           bus_sel_savedwin_data_209_port, curr_proc_regs(208) 
                           => bus_sel_savedwin_data_208_port, 
                           curr_proc_regs(207) => 
                           bus_sel_savedwin_data_207_port, curr_proc_regs(206) 
                           => bus_sel_savedwin_data_206_port, 
                           curr_proc_regs(205) => 
                           bus_sel_savedwin_data_205_port, curr_proc_regs(204) 
                           => bus_sel_savedwin_data_204_port, 
                           curr_proc_regs(203) => 
                           bus_sel_savedwin_data_203_port, curr_proc_regs(202) 
                           => bus_sel_savedwin_data_202_port, 
                           curr_proc_regs(201) => 
                           bus_sel_savedwin_data_201_port, curr_proc_regs(200) 
                           => bus_sel_savedwin_data_200_port, 
                           curr_proc_regs(199) => 
                           bus_sel_savedwin_data_199_port, curr_proc_regs(198) 
                           => bus_sel_savedwin_data_198_port, 
                           curr_proc_regs(197) => 
                           bus_sel_savedwin_data_197_port, curr_proc_regs(196) 
                           => bus_sel_savedwin_data_196_port, 
                           curr_proc_regs(195) => 
                           bus_sel_savedwin_data_195_port, curr_proc_regs(194) 
                           => bus_sel_savedwin_data_194_port, 
                           curr_proc_regs(193) => 
                           bus_sel_savedwin_data_193_port, curr_proc_regs(192) 
                           => bus_sel_savedwin_data_192_port, 
                           curr_proc_regs(191) => 
                           bus_sel_savedwin_data_191_port, curr_proc_regs(190) 
                           => bus_sel_savedwin_data_190_port, 
                           curr_proc_regs(189) => 
                           bus_sel_savedwin_data_189_port, curr_proc_regs(188) 
                           => bus_sel_savedwin_data_188_port, 
                           curr_proc_regs(187) => 
                           bus_sel_savedwin_data_187_port, curr_proc_regs(186) 
                           => bus_sel_savedwin_data_186_port, 
                           curr_proc_regs(185) => 
                           bus_sel_savedwin_data_185_port, curr_proc_regs(184) 
                           => bus_sel_savedwin_data_184_port, 
                           curr_proc_regs(183) => 
                           bus_sel_savedwin_data_183_port, curr_proc_regs(182) 
                           => bus_sel_savedwin_data_182_port, 
                           curr_proc_regs(181) => 
                           bus_sel_savedwin_data_181_port, curr_proc_regs(180) 
                           => bus_sel_savedwin_data_180_port, 
                           curr_proc_regs(179) => 
                           bus_sel_savedwin_data_179_port, curr_proc_regs(178) 
                           => bus_sel_savedwin_data_178_port, 
                           curr_proc_regs(177) => 
                           bus_sel_savedwin_data_177_port, curr_proc_regs(176) 
                           => bus_sel_savedwin_data_176_port, 
                           curr_proc_regs(175) => 
                           bus_sel_savedwin_data_175_port, curr_proc_regs(174) 
                           => bus_sel_savedwin_data_174_port, 
                           curr_proc_regs(173) => 
                           bus_sel_savedwin_data_173_port, curr_proc_regs(172) 
                           => bus_sel_savedwin_data_172_port, 
                           curr_proc_regs(171) => 
                           bus_sel_savedwin_data_171_port, curr_proc_regs(170) 
                           => bus_sel_savedwin_data_170_port, 
                           curr_proc_regs(169) => 
                           bus_sel_savedwin_data_169_port, curr_proc_regs(168) 
                           => bus_sel_savedwin_data_168_port, 
                           curr_proc_regs(167) => 
                           bus_sel_savedwin_data_167_port, curr_proc_regs(166) 
                           => bus_sel_savedwin_data_166_port, 
                           curr_proc_regs(165) => 
                           bus_sel_savedwin_data_165_port, curr_proc_regs(164) 
                           => bus_sel_savedwin_data_164_port, 
                           curr_proc_regs(163) => 
                           bus_sel_savedwin_data_163_port, curr_proc_regs(162) 
                           => bus_sel_savedwin_data_162_port, 
                           curr_proc_regs(161) => 
                           bus_sel_savedwin_data_161_port, curr_proc_regs(160) 
                           => bus_sel_savedwin_data_160_port, 
                           curr_proc_regs(159) => 
                           bus_sel_savedwin_data_159_port, curr_proc_regs(158) 
                           => bus_sel_savedwin_data_158_port, 
                           curr_proc_regs(157) => 
                           bus_sel_savedwin_data_157_port, curr_proc_regs(156) 
                           => bus_sel_savedwin_data_156_port, 
                           curr_proc_regs(155) => 
                           bus_sel_savedwin_data_155_port, curr_proc_regs(154) 
                           => bus_sel_savedwin_data_154_port, 
                           curr_proc_regs(153) => 
                           bus_sel_savedwin_data_153_port, curr_proc_regs(152) 
                           => bus_sel_savedwin_data_152_port, 
                           curr_proc_regs(151) => 
                           bus_sel_savedwin_data_151_port, curr_proc_regs(150) 
                           => bus_sel_savedwin_data_150_port, 
                           curr_proc_regs(149) => 
                           bus_sel_savedwin_data_149_port, curr_proc_regs(148) 
                           => bus_sel_savedwin_data_148_port, 
                           curr_proc_regs(147) => 
                           bus_sel_savedwin_data_147_port, curr_proc_regs(146) 
                           => bus_sel_savedwin_data_146_port, 
                           curr_proc_regs(145) => 
                           bus_sel_savedwin_data_145_port, curr_proc_regs(144) 
                           => bus_sel_savedwin_data_144_port, 
                           curr_proc_regs(143) => 
                           bus_sel_savedwin_data_143_port, curr_proc_regs(142) 
                           => bus_sel_savedwin_data_142_port, 
                           curr_proc_regs(141) => 
                           bus_sel_savedwin_data_141_port, curr_proc_regs(140) 
                           => bus_sel_savedwin_data_140_port, 
                           curr_proc_regs(139) => 
                           bus_sel_savedwin_data_139_port, curr_proc_regs(138) 
                           => bus_sel_savedwin_data_138_port, 
                           curr_proc_regs(137) => 
                           bus_sel_savedwin_data_137_port, curr_proc_regs(136) 
                           => bus_sel_savedwin_data_136_port, 
                           curr_proc_regs(135) => 
                           bus_sel_savedwin_data_135_port, curr_proc_regs(134) 
                           => bus_sel_savedwin_data_134_port, 
                           curr_proc_regs(133) => 
                           bus_sel_savedwin_data_133_port, curr_proc_regs(132) 
                           => bus_sel_savedwin_data_132_port, 
                           curr_proc_regs(131) => 
                           bus_sel_savedwin_data_131_port, curr_proc_regs(130) 
                           => bus_sel_savedwin_data_130_port, 
                           curr_proc_regs(129) => 
                           bus_sel_savedwin_data_129_port, curr_proc_regs(128) 
                           => bus_sel_savedwin_data_128_port, 
                           curr_proc_regs(127) => 
                           bus_sel_savedwin_data_127_port, curr_proc_regs(126) 
                           => bus_sel_savedwin_data_126_port, 
                           curr_proc_regs(125) => 
                           bus_sel_savedwin_data_125_port, curr_proc_regs(124) 
                           => bus_sel_savedwin_data_124_port, 
                           curr_proc_regs(123) => 
                           bus_sel_savedwin_data_123_port, curr_proc_regs(122) 
                           => bus_sel_savedwin_data_122_port, 
                           curr_proc_regs(121) => 
                           bus_sel_savedwin_data_121_port, curr_proc_regs(120) 
                           => bus_sel_savedwin_data_120_port, 
                           curr_proc_regs(119) => 
                           bus_sel_savedwin_data_119_port, curr_proc_regs(118) 
                           => bus_sel_savedwin_data_118_port, 
                           curr_proc_regs(117) => 
                           bus_sel_savedwin_data_117_port, curr_proc_regs(116) 
                           => bus_sel_savedwin_data_116_port, 
                           curr_proc_regs(115) => 
                           bus_sel_savedwin_data_115_port, curr_proc_regs(114) 
                           => bus_sel_savedwin_data_114_port, 
                           curr_proc_regs(113) => 
                           bus_sel_savedwin_data_113_port, curr_proc_regs(112) 
                           => bus_sel_savedwin_data_112_port, 
                           curr_proc_regs(111) => 
                           bus_sel_savedwin_data_111_port, curr_proc_regs(110) 
                           => bus_sel_savedwin_data_110_port, 
                           curr_proc_regs(109) => 
                           bus_sel_savedwin_data_109_port, curr_proc_regs(108) 
                           => bus_sel_savedwin_data_108_port, 
                           curr_proc_regs(107) => 
                           bus_sel_savedwin_data_107_port, curr_proc_regs(106) 
                           => bus_sel_savedwin_data_106_port, 
                           curr_proc_regs(105) => 
                           bus_sel_savedwin_data_105_port, curr_proc_regs(104) 
                           => bus_sel_savedwin_data_104_port, 
                           curr_proc_regs(103) => 
                           bus_sel_savedwin_data_103_port, curr_proc_regs(102) 
                           => bus_sel_savedwin_data_102_port, 
                           curr_proc_regs(101) => 
                           bus_sel_savedwin_data_101_port, curr_proc_regs(100) 
                           => bus_sel_savedwin_data_100_port, 
                           curr_proc_regs(99) => bus_sel_savedwin_data_99_port,
                           curr_proc_regs(98) => bus_sel_savedwin_data_98_port,
                           curr_proc_regs(97) => bus_sel_savedwin_data_97_port,
                           curr_proc_regs(96) => bus_sel_savedwin_data_96_port,
                           curr_proc_regs(95) => bus_sel_savedwin_data_95_port,
                           curr_proc_regs(94) => bus_sel_savedwin_data_94_port,
                           curr_proc_regs(93) => bus_sel_savedwin_data_93_port,
                           curr_proc_regs(92) => bus_sel_savedwin_data_92_port,
                           curr_proc_regs(91) => bus_sel_savedwin_data_91_port,
                           curr_proc_regs(90) => bus_sel_savedwin_data_90_port,
                           curr_proc_regs(89) => bus_sel_savedwin_data_89_port,
                           curr_proc_regs(88) => bus_sel_savedwin_data_88_port,
                           curr_proc_regs(87) => bus_sel_savedwin_data_87_port,
                           curr_proc_regs(86) => bus_sel_savedwin_data_86_port,
                           curr_proc_regs(85) => bus_sel_savedwin_data_85_port,
                           curr_proc_regs(84) => bus_sel_savedwin_data_84_port,
                           curr_proc_regs(83) => bus_sel_savedwin_data_83_port,
                           curr_proc_regs(82) => bus_sel_savedwin_data_82_port,
                           curr_proc_regs(81) => bus_sel_savedwin_data_81_port,
                           curr_proc_regs(80) => bus_sel_savedwin_data_80_port,
                           curr_proc_regs(79) => bus_sel_savedwin_data_79_port,
                           curr_proc_regs(78) => bus_sel_savedwin_data_78_port,
                           curr_proc_regs(77) => bus_sel_savedwin_data_77_port,
                           curr_proc_regs(76) => bus_sel_savedwin_data_76_port,
                           curr_proc_regs(75) => bus_sel_savedwin_data_75_port,
                           curr_proc_regs(74) => bus_sel_savedwin_data_74_port,
                           curr_proc_regs(73) => bus_sel_savedwin_data_73_port,
                           curr_proc_regs(72) => bus_sel_savedwin_data_72_port,
                           curr_proc_regs(71) => bus_sel_savedwin_data_71_port,
                           curr_proc_regs(70) => bus_sel_savedwin_data_70_port,
                           curr_proc_regs(69) => bus_sel_savedwin_data_69_port,
                           curr_proc_regs(68) => bus_sel_savedwin_data_68_port,
                           curr_proc_regs(67) => bus_sel_savedwin_data_67_port,
                           curr_proc_regs(66) => bus_sel_savedwin_data_66_port,
                           curr_proc_regs(65) => bus_sel_savedwin_data_65_port,
                           curr_proc_regs(64) => bus_sel_savedwin_data_64_port,
                           curr_proc_regs(63) => bus_sel_savedwin_data_63_port,
                           curr_proc_regs(62) => bus_sel_savedwin_data_62_port,
                           curr_proc_regs(61) => bus_sel_savedwin_data_61_port,
                           curr_proc_regs(60) => bus_sel_savedwin_data_60_port,
                           curr_proc_regs(59) => bus_sel_savedwin_data_59_port,
                           curr_proc_regs(58) => bus_sel_savedwin_data_58_port,
                           curr_proc_regs(57) => bus_sel_savedwin_data_57_port,
                           curr_proc_regs(56) => bus_sel_savedwin_data_56_port,
                           curr_proc_regs(55) => bus_sel_savedwin_data_55_port,
                           curr_proc_regs(54) => bus_sel_savedwin_data_54_port,
                           curr_proc_regs(53) => bus_sel_savedwin_data_53_port,
                           curr_proc_regs(52) => bus_sel_savedwin_data_52_port,
                           curr_proc_regs(51) => bus_sel_savedwin_data_51_port,
                           curr_proc_regs(50) => bus_sel_savedwin_data_50_port,
                           curr_proc_regs(49) => bus_sel_savedwin_data_49_port,
                           curr_proc_regs(48) => bus_sel_savedwin_data_48_port,
                           curr_proc_regs(47) => bus_sel_savedwin_data_47_port,
                           curr_proc_regs(46) => bus_sel_savedwin_data_46_port,
                           curr_proc_regs(45) => bus_sel_savedwin_data_45_port,
                           curr_proc_regs(44) => bus_sel_savedwin_data_44_port,
                           curr_proc_regs(43) => bus_sel_savedwin_data_43_port,
                           curr_proc_regs(42) => bus_sel_savedwin_data_42_port,
                           curr_proc_regs(41) => bus_sel_savedwin_data_41_port,
                           curr_proc_regs(40) => bus_sel_savedwin_data_40_port,
                           curr_proc_regs(39) => bus_sel_savedwin_data_39_port,
                           curr_proc_regs(38) => bus_sel_savedwin_data_38_port,
                           curr_proc_regs(37) => bus_sel_savedwin_data_37_port,
                           curr_proc_regs(36) => bus_sel_savedwin_data_36_port,
                           curr_proc_regs(35) => bus_sel_savedwin_data_35_port,
                           curr_proc_regs(34) => bus_sel_savedwin_data_34_port,
                           curr_proc_regs(33) => bus_sel_savedwin_data_33_port,
                           curr_proc_regs(32) => bus_sel_savedwin_data_32_port,
                           curr_proc_regs(31) => bus_sel_savedwin_data_31_port,
                           curr_proc_regs(30) => bus_sel_savedwin_data_30_port,
                           curr_proc_regs(29) => bus_sel_savedwin_data_29_port,
                           curr_proc_regs(28) => bus_sel_savedwin_data_28_port,
                           curr_proc_regs(27) => bus_sel_savedwin_data_27_port,
                           curr_proc_regs(26) => bus_sel_savedwin_data_26_port,
                           curr_proc_regs(25) => bus_sel_savedwin_data_25_port,
                           curr_proc_regs(24) => bus_sel_savedwin_data_24_port,
                           curr_proc_regs(23) => bus_sel_savedwin_data_23_port,
                           curr_proc_regs(22) => bus_sel_savedwin_data_22_port,
                           curr_proc_regs(21) => bus_sel_savedwin_data_21_port,
                           curr_proc_regs(20) => bus_sel_savedwin_data_20_port,
                           curr_proc_regs(19) => bus_sel_savedwin_data_19_port,
                           curr_proc_regs(18) => bus_sel_savedwin_data_18_port,
                           curr_proc_regs(17) => bus_sel_savedwin_data_17_port,
                           curr_proc_regs(16) => bus_sel_savedwin_data_16_port,
                           curr_proc_regs(15) => bus_sel_savedwin_data_15_port,
                           curr_proc_regs(14) => bus_sel_savedwin_data_14_port,
                           curr_proc_regs(13) => bus_sel_savedwin_data_13_port,
                           curr_proc_regs(12) => bus_sel_savedwin_data_12_port,
                           curr_proc_regs(11) => bus_sel_savedwin_data_11_port,
                           curr_proc_regs(10) => bus_sel_savedwin_data_10_port,
                           curr_proc_regs(9) => bus_sel_savedwin_data_9_port, 
                           curr_proc_regs(8) => bus_sel_savedwin_data_8_port, 
                           curr_proc_regs(7) => bus_sel_savedwin_data_7_port, 
                           curr_proc_regs(6) => bus_sel_savedwin_data_6_port, 
                           curr_proc_regs(5) => bus_sel_savedwin_data_5_port, 
                           curr_proc_regs(4) => bus_sel_savedwin_data_4_port, 
                           curr_proc_regs(3) => bus_sel_savedwin_data_3_port, 
                           curr_proc_regs(2) => bus_sel_savedwin_data_2_port, 
                           curr_proc_regs(1) => bus_sel_savedwin_data_1_port, 
                           curr_proc_regs(0) => bus_sel_savedwin_data_0_port);
   PUSH_ADDRGEN : address_generator_N16_0 port map( clk => CLK, rst => RESET, 
                           enable => SPILL_port, done => 
                           donespill_donefill_encoding_0_port, working => 
                           working_PUSH, addr(15) => spill_address_ext_15_port,
                           addr(14) => spill_address_ext_14_port, addr(13) => 
                           spill_address_ext_13_port, addr(12) => 
                           spill_address_ext_12_port, addr(11) => 
                           spill_address_ext_11_port, addr(10) => 
                           spill_address_ext_10_port, addr(9) => 
                           spill_address_ext_9_port, addr(8) => 
                           spill_address_ext_8_port, addr(7) => 
                           spill_address_ext_7_port, addr(6) => 
                           spill_address_ext_6_port, addr(5) => 
                           spill_address_ext_5_port, addr(4) => 
                           spill_address_ext_4_port, addr(3) => 
                           spill_address_ext_3_port, addr(2) => 
                           spill_address_ext_2_port, addr(1) => 
                           spill_address_ext_1_port, addr(0) => 
                           spill_address_ext_0_port);
   SPILLADDR_ENC : addr_encoder_N4 port map( Q(15) => spill_address_ext_15_port
                           , Q(14) => spill_address_ext_14_port, Q(13) => 
                           spill_address_ext_13_port, Q(12) => 
                           spill_address_ext_12_port, Q(11) => 
                           spill_address_ext_11_port, Q(10) => 
                           spill_address_ext_10_port, Q(9) => 
                           spill_address_ext_9_port, Q(8) => 
                           spill_address_ext_8_port, Q(7) => 
                           spill_address_ext_7_port, Q(6) => 
                           spill_address_ext_6_port, Q(5) => 
                           spill_address_ext_5_port, Q(4) => 
                           spill_address_ext_4_port, Q(3) => 
                           spill_address_ext_3_port, Q(2) => 
                           spill_address_ext_2_port, Q(1) => 
                           spill_address_ext_1_port, Q(0) => 
                           spill_address_ext_0_port, Y(3) => 
                           spill_address_3_port, Y(2) => spill_address_2_port, 
                           Y(1) => spill_address_1_port, Y(0) => 
                           spill_address_0_port);
   RDPORT_SPILL : mux_N32_M4 port map( S(3) => spill_address_3_port, S(2) => 
                           spill_address_2_port, S(1) => spill_address_1_port, 
                           S(0) => spill_address_0_port, Q(511) => 
                           bus_sel_savedwin_data_511_port, Q(510) => 
                           bus_sel_savedwin_data_510_port, Q(509) => 
                           bus_sel_savedwin_data_509_port, Q(508) => 
                           bus_sel_savedwin_data_508_port, Q(507) => 
                           bus_sel_savedwin_data_507_port, Q(506) => 
                           bus_sel_savedwin_data_506_port, Q(505) => 
                           bus_sel_savedwin_data_505_port, Q(504) => 
                           bus_sel_savedwin_data_504_port, Q(503) => 
                           bus_sel_savedwin_data_503_port, Q(502) => 
                           bus_sel_savedwin_data_502_port, Q(501) => 
                           bus_sel_savedwin_data_501_port, Q(500) => 
                           bus_sel_savedwin_data_500_port, Q(499) => 
                           bus_sel_savedwin_data_499_port, Q(498) => 
                           bus_sel_savedwin_data_498_port, Q(497) => 
                           bus_sel_savedwin_data_497_port, Q(496) => 
                           bus_sel_savedwin_data_496_port, Q(495) => 
                           bus_sel_savedwin_data_495_port, Q(494) => 
                           bus_sel_savedwin_data_494_port, Q(493) => 
                           bus_sel_savedwin_data_493_port, Q(492) => 
                           bus_sel_savedwin_data_492_port, Q(491) => 
                           bus_sel_savedwin_data_491_port, Q(490) => 
                           bus_sel_savedwin_data_490_port, Q(489) => 
                           bus_sel_savedwin_data_489_port, Q(488) => 
                           bus_sel_savedwin_data_488_port, Q(487) => 
                           bus_sel_savedwin_data_487_port, Q(486) => 
                           bus_sel_savedwin_data_486_port, Q(485) => 
                           bus_sel_savedwin_data_485_port, Q(484) => 
                           bus_sel_savedwin_data_484_port, Q(483) => 
                           bus_sel_savedwin_data_483_port, Q(482) => 
                           bus_sel_savedwin_data_482_port, Q(481) => 
                           bus_sel_savedwin_data_481_port, Q(480) => 
                           bus_sel_savedwin_data_480_port, Q(479) => 
                           bus_sel_savedwin_data_479_port, Q(478) => 
                           bus_sel_savedwin_data_478_port, Q(477) => 
                           bus_sel_savedwin_data_477_port, Q(476) => 
                           bus_sel_savedwin_data_476_port, Q(475) => 
                           bus_sel_savedwin_data_475_port, Q(474) => 
                           bus_sel_savedwin_data_474_port, Q(473) => 
                           bus_sel_savedwin_data_473_port, Q(472) => 
                           bus_sel_savedwin_data_472_port, Q(471) => 
                           bus_sel_savedwin_data_471_port, Q(470) => 
                           bus_sel_savedwin_data_470_port, Q(469) => 
                           bus_sel_savedwin_data_469_port, Q(468) => 
                           bus_sel_savedwin_data_468_port, Q(467) => 
                           bus_sel_savedwin_data_467_port, Q(466) => 
                           bus_sel_savedwin_data_466_port, Q(465) => 
                           bus_sel_savedwin_data_465_port, Q(464) => 
                           bus_sel_savedwin_data_464_port, Q(463) => 
                           bus_sel_savedwin_data_463_port, Q(462) => 
                           bus_sel_savedwin_data_462_port, Q(461) => 
                           bus_sel_savedwin_data_461_port, Q(460) => 
                           bus_sel_savedwin_data_460_port, Q(459) => 
                           bus_sel_savedwin_data_459_port, Q(458) => 
                           bus_sel_savedwin_data_458_port, Q(457) => 
                           bus_sel_savedwin_data_457_port, Q(456) => 
                           bus_sel_savedwin_data_456_port, Q(455) => 
                           bus_sel_savedwin_data_455_port, Q(454) => 
                           bus_sel_savedwin_data_454_port, Q(453) => 
                           bus_sel_savedwin_data_453_port, Q(452) => 
                           bus_sel_savedwin_data_452_port, Q(451) => 
                           bus_sel_savedwin_data_451_port, Q(450) => 
                           bus_sel_savedwin_data_450_port, Q(449) => 
                           bus_sel_savedwin_data_449_port, Q(448) => 
                           bus_sel_savedwin_data_448_port, Q(447) => 
                           bus_sel_savedwin_data_447_port, Q(446) => 
                           bus_sel_savedwin_data_446_port, Q(445) => 
                           bus_sel_savedwin_data_445_port, Q(444) => 
                           bus_sel_savedwin_data_444_port, Q(443) => 
                           bus_sel_savedwin_data_443_port, Q(442) => 
                           bus_sel_savedwin_data_442_port, Q(441) => 
                           bus_sel_savedwin_data_441_port, Q(440) => 
                           bus_sel_savedwin_data_440_port, Q(439) => 
                           bus_sel_savedwin_data_439_port, Q(438) => 
                           bus_sel_savedwin_data_438_port, Q(437) => 
                           bus_sel_savedwin_data_437_port, Q(436) => 
                           bus_sel_savedwin_data_436_port, Q(435) => 
                           bus_sel_savedwin_data_435_port, Q(434) => 
                           bus_sel_savedwin_data_434_port, Q(433) => 
                           bus_sel_savedwin_data_433_port, Q(432) => 
                           bus_sel_savedwin_data_432_port, Q(431) => 
                           bus_sel_savedwin_data_431_port, Q(430) => 
                           bus_sel_savedwin_data_430_port, Q(429) => 
                           bus_sel_savedwin_data_429_port, Q(428) => 
                           bus_sel_savedwin_data_428_port, Q(427) => 
                           bus_sel_savedwin_data_427_port, Q(426) => 
                           bus_sel_savedwin_data_426_port, Q(425) => 
                           bus_sel_savedwin_data_425_port, Q(424) => 
                           bus_sel_savedwin_data_424_port, Q(423) => 
                           bus_sel_savedwin_data_423_port, Q(422) => 
                           bus_sel_savedwin_data_422_port, Q(421) => 
                           bus_sel_savedwin_data_421_port, Q(420) => 
                           bus_sel_savedwin_data_420_port, Q(419) => 
                           bus_sel_savedwin_data_419_port, Q(418) => 
                           bus_sel_savedwin_data_418_port, Q(417) => 
                           bus_sel_savedwin_data_417_port, Q(416) => 
                           bus_sel_savedwin_data_416_port, Q(415) => 
                           bus_sel_savedwin_data_415_port, Q(414) => 
                           bus_sel_savedwin_data_414_port, Q(413) => 
                           bus_sel_savedwin_data_413_port, Q(412) => 
                           bus_sel_savedwin_data_412_port, Q(411) => 
                           bus_sel_savedwin_data_411_port, Q(410) => 
                           bus_sel_savedwin_data_410_port, Q(409) => 
                           bus_sel_savedwin_data_409_port, Q(408) => 
                           bus_sel_savedwin_data_408_port, Q(407) => 
                           bus_sel_savedwin_data_407_port, Q(406) => 
                           bus_sel_savedwin_data_406_port, Q(405) => 
                           bus_sel_savedwin_data_405_port, Q(404) => 
                           bus_sel_savedwin_data_404_port, Q(403) => 
                           bus_sel_savedwin_data_403_port, Q(402) => 
                           bus_sel_savedwin_data_402_port, Q(401) => 
                           bus_sel_savedwin_data_401_port, Q(400) => 
                           bus_sel_savedwin_data_400_port, Q(399) => 
                           bus_sel_savedwin_data_399_port, Q(398) => 
                           bus_sel_savedwin_data_398_port, Q(397) => 
                           bus_sel_savedwin_data_397_port, Q(396) => 
                           bus_sel_savedwin_data_396_port, Q(395) => 
                           bus_sel_savedwin_data_395_port, Q(394) => 
                           bus_sel_savedwin_data_394_port, Q(393) => 
                           bus_sel_savedwin_data_393_port, Q(392) => 
                           bus_sel_savedwin_data_392_port, Q(391) => 
                           bus_sel_savedwin_data_391_port, Q(390) => 
                           bus_sel_savedwin_data_390_port, Q(389) => 
                           bus_sel_savedwin_data_389_port, Q(388) => 
                           bus_sel_savedwin_data_388_port, Q(387) => 
                           bus_sel_savedwin_data_387_port, Q(386) => 
                           bus_sel_savedwin_data_386_port, Q(385) => 
                           bus_sel_savedwin_data_385_port, Q(384) => 
                           bus_sel_savedwin_data_384_port, Q(383) => 
                           bus_sel_savedwin_data_383_port, Q(382) => 
                           bus_sel_savedwin_data_382_port, Q(381) => 
                           bus_sel_savedwin_data_381_port, Q(380) => 
                           bus_sel_savedwin_data_380_port, Q(379) => 
                           bus_sel_savedwin_data_379_port, Q(378) => 
                           bus_sel_savedwin_data_378_port, Q(377) => 
                           bus_sel_savedwin_data_377_port, Q(376) => 
                           bus_sel_savedwin_data_376_port, Q(375) => 
                           bus_sel_savedwin_data_375_port, Q(374) => 
                           bus_sel_savedwin_data_374_port, Q(373) => 
                           bus_sel_savedwin_data_373_port, Q(372) => 
                           bus_sel_savedwin_data_372_port, Q(371) => 
                           bus_sel_savedwin_data_371_port, Q(370) => 
                           bus_sel_savedwin_data_370_port, Q(369) => 
                           bus_sel_savedwin_data_369_port, Q(368) => 
                           bus_sel_savedwin_data_368_port, Q(367) => 
                           bus_sel_savedwin_data_367_port, Q(366) => 
                           bus_sel_savedwin_data_366_port, Q(365) => 
                           bus_sel_savedwin_data_365_port, Q(364) => 
                           bus_sel_savedwin_data_364_port, Q(363) => 
                           bus_sel_savedwin_data_363_port, Q(362) => 
                           bus_sel_savedwin_data_362_port, Q(361) => 
                           bus_sel_savedwin_data_361_port, Q(360) => 
                           bus_sel_savedwin_data_360_port, Q(359) => 
                           bus_sel_savedwin_data_359_port, Q(358) => 
                           bus_sel_savedwin_data_358_port, Q(357) => 
                           bus_sel_savedwin_data_357_port, Q(356) => 
                           bus_sel_savedwin_data_356_port, Q(355) => 
                           bus_sel_savedwin_data_355_port, Q(354) => 
                           bus_sel_savedwin_data_354_port, Q(353) => 
                           bus_sel_savedwin_data_353_port, Q(352) => 
                           bus_sel_savedwin_data_352_port, Q(351) => 
                           bus_sel_savedwin_data_351_port, Q(350) => 
                           bus_sel_savedwin_data_350_port, Q(349) => 
                           bus_sel_savedwin_data_349_port, Q(348) => 
                           bus_sel_savedwin_data_348_port, Q(347) => 
                           bus_sel_savedwin_data_347_port, Q(346) => 
                           bus_sel_savedwin_data_346_port, Q(345) => 
                           bus_sel_savedwin_data_345_port, Q(344) => 
                           bus_sel_savedwin_data_344_port, Q(343) => 
                           bus_sel_savedwin_data_343_port, Q(342) => 
                           bus_sel_savedwin_data_342_port, Q(341) => 
                           bus_sel_savedwin_data_341_port, Q(340) => 
                           bus_sel_savedwin_data_340_port, Q(339) => 
                           bus_sel_savedwin_data_339_port, Q(338) => 
                           bus_sel_savedwin_data_338_port, Q(337) => 
                           bus_sel_savedwin_data_337_port, Q(336) => 
                           bus_sel_savedwin_data_336_port, Q(335) => 
                           bus_sel_savedwin_data_335_port, Q(334) => 
                           bus_sel_savedwin_data_334_port, Q(333) => 
                           bus_sel_savedwin_data_333_port, Q(332) => 
                           bus_sel_savedwin_data_332_port, Q(331) => 
                           bus_sel_savedwin_data_331_port, Q(330) => 
                           bus_sel_savedwin_data_330_port, Q(329) => 
                           bus_sel_savedwin_data_329_port, Q(328) => 
                           bus_sel_savedwin_data_328_port, Q(327) => 
                           bus_sel_savedwin_data_327_port, Q(326) => 
                           bus_sel_savedwin_data_326_port, Q(325) => 
                           bus_sel_savedwin_data_325_port, Q(324) => 
                           bus_sel_savedwin_data_324_port, Q(323) => 
                           bus_sel_savedwin_data_323_port, Q(322) => 
                           bus_sel_savedwin_data_322_port, Q(321) => 
                           bus_sel_savedwin_data_321_port, Q(320) => 
                           bus_sel_savedwin_data_320_port, Q(319) => 
                           bus_sel_savedwin_data_319_port, Q(318) => 
                           bus_sel_savedwin_data_318_port, Q(317) => 
                           bus_sel_savedwin_data_317_port, Q(316) => 
                           bus_sel_savedwin_data_316_port, Q(315) => 
                           bus_sel_savedwin_data_315_port, Q(314) => 
                           bus_sel_savedwin_data_314_port, Q(313) => 
                           bus_sel_savedwin_data_313_port, Q(312) => 
                           bus_sel_savedwin_data_312_port, Q(311) => 
                           bus_sel_savedwin_data_311_port, Q(310) => 
                           bus_sel_savedwin_data_310_port, Q(309) => 
                           bus_sel_savedwin_data_309_port, Q(308) => 
                           bus_sel_savedwin_data_308_port, Q(307) => 
                           bus_sel_savedwin_data_307_port, Q(306) => 
                           bus_sel_savedwin_data_306_port, Q(305) => 
                           bus_sel_savedwin_data_305_port, Q(304) => 
                           bus_sel_savedwin_data_304_port, Q(303) => 
                           bus_sel_savedwin_data_303_port, Q(302) => 
                           bus_sel_savedwin_data_302_port, Q(301) => 
                           bus_sel_savedwin_data_301_port, Q(300) => 
                           bus_sel_savedwin_data_300_port, Q(299) => 
                           bus_sel_savedwin_data_299_port, Q(298) => 
                           bus_sel_savedwin_data_298_port, Q(297) => 
                           bus_sel_savedwin_data_297_port, Q(296) => 
                           bus_sel_savedwin_data_296_port, Q(295) => 
                           bus_sel_savedwin_data_295_port, Q(294) => 
                           bus_sel_savedwin_data_294_port, Q(293) => 
                           bus_sel_savedwin_data_293_port, Q(292) => 
                           bus_sel_savedwin_data_292_port, Q(291) => 
                           bus_sel_savedwin_data_291_port, Q(290) => 
                           bus_sel_savedwin_data_290_port, Q(289) => 
                           bus_sel_savedwin_data_289_port, Q(288) => 
                           bus_sel_savedwin_data_288_port, Q(287) => 
                           bus_sel_savedwin_data_287_port, Q(286) => 
                           bus_sel_savedwin_data_286_port, Q(285) => 
                           bus_sel_savedwin_data_285_port, Q(284) => 
                           bus_sel_savedwin_data_284_port, Q(283) => 
                           bus_sel_savedwin_data_283_port, Q(282) => 
                           bus_sel_savedwin_data_282_port, Q(281) => 
                           bus_sel_savedwin_data_281_port, Q(280) => 
                           bus_sel_savedwin_data_280_port, Q(279) => 
                           bus_sel_savedwin_data_279_port, Q(278) => 
                           bus_sel_savedwin_data_278_port, Q(277) => 
                           bus_sel_savedwin_data_277_port, Q(276) => 
                           bus_sel_savedwin_data_276_port, Q(275) => 
                           bus_sel_savedwin_data_275_port, Q(274) => 
                           bus_sel_savedwin_data_274_port, Q(273) => 
                           bus_sel_savedwin_data_273_port, Q(272) => 
                           bus_sel_savedwin_data_272_port, Q(271) => 
                           bus_sel_savedwin_data_271_port, Q(270) => 
                           bus_sel_savedwin_data_270_port, Q(269) => 
                           bus_sel_savedwin_data_269_port, Q(268) => 
                           bus_sel_savedwin_data_268_port, Q(267) => 
                           bus_sel_savedwin_data_267_port, Q(266) => 
                           bus_sel_savedwin_data_266_port, Q(265) => 
                           bus_sel_savedwin_data_265_port, Q(264) => 
                           bus_sel_savedwin_data_264_port, Q(263) => 
                           bus_sel_savedwin_data_263_port, Q(262) => 
                           bus_sel_savedwin_data_262_port, Q(261) => 
                           bus_sel_savedwin_data_261_port, Q(260) => 
                           bus_sel_savedwin_data_260_port, Q(259) => 
                           bus_sel_savedwin_data_259_port, Q(258) => 
                           bus_sel_savedwin_data_258_port, Q(257) => 
                           bus_sel_savedwin_data_257_port, Q(256) => 
                           bus_sel_savedwin_data_256_port, Q(255) => 
                           bus_sel_savedwin_data_255_port, Q(254) => 
                           bus_sel_savedwin_data_254_port, Q(253) => 
                           bus_sel_savedwin_data_253_port, Q(252) => 
                           bus_sel_savedwin_data_252_port, Q(251) => 
                           bus_sel_savedwin_data_251_port, Q(250) => 
                           bus_sel_savedwin_data_250_port, Q(249) => 
                           bus_sel_savedwin_data_249_port, Q(248) => 
                           bus_sel_savedwin_data_248_port, Q(247) => 
                           bus_sel_savedwin_data_247_port, Q(246) => 
                           bus_sel_savedwin_data_246_port, Q(245) => 
                           bus_sel_savedwin_data_245_port, Q(244) => 
                           bus_sel_savedwin_data_244_port, Q(243) => 
                           bus_sel_savedwin_data_243_port, Q(242) => 
                           bus_sel_savedwin_data_242_port, Q(241) => 
                           bus_sel_savedwin_data_241_port, Q(240) => 
                           bus_sel_savedwin_data_240_port, Q(239) => 
                           bus_sel_savedwin_data_239_port, Q(238) => 
                           bus_sel_savedwin_data_238_port, Q(237) => 
                           bus_sel_savedwin_data_237_port, Q(236) => 
                           bus_sel_savedwin_data_236_port, Q(235) => 
                           bus_sel_savedwin_data_235_port, Q(234) => 
                           bus_sel_savedwin_data_234_port, Q(233) => 
                           bus_sel_savedwin_data_233_port, Q(232) => 
                           bus_sel_savedwin_data_232_port, Q(231) => 
                           bus_sel_savedwin_data_231_port, Q(230) => 
                           bus_sel_savedwin_data_230_port, Q(229) => 
                           bus_sel_savedwin_data_229_port, Q(228) => 
                           bus_sel_savedwin_data_228_port, Q(227) => 
                           bus_sel_savedwin_data_227_port, Q(226) => 
                           bus_sel_savedwin_data_226_port, Q(225) => 
                           bus_sel_savedwin_data_225_port, Q(224) => 
                           bus_sel_savedwin_data_224_port, Q(223) => 
                           bus_sel_savedwin_data_223_port, Q(222) => 
                           bus_sel_savedwin_data_222_port, Q(221) => 
                           bus_sel_savedwin_data_221_port, Q(220) => 
                           bus_sel_savedwin_data_220_port, Q(219) => 
                           bus_sel_savedwin_data_219_port, Q(218) => 
                           bus_sel_savedwin_data_218_port, Q(217) => 
                           bus_sel_savedwin_data_217_port, Q(216) => 
                           bus_sel_savedwin_data_216_port, Q(215) => 
                           bus_sel_savedwin_data_215_port, Q(214) => 
                           bus_sel_savedwin_data_214_port, Q(213) => 
                           bus_sel_savedwin_data_213_port, Q(212) => 
                           bus_sel_savedwin_data_212_port, Q(211) => 
                           bus_sel_savedwin_data_211_port, Q(210) => 
                           bus_sel_savedwin_data_210_port, Q(209) => 
                           bus_sel_savedwin_data_209_port, Q(208) => 
                           bus_sel_savedwin_data_208_port, Q(207) => 
                           bus_sel_savedwin_data_207_port, Q(206) => 
                           bus_sel_savedwin_data_206_port, Q(205) => 
                           bus_sel_savedwin_data_205_port, Q(204) => 
                           bus_sel_savedwin_data_204_port, Q(203) => 
                           bus_sel_savedwin_data_203_port, Q(202) => 
                           bus_sel_savedwin_data_202_port, Q(201) => 
                           bus_sel_savedwin_data_201_port, Q(200) => 
                           bus_sel_savedwin_data_200_port, Q(199) => 
                           bus_sel_savedwin_data_199_port, Q(198) => 
                           bus_sel_savedwin_data_198_port, Q(197) => 
                           bus_sel_savedwin_data_197_port, Q(196) => 
                           bus_sel_savedwin_data_196_port, Q(195) => 
                           bus_sel_savedwin_data_195_port, Q(194) => 
                           bus_sel_savedwin_data_194_port, Q(193) => 
                           bus_sel_savedwin_data_193_port, Q(192) => 
                           bus_sel_savedwin_data_192_port, Q(191) => 
                           bus_sel_savedwin_data_191_port, Q(190) => 
                           bus_sel_savedwin_data_190_port, Q(189) => 
                           bus_sel_savedwin_data_189_port, Q(188) => 
                           bus_sel_savedwin_data_188_port, Q(187) => 
                           bus_sel_savedwin_data_187_port, Q(186) => 
                           bus_sel_savedwin_data_186_port, Q(185) => 
                           bus_sel_savedwin_data_185_port, Q(184) => 
                           bus_sel_savedwin_data_184_port, Q(183) => 
                           bus_sel_savedwin_data_183_port, Q(182) => 
                           bus_sel_savedwin_data_182_port, Q(181) => 
                           bus_sel_savedwin_data_181_port, Q(180) => 
                           bus_sel_savedwin_data_180_port, Q(179) => 
                           bus_sel_savedwin_data_179_port, Q(178) => 
                           bus_sel_savedwin_data_178_port, Q(177) => 
                           bus_sel_savedwin_data_177_port, Q(176) => 
                           bus_sel_savedwin_data_176_port, Q(175) => 
                           bus_sel_savedwin_data_175_port, Q(174) => 
                           bus_sel_savedwin_data_174_port, Q(173) => 
                           bus_sel_savedwin_data_173_port, Q(172) => 
                           bus_sel_savedwin_data_172_port, Q(171) => 
                           bus_sel_savedwin_data_171_port, Q(170) => 
                           bus_sel_savedwin_data_170_port, Q(169) => 
                           bus_sel_savedwin_data_169_port, Q(168) => 
                           bus_sel_savedwin_data_168_port, Q(167) => 
                           bus_sel_savedwin_data_167_port, Q(166) => 
                           bus_sel_savedwin_data_166_port, Q(165) => 
                           bus_sel_savedwin_data_165_port, Q(164) => 
                           bus_sel_savedwin_data_164_port, Q(163) => 
                           bus_sel_savedwin_data_163_port, Q(162) => 
                           bus_sel_savedwin_data_162_port, Q(161) => 
                           bus_sel_savedwin_data_161_port, Q(160) => 
                           bus_sel_savedwin_data_160_port, Q(159) => 
                           bus_sel_savedwin_data_159_port, Q(158) => 
                           bus_sel_savedwin_data_158_port, Q(157) => 
                           bus_sel_savedwin_data_157_port, Q(156) => 
                           bus_sel_savedwin_data_156_port, Q(155) => 
                           bus_sel_savedwin_data_155_port, Q(154) => 
                           bus_sel_savedwin_data_154_port, Q(153) => 
                           bus_sel_savedwin_data_153_port, Q(152) => 
                           bus_sel_savedwin_data_152_port, Q(151) => 
                           bus_sel_savedwin_data_151_port, Q(150) => 
                           bus_sel_savedwin_data_150_port, Q(149) => 
                           bus_sel_savedwin_data_149_port, Q(148) => 
                           bus_sel_savedwin_data_148_port, Q(147) => 
                           bus_sel_savedwin_data_147_port, Q(146) => 
                           bus_sel_savedwin_data_146_port, Q(145) => 
                           bus_sel_savedwin_data_145_port, Q(144) => 
                           bus_sel_savedwin_data_144_port, Q(143) => 
                           bus_sel_savedwin_data_143_port, Q(142) => 
                           bus_sel_savedwin_data_142_port, Q(141) => 
                           bus_sel_savedwin_data_141_port, Q(140) => 
                           bus_sel_savedwin_data_140_port, Q(139) => 
                           bus_sel_savedwin_data_139_port, Q(138) => 
                           bus_sel_savedwin_data_138_port, Q(137) => 
                           bus_sel_savedwin_data_137_port, Q(136) => 
                           bus_sel_savedwin_data_136_port, Q(135) => 
                           bus_sel_savedwin_data_135_port, Q(134) => 
                           bus_sel_savedwin_data_134_port, Q(133) => 
                           bus_sel_savedwin_data_133_port, Q(132) => 
                           bus_sel_savedwin_data_132_port, Q(131) => 
                           bus_sel_savedwin_data_131_port, Q(130) => 
                           bus_sel_savedwin_data_130_port, Q(129) => 
                           bus_sel_savedwin_data_129_port, Q(128) => 
                           bus_sel_savedwin_data_128_port, Q(127) => 
                           bus_sel_savedwin_data_127_port, Q(126) => 
                           bus_sel_savedwin_data_126_port, Q(125) => 
                           bus_sel_savedwin_data_125_port, Q(124) => 
                           bus_sel_savedwin_data_124_port, Q(123) => 
                           bus_sel_savedwin_data_123_port, Q(122) => 
                           bus_sel_savedwin_data_122_port, Q(121) => 
                           bus_sel_savedwin_data_121_port, Q(120) => 
                           bus_sel_savedwin_data_120_port, Q(119) => 
                           bus_sel_savedwin_data_119_port, Q(118) => 
                           bus_sel_savedwin_data_118_port, Q(117) => 
                           bus_sel_savedwin_data_117_port, Q(116) => 
                           bus_sel_savedwin_data_116_port, Q(115) => 
                           bus_sel_savedwin_data_115_port, Q(114) => 
                           bus_sel_savedwin_data_114_port, Q(113) => 
                           bus_sel_savedwin_data_113_port, Q(112) => 
                           bus_sel_savedwin_data_112_port, Q(111) => 
                           bus_sel_savedwin_data_111_port, Q(110) => 
                           bus_sel_savedwin_data_110_port, Q(109) => 
                           bus_sel_savedwin_data_109_port, Q(108) => 
                           bus_sel_savedwin_data_108_port, Q(107) => 
                           bus_sel_savedwin_data_107_port, Q(106) => 
                           bus_sel_savedwin_data_106_port, Q(105) => 
                           bus_sel_savedwin_data_105_port, Q(104) => 
                           bus_sel_savedwin_data_104_port, Q(103) => 
                           bus_sel_savedwin_data_103_port, Q(102) => 
                           bus_sel_savedwin_data_102_port, Q(101) => 
                           bus_sel_savedwin_data_101_port, Q(100) => 
                           bus_sel_savedwin_data_100_port, Q(99) => 
                           bus_sel_savedwin_data_99_port, Q(98) => 
                           bus_sel_savedwin_data_98_port, Q(97) => 
                           bus_sel_savedwin_data_97_port, Q(96) => 
                           bus_sel_savedwin_data_96_port, Q(95) => 
                           bus_sel_savedwin_data_95_port, Q(94) => 
                           bus_sel_savedwin_data_94_port, Q(93) => 
                           bus_sel_savedwin_data_93_port, Q(92) => 
                           bus_sel_savedwin_data_92_port, Q(91) => 
                           bus_sel_savedwin_data_91_port, Q(90) => 
                           bus_sel_savedwin_data_90_port, Q(89) => 
                           bus_sel_savedwin_data_89_port, Q(88) => 
                           bus_sel_savedwin_data_88_port, Q(87) => 
                           bus_sel_savedwin_data_87_port, Q(86) => 
                           bus_sel_savedwin_data_86_port, Q(85) => 
                           bus_sel_savedwin_data_85_port, Q(84) => 
                           bus_sel_savedwin_data_84_port, Q(83) => 
                           bus_sel_savedwin_data_83_port, Q(82) => 
                           bus_sel_savedwin_data_82_port, Q(81) => 
                           bus_sel_savedwin_data_81_port, Q(80) => 
                           bus_sel_savedwin_data_80_port, Q(79) => 
                           bus_sel_savedwin_data_79_port, Q(78) => 
                           bus_sel_savedwin_data_78_port, Q(77) => 
                           bus_sel_savedwin_data_77_port, Q(76) => 
                           bus_sel_savedwin_data_76_port, Q(75) => 
                           bus_sel_savedwin_data_75_port, Q(74) => 
                           bus_sel_savedwin_data_74_port, Q(73) => 
                           bus_sel_savedwin_data_73_port, Q(72) => 
                           bus_sel_savedwin_data_72_port, Q(71) => 
                           bus_sel_savedwin_data_71_port, Q(70) => 
                           bus_sel_savedwin_data_70_port, Q(69) => 
                           bus_sel_savedwin_data_69_port, Q(68) => 
                           bus_sel_savedwin_data_68_port, Q(67) => 
                           bus_sel_savedwin_data_67_port, Q(66) => 
                           bus_sel_savedwin_data_66_port, Q(65) => 
                           bus_sel_savedwin_data_65_port, Q(64) => 
                           bus_sel_savedwin_data_64_port, Q(63) => 
                           bus_sel_savedwin_data_63_port, Q(62) => 
                           bus_sel_savedwin_data_62_port, Q(61) => 
                           bus_sel_savedwin_data_61_port, Q(60) => 
                           bus_sel_savedwin_data_60_port, Q(59) => 
                           bus_sel_savedwin_data_59_port, Q(58) => 
                           bus_sel_savedwin_data_58_port, Q(57) => 
                           bus_sel_savedwin_data_57_port, Q(56) => 
                           bus_sel_savedwin_data_56_port, Q(55) => 
                           bus_sel_savedwin_data_55_port, Q(54) => 
                           bus_sel_savedwin_data_54_port, Q(53) => 
                           bus_sel_savedwin_data_53_port, Q(52) => 
                           bus_sel_savedwin_data_52_port, Q(51) => 
                           bus_sel_savedwin_data_51_port, Q(50) => 
                           bus_sel_savedwin_data_50_port, Q(49) => 
                           bus_sel_savedwin_data_49_port, Q(48) => 
                           bus_sel_savedwin_data_48_port, Q(47) => 
                           bus_sel_savedwin_data_47_port, Q(46) => 
                           bus_sel_savedwin_data_46_port, Q(45) => 
                           bus_sel_savedwin_data_45_port, Q(44) => 
                           bus_sel_savedwin_data_44_port, Q(43) => 
                           bus_sel_savedwin_data_43_port, Q(42) => 
                           bus_sel_savedwin_data_42_port, Q(41) => 
                           bus_sel_savedwin_data_41_port, Q(40) => 
                           bus_sel_savedwin_data_40_port, Q(39) => 
                           bus_sel_savedwin_data_39_port, Q(38) => 
                           bus_sel_savedwin_data_38_port, Q(37) => 
                           bus_sel_savedwin_data_37_port, Q(36) => 
                           bus_sel_savedwin_data_36_port, Q(35) => 
                           bus_sel_savedwin_data_35_port, Q(34) => 
                           bus_sel_savedwin_data_34_port, Q(33) => 
                           bus_sel_savedwin_data_33_port, Q(32) => 
                           bus_sel_savedwin_data_32_port, Q(31) => 
                           bus_sel_savedwin_data_31_port, Q(30) => 
                           bus_sel_savedwin_data_30_port, Q(29) => 
                           bus_sel_savedwin_data_29_port, Q(28) => 
                           bus_sel_savedwin_data_28_port, Q(27) => 
                           bus_sel_savedwin_data_27_port, Q(26) => 
                           bus_sel_savedwin_data_26_port, Q(25) => 
                           bus_sel_savedwin_data_25_port, Q(24) => 
                           bus_sel_savedwin_data_24_port, Q(23) => 
                           bus_sel_savedwin_data_23_port, Q(22) => 
                           bus_sel_savedwin_data_22_port, Q(21) => 
                           bus_sel_savedwin_data_21_port, Q(20) => 
                           bus_sel_savedwin_data_20_port, Q(19) => 
                           bus_sel_savedwin_data_19_port, Q(18) => 
                           bus_sel_savedwin_data_18_port, Q(17) => 
                           bus_sel_savedwin_data_17_port, Q(16) => 
                           bus_sel_savedwin_data_16_port, Q(15) => 
                           bus_sel_savedwin_data_15_port, Q(14) => 
                           bus_sel_savedwin_data_14_port, Q(13) => 
                           bus_sel_savedwin_data_13_port, Q(12) => 
                           bus_sel_savedwin_data_12_port, Q(11) => 
                           bus_sel_savedwin_data_11_port, Q(10) => 
                           bus_sel_savedwin_data_10_port, Q(9) => 
                           bus_sel_savedwin_data_9_port, Q(8) => 
                           bus_sel_savedwin_data_8_port, Q(7) => 
                           bus_sel_savedwin_data_7_port, Q(6) => 
                           bus_sel_savedwin_data_6_port, Q(5) => 
                           bus_sel_savedwin_data_5_port, Q(4) => 
                           bus_sel_savedwin_data_4_port, Q(3) => 
                           bus_sel_savedwin_data_3_port, Q(2) => 
                           bus_sel_savedwin_data_2_port, Q(1) => 
                           bus_sel_savedwin_data_1_port, Q(0) => 
                           bus_sel_savedwin_data_0_port, Y(31) => BUS_TOMEM(31)
                           , Y(30) => BUS_TOMEM(30), Y(29) => BUS_TOMEM(29), 
                           Y(28) => BUS_TOMEM(28), Y(27) => BUS_TOMEM(27), 
                           Y(26) => BUS_TOMEM(26), Y(25) => BUS_TOMEM(25), 
                           Y(24) => BUS_TOMEM(24), Y(23) => BUS_TOMEM(23), 
                           Y(22) => BUS_TOMEM(22), Y(21) => BUS_TOMEM(21), 
                           Y(20) => BUS_TOMEM(20), Y(19) => BUS_TOMEM(19), 
                           Y(18) => BUS_TOMEM(18), Y(17) => BUS_TOMEM(17), 
                           Y(16) => BUS_TOMEM(16), Y(15) => BUS_TOMEM(15), 
                           Y(14) => BUS_TOMEM(14), Y(13) => BUS_TOMEM(13), 
                           Y(12) => BUS_TOMEM(12), Y(11) => BUS_TOMEM(11), 
                           Y(10) => BUS_TOMEM(10), Y(9) => BUS_TOMEM(9), Y(8) 
                           => BUS_TOMEM(8), Y(7) => BUS_TOMEM(7), Y(6) => 
                           BUS_TOMEM(6), Y(5) => BUS_TOMEM(5), Y(4) => 
                           BUS_TOMEM(4), Y(3) => BUS_TOMEM(3), Y(2) => 
                           BUS_TOMEM(2), Y(1) => BUS_TOMEM(1), Y(0) => 
                           BUS_TOMEM(0));
   EQ_CHECK_POP : equal_check_N5_1 port map( A(4) => c_win_4_port, A(3) => 
                           c_win_3_port, A(2) => c_win_2_port, A(1) => 
                           c_win_1_port, A(0) => c_win_0_port, B(4) => 
                           c_swin_4_port, B(3) => c_swin_3_port, B(2) => 
                           c_swin_2_port, B(1) => c_swin_1_port, B(0) => 
                           c_swin_0_port, EQUAL => filleq);
   POP_ADDRGEN : address_generator_N16_1 port map( clk => CLK, rst => RESET, 
                           enable => FILL_port, done => 
                           donespill_donefill_encoding_1_port, working => 
                           working_POP, addr(15) => fill_address_ext_15_port, 
                           addr(14) => fill_address_ext_14_port, addr(13) => 
                           fill_address_ext_13_port, addr(12) => 
                           fill_address_ext_12_port, addr(11) => 
                           fill_address_ext_11_port, addr(10) => 
                           fill_address_ext_10_port, addr(9) => 
                           fill_address_ext_9_port, addr(8) => 
                           fill_address_ext_8_port, addr(7) => 
                           fill_address_ext_7_port, addr(6) => 
                           fill_address_ext_6_port, addr(5) => 
                           fill_address_ext_5_port, addr(4) => 
                           fill_address_ext_4_port, addr(3) => 
                           fill_address_ext_3_port, addr(2) => 
                           fill_address_ext_2_port, addr(1) => 
                           fill_address_ext_1_port, addr(0) => 
                           fill_address_ext_0_port);
   U52 : NOR2_X2 port map( A1 => n37, A2 => n38, ZN => 
                           internal_inloc_data_4_29_port);
   U53 : NOR2_X2 port map( A1 => n41, A2 => n42, ZN => 
                           internal_inloc_data_4_27_port);
   U54 : NOR2_X2 port map( A1 => n43, A2 => n44, ZN => 
                           internal_inloc_data_4_26_port);
   U55 : NOR2_X2 port map( A1 => n45, A2 => n46, ZN => 
                           internal_inloc_data_4_25_port);
   U56 : NOR2_X2 port map( A1 => n95, A2 => n96, ZN => 
                           internal_inloc_data_3_31_port);
   U57 : NOR2_X2 port map( A1 => n97, A2 => n98, ZN => 
                           internal_inloc_data_3_30_port);
   U58 : NOR2_X2 port map( A1 => n101, A2 => n102, ZN => 
                           internal_inloc_data_3_29_port);
   U59 : NOR2_X2 port map( A1 => n105, A2 => n106, ZN => 
                           internal_inloc_data_3_27_port);
   U60 : NOR2_X2 port map( A1 => n107, A2 => n108, ZN => 
                           internal_inloc_data_3_26_port);
   U61 : NOR2_X2 port map( A1 => n109, A2 => n110, ZN => 
                           internal_inloc_data_3_25_port);
   U62 : NOR2_X2 port map( A1 => n159, A2 => n160, ZN => 
                           internal_inloc_data_2_31_port);
   U63 : NOR2_X2 port map( A1 => n161, A2 => n162, ZN => 
                           internal_inloc_data_2_30_port);
   U64 : NOR2_X2 port map( A1 => n165, A2 => n166, ZN => 
                           internal_inloc_data_2_29_port);
   U65 : NOR2_X2 port map( A1 => n169, A2 => n170, ZN => 
                           internal_inloc_data_2_27_port);
   U66 : NOR2_X2 port map( A1 => n171, A2 => n172, ZN => 
                           internal_inloc_data_2_26_port);
   U67 : NOR2_X2 port map( A1 => n173, A2 => n174, ZN => 
                           internal_inloc_data_2_25_port);
   U68 : NOR2_X2 port map( A1 => n223, A2 => n224, ZN => 
                           internal_inloc_data_1_31_port);
   U69 : NOR2_X2 port map( A1 => n225, A2 => n226, ZN => 
                           internal_inloc_data_1_30_port);
   U70 : NOR2_X2 port map( A1 => n229, A2 => n230, ZN => 
                           internal_inloc_data_1_29_port);
   U71 : NOR2_X2 port map( A1 => n233, A2 => n234, ZN => 
                           internal_inloc_data_1_27_port);
   U72 : NOR2_X2 port map( A1 => n235, A2 => n236, ZN => 
                           internal_inloc_data_1_26_port);
   U73 : NOR2_X2 port map( A1 => n237, A2 => n238, ZN => 
                           internal_inloc_data_1_25_port);
   U74 : NOR2_X2 port map( A1 => n287, A2 => n288, ZN => 
                           internal_inloc_data_0_31_port);
   U75 : NOR2_X2 port map( A1 => n289, A2 => n290, ZN => 
                           internal_inloc_data_0_30_port);
   U76 : NOR2_X2 port map( A1 => n293, A2 => n294, ZN => 
                           internal_inloc_data_0_29_port);
   U77 : NOR2_X2 port map( A1 => n297, A2 => n298, ZN => 
                           internal_inloc_data_0_27_port);
   U78 : NOR2_X2 port map( A1 => n299, A2 => n300, ZN => 
                           internal_inloc_data_0_26_port);
   U79 : NOR2_X2 port map( A1 => n301, A2 => n302, ZN => 
                           internal_inloc_data_0_25_port);
   U80 : NOR2_X2 port map( A1 => n31, A2 => n32, ZN => 
                           internal_inloc_data_4_31_port);
   U81 : NOR2_X2 port map( A1 => n33, A2 => n34, ZN => 
                           internal_inloc_data_4_30_port);
   U82 : NOR2_X2 port map( A1 => n39, A2 => n40, ZN => 
                           internal_inloc_data_4_28_port);
   U83 : NOR2_X2 port map( A1 => n47, A2 => n48, ZN => 
                           internal_inloc_data_4_24_port);
   U84 : NOR2_X2 port map( A1 => n103, A2 => n104, ZN => 
                           internal_inloc_data_3_28_port);
   U85 : NOR2_X2 port map( A1 => n111, A2 => n112, ZN => 
                           internal_inloc_data_3_24_port);
   U86 : NOR2_X2 port map( A1 => n167, A2 => n168, ZN => 
                           internal_inloc_data_2_28_port);
   U87 : NOR2_X2 port map( A1 => n175, A2 => n176, ZN => 
                           internal_inloc_data_2_24_port);
   U88 : NOR2_X2 port map( A1 => n231, A2 => n232, ZN => 
                           internal_inloc_data_1_28_port);
   U89 : NOR2_X2 port map( A1 => n239, A2 => n240, ZN => 
                           internal_inloc_data_1_24_port);
   U90 : NOR2_X2 port map( A1 => n295, A2 => n296, ZN => 
                           internal_inloc_data_0_28_port);
   U91 : NOR2_X2 port map( A1 => n303, A2 => n304, ZN => 
                           internal_inloc_data_0_24_port);
   U92 : NOR2_X2 port map( A1 => n49, A2 => n50, ZN => 
                           internal_inloc_data_4_23_port);
   U93 : NOR2_X2 port map( A1 => n65, A2 => n66, ZN => 
                           internal_inloc_data_4_16_port);
   U94 : NOR2_X2 port map( A1 => n17, A2 => n18, ZN => 
                           internal_inloc_data_4_9_port);
   U95 : NOR2_X2 port map( A1 => n113, A2 => n114, ZN => 
                           internal_inloc_data_3_23_port);
   U96 : NOR2_X2 port map( A1 => n129, A2 => n130, ZN => 
                           internal_inloc_data_3_16_port);
   U97 : NOR2_X2 port map( A1 => n81, A2 => n82, ZN => 
                           internal_inloc_data_3_9_port);
   U98 : NOR2_X2 port map( A1 => n177, A2 => n178, ZN => 
                           internal_inloc_data_2_23_port);
   U99 : NOR2_X2 port map( A1 => n193, A2 => n194, ZN => 
                           internal_inloc_data_2_16_port);
   U100 : NOR2_X2 port map( A1 => n145, A2 => n146, ZN => 
                           internal_inloc_data_2_9_port);
   U101 : NOR2_X2 port map( A1 => n241, A2 => n242, ZN => 
                           internal_inloc_data_1_23_port);
   U102 : NOR2_X2 port map( A1 => n257, A2 => n258, ZN => 
                           internal_inloc_data_1_16_port);
   U103 : NOR2_X2 port map( A1 => n209, A2 => n210, ZN => 
                           internal_inloc_data_1_9_port);
   U104 : NOR2_X2 port map( A1 => n305, A2 => n306, ZN => 
                           internal_inloc_data_0_23_port);
   U105 : NOR2_X2 port map( A1 => n321, A2 => n322, ZN => 
                           internal_inloc_data_0_16_port);
   U106 : NOR2_X2 port map( A1 => n273, A2 => n274, ZN => 
                           internal_inloc_data_0_9_port);
   U107 : NOR2_X2 port map( A1 => n51, A2 => n52, ZN => 
                           internal_inloc_data_4_22_port);
   U108 : NOR2_X2 port map( A1 => n67, A2 => n68, ZN => 
                           internal_inloc_data_4_15_port);
   U109 : NOR2_X2 port map( A1 => n19, A2 => n20, ZN => 
                           internal_inloc_data_4_8_port);
   U110 : NOR2_X2 port map( A1 => n115, A2 => n116, ZN => 
                           internal_inloc_data_3_22_port);
   U111 : NOR2_X2 port map( A1 => n131, A2 => n132, ZN => 
                           internal_inloc_data_3_15_port);
   U112 : NOR2_X2 port map( A1 => n83, A2 => n84, ZN => 
                           internal_inloc_data_3_8_port);
   U113 : NOR2_X2 port map( A1 => n179, A2 => n180, ZN => 
                           internal_inloc_data_2_22_port);
   U114 : NOR2_X2 port map( A1 => n195, A2 => n196, ZN => 
                           internal_inloc_data_2_15_port);
   U115 : NOR2_X2 port map( A1 => n147, A2 => n148, ZN => 
                           internal_inloc_data_2_8_port);
   U116 : NOR2_X2 port map( A1 => n243, A2 => n244, ZN => 
                           internal_inloc_data_1_22_port);
   U117 : NOR2_X2 port map( A1 => n259, A2 => n260, ZN => 
                           internal_inloc_data_1_15_port);
   U118 : NOR2_X2 port map( A1 => n211, A2 => n212, ZN => 
                           internal_inloc_data_1_8_port);
   U119 : NOR2_X2 port map( A1 => n307, A2 => n308, ZN => 
                           internal_inloc_data_0_22_port);
   U120 : NOR2_X2 port map( A1 => n323, A2 => n324, ZN => 
                           internal_inloc_data_0_15_port);
   U121 : NOR2_X2 port map( A1 => n275, A2 => n276, ZN => 
                           internal_inloc_data_0_8_port);
   U122 : NOR2_X2 port map( A1 => n53, A2 => n54, ZN => 
                           internal_inloc_data_4_21_port);
   U123 : NOR2_X2 port map( A1 => n69, A2 => n70, ZN => 
                           internal_inloc_data_4_14_port);
   U124 : NOR2_X2 port map( A1 => n21, A2 => n22, ZN => 
                           internal_inloc_data_4_7_port);
   U125 : NOR2_X2 port map( A1 => n117, A2 => n118, ZN => 
                           internal_inloc_data_3_21_port);
   U126 : NOR2_X2 port map( A1 => n133, A2 => n134, ZN => 
                           internal_inloc_data_3_14_port);
   U127 : NOR2_X2 port map( A1 => n85, A2 => n86, ZN => 
                           internal_inloc_data_3_7_port);
   U128 : NOR2_X2 port map( A1 => n181, A2 => n182, ZN => 
                           internal_inloc_data_2_21_port);
   U129 : NOR2_X2 port map( A1 => n197, A2 => n198, ZN => 
                           internal_inloc_data_2_14_port);
   U130 : NOR2_X2 port map( A1 => n149, A2 => n150, ZN => 
                           internal_inloc_data_2_7_port);
   U131 : NOR2_X2 port map( A1 => n245, A2 => n246, ZN => 
                           internal_inloc_data_1_21_port);
   U132 : NOR2_X2 port map( A1 => n261, A2 => n262, ZN => 
                           internal_inloc_data_1_14_port);
   U133 : NOR2_X2 port map( A1 => n213, A2 => n214, ZN => 
                           internal_inloc_data_1_7_port);
   U134 : NOR2_X2 port map( A1 => n309, A2 => n310, ZN => 
                           internal_inloc_data_0_21_port);
   U135 : NOR2_X2 port map( A1 => n325, A2 => n326, ZN => 
                           internal_inloc_data_0_14_port);
   U136 : NOR2_X2 port map( A1 => n277, A2 => n278, ZN => 
                           internal_inloc_data_0_7_port);
   U137 : NOR2_X2 port map( A1 => n55, A2 => n56, ZN => 
                           internal_inloc_data_4_20_port);
   U138 : NOR2_X2 port map( A1 => n71, A2 => n72, ZN => 
                           internal_inloc_data_4_13_port);
   U139 : NOR2_X2 port map( A1 => n23, A2 => n24, ZN => 
                           internal_inloc_data_4_6_port);
   U140 : NOR2_X2 port map( A1 => n119, A2 => n120, ZN => 
                           internal_inloc_data_3_20_port);
   U141 : NOR2_X2 port map( A1 => n135, A2 => n136, ZN => 
                           internal_inloc_data_3_13_port);
   U142 : NOR2_X2 port map( A1 => n87, A2 => n88, ZN => 
                           internal_inloc_data_3_6_port);
   U143 : NOR2_X2 port map( A1 => n183, A2 => n184, ZN => 
                           internal_inloc_data_2_20_port);
   U144 : NOR2_X2 port map( A1 => n199, A2 => n200, ZN => 
                           internal_inloc_data_2_13_port);
   U145 : NOR2_X2 port map( A1 => n151, A2 => n152, ZN => 
                           internal_inloc_data_2_6_port);
   U146 : NOR2_X2 port map( A1 => n247, A2 => n248, ZN => 
                           internal_inloc_data_1_20_port);
   U147 : NOR2_X2 port map( A1 => n263, A2 => n264, ZN => 
                           internal_inloc_data_1_13_port);
   U148 : NOR2_X2 port map( A1 => n215, A2 => n216, ZN => 
                           internal_inloc_data_1_6_port);
   U149 : NOR2_X2 port map( A1 => n311, A2 => n312, ZN => 
                           internal_inloc_data_0_20_port);
   U150 : NOR2_X2 port map( A1 => n327, A2 => n328, ZN => 
                           internal_inloc_data_0_13_port);
   U151 : NOR2_X2 port map( A1 => n279, A2 => n280, ZN => 
                           internal_inloc_data_0_6_port);
   U152 : NOR2_X2 port map( A1 => n59, A2 => n60, ZN => 
                           internal_inloc_data_4_19_port);
   U153 : NOR2_X2 port map( A1 => n73, A2 => n74, ZN => 
                           internal_inloc_data_4_12_port);
   U154 : NOR2_X2 port map( A1 => n25, A2 => n26, ZN => 
                           internal_inloc_data_4_5_port);
   U155 : NOR2_X2 port map( A1 => n123, A2 => n124, ZN => 
                           internal_inloc_data_3_19_port);
   U156 : NOR2_X2 port map( A1 => n137, A2 => n138, ZN => 
                           internal_inloc_data_3_12_port);
   U157 : NOR2_X2 port map( A1 => n89, A2 => n90, ZN => 
                           internal_inloc_data_3_5_port);
   U158 : NOR2_X2 port map( A1 => n187, A2 => n188, ZN => 
                           internal_inloc_data_2_19_port);
   U159 : NOR2_X2 port map( A1 => n201, A2 => n202, ZN => 
                           internal_inloc_data_2_12_port);
   U160 : NOR2_X2 port map( A1 => n153, A2 => n154, ZN => 
                           internal_inloc_data_2_5_port);
   U161 : NOR2_X2 port map( A1 => n251, A2 => n252, ZN => 
                           internal_inloc_data_1_19_port);
   U162 : NOR2_X2 port map( A1 => n265, A2 => n266, ZN => 
                           internal_inloc_data_1_12_port);
   U163 : NOR2_X2 port map( A1 => n217, A2 => n218, ZN => 
                           internal_inloc_data_1_5_port);
   U164 : NOR2_X2 port map( A1 => n315, A2 => n316, ZN => 
                           internal_inloc_data_0_19_port);
   U165 : NOR2_X2 port map( A1 => n329, A2 => n330, ZN => 
                           internal_inloc_data_0_12_port);
   U166 : NOR2_X2 port map( A1 => n281, A2 => n282, ZN => 
                           internal_inloc_data_0_5_port);
   U167 : NOR2_X2 port map( A1 => n61, A2 => n62, ZN => 
                           internal_inloc_data_4_18_port);
   U168 : NOR2_X2 port map( A1 => n75, A2 => n76, ZN => 
                           internal_inloc_data_4_11_port);
   U169 : NOR2_X2 port map( A1 => n27, A2 => n28, ZN => 
                           internal_inloc_data_4_4_port);
   U170 : NOR2_X2 port map( A1 => n125, A2 => n126, ZN => 
                           internal_inloc_data_3_18_port);
   U171 : NOR2_X2 port map( A1 => n139, A2 => n140, ZN => 
                           internal_inloc_data_3_11_port);
   U172 : NOR2_X2 port map( A1 => n91, A2 => n92, ZN => 
                           internal_inloc_data_3_4_port);
   U173 : NOR2_X2 port map( A1 => n189, A2 => n190, ZN => 
                           internal_inloc_data_2_18_port);
   U174 : NOR2_X2 port map( A1 => n203, A2 => n204, ZN => 
                           internal_inloc_data_2_11_port);
   U175 : NOR2_X2 port map( A1 => n155, A2 => n156, ZN => 
                           internal_inloc_data_2_4_port);
   U176 : NOR2_X2 port map( A1 => n253, A2 => n254, ZN => 
                           internal_inloc_data_1_18_port);
   U177 : NOR2_X2 port map( A1 => n267, A2 => n268, ZN => 
                           internal_inloc_data_1_11_port);
   U178 : NOR2_X2 port map( A1 => n219, A2 => n220, ZN => 
                           internal_inloc_data_1_4_port);
   U179 : NOR2_X2 port map( A1 => n317, A2 => n318, ZN => 
                           internal_inloc_data_0_18_port);
   U180 : NOR2_X2 port map( A1 => n331, A2 => n332, ZN => 
                           internal_inloc_data_0_11_port);
   U181 : NOR2_X2 port map( A1 => n283, A2 => n284, ZN => 
                           internal_inloc_data_0_4_port);
   U182 : NOR2_X2 port map( A1 => n63, A2 => n64, ZN => 
                           internal_inloc_data_4_17_port);
   U183 : NOR2_X2 port map( A1 => n77, A2 => n78, ZN => 
                           internal_inloc_data_4_10_port);
   U184 : NOR2_X2 port map( A1 => n29, A2 => n30, ZN => 
                           internal_inloc_data_4_3_port);
   U185 : NOR2_X2 port map( A1 => n127, A2 => n128, ZN => 
                           internal_inloc_data_3_17_port);
   U186 : NOR2_X2 port map( A1 => n141, A2 => n142, ZN => 
                           internal_inloc_data_3_10_port);
   U187 : NOR2_X2 port map( A1 => n93, A2 => n94, ZN => 
                           internal_inloc_data_3_3_port);
   U188 : NOR2_X2 port map( A1 => n191, A2 => n192, ZN => 
                           internal_inloc_data_2_17_port);
   U189 : NOR2_X2 port map( A1 => n205, A2 => n206, ZN => 
                           internal_inloc_data_2_10_port);
   U190 : NOR2_X2 port map( A1 => n157, A2 => n158, ZN => 
                           internal_inloc_data_2_3_port);
   U191 : NOR2_X2 port map( A1 => n255, A2 => n256, ZN => 
                           internal_inloc_data_1_17_port);
   U192 : NOR2_X2 port map( A1 => n269, A2 => n270, ZN => 
                           internal_inloc_data_1_10_port);
   U193 : NOR2_X2 port map( A1 => n221, A2 => n222, ZN => 
                           internal_inloc_data_1_3_port);
   U194 : NOR2_X2 port map( A1 => n319, A2 => n320, ZN => 
                           internal_inloc_data_0_17_port);
   U195 : NOR2_X2 port map( A1 => n333, A2 => n334, ZN => 
                           internal_inloc_data_0_10_port);
   U196 : NOR2_X2 port map( A1 => n285, A2 => n286, ZN => 
                           internal_inloc_data_0_3_port);
   U197 : NOR2_X2 port map( A1 => n35, A2 => n36, ZN => 
                           internal_inloc_data_4_2_port);
   U198 : NOR2_X2 port map( A1 => n57, A2 => n58, ZN => 
                           internal_inloc_data_4_1_port);
   U199 : NOR2_X2 port map( A1 => n79, A2 => n80, ZN => 
                           internal_inloc_data_4_0_port);
   U200 : NOR2_X2 port map( A1 => n99, A2 => n100, ZN => 
                           internal_inloc_data_3_2_port);
   U201 : NOR2_X2 port map( A1 => n121, A2 => n122, ZN => 
                           internal_inloc_data_3_1_port);
   U202 : NOR2_X2 port map( A1 => n143, A2 => n144, ZN => 
                           internal_inloc_data_3_0_port);
   U203 : NOR2_X2 port map( A1 => n163, A2 => n164, ZN => 
                           internal_inloc_data_2_2_port);
   U204 : NOR2_X2 port map( A1 => n185, A2 => n186, ZN => 
                           internal_inloc_data_2_1_port);
   U205 : NOR2_X2 port map( A1 => n207, A2 => n208, ZN => 
                           internal_inloc_data_2_0_port);
   U206 : NOR2_X2 port map( A1 => n227, A2 => n228, ZN => 
                           internal_inloc_data_1_2_port);
   U207 : NOR2_X2 port map( A1 => n249, A2 => n250, ZN => 
                           internal_inloc_data_1_1_port);
   U208 : NOR2_X2 port map( A1 => n271, A2 => n272, ZN => 
                           internal_inloc_data_1_0_port);
   U209 : NOR2_X2 port map( A1 => n291, A2 => n292, ZN => 
                           internal_inloc_data_0_2_port);
   U210 : NOR2_X2 port map( A1 => n313, A2 => n314, ZN => 
                           internal_inloc_data_0_1_port);
   U211 : NOR2_X2 port map( A1 => n335, A2 => n336, ZN => 
                           internal_inloc_data_0_0_port);
   U212 : INV_X1 port map( A => n12, ZN => n340);
   U213 : AOI21_X1 port map( B1 => n13, B2 => RET, A => 
                           fill_address_ext_15_port, ZN => n12);
   U214 : INV_X1 port map( A => n14, ZN => n341);
   U215 : AOI21_X1 port map( B1 => n15, B2 => CALL, A => 
                           spill_address_ext_15_port, ZN => n14);
   U216 : OAI21_X1 port map( B1 => n16, B2 => n15, A => 
                           spill_address_ext_0_port, ZN => SPILL_port);
   U217 : INV_X1 port map( A => spilleq, ZN => n15);
   U218 : INV_X1 port map( A => CALL, ZN => n16);
   U219 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => n18);
   U220 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => n17);
   U221 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => n20);
   U222 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => n19);
   U223 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => n22);
   U224 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => n21);
   U225 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => n24);
   U226 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => n23);
   U227 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => n26);
   U228 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => n25);
   U229 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => n28);
   U230 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => n27);
   U231 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => n30);
   U232 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => n29);
   U233 : NAND4_X1 port map( A1 => n598, A2 => n597, A3 => n596, A4 => n595, ZN
                           => n32);
   U234 : NAND4_X1 port map( A1 => n594, A2 => n593, A3 => n592, A4 => n591, ZN
                           => n31);
   U235 : NAND4_X1 port map( A1 => n590, A2 => n589, A3 => n588, A4 => n587, ZN
                           => n34);
   U236 : NAND4_X1 port map( A1 => n586, A2 => n585, A3 => n584, A4 => n583, ZN
                           => n33);
   U237 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => n36);
   U238 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => n35);
   U239 : NAND4_X1 port map( A1 => n582, A2 => n581, A3 => n580, A4 => n579, ZN
                           => n38);
   U240 : NAND4_X1 port map( A1 => n578, A2 => n577, A3 => n576, A4 => n575, ZN
                           => n37);
   U241 : NAND4_X1 port map( A1 => n574, A2 => n573, A3 => n572, A4 => n571, ZN
                           => n40);
   U242 : NAND4_X1 port map( A1 => n570, A2 => n569, A3 => n568, A4 => n567, ZN
                           => n39);
   U243 : NAND4_X1 port map( A1 => n566, A2 => n565, A3 => n564, A4 => n563, ZN
                           => n42);
   U244 : NAND4_X1 port map( A1 => n562, A2 => n561, A3 => n560, A4 => n559, ZN
                           => n41);
   U245 : NAND4_X1 port map( A1 => n558, A2 => n557, A3 => n556, A4 => n555, ZN
                           => n44);
   U246 : NAND4_X1 port map( A1 => n554, A2 => n553, A3 => n552, A4 => n551, ZN
                           => n43);
   U247 : NAND4_X1 port map( A1 => n550, A2 => n549, A3 => n548, A4 => n547, ZN
                           => n46);
   U248 : NAND4_X1 port map( A1 => n546, A2 => n545, A3 => n544, A4 => n543, ZN
                           => n45);
   U249 : NAND4_X1 port map( A1 => n542, A2 => n541, A3 => n540, A4 => n539, ZN
                           => n48);
   U250 : NAND4_X1 port map( A1 => n538, A2 => n537, A3 => n536, A4 => n535, ZN
                           => n47);
   U251 : NAND4_X1 port map( A1 => n534, A2 => n533, A3 => n532, A4 => n531, ZN
                           => n50);
   U252 : NAND4_X1 port map( A1 => n530, A2 => n529, A3 => n528, A4 => n527, ZN
                           => n49);
   U253 : NAND4_X1 port map( A1 => n526, A2 => n525, A3 => n524, A4 => n523, ZN
                           => n52);
   U254 : NAND4_X1 port map( A1 => n522, A2 => n521, A3 => n520, A4 => n519, ZN
                           => n51);
   U255 : NAND4_X1 port map( A1 => n518, A2 => n517, A3 => n516, A4 => n515, ZN
                           => n54);
   U256 : NAND4_X1 port map( A1 => n514, A2 => n513, A3 => n512, A4 => n511, ZN
                           => n53);
   U257 : NAND4_X1 port map( A1 => n510, A2 => n509, A3 => n508, A4 => n507, ZN
                           => n56);
   U258 : NAND4_X1 port map( A1 => n506, A2 => n505, A3 => n504, A4 => n503, ZN
                           => n55);
   U259 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => n58);
   U260 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => n57);
   U261 : NAND4_X1 port map( A1 => n502, A2 => n501, A3 => n500, A4 => n499, ZN
                           => n60);
   U262 : NAND4_X1 port map( A1 => n498, A2 => n497, A3 => n496, A4 => n495, ZN
                           => n59);
   U263 : NAND4_X1 port map( A1 => n494, A2 => n493, A3 => n492, A4 => n491, ZN
                           => n62);
   U264 : NAND4_X1 port map( A1 => n490, A2 => n489, A3 => n488, A4 => n487, ZN
                           => n61);
   U265 : NAND4_X1 port map( A1 => n486, A2 => n485, A3 => n484, A4 => n483, ZN
                           => n64);
   U266 : NAND4_X1 port map( A1 => n482, A2 => n481, A3 => n480, A4 => n479, ZN
                           => n63);
   U267 : NAND4_X1 port map( A1 => n478, A2 => n477, A3 => n476, A4 => n475, ZN
                           => n66);
   U268 : NAND4_X1 port map( A1 => n474, A2 => n473, A3 => n472, A4 => n471, ZN
                           => n65);
   U269 : NAND4_X1 port map( A1 => n470, A2 => n469, A3 => n468, A4 => n467, ZN
                           => n68);
   U270 : NAND4_X1 port map( A1 => n466, A2 => n465, A3 => n464, A4 => n463, ZN
                           => n67);
   U271 : NAND4_X1 port map( A1 => n462, A2 => n461, A3 => n460, A4 => n459, ZN
                           => n70);
   U272 : NAND4_X1 port map( A1 => n458, A2 => n457, A3 => n456, A4 => n455, ZN
                           => n69);
   U273 : NAND4_X1 port map( A1 => n454, A2 => n453, A3 => n452, A4 => n451, ZN
                           => n72);
   U274 : NAND4_X1 port map( A1 => n450, A2 => n449, A3 => n448, A4 => n447, ZN
                           => n71);
   U275 : NAND4_X1 port map( A1 => n446, A2 => n445, A3 => n444, A4 => n443, ZN
                           => n74);
   U276 : NAND4_X1 port map( A1 => n442, A2 => n441, A3 => n440, A4 => n439, ZN
                           => n73);
   U277 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => n76);
   U278 : NAND4_X1 port map( A1 => n434, A2 => n433, A3 => n432, A4 => n431, ZN
                           => n75);
   U279 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => n78);
   U280 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => n77);
   U281 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => n80);
   U282 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => n79);
   U283 : NAND4_X1 port map( A1 => n678, A2 => n677, A3 => n676, A4 => n675, ZN
                           => n82);
   U284 : NAND4_X1 port map( A1 => n674, A2 => n673, A3 => n672, A4 => n671, ZN
                           => n81);
   U285 : NAND4_X1 port map( A1 => n670, A2 => n669, A3 => n668, A4 => n667, ZN
                           => n84);
   U286 : NAND4_X1 port map( A1 => n666, A2 => n665, A3 => n664, A4 => n663, ZN
                           => n83);
   U287 : NAND4_X1 port map( A1 => n662, A2 => n661, A3 => n660, A4 => n659, ZN
                           => n86);
   U288 : NAND4_X1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, ZN
                           => n85);
   U289 : NAND4_X1 port map( A1 => n654, A2 => n653, A3 => n652, A4 => n651, ZN
                           => n88);
   U290 : NAND4_X1 port map( A1 => n650, A2 => n649, A3 => n648, A4 => n647, ZN
                           => n87);
   U291 : NAND4_X1 port map( A1 => n646, A2 => n645, A3 => n644, A4 => n643, ZN
                           => n90);
   U292 : NAND4_X1 port map( A1 => n642, A2 => n641, A3 => n640, A4 => n639, ZN
                           => n89);
   U293 : NAND4_X1 port map( A1 => n638, A2 => n637, A3 => n636, A4 => n635, ZN
                           => n92);
   U294 : NAND4_X1 port map( A1 => n634, A2 => n633, A3 => n632, A4 => n631, ZN
                           => n91);
   U295 : NAND4_X1 port map( A1 => n630, A2 => n629, A3 => n628, A4 => n627, ZN
                           => n94);
   U296 : NAND4_X1 port map( A1 => n626, A2 => n625, A3 => n624, A4 => n623, ZN
                           => n93);
   U297 : NAND4_X1 port map( A1 => n854, A2 => n853, A3 => n852, A4 => n851, ZN
                           => n96);
   U298 : NAND4_X1 port map( A1 => n850, A2 => n849, A3 => n848, A4 => n847, ZN
                           => n95);
   U299 : NAND4_X1 port map( A1 => n846, A2 => n845, A3 => n844, A4 => n843, ZN
                           => n98);
   U300 : NAND4_X1 port map( A1 => n842, A2 => n841, A3 => n840, A4 => n839, ZN
                           => n97);
   U301 : NAND4_X1 port map( A1 => n622, A2 => n621, A3 => n620, A4 => n619, ZN
                           => n100);
   U302 : NAND4_X1 port map( A1 => n618, A2 => n617, A3 => n616, A4 => n615, ZN
                           => n99);
   U303 : NAND4_X1 port map( A1 => n838, A2 => n837, A3 => n836, A4 => n835, ZN
                           => n102);
   U304 : NAND4_X1 port map( A1 => n834, A2 => n833, A3 => n832, A4 => n831, ZN
                           => n101);
   U305 : NAND4_X1 port map( A1 => n830, A2 => n829, A3 => n828, A4 => n827, ZN
                           => n104);
   U306 : NAND4_X1 port map( A1 => n826, A2 => n825, A3 => n824, A4 => n823, ZN
                           => n103);
   U307 : NAND4_X1 port map( A1 => n822, A2 => n821, A3 => n820, A4 => n819, ZN
                           => n106);
   U308 : NAND4_X1 port map( A1 => n818, A2 => n817, A3 => n816, A4 => n815, ZN
                           => n105);
   U309 : NAND4_X1 port map( A1 => n814, A2 => n813, A3 => n812, A4 => n811, ZN
                           => n108);
   U310 : NAND4_X1 port map( A1 => n810, A2 => n809, A3 => n808, A4 => n807, ZN
                           => n107);
   U311 : NAND4_X1 port map( A1 => n806, A2 => n805, A3 => n804, A4 => n803, ZN
                           => n110);
   U312 : NAND4_X1 port map( A1 => n802, A2 => n801, A3 => n800, A4 => n799, ZN
                           => n109);
   U313 : NAND4_X1 port map( A1 => n798, A2 => n797, A3 => n796, A4 => n795, ZN
                           => n112);
   U314 : NAND4_X1 port map( A1 => n794, A2 => n793, A3 => n792, A4 => n791, ZN
                           => n111);
   U315 : NAND4_X1 port map( A1 => n790, A2 => n789, A3 => n788, A4 => n787, ZN
                           => n114);
   U316 : NAND4_X1 port map( A1 => n786, A2 => n785, A3 => n784, A4 => n783, ZN
                           => n113);
   U317 : NAND4_X1 port map( A1 => n782, A2 => n781, A3 => n780, A4 => n779, ZN
                           => n116);
   U318 : NAND4_X1 port map( A1 => n778, A2 => n777, A3 => n776, A4 => n775, ZN
                           => n115);
   U319 : NAND4_X1 port map( A1 => n774, A2 => n773, A3 => n772, A4 => n771, ZN
                           => n118);
   U320 : NAND4_X1 port map( A1 => n770, A2 => n769, A3 => n768, A4 => n767, ZN
                           => n117);
   U321 : NAND4_X1 port map( A1 => n766, A2 => n765, A3 => n764, A4 => n763, ZN
                           => n120);
   U322 : NAND4_X1 port map( A1 => n762, A2 => n761, A3 => n760, A4 => n759, ZN
                           => n119);
   U323 : NAND4_X1 port map( A1 => n614, A2 => n613, A3 => n612, A4 => n611, ZN
                           => n122);
   U324 : NAND4_X1 port map( A1 => n610, A2 => n609, A3 => n608, A4 => n607, ZN
                           => n121);
   U325 : NAND4_X1 port map( A1 => n758, A2 => n757, A3 => n756, A4 => n755, ZN
                           => n124);
   U326 : NAND4_X1 port map( A1 => n754, A2 => n753, A3 => n752, A4 => n751, ZN
                           => n123);
   U327 : NAND4_X1 port map( A1 => n750, A2 => n749, A3 => n748, A4 => n747, ZN
                           => n126);
   U328 : NAND4_X1 port map( A1 => n746, A2 => n745, A3 => n744, A4 => n743, ZN
                           => n125);
   U329 : NAND4_X1 port map( A1 => n742, A2 => n741, A3 => n740, A4 => n739, ZN
                           => n128);
   U330 : NAND4_X1 port map( A1 => n738, A2 => n737, A3 => n736, A4 => n735, ZN
                           => n127);
   U331 : NAND4_X1 port map( A1 => n734, A2 => n733, A3 => n732, A4 => n731, ZN
                           => n130);
   U332 : NAND4_X1 port map( A1 => n730, A2 => n729, A3 => n728, A4 => n727, ZN
                           => n129);
   U333 : NAND4_X1 port map( A1 => n726, A2 => n725, A3 => n724, A4 => n723, ZN
                           => n132);
   U334 : NAND4_X1 port map( A1 => n722, A2 => n721, A3 => n720, A4 => n719, ZN
                           => n131);
   U335 : NAND4_X1 port map( A1 => n718, A2 => n717, A3 => n716, A4 => n715, ZN
                           => n134);
   U336 : NAND4_X1 port map( A1 => n714, A2 => n713, A3 => n712, A4 => n711, ZN
                           => n133);
   U337 : NAND4_X1 port map( A1 => n710, A2 => n709, A3 => n708, A4 => n707, ZN
                           => n136);
   U338 : NAND4_X1 port map( A1 => n706, A2 => n705, A3 => n704, A4 => n703, ZN
                           => n135);
   U339 : NAND4_X1 port map( A1 => n702, A2 => n701, A3 => n700, A4 => n699, ZN
                           => n138);
   U340 : NAND4_X1 port map( A1 => n698, A2 => n697, A3 => n696, A4 => n695, ZN
                           => n137);
   U341 : NAND4_X1 port map( A1 => n694, A2 => n693, A3 => n692, A4 => n691, ZN
                           => n140);
   U342 : NAND4_X1 port map( A1 => n690, A2 => n689, A3 => n688, A4 => n687, ZN
                           => n139);
   U343 : NAND4_X1 port map( A1 => n686, A2 => n685, A3 => n684, A4 => n683, ZN
                           => n142);
   U344 : NAND4_X1 port map( A1 => n682, A2 => n681, A3 => n680, A4 => n679, ZN
                           => n141);
   U345 : NAND4_X1 port map( A1 => n606, A2 => n605, A3 => n604, A4 => n603, ZN
                           => n144);
   U346 : NAND4_X1 port map( A1 => n602, A2 => n601, A3 => n600, A4 => n599, ZN
                           => n143);
   U347 : NAND4_X1 port map( A1 => n934, A2 => n933, A3 => n932, A4 => n931, ZN
                           => n146);
   U348 : NAND4_X1 port map( A1 => n930, A2 => n929, A3 => n928, A4 => n927, ZN
                           => n145);
   U349 : NAND4_X1 port map( A1 => n926, A2 => n925, A3 => n924, A4 => n923, ZN
                           => n148);
   U350 : NAND4_X1 port map( A1 => n922, A2 => n921, A3 => n920, A4 => n919, ZN
                           => n147);
   U351 : NAND4_X1 port map( A1 => n918, A2 => n917, A3 => n916, A4 => n915, ZN
                           => n150);
   U352 : NAND4_X1 port map( A1 => n914, A2 => n913, A3 => n912, A4 => n911, ZN
                           => n149);
   U353 : NAND4_X1 port map( A1 => n910, A2 => n909, A3 => n908, A4 => n907, ZN
                           => n152);
   U354 : NAND4_X1 port map( A1 => n906, A2 => n905, A3 => n904, A4 => n903, ZN
                           => n151);
   U355 : NAND4_X1 port map( A1 => n902, A2 => n901, A3 => n900, A4 => n899, ZN
                           => n154);
   U356 : NAND4_X1 port map( A1 => n898, A2 => n897, A3 => n896, A4 => n895, ZN
                           => n153);
   U357 : NAND4_X1 port map( A1 => n894, A2 => n893, A3 => n892, A4 => n891, ZN
                           => n156);
   U358 : NAND4_X1 port map( A1 => n890, A2 => n889, A3 => n888, A4 => n887, ZN
                           => n155);
   U359 : NAND4_X1 port map( A1 => n886, A2 => n885, A3 => n884, A4 => n883, ZN
                           => n158);
   U360 : NAND4_X1 port map( A1 => n882, A2 => n881, A3 => n880, A4 => n879, ZN
                           => n157);
   U361 : NAND4_X1 port map( A1 => n1110, A2 => n1109, A3 => n1108, A4 => n1107
                           , ZN => n160);
   U362 : NAND4_X1 port map( A1 => n1106, A2 => n1105, A3 => n1104, A4 => n1103
                           , ZN => n159);
   U363 : NAND4_X1 port map( A1 => n1102, A2 => n1101, A3 => n1100, A4 => n1099
                           , ZN => n162);
   U364 : NAND4_X1 port map( A1 => n1098, A2 => n1097, A3 => n1096, A4 => n1095
                           , ZN => n161);
   U365 : NAND4_X1 port map( A1 => n878, A2 => n877, A3 => n876, A4 => n875, ZN
                           => n164);
   U366 : NAND4_X1 port map( A1 => n874, A2 => n873, A3 => n872, A4 => n871, ZN
                           => n163);
   U367 : NAND4_X1 port map( A1 => n1094, A2 => n1093, A3 => n1092, A4 => n1091
                           , ZN => n166);
   U368 : NAND4_X1 port map( A1 => n1090, A2 => n1089, A3 => n1088, A4 => n1087
                           , ZN => n165);
   U369 : NAND4_X1 port map( A1 => n1086, A2 => n1085, A3 => n1084, A4 => n1083
                           , ZN => n168);
   U370 : NAND4_X1 port map( A1 => n1082, A2 => n1081, A3 => n1080, A4 => n1079
                           , ZN => n167);
   U371 : NAND4_X1 port map( A1 => n1078, A2 => n1077, A3 => n1076, A4 => n1075
                           , ZN => n170);
   U372 : NAND4_X1 port map( A1 => n1074, A2 => n1073, A3 => n1072, A4 => n1071
                           , ZN => n169);
   U373 : NAND4_X1 port map( A1 => n1070, A2 => n1069, A3 => n1068, A4 => n1067
                           , ZN => n172);
   U374 : NAND4_X1 port map( A1 => n1066, A2 => n1065, A3 => n1064, A4 => n1063
                           , ZN => n171);
   U375 : NAND4_X1 port map( A1 => n1062, A2 => n1061, A3 => n1060, A4 => n1059
                           , ZN => n174);
   U376 : NAND4_X1 port map( A1 => n1058, A2 => n1057, A3 => n1056, A4 => n1055
                           , ZN => n173);
   U377 : NAND4_X1 port map( A1 => n1054, A2 => n1053, A3 => n1052, A4 => n1051
                           , ZN => n176);
   U378 : NAND4_X1 port map( A1 => n1050, A2 => n1049, A3 => n1048, A4 => n1047
                           , ZN => n175);
   U379 : NAND4_X1 port map( A1 => n1046, A2 => n1045, A3 => n1044, A4 => n1043
                           , ZN => n178);
   U380 : NAND4_X1 port map( A1 => n1042, A2 => n1041, A3 => n1040, A4 => n1039
                           , ZN => n177);
   U381 : NAND4_X1 port map( A1 => n1038, A2 => n1037, A3 => n1036, A4 => n1035
                           , ZN => n180);
   U382 : NAND4_X1 port map( A1 => n1034, A2 => n1033, A3 => n1032, A4 => n1031
                           , ZN => n179);
   U383 : NAND4_X1 port map( A1 => n1030, A2 => n1029, A3 => n1028, A4 => n1027
                           , ZN => n182);
   U384 : NAND4_X1 port map( A1 => n1026, A2 => n1025, A3 => n1024, A4 => n1023
                           , ZN => n181);
   U385 : NAND4_X1 port map( A1 => n1022, A2 => n1021, A3 => n1020, A4 => n1019
                           , ZN => n184);
   U386 : NAND4_X1 port map( A1 => n1018, A2 => n1017, A3 => n1016, A4 => n1015
                           , ZN => n183);
   U387 : NAND4_X1 port map( A1 => n870, A2 => n869, A3 => n868, A4 => n867, ZN
                           => n186);
   U388 : NAND4_X1 port map( A1 => n866, A2 => n865, A3 => n864, A4 => n863, ZN
                           => n185);
   U389 : NAND4_X1 port map( A1 => n1014, A2 => n1013, A3 => n1012, A4 => n1011
                           , ZN => n188);
   U390 : NAND4_X1 port map( A1 => n1010, A2 => n1009, A3 => n1008, A4 => n1007
                           , ZN => n187);
   U391 : NAND4_X1 port map( A1 => n1006, A2 => n1005, A3 => n1004, A4 => n1003
                           , ZN => n190);
   U392 : NAND4_X1 port map( A1 => n1002, A2 => n1001, A3 => n1000, A4 => n999,
                           ZN => n189);
   U393 : NAND4_X1 port map( A1 => n998, A2 => n997, A3 => n996, A4 => n995, ZN
                           => n192);
   U394 : NAND4_X1 port map( A1 => n994, A2 => n993, A3 => n992, A4 => n991, ZN
                           => n191);
   U395 : NAND4_X1 port map( A1 => n990, A2 => n989, A3 => n988, A4 => n987, ZN
                           => n194);
   U396 : NAND4_X1 port map( A1 => n986, A2 => n985, A3 => n984, A4 => n983, ZN
                           => n193);
   U397 : NAND4_X1 port map( A1 => n982, A2 => n981, A3 => n980, A4 => n979, ZN
                           => n196);
   U398 : NAND4_X1 port map( A1 => n978, A2 => n977, A3 => n976, A4 => n975, ZN
                           => n195);
   U399 : NAND4_X1 port map( A1 => n974, A2 => n973, A3 => n972, A4 => n971, ZN
                           => n198);
   U400 : NAND4_X1 port map( A1 => n970, A2 => n969, A3 => n968, A4 => n967, ZN
                           => n197);
   U401 : NAND4_X1 port map( A1 => n966, A2 => n965, A3 => n964, A4 => n963, ZN
                           => n200);
   U402 : NAND4_X1 port map( A1 => n962, A2 => n961, A3 => n960, A4 => n959, ZN
                           => n199);
   U403 : NAND4_X1 port map( A1 => n958, A2 => n957, A3 => n956, A4 => n955, ZN
                           => n202);
   U404 : NAND4_X1 port map( A1 => n954, A2 => n953, A3 => n952, A4 => n951, ZN
                           => n201);
   U405 : NAND4_X1 port map( A1 => n950, A2 => n949, A3 => n948, A4 => n947, ZN
                           => n204);
   U406 : NAND4_X1 port map( A1 => n946, A2 => n945, A3 => n944, A4 => n943, ZN
                           => n203);
   U407 : NAND4_X1 port map( A1 => n942, A2 => n941, A3 => n940, A4 => n939, ZN
                           => n206);
   U408 : NAND4_X1 port map( A1 => n938, A2 => n937, A3 => n936, A4 => n935, ZN
                           => n205);
   U409 : NAND4_X1 port map( A1 => n862, A2 => n861, A3 => n860, A4 => n859, ZN
                           => n208);
   U410 : NAND4_X1 port map( A1 => n858, A2 => n857, A3 => n856, A4 => n855, ZN
                           => n207);
   U411 : NAND4_X1 port map( A1 => n1190, A2 => n1189, A3 => n1188, A4 => n1187
                           , ZN => n210);
   U412 : NAND4_X1 port map( A1 => n1186, A2 => n1185, A3 => n1184, A4 => n1183
                           , ZN => n209);
   U413 : NAND4_X1 port map( A1 => n1182, A2 => n1181, A3 => n1180, A4 => n1179
                           , ZN => n212);
   U414 : NAND4_X1 port map( A1 => n1178, A2 => n1177, A3 => n1176, A4 => n1175
                           , ZN => n211);
   U415 : NAND4_X1 port map( A1 => n1174, A2 => n1173, A3 => n1172, A4 => n1171
                           , ZN => n214);
   U416 : NAND4_X1 port map( A1 => n1170, A2 => n1169, A3 => n1168, A4 => n1167
                           , ZN => n213);
   U417 : NAND4_X1 port map( A1 => n1166, A2 => n1165, A3 => n1164, A4 => n1163
                           , ZN => n216);
   U418 : NAND4_X1 port map( A1 => n1162, A2 => n1161, A3 => n1160, A4 => n1159
                           , ZN => n215);
   U419 : NAND4_X1 port map( A1 => n1158, A2 => n1157, A3 => n1156, A4 => n1155
                           , ZN => n218);
   U420 : NAND4_X1 port map( A1 => n1154, A2 => n1153, A3 => n1152, A4 => n1151
                           , ZN => n217);
   U421 : NAND4_X1 port map( A1 => n1150, A2 => n1149, A3 => n1148, A4 => n1147
                           , ZN => n220);
   U422 : NAND4_X1 port map( A1 => n1146, A2 => n1145, A3 => n1144, A4 => n1143
                           , ZN => n219);
   U423 : NAND4_X1 port map( A1 => n1142, A2 => n1141, A3 => n1140, A4 => n1139
                           , ZN => n222);
   U424 : NAND4_X1 port map( A1 => n1138, A2 => n1137, A3 => n1136, A4 => n1135
                           , ZN => n221);
   U425 : NAND4_X1 port map( A1 => n1366, A2 => n1365, A3 => n1364, A4 => n1363
                           , ZN => n224);
   U426 : NAND4_X1 port map( A1 => n1362, A2 => n1361, A3 => n1360, A4 => n1359
                           , ZN => n223);
   U427 : NAND4_X1 port map( A1 => n1358, A2 => n1357, A3 => n1356, A4 => n1355
                           , ZN => n226);
   U428 : NAND4_X1 port map( A1 => n1354, A2 => n1353, A3 => n1352, A4 => n1351
                           , ZN => n225);
   U429 : NAND4_X1 port map( A1 => n1134, A2 => n1133, A3 => n1132, A4 => n1131
                           , ZN => n228);
   U430 : NAND4_X1 port map( A1 => n1130, A2 => n1129, A3 => n1128, A4 => n1127
                           , ZN => n227);
   U431 : NAND4_X1 port map( A1 => n1350, A2 => n1349, A3 => n1348, A4 => n1347
                           , ZN => n230);
   U432 : NAND4_X1 port map( A1 => n1346, A2 => n1345, A3 => n1344, A4 => n1343
                           , ZN => n229);
   U433 : NAND4_X1 port map( A1 => n1342, A2 => n1341, A3 => n1340, A4 => n1339
                           , ZN => n232);
   U434 : NAND4_X1 port map( A1 => n1338, A2 => n1337, A3 => n1336, A4 => n1335
                           , ZN => n231);
   U435 : NAND4_X1 port map( A1 => n1334, A2 => n1333, A3 => n1332, A4 => n1331
                           , ZN => n234);
   U436 : NAND4_X1 port map( A1 => n1330, A2 => n1329, A3 => n1328, A4 => n1327
                           , ZN => n233);
   U437 : NAND4_X1 port map( A1 => n1326, A2 => n1325, A3 => n1324, A4 => n1323
                           , ZN => n236);
   U438 : NAND4_X1 port map( A1 => n1322, A2 => n1321, A3 => n1320, A4 => n1319
                           , ZN => n235);
   U439 : NAND4_X1 port map( A1 => n1318, A2 => n1317, A3 => n1316, A4 => n1315
                           , ZN => n238);
   U440 : NAND4_X1 port map( A1 => n1314, A2 => n1313, A3 => n1312, A4 => n1311
                           , ZN => n237);
   U441 : NAND4_X1 port map( A1 => n1310, A2 => n1309, A3 => n1308, A4 => n1307
                           , ZN => n240);
   U442 : NAND4_X1 port map( A1 => n1306, A2 => n1305, A3 => n1304, A4 => n1303
                           , ZN => n239);
   U443 : NAND4_X1 port map( A1 => n1302, A2 => n1301, A3 => n1300, A4 => n1299
                           , ZN => n242);
   U444 : NAND4_X1 port map( A1 => n1298, A2 => n1297, A3 => n1296, A4 => n1295
                           , ZN => n241);
   U445 : NAND4_X1 port map( A1 => n1294, A2 => n1293, A3 => n1292, A4 => n1291
                           , ZN => n244);
   U446 : NAND4_X1 port map( A1 => n1290, A2 => n1289, A3 => n1288, A4 => n1287
                           , ZN => n243);
   U447 : NAND4_X1 port map( A1 => n1286, A2 => n1285, A3 => n1284, A4 => n1283
                           , ZN => n246);
   U448 : NAND4_X1 port map( A1 => n1282, A2 => n1281, A3 => n1280, A4 => n1279
                           , ZN => n245);
   U449 : NAND4_X1 port map( A1 => n1278, A2 => n1277, A3 => n1276, A4 => n1275
                           , ZN => n248);
   U450 : NAND4_X1 port map( A1 => n1274, A2 => n1273, A3 => n1272, A4 => n1271
                           , ZN => n247);
   U451 : NAND4_X1 port map( A1 => n1126, A2 => n1125, A3 => n1124, A4 => n1123
                           , ZN => n250);
   U452 : NAND4_X1 port map( A1 => n1122, A2 => n1121, A3 => n1120, A4 => n1119
                           , ZN => n249);
   U453 : NAND4_X1 port map( A1 => n1270, A2 => n1269, A3 => n1268, A4 => n1267
                           , ZN => n252);
   U454 : NAND4_X1 port map( A1 => n1266, A2 => n1265, A3 => n1264, A4 => n1263
                           , ZN => n251);
   U455 : NAND4_X1 port map( A1 => n1262, A2 => n1261, A3 => n1260, A4 => n1259
                           , ZN => n254);
   U456 : NAND4_X1 port map( A1 => n1258, A2 => n1257, A3 => n1256, A4 => n1255
                           , ZN => n253);
   U457 : NAND4_X1 port map( A1 => n1254, A2 => n1253, A3 => n1252, A4 => n1251
                           , ZN => n256);
   U458 : NAND4_X1 port map( A1 => n1250, A2 => n1249, A3 => n1248, A4 => n1247
                           , ZN => n255);
   U459 : NAND4_X1 port map( A1 => n1246, A2 => n1245, A3 => n1244, A4 => n1243
                           , ZN => n258);
   U460 : NAND4_X1 port map( A1 => n1242, A2 => n1241, A3 => n1240, A4 => n1239
                           , ZN => n257);
   U461 : NAND4_X1 port map( A1 => n1238, A2 => n1237, A3 => n1236, A4 => n1235
                           , ZN => n260);
   U462 : NAND4_X1 port map( A1 => n1234, A2 => n1233, A3 => n1232, A4 => n1231
                           , ZN => n259);
   U463 : NAND4_X1 port map( A1 => n1230, A2 => n1229, A3 => n1228, A4 => n1227
                           , ZN => n262);
   U464 : NAND4_X1 port map( A1 => n1226, A2 => n1225, A3 => n1224, A4 => n1223
                           , ZN => n261);
   U465 : NAND4_X1 port map( A1 => n1222, A2 => n1221, A3 => n1220, A4 => n1219
                           , ZN => n264);
   U466 : NAND4_X1 port map( A1 => n1218, A2 => n1217, A3 => n1216, A4 => n1215
                           , ZN => n263);
   U467 : NAND4_X1 port map( A1 => n1214, A2 => n1213, A3 => n1212, A4 => n1211
                           , ZN => n266);
   U468 : NAND4_X1 port map( A1 => n1210, A2 => n1209, A3 => n1208, A4 => n1207
                           , ZN => n265);
   U469 : NAND4_X1 port map( A1 => n1206, A2 => n1205, A3 => n1204, A4 => n1203
                           , ZN => n268);
   U470 : NAND4_X1 port map( A1 => n1202, A2 => n1201, A3 => n1200, A4 => n1199
                           , ZN => n267);
   U471 : NAND4_X1 port map( A1 => n1198, A2 => n1197, A3 => n1196, A4 => n1195
                           , ZN => n270);
   U472 : NAND4_X1 port map( A1 => n1194, A2 => n1193, A3 => n1192, A4 => n1191
                           , ZN => n269);
   U473 : NAND4_X1 port map( A1 => n1118, A2 => n1117, A3 => n1116, A4 => n1115
                           , ZN => n272);
   U474 : NAND4_X1 port map( A1 => n1114, A2 => n1113, A3 => n1112, A4 => n1111
                           , ZN => n271);
   U475 : NAND4_X1 port map( A1 => n1446, A2 => n1445, A3 => n1444, A4 => n1443
                           , ZN => n274);
   U476 : NAND4_X1 port map( A1 => n1442, A2 => n1441, A3 => n1440, A4 => n1439
                           , ZN => n273);
   U477 : NAND4_X1 port map( A1 => n1438, A2 => n1437, A3 => n1436, A4 => n1435
                           , ZN => n276);
   U478 : NAND4_X1 port map( A1 => n1434, A2 => n1433, A3 => n1432, A4 => n1431
                           , ZN => n275);
   U479 : NAND4_X1 port map( A1 => n1430, A2 => n1429, A3 => n1428, A4 => n1427
                           , ZN => n278);
   U480 : NAND4_X1 port map( A1 => n1426, A2 => n1425, A3 => n1424, A4 => n1423
                           , ZN => n277);
   U481 : NAND4_X1 port map( A1 => n1422, A2 => n1421, A3 => n1420, A4 => n1419
                           , ZN => n280);
   U482 : NAND4_X1 port map( A1 => n1418, A2 => n1417, A3 => n1416, A4 => n1415
                           , ZN => n279);
   U483 : NAND4_X1 port map( A1 => n1414, A2 => n1413, A3 => n1412, A4 => n1411
                           , ZN => n282);
   U484 : NAND4_X1 port map( A1 => n1410, A2 => n1409, A3 => n1408, A4 => n1407
                           , ZN => n281);
   U485 : NAND4_X1 port map( A1 => n1406, A2 => n1405, A3 => n1404, A4 => n1403
                           , ZN => n284);
   U486 : NAND4_X1 port map( A1 => n1402, A2 => n1401, A3 => n1400, A4 => n1399
                           , ZN => n283);
   U487 : NAND4_X1 port map( A1 => n1398, A2 => n1397, A3 => n1396, A4 => n1395
                           , ZN => n286);
   U488 : NAND4_X1 port map( A1 => n1394, A2 => n1393, A3 => n1392, A4 => n1391
                           , ZN => n285);
   U489 : NAND4_X1 port map( A1 => n1622, A2 => n1621, A3 => n1620, A4 => n1619
                           , ZN => n288);
   U490 : NAND4_X1 port map( A1 => n1618, A2 => n1617, A3 => n1616, A4 => n1615
                           , ZN => n287);
   U491 : NAND4_X1 port map( A1 => n1614, A2 => n1613, A3 => n1612, A4 => n1611
                           , ZN => n290);
   U492 : NAND4_X1 port map( A1 => n1610, A2 => n1609, A3 => n1608, A4 => n1607
                           , ZN => n289);
   U493 : NAND4_X1 port map( A1 => n1390, A2 => n1389, A3 => n1388, A4 => n1387
                           , ZN => n292);
   U494 : NAND4_X1 port map( A1 => n1386, A2 => n1385, A3 => n1384, A4 => n1383
                           , ZN => n291);
   U495 : NAND4_X1 port map( A1 => n1606, A2 => n1605, A3 => n1604, A4 => n1603
                           , ZN => n294);
   U496 : NAND4_X1 port map( A1 => n1602, A2 => n1601, A3 => n1600, A4 => n1599
                           , ZN => n293);
   U497 : NAND4_X1 port map( A1 => n1598, A2 => n1597, A3 => n1596, A4 => n1595
                           , ZN => n296);
   U498 : NAND4_X1 port map( A1 => n1594, A2 => n1593, A3 => n1592, A4 => n1591
                           , ZN => n295);
   U499 : NAND4_X1 port map( A1 => n1590, A2 => n1589, A3 => n1588, A4 => n1587
                           , ZN => n298);
   U500 : NAND4_X1 port map( A1 => n1586, A2 => n1585, A3 => n1584, A4 => n1583
                           , ZN => n297);
   U501 : NAND4_X1 port map( A1 => n1582, A2 => n1581, A3 => n1580, A4 => n1579
                           , ZN => n300);
   U502 : NAND4_X1 port map( A1 => n1578, A2 => n1577, A3 => n1576, A4 => n1575
                           , ZN => n299);
   U503 : NAND4_X1 port map( A1 => n1574, A2 => n1573, A3 => n1572, A4 => n1571
                           , ZN => n302);
   U504 : NAND4_X1 port map( A1 => n1570, A2 => n1569, A3 => n1568, A4 => n1567
                           , ZN => n301);
   U505 : NAND4_X1 port map( A1 => n1566, A2 => n1565, A3 => n1564, A4 => n1563
                           , ZN => n304);
   U506 : NAND4_X1 port map( A1 => n1562, A2 => n1561, A3 => n1560, A4 => n1559
                           , ZN => n303);
   U507 : NAND4_X1 port map( A1 => n1558, A2 => n1557, A3 => n1556, A4 => n1555
                           , ZN => n306);
   U508 : NAND4_X1 port map( A1 => n1554, A2 => n1553, A3 => n1552, A4 => n1551
                           , ZN => n305);
   U509 : NAND4_X1 port map( A1 => n1550, A2 => n1549, A3 => n1548, A4 => n1547
                           , ZN => n308);
   U510 : NAND4_X1 port map( A1 => n1546, A2 => n1545, A3 => n1544, A4 => n1543
                           , ZN => n307);
   U511 : NAND4_X1 port map( A1 => n1542, A2 => n1541, A3 => n1540, A4 => n1539
                           , ZN => n310);
   U512 : NAND4_X1 port map( A1 => n1538, A2 => n1537, A3 => n1536, A4 => n1535
                           , ZN => n309);
   U513 : NAND4_X1 port map( A1 => n1534, A2 => n1533, A3 => n1532, A4 => n1531
                           , ZN => n312);
   U514 : NAND4_X1 port map( A1 => n1530, A2 => n1529, A3 => n1528, A4 => n1527
                           , ZN => n311);
   U515 : NAND4_X1 port map( A1 => n1382, A2 => n1381, A3 => n1380, A4 => n1379
                           , ZN => n314);
   U516 : NAND4_X1 port map( A1 => n1378, A2 => n1377, A3 => n1376, A4 => n1375
                           , ZN => n313);
   U517 : NAND4_X1 port map( A1 => n1526, A2 => n1525, A3 => n1524, A4 => n1523
                           , ZN => n316);
   U518 : NAND4_X1 port map( A1 => n1522, A2 => n1521, A3 => n1520, A4 => n1519
                           , ZN => n315);
   U519 : NAND4_X1 port map( A1 => n1518, A2 => n1517, A3 => n1516, A4 => n1515
                           , ZN => n318);
   U520 : NAND4_X1 port map( A1 => n1514, A2 => n1513, A3 => n1512, A4 => n1511
                           , ZN => n317);
   U521 : NAND4_X1 port map( A1 => n1510, A2 => n1509, A3 => n1508, A4 => n1507
                           , ZN => n320);
   U522 : NAND4_X1 port map( A1 => n1506, A2 => n1505, A3 => n1504, A4 => n1503
                           , ZN => n319);
   U523 : NAND4_X1 port map( A1 => n1502, A2 => n1501, A3 => n1500, A4 => n1499
                           , ZN => n322);
   U524 : NAND4_X1 port map( A1 => n1498, A2 => n1497, A3 => n1496, A4 => n1495
                           , ZN => n321);
   U525 : NAND4_X1 port map( A1 => n1494, A2 => n1493, A3 => n1492, A4 => n1491
                           , ZN => n324);
   U526 : NAND4_X1 port map( A1 => n1490, A2 => n1489, A3 => n1488, A4 => n1487
                           , ZN => n323);
   U527 : NAND4_X1 port map( A1 => n1486, A2 => n1485, A3 => n1484, A4 => n1483
                           , ZN => n326);
   U528 : NAND4_X1 port map( A1 => n1482, A2 => n1481, A3 => n1480, A4 => n1479
                           , ZN => n325);
   U529 : NAND4_X1 port map( A1 => n1478, A2 => n1477, A3 => n1476, A4 => n1475
                           , ZN => n328);
   U530 : NAND4_X1 port map( A1 => n1474, A2 => n1473, A3 => n1472, A4 => n1471
                           , ZN => n327);
   U531 : NAND4_X1 port map( A1 => n1470, A2 => n1469, A3 => n1468, A4 => n1467
                           , ZN => n330);
   U532 : NAND4_X1 port map( A1 => n1466, A2 => n1465, A3 => n1464, A4 => n1463
                           , ZN => n329);
   U533 : NAND4_X1 port map( A1 => n1462, A2 => n1461, A3 => n1460, A4 => n1459
                           , ZN => n332);
   U534 : NAND4_X1 port map( A1 => n1458, A2 => n1457, A3 => n1456, A4 => n1455
                           , ZN => n331);
   U535 : NAND4_X1 port map( A1 => n1454, A2 => n1453, A3 => n1452, A4 => n1451
                           , ZN => n334);
   U536 : NAND4_X1 port map( A1 => n1450, A2 => n1449, A3 => n1448, A4 => n1447
                           , ZN => n333);
   U537 : NAND4_X1 port map( A1 => n1374, A2 => n1373, A3 => n1372, A4 => n1371
                           , ZN => n336);
   U538 : NAND4_X1 port map( A1 => n1370, A2 => n1369, A3 => n1368, A4 => n1367
                           , ZN => n335);
   U539 : AND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => int_RD2);
   U540 : AND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => int_RD1);
   U541 : AND2_X1 port map( A1 => dec_output_9_port, A2 => n337, ZN => 
                           dec_out_with_wen_9_port);
   U542 : AND2_X1 port map( A1 => dec_output_8_port, A2 => n337, ZN => 
                           dec_out_with_wen_8_port);
   U543 : AND2_X1 port map( A1 => dec_output_7_port, A2 => n337, ZN => 
                           dec_out_with_wen_7_port);
   U544 : AND2_X1 port map( A1 => dec_output_6_port, A2 => n337, ZN => 
                           dec_out_with_wen_6_port);
   U545 : AND2_X1 port map( A1 => dec_output_5_port, A2 => n337, ZN => 
                           dec_out_with_wen_5_port);
   U546 : AND2_X1 port map( A1 => dec_output_4_port, A2 => n337, ZN => 
                           dec_out_with_wen_4_port);
   U547 : AND2_X1 port map( A1 => dec_output_3_port, A2 => n337, ZN => 
                           dec_out_with_wen_3_port);
   U548 : AND2_X1 port map( A1 => dec_output_31_port, A2 => n337, ZN => 
                           dec_out_with_wen_31_port);
   U549 : AND2_X1 port map( A1 => dec_output_30_port, A2 => n337, ZN => 
                           dec_out_with_wen_30_port);
   U550 : AND2_X1 port map( A1 => dec_output_2_port, A2 => n337, ZN => 
                           dec_out_with_wen_2_port);
   U551 : AND2_X1 port map( A1 => dec_output_29_port, A2 => n337, ZN => 
                           dec_out_with_wen_29_port);
   U552 : AND2_X1 port map( A1 => dec_output_28_port, A2 => n337, ZN => 
                           dec_out_with_wen_28_port);
   U553 : AND2_X1 port map( A1 => dec_output_27_port, A2 => n337, ZN => 
                           dec_out_with_wen_27_port);
   U554 : AND2_X1 port map( A1 => dec_output_26_port, A2 => n337, ZN => 
                           dec_out_with_wen_26_port);
   U555 : AND2_X1 port map( A1 => dec_output_25_port, A2 => n337, ZN => 
                           dec_out_with_wen_25_port);
   U556 : AND2_X1 port map( A1 => dec_output_24_port, A2 => n337, ZN => 
                           dec_out_with_wen_24_port);
   U557 : AND2_X1 port map( A1 => dec_output_23_port, A2 => n337, ZN => 
                           dec_out_with_wen_23_port);
   U558 : AND2_X1 port map( A1 => dec_output_22_port, A2 => n337, ZN => 
                           dec_out_with_wen_22_port);
   U559 : AND2_X1 port map( A1 => dec_output_21_port, A2 => n337, ZN => 
                           dec_out_with_wen_21_port);
   U560 : AND2_X1 port map( A1 => dec_output_20_port, A2 => n337, ZN => 
                           dec_out_with_wen_20_port);
   U561 : AND2_X1 port map( A1 => dec_output_1_port, A2 => n337, ZN => 
                           dec_out_with_wen_1_port);
   U562 : AND2_X1 port map( A1 => dec_output_19_port, A2 => n337, ZN => 
                           dec_out_with_wen_19_port);
   U563 : AND2_X1 port map( A1 => dec_output_18_port, A2 => n337, ZN => 
                           dec_out_with_wen_18_port);
   U564 : AND2_X1 port map( A1 => dec_output_17_port, A2 => n337, ZN => 
                           dec_out_with_wen_17_port);
   U565 : AND2_X1 port map( A1 => dec_output_16_port, A2 => n337, ZN => 
                           dec_out_with_wen_16_port);
   U566 : AND2_X1 port map( A1 => dec_output_15_port, A2 => n337, ZN => 
                           dec_out_with_wen_15_port);
   U567 : AND2_X1 port map( A1 => dec_output_14_port, A2 => n337, ZN => 
                           dec_out_with_wen_14_port);
   U568 : AND2_X1 port map( A1 => dec_output_13_port, A2 => n337, ZN => 
                           dec_out_with_wen_13_port);
   U569 : AND2_X1 port map( A1 => dec_output_12_port, A2 => n337, ZN => 
                           dec_out_with_wen_12_port);
   U570 : AND2_X1 port map( A1 => dec_output_11_port, A2 => n337, ZN => 
                           dec_out_with_wen_11_port);
   U571 : AND2_X1 port map( A1 => dec_output_10_port, A2 => n337, ZN => 
                           dec_out_with_wen_10_port);
   U572 : AND2_X1 port map( A1 => dec_output_0_port, A2 => n337, ZN => 
                           dec_out_with_wen_0_port);
   U573 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n337);
   U574 : AND2_X1 port map( A1 => c_swin_0_port, A2 => FILL_port, ZN => 
                           c_swin_masked_1bit_4_0_port);
   U575 : AND2_X1 port map( A1 => c_swin_4_port, A2 => FILL_port, ZN => 
                           c_swin_masked_1bit_3_0_port);
   U576 : AND2_X1 port map( A1 => c_swin_3_port, A2 => FILL_port, ZN => 
                           c_swin_masked_1bit_2_0_port);
   U577 : AND2_X1 port map( A1 => c_swin_2_port, A2 => FILL_port, ZN => 
                           c_swin_masked_1bit_1_0_port);
   U578 : AND2_X1 port map( A1 => c_swin_1_port, A2 => FILL_port, ZN => 
                           c_swin_masked_1bit_0_0_port);
   U579 : OAI21_X1 port map( B1 => n338, B2 => n13, A => 
                           fill_address_ext_0_port, ZN => FILL_port);
   U580 : INV_X1 port map( A => filleq, ZN => n13);
   U581 : INV_X1 port map( A => RET, ZN => n338);

end SYN_mix;
